-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
TKKoLN1qdRKFrJVMhU/GhY49huWWv5YhI9K3i5Cxhrc3SMMbHtoag9m24fI6F1Mg
enx+LET/0hYfHO+e6kG3FMhhDeWU0rAC2tPySBLxuy41qh0oNLjgjyYdsDch5dZS
Dq6Bd6e/WxmP04ECXMM2am7sNjJEdhGrJa83G3qfKwU=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 11535)

`protect DATA_BLOCK
uF2/xHskxjw9eEPN8XuFbdSbB70YhdaYw54z3dY0kPQvJzDvuLRtxYkq24Z+klDy
2dKlxtoUVIs6tud7X92rfDAXQUBkSu2cMj7MR9X1GFpDJXIKhJn7NOnYBVYDSuGg
jGbVsXY1YGhNcb9i99dshbaRO/EDTLRa1l5RQc1wvjwnZHkpQexgPGuHvYjbwHi7
zwRsow0stQUpQAKWYRtF5bdaKAEjy/N3TK8L5atLJsOkyZ6fS+tvWzIwxf+UdNNZ
WnPKWgzSREmr4LlWkEKmHplA8Z6PDx7qHxJ7YXuYcn2qnI2vHZCt7XQ/4F86C4Tw
UOvex9v/y4lf5Bl3wHYs97hdexmqOIOXfFthHjQngbbFn6onenESiXZxroHj5Rm9
gsKyWQqjIjncfIH3rvJrDM5TmRbuCTdoxQEzC27YYQLMh0p3o9WgAT91Nzr3bZQY
qyhZgirk5e4Da51S72SFtCjNbshbXJLmn6tadJiHI9hX6N2sKk4Pt3T/KMXw+W4w
RqKZrRdKZR9HlBkbYSUCmPzrLlhPNQHX0TinTTKr1ScZOjyk90vPkx3jKi/xt7wb
pyx9l8r2jTmoB1R2/TvL3VlDD/p6rmfCFbhz2mfXrdkgGPaDLYImpgjvaDJPSRSi
nFec+NTR80ORUt4wnghziaD/g0CbmHYG9x6BALT25lx9uLwjpS7HXN+zsEpZsCeA
o+OhrOWcpAGh/U8XEHnnAIbK9irWGE4vLT89bHjiqO/V/OQDwtGTLfI00dVbSCFn
BcncLt7C0i2532rHTRzjB9KrAwPTS6W/nH8GJ17tql0cpvri9Jh+ctTfHBbF5p2T
gLlcEXsAZM0sagEN61Kib9H/ZD6B27ESYldl12sRFNabcvJLLiNiFXSTuQj/1WJg
d39y9qDzqbJLpcuUxfQ5BLRwdttAMFEwgVyRHY1mtT6aeZtzKYF9pzOYNmcMXUsu
HZP9ZNZaC8Cqp+eU43ZrcnK6Ih2jDewxy/FmMe8kfueFfvHMjgdu1Ttj8jyim2OX
FDxCLOwwDllteQ31bCOtG0j8sxndVKpwEpg7D2EKaIr/lo1s1O8lUm9sCCFJ5gjF
WRcqj1dRshwkoTlh7NwTxJD2jUq0KhoPQagNlgSli47J5k3TpuOFwYGON5ttsLCx
96z3Iqcrlf/BIJnzprojk/pFO6+Ak80n0wsbmZewSWA3O1hRARKMhUw1x6SCM6Me
fwGS2FrE0JiusFbsUYl5fNRchQ+M2Y21x0knZSMmFtW6FYxqHHE7KAzEPDIK61cF
2PS7cBoUiQ1B0M7Y8hcJjcIACyztdgPu3dQGBNQkOIROU9pt+r6Nfcop+TT+juLD
jN+sLimgjewIA5xvs3NKwo+tmidLMYSXIPLWCeYGKUPPIFSQfvO9lczL6NKHYz93
k08ng6Y0quL+ECMZKhBge4Y8GODibvyTY9wwVtYWfjAadobF2WPsqcgBbAcPrEcx
nDJzG4opiRf3io18FYwSG4388XvhM2fUF0Mr5dlueaLjuQu5h68i3QoVyx1CxZV1
RXhOxWxWPiKjRml5DeuyCPfVoc5itorbiFerVXqER61Y5YohA1HizHQnyrRVsXcb
NAYP+FBTkJnbdhQdWXwdzpYQZq27QYWH8baVbDsKUVuSz8G2i8AOJ1SkLR5CY0RO
S4tJQE0MfHLvqIczsa36EOp0akuuMWc1N1B30VSyxAWMXlp/jfRDf1xgdhk61v8+
WLj7XzMx9KGyVucSukzwMKyTEUVVkUkeqQWnUEvetZ+9o7OPqR06gFbxzaPcRiBI
/89RHnmFD9dLY+O+FS69hVWLIhJflI/a+NQqfQ+9p8VHK5L9C75PT/rUMUg/rjt6
bTJ0IC/gWsFtJ+YwnPh+UZmfbi9Swd3Gut5mRzBdp+aHPTddlsy/65NQZJa5XfBM
WaFf4jzsc3rlGSPvGXJDUFgAzhEiCEaufvDI3GRP6N53/j+VaJ0wtHzyt+UvDLVs
kmm3Oi3iA5l0r1EG65KchmPL1E0i+5lrVv5Ii7XHSpZDgk07OuXDFv4klOb3CZXx
9+Zs5hDMQn4dMxhtGlaev+HrnwssuYynvoyFoiTKg5+JTLlu/4x25bwBoJVBBk7r
rluzSXO++ksu/nEL2DZnQoIGHVw4/fJV48Gt3ccLPpq5izDkzfjqRhdMx5MModiu
r94SSy+4l6wfuPQ1lvYA6H055eHVyxwITZK34So3teyU6O7avMyEliTe/YDHhb76
CoOUXBAQwrZJxSSg51fRu4gTsAzKOzTV2DFg9EqXJYVYYbshcMk0/vdpBOIlKyn6
pLOJl4W+VkR5rVAvV9rBSIiABr/V9yyViDO/25Be6LL5LKahHhES6ROVPd8Kmc8+
5BqBD4FXC3gY8f9E1yo1/dZv8Ov95f4FElqmOAdsQxUlwSU9UvIPY2E6xShb+lhp
hcMuDTFCmZjRX0HwsZSArNok+aJAQgAVCH6pA93hPYEiIwXPhmS19S/hCuk2m0Nd
Vhe54Q6Dg2Gi9+wkZKSyw6E8FHbf6AR2wZJ2bzMvCXslZnfgwVC6CYk7z4LCpNRP
/ofSVZQX4YrAndppIwnzAIt+NjdOXq7ODJZ3Pxy+lFNAUeJ/IVDzgBAtdspLQMnS
TYbVsXJZvE4lILLbliLO8snCqgakrRXlg8PcSIeGu1tEWtCPnWAXWkqq9RhvOxFO
DFoGoCqP6nwlR7zFAUY+bmWpCtOaToDn3PXGTjjRB2+OLM0aG6MFlDGp5CF7F1to
Z4dq+2AOaSmMLi8+VlS4BRSdP1gcVR3kTnwY1f/r4A0vUVaqBsRAoyoK3mtg8Oy9
2IQXJaaoun//Aq6QkHKcBwo5mbT3mG4LrtbpBEk1/8JXOyq8BS3Bq/5B2o50don9
xo01haZa+buuAV0dTPvM5G2xEejfn902mHOmPDVc5kl4ip0x+94OcnL6L3OPQE7c
7igdWNlaTGgl3KSy/Hfhbn1KKUPBF6rpadEO070q/YR3vfy25kB5Y91Br9OB4vRY
3pvk+S1eGs1B2d1pCkamGgkuSldy9u1dWU2VVGTa0N3YErNwXELyfG6V7hTRtl41
U2fJB5fw76j5YjPuRAJ3OmmJ3OckcfHqzBqEQmpphplFc2j+YvQLqW5LVNakawtf
6Wl0/9+YnwH096hYqR3igCSFCAY7arBzPc0GcLCWppdOTjjLVkUaL0BY/JtmEfo7
SUpxVUQKrX01VPD4qJnHgx5SoJ+PVuPoCF1wkAYSoRDWJpKqtj1LbCt/neNrDBDE
d7Sesf0wCl8fkZGcd+ELe8L6NS/6GimcQblzfR00A98tereHLvX/8owAnKY3LKDJ
/zazilam1IAAMe2H9WfHhVnbt7JWLEobBVr/AEDHgMhdcygBvutelpek4vS4vX5W
4qrmrl8oJ2E7gZZWxedjIyWwh53O5XxhUUszxBEe3DZepZEGJJC6sfVGL0kZi3b0
GgCaL+no9e8Zcvkl/b5nvHtae9ivoM7WpdNnzz8D5SZ+Ox1McCB0yT71a0bjfqH4
ECJ/vxkAdZGfVlnvVT1lUhNIQLfD2Xq9mnxiuhZ5Mb21/Ds1b4dQyiDsCim7qS08
JZdNrm3XS/P5U2v5wuray68iF5qJihG8pfiyZF1+5U44mg2vxvZeruCpSRvvd6JQ
FSiPftYpN74aq2SR9BsBJkXRskOhPmwajQHcn7GnOyDcMIF+Z92x8R7YFkV6lPJ7
7CSH8pKfWBQ/3mf72JdbXNHk3GqTywxM6hW0JDgdyAJXqwzCbNX4SXh8sJnG6ISO
s3MebNLIVyK/09vI4scijj4WAs0ayGrAloR73ku9tQJFVJDbjdBixhytpppXWnfy
w5dDxtWtJq5caFygaqhLBM8WahY2a+vJV2q5CssjyNb+WKeckV2wSL53Pa1VXjP7
DTSpGxgE0dDv1U4+B8mCA3BkCL4rPs7cU9xJlhpF4dxBWBD8EVcyAVbo0P9TjOZ/
K9BOze9LAdigUcLYL3+mPS7GkZarqKzKcDHaJkq1/kgIaz4fakhR3YE3zx2mlqLW
3O8RxYSbOyyex7KTYn5OX0kz72zmvhZbeSbjp961KH4hAz4z3ksQcVfm6R+ZWHIL
hz0oiGxv1vSC9XhDKAYOiKvjskUgGfHbtjinYFKBFRGXz2IiIn2y7qlMGBCOB306
/Hpvjtt4RuHCQyymIV+szTWb2uWf78j+PhBs0ngWrkRiuJJXwup4PuPmiUIIu3ie
WSq+zC6DUm6Z5YMyb+0DfHyUErA4lTfDdZUg/J69a/tk2NZGmhAEdPtKnGoCxtFW
51yNSJzdIHqcIZXGrLvKGJbPVsVAC+OLru3SjeqZA8miipqdx2U9w2rN3a+UNpUN
LYnhtZAW8yjAwpc3MNEEKahoenM7eEAgVpXnjGTX/bMnll+GlW+2HLl5+yDmH30H
O/VklLrdg5DlRF8VOwd22O789tTThqy5AV1JcsGnmzVgYkY/3V0i/42T/QVs1Q1k
1VQoBo3t3RFC8GxU0C5cvdD2EWV3YmtwZfRmLuKDLA1lGQf12VmwgNEQ0dIkC7ne
TzpfbyZalXFaaFEZusJSF1eg370TowWZLG9isEzdT4h6dYHhA3cFaekNADb/Dqqo
ECu2zNRyMd80FW4Pmi3A2JFbWY/59qkLWgRzdrLNtZwIMWJLcVNoypysnEIpTeVx
a+Qt9nWH/0Zo3aDR3mrwYxzCwBAIOS7f9+/DNa1pXi+VDivK+jwZm8pqsgsNiUFP
jdndOQg5RlRhA+et1PAjWurqZnABBWBV7ic/t5/h6GNp/0W3uAl3wHXlpbbnWXUi
Uj41LsecWEI3x4cNB+bsleHlCAo6BTwQECSU/zzncygdD0m9dsNcMFPlVvxTBIKf
ewUrCtFy8APxR2cfe45mnWNDavAlBKiZuI0AtOnx2f4m+VVyHypOxKbvCYJU5rbs
78DTVc850flbAsgxa675oMFMxXwrjp0OERY2DbGcWbf+GJV3wv4pP/Ijq5XnTMJy
v24AyggpkzUqSKAMZzkQ/2TQGPUIU8/I/pKXfbP9p3t8c31Q4UUi+im3FQCKrY4J
YrEmoOwlu8gsWrA2yKYyCvQxNVw7jVZguxS2yMvHbKcPmtJpgfjXKwmjIBOyQ8BT
gPPJR8gVtbU11JREve4KbVTzVWsOjGo7p4LVpq6nveEw3kJbRDQWTU7qPNNBG0+W
ZPBpYjnUTvSTQ+XCxhPp8fO6DLWo61Te0ub+ChSwsgflz7fjIJ76grLjQBQ38/PT
UaparoBa5EB4FGl5JGewuXuYS9C4nLuV38zaBXpeouXx5Y7Xez1dkSh6PMcMGMHt
vv20/MyiH0gZbVf9BsxHvLUpVvTlKIWKKWl1MSCOwVUPwg5PlQDS+UmZRXqjfjCK
WF6n/7ailZjc62efEBJNCRxfDZZiY0fGgtGBGNaM1/Ayx0A7MFX15BPEdNcyRaNd
dIjP20r4KcmSXCni1/AD0ztUn5EEUJRyqWBMokJzbOanilI3Pjpgw8eHvf3t4nAu
bBDfrN3+BrXCY/dS9ta0LUkBrMw5poqotC9rw6aldrcciruWbNf2xV1gkTuEyZXh
qEkkeG4q3eyPFtAPt5Twr9Df4oeuOP3kxWmW6SsOdSbdiaZptn3v4R99O+Lbx3H6
EBJjEvL+rZhAaG5tzZrsfebbWK8c05sF/P50toU/tL/XNVSQtcAlLIEKcVkm9RLt
xTUP7gzduQX9eK6m65rEL7hvMao6fmK2UCyH3IS2SBGRkzh0gqzmAL56ZNfes1ic
R6J1GO4cbKTT7WkkxGL3RVaQJmq1T5UFdTmuWeR6AsYt5LKZsvTMQHRqUq0tbnWl
Ump+JoLza63xEePSzujj6gx/yWVIArDPvkx7oFrk168WkUbHu3gV4km0ZVtAsPVB
Zp39JxMrwh778+xqDEFeBDuCzhiUrDTjIf4nr5qvE9KvK7rzoUxXLCMkXHI62cmo
KM/jp9UqAuobX9Oeqo/my4SN6JZoVXMm9RBZrsXZAY0dmy25QxZGnx/cLOBvFx0I
4bpttuZXc8bbleTLH9an6Osb3Vn5FoEg8V39+mz+/BxO6xREpjPJt9J/njZKrc9O
WkqNuiYAkwlYGpFLNE5PsdqmkPmr9OSQ7w1Uj4TRwckBIZ/3qQONMDz3TSzMehRt
fX1oen3iR5QOokNaeB4ab4ugKTq3qmRWUy3FrN7/IhpMs/GDuajUgI//PRgcFhDd
CLwFu0/PN8fMEsEKzHr3VIG7d9RYpsffkwnOysSCay3anH4vxubG2NK3qChrSQ22
tLGR/LE9EMjD5LHe+tAep+1gq4kr+uKvEw1JnBcMiYNdHLohL82suoztHaTJdMJ7
MelGFNPDd8vbahh5TzfuIV2uBGXkDuxfGoctQOT8I5VyNiQS3FRq3cp2MI+tBkuu
E+ylQ6TqfucvqDQ6LTiplEGhHJhfcIrf+bQqqPGBK/gwkvMuTpp6hlsrrt8xaqce
xClRlSJpojd5rxFVCemDiDHkKKjaX+y7vuguITHEaY32DZJkcoPU5QYhE8qP5v2s
wK6mS/a3Z4xpGUINAsMfjo3NooiaD3mVJwSojwh0q42PB3jaYSOYw0++wIPeQmwr
xqtqoq4h1nL5WM3/iKZAlEa6eH1VXBL5bOXdPABI5AFHAgBZFis0hel20GnNAyO9
F+xKZBfrEUXf6LamEutA6Y0Qq7W86o/+paXqiPmBszf8FI//7zvnUpjCH1wLxPAi
wwwESuoas5WJxaREWLAN/MbrJXJPdo+rbJWXMk2+RKYZJacBzPa61zxVpJXTxRcw
udMGgrHyDASyn7VKr/hRWQq4HPO0f4C26tpABfnBSW64GrTrMYzMavnDuNEakMyJ
lZVs2JAO3N/OShyet+VJ5xt+v7w5sMQlFoNoC/l/D4X8sBRS/4bp8u3MHTMYw0dI
pctNMg91AejMLc8XNHrtJFPDpZKHLGxKcxNCwmgWn3c6aN7oYexr4FjKpg/F26DF
7rGFEroddSj/0nJfr5WyyjMtQ3huEGAFg7R6KBKaol+6Imvue5M3XP9WMR3szHKt
w8tj6gyEHVd+1Ni2HG3pVRev1DXhDFLgApTmz+jT1432pSKaUXJBSdxFzfOQnvgD
SW9cxnclkKlo4TtFCWQD0Rg2xK52gUW2uNZ0pSYNcaVj+S7PIEKz2FWzOIDNrhpB
oUm+VD//mWkh/J07kcdm2P/fLpkYMwy6RLULWk736vJ+IVcJVh7q1PqkLDNlMQCl
rtYunYPQfO/UJtZiK5BiwyoivpgPLYLhU9iq29mzYVt7PkIH/qipTk8LbeExS3Cy
p6mUGurDDXtKO/0eZ3s/DN7ruLH5yQD4WsTOwDum+kAUuyv5l9LgzP9rlO2f2l1J
I/e4oNo902EJbM9dg1a2Zr8+xoUVLv2+6n//FSDZmWANi9I8Ux04uW/seKsBqb8S
5qqQHeIoNDNvHJ5QwdlMGuC7cn/iivo3OB0iVk9vbRgYXdaSANdpdJPs7FWGyUXB
5IhdXNaZ5+JGmuOeLmNQ52AbrRxsREduXA/h9t2CTengUJ0Vhyic5Pw3+T5ZQNJA
vr88svDahFOOreMAQlYmh6prN4Q1KBaew646zgkWDlZoz0CGMWrnbLcBDe8p4NNL
YyzFATdAbVrpaOvpnqc+nF2tQIcOXArYiZ7+YnLjefJcvZg4vslHExFJb0/Tf8Je
bXfG755Q2goCHZ3gRe3KGCaRHdfdaZoPdgHde7W4jhSob8plO9j5NpvVNYpi57kE
KdMBQJRTH1ArvbmcbWGltPk3QFrUnckD60TOqN2xmA2/JGj9PldhDlnd4huNIKq2
FMWTAz3fRdBut+crJWIZwyKPSHvudch/2es20DgD95S9WgSmjvS4Cc6bH5PLuzVx
w4X/7YwHue6GOzlchoVdlSBjMuy74GqLAejj503V1NGO2M85F8IDUxL6XhLCZuBh
C2wpjBeKEk33+mq1FUNnWSzfpqdlKm6whr1ruG75b6MLF9gU0yqK5JIpGraFNGup
1uD3ojz9gnt1lBZqy0JIvmpHdmv8MbNyD/ozbx9NNotkTNz0ZoUcGYdnQGAqc9rO
Q2FLbsgAK4CM/8ANdMuuvlB3yDf0ZITmtrYFjoJuSXF8WkqyNmHg5Ndw8vBLjyR8
hdSs0UQ4GQx5keGOAyRdsxCV/7dAzU7I15UEWguQno9KX+fY/KA0lZp/cPBSpFjx
9EzJLnJOJ2YC9ofCzC6ba2oWSXbGZ1f2tJcDywbHB9+PrLQhW8peKBUz0ZfXE8bJ
A9j79oQ7D5dhbbOd8QN3aMZ840OAvh47zj8pLux/1UZWX/pJqCDYFBSd14h8cXgs
YHUvbvT/PpgRattknQHp+3KOsRW8Ychrv7SPLb8sbYVjP7yX97grha70QzT1rNfH
oWyB0G1P+LvOvKqScI6vEj1R3Ew/HYsEMiUj0WDrLfVGGZJ1FdxAueuCHdthXs+B
OVM41DFzELfMeV/DevkYWrHvwGBumMp5siE6I8FPg3/uRH+RN9C6tFtshp71/opI
o7vgKWuk4eEr4/rVuvE0p2g/PTmw8oI1N5/3fBjS16ENcWU+ftZ1esnaz251KsYL
HJus7HE1NkQsIOQ+XRQ8hTK3irlaC05nAHyk3RmG1Y6f8ngiuHsie2YY2zXXonmk
hC2klN5+gEbgRIcK3c0lbC4XoI7c2kx7/qMbvpaY/YDDRShik4KXDVSXxGBgviJs
c6//dL1cqFxKFSZznRgOqT2FCoPTvEJrft9oJDppKTGeL23xNvI5EnpJk4FawEe/
qc39TR7hTo5w6KdyJQJo+4vUZpAnF9uKNXVq9OJ5I1F3JEBpOkjugohjSnNkbwnz
3pKcWYI2R/k3D4igSh+CgjhIQYouu+AZ6eoAq1rF0tB5bzJhwFq16S8BW6O/hp5U
wWsUBNJkN/hcaIAoysWgcNTAF3AT6XauJrBOVo5i99Y+0wiIQ8/qxnB+Q8f6poDZ
y45+IAhMNwF7E+l8G8NkTuKDhcdvhBry1rCU45HP/i4BoNCG+6FSGdhbEmJE7jL1
AYVTPWOofjlD6A2HDUj6PdCtoqBfq7bhz+BQzLKJNl+D7oGf8zVLG3Ol6B/urerZ
wf8IV+7ShA/YwGefZS5rfPuj4plzuLTRsHtIKkNSLSaK80b3j9p9TvnH7btiW/Ii
xzCnmasBRBSLkik0NhiGbQTZnaZbFGaIMCOFAKUv+4lKBRHz2rpGGvGOXhkwdGgt
XLP4VSyja/zLHJjsIn2ELEYQHnD7MpgiPnu0BXbRTiMibwI+auKI9ESo+T5ypMMV
oSgaOhZ8oseRlX70yuY/hslVKf1xGbG9g+/EY6V7xlle7gsg0BInKK1UZA4t7Uqo
KpMRFMJbkNGKRJltcGm4QtguAfPqd68Vu4FhUEhbToTxk8vEetm5SqkFQ9hgg7cG
yBrTPRo+OA2Nj3klW5We7FF/O6gfRHGRzDu6KNXjSss1IVXYjKSVXE+86MUfjk5a
HxlHQv1eiGBXw+C0vtzOHoCOSIMAYhSwffNwzYsZ/B4CVtXWPQfYV0XLOLv2z3OI
W1yagEFBEUHbDoKSwwn8PGiB79+PjaN/iTHYhuKfTTCd9f4zPXDhbe7ipDvnJyg/
J+c6dmBstGMIwAsuSYDZZ7z6VsuZBbAKJvScvIqCRrTdzYM89s2QK7AkAb1xM83l
GL+HUUwsBN/t7nRnE2y9klUcDmWQv8cNZPIWWafj066C9fMOYz82xSvSFHEq4eZI
8Zlm9kLAxLymRLcqm2mB3R5tTu3SiiY4ddglBdjkXxqyfEed4Qzpj4U3fQJf7b5X
OxKmKlAmiaOUDcYjvelkT4wc5RmnLeez54irUTgo+gNX5BlslDcb2pV2IgZwbuS7
UEsyQRpZ2vvyKV6idqklHi507xwGv+LGpwcez0mWNoAcytiVIE2DsuMCK55brTab
KQydS0+wnZ9ttlYRfNpbyiAfvi/2SMKHXSBXIzGInGUiCAMdCEYxIVTZotvmPdX1
Oql/roHD3bKvFyTRNtP5xCCuqqUry8fx0j4ro3lBy4ZRbeNTWk3T0ud5qVadbYX9
WCnoyq4D6iNOxamosXo01vxckurM5bnHxyTd3ewoh5Yub1jBxmkD10C2cxh9ZY7t
Nl5RvMDDEcaDUy6dm6Lihiedav7TPbjA9XdTwXCI2dOQzsSxQR9iKTeglTaMCQ7v
AdwXxUSWBP+9gB8+Un4J3g1DnSSKSGvX8b2rVQ4/TQ/pbhGN4HKkU3rUjschKP/y
TgWSv7b53i9vZkjgR/kagY/hFLCIS4J0nC1Wi5c8xVy/H74dTcn53R+t4921R+1t
TPs6RsxM/jPdl5vKW7JF/BO1MQvsomrI/7IQoGLjtIHANtJeF0w9keMpx9BEk6e7
dyXKyH6yzXavIWxgfTR4+zuPhSrm5w7K9jvzig2TBQwmgMjA7titG62nb+dVew65
5+Jx7VIqE2R2RTCO5ruhJd/gx4fLqK7EIgBPAU1CdXaxWn9Bb6b+yDDXMJ57JJyh
We5v1P5r/9cSd3cDMU2D3Buu+gO1JbJLXnxLTtqw5EUL4g9rF/rApuAk0wcYcHu/
Bk3dnlNTnGRn1F/VRqnoMiAO2dM36Mdfvqin0PJxl1tJ7t2wWj8V3yZL5iuSqTB9
QxcG6sGVJZNdwZKYQa5deztjXAgmV1cpEtbzi7/wFLugZuqjmO1NSt+cBg6p5Sat
XRr4fUMirVwutJ0xWNtRrTdbTRtu7bY+DTKoLCB1D9vWiQ/PZoJezN2mEQ46yRLv
XLvVBLO+ER4Kr10Su9FgQXahyquwF0IBVcckgAnNO82JFyB80UKZ9P2vBBOcmzHw
rRNDrzUEV3xa9sYRgyd1RXKL3qvkkOAGaKRSO5o2xZqLa2A0rfNCdrthQl+J5CXo
9TkTzDg7YMvAJglqUP62+t7Vr4QMXYHe9N84WjTQg40lLjhW3lWti8gGKdWR1l8K
1hjNC9tzhTBqtrUj8nRZZlHvYBqwsUeYZdi3pW9eTRdeAXANy38lDzuShsQ4WtJs
V7DnoynDRCUCwXacAgtk4mvZj1kEfQXJrtHxg+iQjf5WJxluJK16XQ0b/StWMZuT
A3xgMDnNdtNHfNERS4RqE6pRu8RFxzfqdlXPimKZl+aIcELXDHPjXKIQ0k8lAFwe
/8tVOing+ZXNgHmr8P+jDsnhYMO/i+4T3gnHX0dkTdJPyuCrnf2za6ajF3Mpu6N5
/F42M1yA4b7hLPQKyjv32np/LFafvEPNh0/I1UKYAepnMoaEHIFpMaAskQzycjCl
H5I9Sht9Cdvg32lplfc1XO9m7H0Tp+cjO2wEZoViXDz9CtO54us7iv7AxQO8ia2d
ng8+lEi20IPJKh90ZHmUMLSUVfj/mspJgxEXjfmQPanytTcUEbBDDAfsvfS4MnWA
Ue+p407h/UQz6qfQZHd5z0kekL8yBq2Gr+oCJ5LdSYvhWrxQTljurzv90djC+5TN
3KVwR58hvot8M3kO9YgTbLztEn7NBFEFGpzZhO18HUA3u3z6LrXOQczrBXUc9foA
p27U66vwHCg09Myy+Slaj2ppfK4fz5SKoovLh+a/IqagAjZi/DYPDhhG7VSPE36t
Cf6NovzBGRrglDACE/eG6FgsGBeULIWy01PJDN/Zr/q1+LS17tQ4WO5+EI1VwHPj
/Wl5kPk/Yx1OMYPc49NT19939CnFsJ6w1JdxO9oJ3az9wnsA8GVESH38GzDHBDSM
Fkj7581/OKOKzgDrMhHAF24JM2TTNQi9NCSBEz40wAElumBYDrasrcrKXWhohCab
HDnsyTeM/IWZ1/moSmTlBhH062Ft/SDrXq8hBYfg6LzhTTLtu9wv8i+60Y1kkmBM
JO6cyEoW1k0OmLiAOOokfpFkkdOnszp5ho+c158DLCV+s7OmgHDu0X0g+g1YEy1E
tnVLRqHDkt7Zq6Snm3Cx5ry0+m2dozp+gOa5Y9tjA/iB1pn91m12ueJ0iIw7NvXz
7875bmGKE7C2e2PYqT+p5ygIuygUzaOChYRaeNQ7nfq31f6fPQpC09wW9CkV/Gg1
8P3Qmp9AdfvFz5KnxwUf6TA+ZVg9Guaj/splweiywVFrm8q7A0kvfcbr1JOG9Nxf
xCgkWxoUngv3RTQpVDGgAC47SycCgJLlz+/MuOJbeUlJA3FUId4Yo32JsUvzkLhd
X2/iEBCZ6ww83D9wYcOJg8ekUQSFiXQeLMOHoo01cuytwNNaPHxJ4TLqVxm5MIOs
pbOyvUJoaD6uqbtxemIhTAl/8sIpWOx7osTpcn5w5i1HcfHr7zb/yFPTxXCyEv9+
Q7G4CXfWWhZh+Vyv3ZQ3TOIP2qRqM91+9bCAB0BmJ3L/ZHR3kzkKHIrqjvVYTepq
Foev45n2so9z42vScfrh1OYSRQnBwD/8/TjxhiarRSnifiN1CGCiNcLldhNhBZLu
CzPngLqCA+VRjMN3K5TXiBwryyaLsQqoXRoTOUpBoOGBK7TFlCD1/XcHgCv2Lcx1
tKrZTFEMrSD2ztJ93/w5Ca3S3f//ysxBoYTQ3qE9a9CcaMbwLn6rnEpXFQKMHBZe
7d0GKbNqsxoh/p5y3GCfu34iBdNF6Qwn4WS8223LXda5XfOyc46hZAroHajq8uKS
CB81dorVeRt4vwVYhYLEfJQBZFkXmV3jH5tMWoI5lVRVRai6XnAnErcJ+dYC8T4+
wWvPCTBU6unuO3ILGJg4Al0hR2LqI2BBHap5xLTs7JxSNaddTQeh3Z23eSbU5oq7
uRhVJhe6b1YJg8A0m2WDb8Iu037cOOWkq0rlCyTd+4uJ4WVa9PUcneUfPQ6RXccF
LvxRIt1C7Z7rDQ1gxA7C/tMgPk1u2wHeG1BZKubX6TGs39m2Ev1TD41dlDN4lH1n
lnzJ2YwG3SiuyyQ24OwTv0hDm74Z7URSaZcRMhJfjtR+LRHVVtQ2p1yxyFHOo+un
L6wa9Z107YPWhOW/cMoUS2CBKwGjSxn+HfrOp3Wh6KHKOuPzidqi5vp+5XjkQHMG
LaGFcPY1yZlK/DOl65yY+dW/7737G63vQpCxXMWGSRpO4NTRDro8olDOuyyoX3R6
ObiXYPpcMJeNS3be6yYft63bkcHh/LA/lcYFMa6Zvp4o6qOJx4q+pFpGDIM4LqCL
ti56nGwjiLJferd+/ED/gdRf/r8J/tBYtGPmcy9S4v4KD/+IBFOa5HIDG9XeriQW
dDDS5tNCvFeO8hhXdGKsEaMz8mY4l00lN91jTCEi9e6ymeFArNp/CFKfNMLQwI9D
r0Qk2jP0IJRgvN9817FXyx9oms2GyPUwpeRQDjYAq1krLSiqzxNgACByuC3N5h1I
LMReMu/zWAwO87Ds3WPsR6gSt4CKlKSRNIX4uI7XjA5ZTnoMbqiwEihFw5an1yVI
XTyathL/UmUHekg7RaaIGl49/DWbPmnRruyNhPvlwHDJLU30UzwKKQP4PsH8ip1s
xlrB8tqAtO5SpA3Hr+vJxLHUyjiyld4B/tUkR632h9m0D1oS0Aal2fkgCxbhmlYa
OFs9rfCnmVX/nm+Dlf7fPE3wWNFMHjRG2P4oy4MTxdDCi5Ii4YIr2MdvcGgqsJN4
2RTqm5A08hToegEqAAAV8n3hn6lp3Df33LinaZatP6Tg0wFwBb0fFXavmqwRSiQn
jE4kOToIyjjc3HW4RFr0YoPYj8eLMemFNj/tS11X4pMJxGKq23KlpRur5d2wwOwU
AriU29cqBQ5om8eKS0MgtbMbzUUXTGYu0Dl7nqYyomAIp6w/1u8PfgXgv22Qm23c
Z+I/nF/XBWWH1g00D3/8bXNxDvpp3Q+f0JUC/lWEFoi9ApoTdEH569qyQlkwccJ2
TimR+wMZbpe0MYJTNul3/G1dE3o5VtLPPHpkz3IXuTrIuvlxE2GlEWfifgioVI2P
t1NYcHI/Yzw1hA2BBMBcYazgXVWhbgKbveAQz00Y29QPPIuZ1YA8vD98MvfYyVPE
zvumh9OlrfSNo6scGjKoHERlx+gGR0iEdV3yyq9D6Dft6hwiX/LpF3IOb3voP8WE
XKTAHa4aU9/oTlDjB48C3PmUYkcPuk1HDLcDdMXb9kAjLkZ0N5on68XQLd5NNJcl
53C3Gmjf8Z85zwDh9zYLyJQs7jSn/NhGCMJVg/NScxDN0QmgNjn/TWjK0SfckhRm
VtYuPEKG2U2DhrLZ0HUMwU45LLzbobzwWecIxyFljGCeICh82d3FEYxAmip81+d8
51tDei/votkqcUII7UKsNWekYXnUOy4QGXNKNEje+rVWAgkole2N+7Pl/sc37coU
m3et4S8KDO39yNbqcedouIy0AJnUdDe3Y/0XiWgJjAQJGQdv2934+hhO7VEfWGJ8
XaXAmrLaHNcObi8j7G2Lce1R0JTKXiX4vmZqsYldP0zs0CqP26o7vgFfS5DGSPQX
GKk6epszrgqFxwifCOjdF8K4ZsJuFw7za9T2RSnby9I7tNjMtZ1f6SjAT0ukgq4W
uzra80dlOlKF+lDSsRE6CmBgv/oGuQpiie+v4Xec/P5eu3U7tTpCa22Oy8zD0UcM
GzlGhx53NdvvBpBWBVJpBTLQzL1i8AhUa+u+AtJu0kO/005F7sG12Qdbo2TvTtxO
2841EXEOJp3rVVvE9MDegeFpXCMcB5xxOBumnZ1LK0jlGaJlG7NpjcbjSfbNpAfn
ctyTELb4n7PY1HFuN7fTJnT9rW/1pAOem9wf28yOwTY03G8ygzvEuNFT8JCwRext
ntCXW9/HIGA/9kMhyKXFfk3ZcLk1BRDLJhYRUJLkFohBlZnLZB1n9T4OpgQaO9QF
aqgzr5xeNgYkTPDqxjGjWERR/wUnm5W0IB0Q819uLsj22HKcBtbtcLUjPbsEHe9z
C+XHZ7qEKQj9vSnTQUk3+6XTaGPIssFw9KUPUp+9I0sPS5McWfR6LzWnQtNo8tCb
34auX6y95Eco7B1oIRsX59j98Ds+KXNd1FBN6YrYXPS5MfuItLpm94HWhg3FfAXF
NnLKPsaXXUTowH5bA+3g3s/Z9C9wHraBQSl+aaSr03ZoGjElvPo92wS5J/8DG38y
XoKqE34mFjco4yAa6bi8Xo8aGF7CxhnWGnPAdvKQHsWwYgrODYtT4lMvj/aUTUa4
e7bA+lpmoMzTx6soyEWdNobt/LcwGCr8QHMmOdDpW4cDVQsCExYamW9JbVcQ3J6V
jeB9g1l2w9d+dI79l76y35bGR6oH9eItBcn9I6pOrbovaBtjvd0fjI002WPj8LGn
2TQess3OMCLL3wEupwmBRnWzmAE3mwDsygCMIMILgb8ro1gFx6vg+gY5mLJ+sy5h
/S6L87eXAxrACISZkgeDC+X+doidJ3feOVKw6Z1vmEH2IxogDrmQ+XENGQeHM3XQ
agr9FGNF1g0Kmgx5vW+1pgmqBw3WAiESbSruM/1LNz4=
`protect END_PROTECTED