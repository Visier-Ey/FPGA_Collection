��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F����Z4��#����m�ǵp��}��a��1��qh8��ɞq�t�m$��?�Y�¤.��i̓X�☾�}ד�^
*4FFx��:�o�""�k@�n�H�����s����F #ʨ���~\��-X�����[��Mm-;>�B0U�s�Z|;�N��I)4�][8x;�Ȇ]�i�?�@%+�"q���#\֢���
�3���ۻ�έԲ���L�y����tV��fw٭P�NKQ��7m�k�|��/���+�,��h	��#}ǂ�	;\=���W�j��"`!	"��N�s�$�'��z�X��̝J���+)|�7c ��t2M@Jw�[�)Q��A�R��p�������
��O��>é�}I*�7A1X�;�X�hk��tb���]�"oG��]j�4<�^�`�5���S �.]d��E�������Ym%��7��	�<�5�G��{Iu�~��a�e�z�Q�/��;P�0�F��{�"�7��,��ړ-	
ُ�k�>&.2�f�%$p��4�V ��]ͱ?~��т-��˴��&ͬ1,q5�L�l��jR�"h�����R��Z���P�a�F�E��A��7���w�+�'���O���3�K�j:7�Gl�f�&���$�����6��nhr?���/B�]q�NO6a����#Fwu�*i'�Q���-á_p�F��{���H�|���a���~%�� Kf���+���ke+
��4�1���]�OO.�� #ʺ�^���~��[f� ���5�l�4k�J��v0�o�(m�2�� ���1�-�;��Y�njT�k��-jL�T�T�����Ӽ�����y�>�%�F��`�G�z�ߍ��xuo�Bw��|��;�hR�b���w�-8}�9J�����G��B{�ܺnw�����j� ��u7&�����Y���|��&���:��D�E��-G��Or���j��޻��Oe8��t����s��� �pnVW:WrS"����!9��!����

�M��Ë�NE�~�:��u� ��\Bf����9��\���`>�Ȧ����Ns��D� ����Lv.}���	`]���O5��t�`��0���� l.x�I�T�?�wu�k�!��+O�f3Co����4$�|����|�Gul�C�xu��V����N00�C BO��\=aQam=�M\%�Ř����	�|$���(�gB����'��&��-�e���h^���JܡH��i`]��j���rR5��U�L��iE����rS1zu����b�#.1�IK��o�j��: ���{�^YÙr�:p��J�3aI,��D�I���3�M��
(��c�艓��
Mʧ�S�� ���m��	M��������:e�RK!�c7���ˇm���^�SP?G�H�-{������y�֏�Pb
"���� q��;C��k��}�����/	=-��T�O&��Q"���G�d�J�+���@�
G.4� �n���}{W���}�P��:i���R"�Er�.��`�����#��~�S�&1�ŅeF^�	�e3f���:���K��E�$O.��w���'�R�i�VMO�Qg��İyƂƇ�9*��hE�@҉�ru�RD����?�'�o�,vQJ9�G����I=�T��!6��ڣ�U�ӻ���-���j�Б�Q�`�S'���^A��Esc��c��ۅ�~gz'I6�wl� ^��	\(@������̃@B%���5
W��x�U{8-��`�E'��`�Z�7�����z7J��I)ԩo9�gP�	���3��t�'
v����~��/�ٍ]tŏWPݖ�.ȷ�9�J��B\Ї� #����a�Š�Jk ��e����m��A�R8v��JR��(�Ts×2`rՀ6����eq�#�@U�J ���K�Q�:l�5=
!�=Խ(�� r�_����U[˹��Lca_F;{5I�i���0	�������5��[�y^Ź�3�gl���b��#"����!׆Ҧjr	�>�
�ܡ�&F��3#�?����Cw�����%�*����G��j6l��â����"�|L�:������<���x��De�h�7�x}
b���V�z������U>��Y�<��!�=��f���ޢ�li�A%V(�֗ғ��L��
>l����=cxk�~��K7T~�,6��D�J�˓yI+��v�k^�<RD�m���0sqL\�(W����z�@� h)숬D�\��>�����,���Xe��*���=�7����4f=)��s��c;Hl�
����k�r,I��b1x/{[&4�\��b,���gy�"Q2|�[n��lH�O^�̩Cu��X��HKU�4a���]���=�~��U�L���J�0!�*��o:{S-�����9��Z>�|�~��z���b����y�Ce9�i���І��00�ص�/q��4ri�D!�lpK�A�[Y^5�=�Bf�k�Q��O�ɂ���U(͝%��T%�U�A�����N����AF����&��0��1S'�R]��Ld$�9R]��.�ʨD��<&F#�����(/*`�,t�^��nU���#2Ӎ�c�taL�;��`�JvɜS��Yc�	0��O���{CT�>�E�\�"�zS�nN��xl��m$�m����>sE9���{��dU���:��&o�xy��R\�ݤOĂцQ��q��`�T�鳍��q[^��ߘQ��^�+��U)�����5@��;i����?��(�h��+���R���҆���W�l��L�(|�QH��|�c��ەI�_�:�qq 2n�=��mA�������\�,F����s�C.vf��aT�Gg83Q���Ǫ�S�3�)��PȤ�6 R(��t�ܿ]��wWJ��[n
N|I���޿J�����'��5�BP��&�z��-�R���>��7kF���o��f�{��~>�s���@Hׂ���-���������ң�}�j���a��p3�r#�J09k?^H0s�U�/�Q��:��8rDO'V8�of��i�K#N���O`��b]L7%�߮ �^<�勮k���&���gv�I��$�ۋ'�����߿�0D�o���Ⱥ�gQ�+y���A���.&#��𳆀y���n?���BJ���~�8�v8s�#�<��C(���s���u�HbQ..����;�dX���	�?�<��F�v���Ҙ8	Ǧ�)��8��)�!֕+��<��7��\轌�� 52�I�v�m�Q��3ߵ�{����;�E��>�o��y�*�J��k���L��Q�
O�5���6���4��#@Us,�1��f�%�P�8�l�3�%z��'�s{�(������YD���s 
(@�jІ�a����U�S;yͽ�$��2D!W5En�g��܉���(���I?����w
v�O�F�^C���HP"@s���e/��d'�~XA�!`���o��"����A�W�/4W�ܳ`����
�?vA�;a��[�A��o��ɺ�e��b����l�*z�v&����E��j������U��2�]�8c�}z�o�(��w�}r����Q�&���q5@h!�Ii��
��Z$R��*�=�Vv$��-�n�@1���-#�@�����#���*�p�N�m����,��c�&�m�ѿ�ʂZ���Z\ܟ��%Z��^D���'��Y�pu��]^���p�)�����q�NL��۟+�^^u=�Q�_}���G�ru_E܃���Ä��.���.��l�˱j�FP!��'��[����C��P�Xs��o��&W����Q1�"I���R�qV��q��}��@�1~��woZ�e�g'7; VS�8�g}y�(Fb�;�X�r�8Q��@)�����q2R��C{\$�ޫ֗�Ud6�@�� F��K �X���=b=�IX�P��ӊ��<�x�BZ �$��Ry�H?R^{$��S@P�q�<������	�7V
��B�Nͨ�Ke��O;@Z=�2њ���Bb)J=�Ȃ���liz���(�	�bG0�?ǂ�G��Iz�8䪨=,*���B�M�������?B��#M��|p"a��r�
�B�Y��d�8�0�V�%���P��nО�ǿITZ}L8-�%l����xz��4���͚A堘���G�����c�=jq��_�6 ��N�eG�H.R�:A<��Y%V�A�D���b�S/$�O�:����I��˴Ms�7>'�u�QZ�}z�I�)z�WH�V,b��6&
�X�彘�;�o,�ѕ�dh�|��jk�9W�^�:�t3.�\q�0�'��l��1t����J��
�QL�*���N�^�!�z��ޞ��7��W��E'�;�e�H�2@���3&7T�
�]��j�]L������m�^��?6��2.hl76o�Ѳ��V[����G����&Fy�[�yq��s]��a$�����U3j�_���/��$JWQ��W�wƵ�ٹL��Z��Y�����m�U!�c��p~$I3��<��>r������$ߎ2mf�vd8]��$uWcę�V��Yp��A�!���EZ3�8��,ȵ����ё��"������&�����Zc{�����������y��<��-�����;:&��>��D�eN���vru�h�D�ܸ_�j��Ƿ���i�ot���iD���ءMD���v1ϒ�L����S��C��t��+��������U[7��Q(�W�����)]���a
�Nf����닠�װ�w�b���rϤⅰ���d�ܓ�A;����r)��Z_��?p��`:&>��7����D��F�M21� �ߺ{���X��(u���P��dMenϘ��k���{��X�Ѭ�e�f;��� �`�&j8��]o9���ٞ�7?:��E^���#���G�H�N��r�82�S8�c�:�{�ŎTR�؅u.���<��vkEz�Ϳ�|#��g���xӉ	t@g��jD�Y��������ϩ�0���Xs�2��h5���n�#��T��p��w�e��V�Y�Ix��^䂝m�얿�e�9�������6Q���9����I]�V���-s���͎eN������q�v�|��Jqu�Sj�c�����Y��Q�j��� �˔�����J�u��J�i��W��q���5���tn~-c�Cj