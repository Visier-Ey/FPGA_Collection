-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
0S+ZRpbNOah1cDplnB7yo7UNFYPg0tNHYcWaLA9l/F8/DXG8/MinhpcX9DdPxjshisZQ26zSGGcP
LEpDlux0CPHN8/1d5RNgJ64AvH5pui3eKjSJi5FVXiGbWxVFEUrLRPbDymEjBPdepIHb3WKynTLI
Uz0/5CUyB1vvY/8orIqzfzPnkcgsWeaY4PtAtdWFhE/tLMrCkG6LlG8YCL5jiADTvm9idGg7CPvc
gcVPE4EeBv9CHcebhtJCyFfkSG8i6ZnSD8YHNnQa/mlFywSiSvbtZnr+FDYuOWgqDXXIPcHBzW7b
MvuOe52Svwbvb9mpmlynz+OcLfXDBYM97voqUQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6336)
`protect data_block
mYw7nN1Lk+F/C5LdN1BG3y15jRcuV0fNNiuj4w3+YVVBgNKZhMD8VtkaZdXcwk7bWArKbAPA5I4a
gUuRSY2G/TLeh74Tm9JpStpCk0VJxUHOkbJviFtTy6PIEQbP39GOSwtz642lPYemG+ZhYX4gXgnL
AXnZUO6F/8CulbtkVgkyNKE1ifhmm6aZO+hZ6yNGNuNtdc7cZ4dYulAstleqpfP+WVo5durTD0ba
yZKyDXxJymWO0t2vuerLJiJX86+0NjU2KjjCLQTUCpp7qQyTkrYhs95S39AKSVFOcE35S2bM59hC
luJZ2EHBYsS6nZZgNwYaddnkWwlmI88CGFIv7zy+hSp0AYbyR08ELl6bKnF1rQcj0nS5v4J7Qyl7
U53qvNWTaFIfu0jqtT8BAvGmCRKq+LzaPzisAMARqWqXg2AjtVR+3z7WPVoM+bhQGyrE3vxLdY83
JRRezP6pAvCG1ejk8Qezf8J+CeTNp/GXTVAEuBc2poFsZ4FrIhz9wzpOTtGMLLjrqkWmyHBve5MM
YPxfXME1dMjX62B80XyD8KsrM8W3BIDdd/qSet4sW4LPaghWKwx8LKiAsuwrhnxpULLUPydwn3r3
KFIyN7YksPMUQkHODFcAHGaybO2yi7a3M3jxwVvmprmFEqFWcGDCOsAl1wOv/sXzwswd/GFraAOP
SEeyVajLDCGAnnQ1VSzImb3GxxPiQqZnG/cLzDyWPqGkL2JzYTd/oHZ5zMftM5nyCHcJZ0+sIS7y
LxLQVQ8MseP265BjzglGRhTQH3h1IThQ79ldO0MsovseEXLh+UF8r9SGnb+ETmNZc/fyXFanG+b4
YRd/yhPJxk4DuhbWKfXIYnD8XcQ8CdPL7bjiidJ/wPu5LwxiY62F/NWu0jeOPa6fCLR8FrbfegvB
nj6Xts5LOP2EZ9OMnYBSh6HFUPA/e1rZ0mUBumBDj9pB+/Qlc01lYRHK6w3mLAomke9Y1jX9vBad
c3nKNOf+rxR0RU0Wa2QruueKbWYPlevKV9YupBpu/EuUzDpwDPmITPzx66O4KwQvkAX1Db3veh7u
PsEBSQSWyN21Bj20ivMvh2TfYmVm0yieOlGUdqRzlr+R2n7xUgrKQ5FELXGabNc82fHigTuCUecQ
hABhfy4uqvf/Faq9qLdAWCk00TFK3JEZGWW2mDK4akpCaFxNjFh2v9eFiVtd4r8Cd/FwAzLR6hFP
rJWGSZfRqyTTEoGReioJFZ/ko6THlO+IDFpAiDp1judeE4yLb2wFTbEiD3lbh/P19qSvjOORUC18
d4SCsaW36O9MA6yuK+IctR+YTw47r7TA1rOfKPVP9szkcT5ynLBwWoqyLKfJQUfMhyGHlMTAub3G
kg7vHZzHwSEn2lwvRg/lX9KTYZaYKXSg4DoOk+HDLKkcME46whb7PxK+RqfkcszUlgJUyFLnCuL0
KKm9zy99u3y/nWoxezWkSxKRsP/4WeihskBKV4nFN/1RZZyc7vMVX5oEZeaX2eJbVdvOmq3K9K9z
FAAhcWGMXY0yTt0ZMIWCWnvmZCPWtHFJB3UhtxlhVnln8j24pFn0mLKebYHdVAq2HBWuA2g9AR1L
BikFoJ/4N0qvMDw9DiQMfz8m0OHtoNPbWyLzu8ih961djeV/gaiwosOWgEBzxjskjWYYjj20Oyik
3Ha/d3wR3iOwxQW1heexHXJGG+4SBl5WNOkK/zyjSLGBiJF76I+08QojjmSIVLbwp13cLMENfaLQ
2B/TcBJQS+rSwAucFfYHsFigZ/qtv28ainKn3liHW6lin/41G4A85UgsYdVh1On95AhLqO2AQWsz
KdnxdwE9y1/Wnd4LjKsT/J1SFeAqgORh33VphY879e7JWHcNp4huajE384LJx7RJ1oASs6VTD6Th
uLilI/0a4eTSYIITRcF77t8LMALb/jpuVnevjCCUGHOSJ9CCKYWd14jIS1t7SFlY8d1s3jFJd8fn
4OFARgUvE+DqfzLyghYvb8Fll+DXbQjd8HFmBBu3jKrghfeiz5qEMOkYm1AA8wXXTEqz78eFQfSu
wEZk1fYpV5Kf27mzIJFzA/oqnPJjrWseoGfa4jfxOEv7uKaWuZy8JoSqkMBGQxGE8zHk8Ei7Jr74
+SIH+xxC2V2hChmK+XaVGSKSVNio2C//r0koFdf9oQF34GS4patbzvR9/pTnpdvLvz1G91wSfvGc
eMpvIBdgrK26JxZC4UI4jro1Py8l3sXQKgxz/46JuSYs2OIqPG5Lxiqzn0iG/o63nTXrtWIGJhw0
H9lYgE6muLUdVS3iPB9ax7TpRt/bPI5Mu+JQwnob3R81Kwamjly1b1SBcdS89UHsg3VfzI7vNIKr
VHUj/+n/sxOySuKPADBxC1yKgY/UN5h5T7GBw1n58dzEBgH1iqF3I0S7TGJJxA9gGPXzdxgbADq1
JrUAYf49z7tNH0rabqlCdKpMfcCMP0jrfLaMvj83vHQSCKAh6+O2Ylq/77wWniEd+fBlbkKf8y09
lq3cMGIn342GkMrDzQy8HCZmH3VqSNoL/PoMfRAtdqnMH+7yMrPdKw6PBivuHNlGpb/FsXyudZIe
x/QgR8t/Qt2BBxC+96vfDfFOvr5Pyfh1/wlYdAq9ivgI0gPj11uPXQ65SOkG3ZwSqJbLHmvtAd31
65QQacOehVtj8cE9vh6XI5qo6CEq6uVPaHNagVACvr8TJr4Q6XWBfa0yXcI/BMC1wJCRiG4XCjc0
CmyLK82RD3OvV5/AR+ZIAnx+KOrskPwS8q1gRXs9HiJtwRUw04DCr6GC2xuuNKT/Yn35/cRuIGDD
BifK1c3FuzO/DpFIi/c5uQyouJJX8GOaaEhmEfL3qTH45jF0NLj1/sZiockAXz87A1cl8IxSLb7n
cOfFqzKdHIuYOtPFFARssDBgaEhHOH1d4jgURTepxIxRPNIjXc/xSHZ9g4PFjg+6X+f4AVOuwtXA
0ysiLJCJhRbxxhxuBl9M+h4e99wC7u4Nf3qnYQkHcboGB/69KnNbtEy1roO2+1RW8TSvGUE3DkBf
l5tskxSwONrF4oYNMM5TUSS5f7pKPQAVtIYgnpqysOo6wRlc84A0SCqeVQJKPtgXbNz+y9Tb0MBX
Vh775MGTb5+w4yPfufs29P/KueJdMS+Gcoj6oXZ6Egi04RA9Cu8YhO/Z3H513kXsQi8Cm+4t+f7I
KduTJ9yXvj63zvxaFEBgKhdQZ6Yrg/GILb+1B10QBBBGImWihuG8UL4EmabpSOOptnnY6gOsfXIi
sJvxCypyKsRXHRN8t2AqZqU3PMBE4O2eXkpestLNe/9G6iVALO4+U8+U029P5UmkM/lk+MpOwTCG
hW4vlmaPMYDmXTcbXd3sYNIiSAKoINQ+3oMAO51JNw2l8bxuS9dodjrPC+Yajh3iOfGKiPHIfb/A
TdoA4UzaqY7aqdZtnRKSnfRKMCmdxKySEOvtnXS4rsAbwFEq8OrOjVRWlO8sz27zGsMEuYXKRkos
lNOzpj7pQ7OmuwM95nMhUp93MvSoACFb+TQ8mrk3VKMQxxPsG+Y72LofnuaqSwDdQs3947cGZhmU
VdM+F3ZOfGeTPmjYHPcwRrIU9RgLyTj0uliIePcu1YyfKzdMXVcrnUKZfD+V4kB9bquOmZ+gzjwD
rOhGYyT2swwzGbePBGFyA4uShS1F/CCXaPxEpHaRhwgZ3hHf3eO/cGHGpyOsvgxg/7VKBPF9IzaH
48HIIHMtUWwH9BOHk6dXhCRx/qs77bg3y6XnQVWUe/osv9J51SH+yrPqRCXPEA+jDk8bEmdpC91n
+rdjoBbkHD7cUpZnz3QQgH+ZqZkZ41v+GoD/x9IuoYSpmgPQ3EJXTIM2ACUwQkZ2fQXybWO/eZ6T
LO55EvHIth3FjpwWvTUu3ehGlkhRuEjUCVHRjSUVfwA4gO/ukAz+Qoq/d8LzIOjMpP9y8YVt/WKM
uoXav6uTCnM1egqB+B7JQBnCdj3G6hCOng8geSBorLPZCZhF3aaw3K6+dhedjZoEhfwg3PuD8V6N
ffb/1D5fdemsqtgDgm5uQclvfmHraEEMbkusbwkJyEidcg3VxDXPF+NXnzB4ryQNCXlkT+yRQAuh
7xYqddJWB1VDFCn85XyZIGkHF9W23OKFRq/taejmFXpZaeyvjJLtcU2AcdaJg/AI5p/JZH9M77hw
ErdWau6ulwnWc+O4OLW5crMFJnvabHlXWZYUbnoesE6k7gRAYof/8dBbxfAw2yhtgWVOeG/pUIEa
O4Bj/C9NGkdwwdH7jgdgs1IotLcvBk1soNIkyLS8RhWNHDNIeSZ092QXo6/Gb+1bqG6fPBdx2FKH
jhCHZwXx7EPbjCNA1JDp+RgGL4W2sy9pR0CsVVyWfmNnCgxpge097UOSEjBNhTltwT3lP4TBiG+m
l/sK3JwPuE+pOqaA9QBSZTEUK+do29kboJtgjhfSDMeWWn+kzLyDIQy8gskyGgkMi84T3k5AH6s4
x4QpopZnTVSK1pLRYxZRW+Tm6sWPmrQ3h91ORi68K8NkY2VRrN6WLgtlrAoAfDjG3HYNSu8BRQJh
nJ4WZKXHFYParVRPTU5q70F/gXJB46ZRGMXqyTKTmwv7eiUzXHWRxL4W9tKDz4F84fc0dL+EIROV
tDUxHegMNjq4hpWpHsmDlml5tYqWSf1bfq7U9MuvxopptQYP4W4CadRM/cEqEzeGvjmvyqU1pJCE
nML9KIPhFjy7pq7NjsqBr/lg9+8QPgqrcurv/bIvzzEv9Nuoa8JCRKhJIAMc7LAukvSdQUK6YWiE
OnUBuoA+JHJZo6jV1N79Iw/CtK6fobY3qrmlOMRJLxRiP6mvL3sB1m04rR8jOpsbPA0jMElYypZ0
ZWSwgLknx2q6B54BI9slBxNOeX+tBOZ8hVxgnRcq0Mvmzrs0yXWc6ON9CAIUsMC17SlmLgKvoQGi
2a4UHSIYadoYhLq4Oi8GUTxC1Py7bDBLgEbwXbSjfMdydbr+MBPfZbJ2TpjvDkluyM9h9fLsEn6A
et1JvmCD+kBtF80jxZSXNsiixWNbR9EQMQEEePh2ANhnq0ECDujsPQXOC+t5bPbw+7fR6VtLaqw8
A4GRHGcAcT9gAoOmasCzWm4YdOvAm8qI7Exrq3msUQ5e4MYftNRNN/3bdne/G+9q3H8bFO+w2UPh
DwUsfI7Pes3Zk/HvgCCS2u1kz8cpar5ZbuBw617LCPC2tIQlYaYls7wzhM+6T4UcXkDr8k9cJ1ug
qRtCI859sZj5CROwSzlmR11nolMxdvL20DTJY/aKHGQm08nbuLaDlBDkRMAYarLy5bEtGpHklepU
/JQO4vucJxAjMNAgkdc6kYnPyDCVzI0FYcMJasiC5dE3P5KX+DsrownpbSUJBlyM6jeNjsvQlf2+
aU3/QOGQ2R5QoKfcMdyIYnESXPb0IqgVYt1VWsCdbpRyScH/nzS4FDVZiEl9AdTJ8J43hq70cT4f
bxEyaHtJa5h2sumaEP8u6iiLjOwtYg/bUyLDozHZ296o7Q1rHl9p6C/ZWAr+44VMtqB8ZqX2ZQXu
/ktvD++9xpYk/78ZPdXEbaCZIpis2hnqkLZr1pJJV2NFBd0XMwDWJTY+3FLO9y/w35q78lHe7Ti5
zYnokEt7527ea2MUjxpCPkV6TLCaW3Rumw898R3XjKNyLbghRcrSq98XrwSUgh4Shr8/BYAEsSWX
X54rVbdvl7tzDFx30BftMnfC5xGwkNmqEyTVdCmBmDG633PC2DVeuQT+iox05UnV/pAW1Eczyfrh
m3HnsT4z2gpR33E44Lger5SFsYQ9cnXWG7/lN7jmrbOAoihBW92KHPzTmRNzjURxL5hW6RMGk8NA
U/4oYrDnG71I5Dn3fEVa52OZ53X2aIEHb2IHn6bofDokR1B3UVwnjZDbIqdmBKyC78fE8xZg3pb7
VxibED8MBZsoZVBWKt1cUSJaDGJNWNsWgPc6cq7qqMrtIf7m/bO38tnz9AgQDxXx9GxuooJb/vxh
QLaakf6/mgipuOER9EooC4EE1SmwPUHJkIXzA3uqIlUQTzuKetwYgeEgVE+OzFfDGfJ4UwlWq1fd
B8x9p8xMO4pxDpw9TgkFcN0ppbOvvYSa/RFacxPJwrkFJFvHLGCz2BwpVoN7I98OmpZt+A3qC7KR
5J5kZWSZ/ibAMag1ySvTpsRHPwKU46c915AuXFUKI2TKAAvquf41u/lUvzlRGNA0bmclbnnS2axt
oMOG98acel8LOM0h57TqHtV55xG+KgQJloukwrHsM8y3Mgc0j57+BfV782ElSIXbsNEpx4Fsq8DA
cSyxFdqN17NMVY488V2oZe9uCHnr1EzhRaywBjLKwYUqupiKY9IaJL6NRRAtLNB0PCnFv0BVQg1b
owGCC8YSvKfH9s8t7L8he3zuTsYF73ubBWXUvtQYDFCvs+Pecqd9KepaZsJS5L7re50RYq1THKvS
z49UbN6e774gkOUUA7YAS091W+IVUvm2jmq2WtJuUk32cJHeJXoafePvVEMbPECWQNylcChPUSRd
4gYFVPqTYTjfPkxftxQ7gkGJC1TEsT2zq6RJZuxDDPziPwVNAx6PqnISFFQ+N4h76ubXVKc31bAs
QzPfW3Hvvk8kxQkbzhPNzpAd0PA1n6kU/ABuyaLkWKEqikcX5tSyVQarS+FST52R/xBEqy689icv
sYNbGe1i7GQ95xM3OJEKM7+iw85CR/wWbmci5epj1L+xluNuTQyl1xmsU70cCByH151EIbNjUw6v
KcJDzREu8TRG0aoU3aICkRE6IpXZVWWEY0s8hSh9/M2OAHz8plaadbPDjKkUhBXPBPLDwJyRSCjG
7lXmVwbrF8+9+QFylkq8MFUQjs1aOBf8a4LjVEuUL+USonDPvvsCCp5r+9jNaow+r79KsdkS55Bs
CdPy7uP1wjbOGd4gFOIIKJJxVNZnNwEqwfFM439uGRIgIs34KYewHY4uhz2dEqBeMlgEmHORF0TL
D5ZsTmzl3wEGrAyJ2QTl1lAcc8FRF+3w59KB6W0B/HPY2nWOzc5DQltE/CPj4whFRSSt6VZDOf7v
y3Ow0EujmaS3xmi9YL+EM/XmVHLFUeariON8fKn1gIvtncCkaMnHPhOKZqQhqpRq/ZbISOOjGvvd
tyO3PNRsdivwUwIOO1rUOS34Ql7hN4lDTjHcrzFuDQv2XkvD/fjoXud6jzFfOqFL+SiRSZU9nijB
MWVbayW/tC/FPInofGSKekJyLzQn/VzMbq+RA35QSREjgRHyk3ewTqo2X4R5t1tZh0I71l3wgEHa
tAFbhctk5pxOZIxsWt7ZZH/DOi/gr/YXmTwXWI9JlvR8hElZ/ZzON5Mqu0q5KO0s5ccEhkt8jk80
KuvRSzD/HNzUpAu8/KS4e+098XQUj+U7uibJmFCsviDqGCEoKqEzcp1/k6HpXYrWn98Wg9rLeUj5
4Qjzunm8L7CaGal/RmDUdT9yV2j/YN5zkyiejjyMrzM7kLkyykydTMW3qcYjnJWIJkb6F9+QSKcr
3dguKicSgzGZGMTlGvv8Ez8bMDcQEmK5nRgjC0opKtUVFXDGQS4XTpIaRXSbOqvvXegjcfBWKT91
/Etz+vhLh/YchQyFh+UxZVobuRDN9BqKzr+6MFPcLpuPv7MFWK6Kcgj43gObrBAPjIB52XGiL0rQ
rkSq9s0UybNud9vRhxR/SnZeUoUovGQ83NKH3F4rMxuZsU1mbj/rjISZoRUxZm/wCNlulFqk/45C
9W+ViQ3DeJHVkUHzUUGpk6ADAoDj1/wzmjWlN0XxwlUOmV3goyXdVThXQ8OAaaz5qf72y0IzFJf2
k/9IIHlCJjCKxxuAJl/Brr7SacrqkoYrGEOd/sOm3vitdg7qoALSPgBp6uTY/u0t3n3yaLvfWKLV
889r4rl6FItaA/c6PAMj+IoCcr1RV1Q0mcWeJ01K+zrNZhCg9ZfzhYvEU1y5NOpHQ7TsvNbD1Ei0
CioYfl1danWEKwaXepPkJSnULlNix1YX8h2ia7u+BmV2tenoS9WHoxbTvKaWOgrgi67rjoXnZOT2
GUhG6HgVwoa22VqaYHym9qIZnouRmTBTRIMMzymE7GqAQYrHr+KlmYcULMqJK2sTgO/BoMnSZa66
xO/axy8Xog9vopTvW7VYbJ447x+/uKlRFeO+iEuFFaANBRmhVC8hQgECxlzfZjO/lkcKLEfv/JGD
feAlJFcWVVQhczc3HG60MGwEhjz4ScpHl7c0KGMC1eu6q08YaJ8m8JZ8px96gIjgeBu9CuAxT517
U7pCiEs4+5NKcFgAdQxhuDzfWlYS01sCG0XVYBOEOWlMVww/HFVY7UvRAOBzJ9rxnB+hLdTPTjY0
yD8qDA48q69hWzj2gpVh8XpQOR/9bQ+te2SbGc/YqM2ftNzNrLyvuZc4QMJ6ycucUVam40nFM6jP
7lAuPPj8oH0r
`protect end_protected
