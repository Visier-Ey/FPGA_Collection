-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
cIBsaEegKEX/0dx/QggVzcyFlXWsTOIDqYpkQKFo8eGizbgdsNaHQeCa8TPs7x+w
Chk2iGaFqNUH/u+JR5TdNDnwMYiTdd/BOa+QBBlnEmQOqeAe9krazq9gheAPl9zP
jx9SjYGkWVgL84DI65Oong/ja/qRxy/WTEB2Tj3FDIA=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 1013)

`protect DATA_BLOCK
wNzuk1rGQ2X6lJvSKzDFjewMCKOls/ENJlWQXYrMsgf6dAOaynMlhUdxBLLYW/1r
t4Kk7SmLc+wlMGg5nMvpqzTMq8MkjReWo9kTcAX9fWGpuKj64y0qAsPoAj7U25kh
FxztOiHXVqG5YoZ6LMRpH1qW8kbqf/az/DDfK48ROEi3JRVMKEmCkd/toSRxQR0f
GTBnfaz0humOM7hU+ecLGju3PFje7XFePriBFgu7ZwCRmlOep68C8o33gdEuqXYd
plVEaXiM14l4PKZ5IDsQlly8SVipAh4qnKhw9ZtmiRqDSTi0CPB9lmYtvF8Jw/XL
fmESsrFA6YXWbsVN2D/orN3u6NeVnrqULd7yyGuhi1U9GYnV0v6Y5L+aC1pi4mlP
y4j3NnAKPPOd2f/z670d/SwnLpFOED4JUHkr3iXKkeLX4ZgESa3jkunvVqbXsOYa
usCrdBmmLphfzXbz999WIVUzTTtMyN3o73sFEkFK/X2JTF5wpi4nZ40272qZ85Xz
/TtB6IWfxpDp0sDUraL89CAH7x3TrIk1miSBj/cIV3lPmA8z+u4/Lykn6N83vurs
etw3bVOvzI8t+zalSjOTa9TMfS+3IfetxvHqCNISk/aFhH2qz/L54aWDyIIqKohr
bCgG+M9ICbkVoVHpGW0DgVRUu3SJ3azV563XTYF1c4wmxmBvn/AQJPydBO0ntOw5
SrLAJXThuA7yoYvR+lQaB6742JDLc9XSzGR5iNxKPKLaeq/EtxE4uTMav6H7DdNp
G2L41HWxdGcd0HMURjqEzyx7/r6VM2P90qWfQEPk19QZjn+PP5Ys+AmUOLv+66U3
CWXx7PrE7W36RHKDHXHgV/m6noyioutsU44O83mKsYiwm1Wx/ZRteYqhLzFL8trF
BRunon2FoiZ5LO/lykNOTjHAB3vyB7W0ARJJ1r+bOPAMj4jbmHH8SQtUm08T7O4S
aIljmcb3p2OgFKfyUN/vil7j+6gDQ5NG2XpI6DnJUUwQPnJxgmAN8Wieq+dUgeRl
6D5g6BrZDD1Z4XcgI+1zLAsiztSgLFOUC0/A63qmQ28xLg5Wbp4np7jtWlKwSCUJ
LbGPQxiGzg1RQ3PUk8cP9BzDM6XRCItjOERpXq0zLwUgq4hFMKtC31iUUrgx5J61
9uF8CUdf0ayZDFQXEIwyQdjdOEhbgaCOwqv68zd6yyBgeZJuw6QboNiWQWp9qA7+
6VdAPrw1lktLMLsU8ighuiu7u2VkXXiP36KUGm0PST9fJEuobm+OFD0xtSMlinBQ
ZcJeyo3Bb1hASm96Cr1W8opN5rWB3+POoo7jgT0hFpdYWHIRX++X23sPS/EnEl9C
DGpYGyZwhqR7ED/k6N5XGx833TMXqOfzCFau6fXLGZ0=
`protect END_PROTECTED