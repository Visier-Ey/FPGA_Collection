-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
U7PzwgsX8y/Z7lXoZAmg7cOPng/OksdpjGT/v/4I1QKIgL4JI1VJDa/y3vGsPcTU
rNb6wIRNFy/gibYfCFLE60pV6/4IboXs/W2C2m6UDdg+gwRbmcBYgCBq8wqUJOFV
D0BqkYyLmb8CZVvrKBRg5or43evXdeJwRRoaCXQeSgg=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 27995)

`protect DATA_BLOCK
8RgoX7mlTAwRGuYbIZVI3aGgBilKyx60TkF/BIMLnijNaktH3z5vC67ihOI17v2h
xDUWVtCXL/pPRJNRHqFN7Esieuj4wvUEDRGd/ubYdsuTqjy7t5skGzbGlhFEpCdZ
X2Sa//joMczls/LZ+Ts2gvqJdRPoWWnejkqILdVnzKbiCntz9bpyEbfAU8xvT9CF
yRDs+3KI/DR7tHyhvGy++w76qjGykm6hlDJHArHl0t4SV0O6uIS4FKa7ImKLZJDK
hsLquIrak77t0wnzCEfJ2nKj82abBSho87+JbC/yHxhx77cGaKhxItk286flmbBw
H7VkP03UJpCg/BtbP9YyL9SGsP7NZfenHl4oYRLbRpHf0lI64TYgWYAYKCJ7kTim
wT88nT/6VdmBsKWZgQATuX5iwgpC9y5AZi4yT9lolAFC3KQtupZJNlddTrOhA0Sd
huIWEzaVmosr9svdQ/hN5gw1EJ265dVAQfOfT5NlKTebGOB1/UKx7JnPV6rsTkCu
suPSvucKVjwYTIWqvh6wKx0aE9ajLa0SCIiSLjac3UCNW0g5T4Mw5oBr93TXVT1H
N6lNng8aM0fNFNOsiJ4+zDtome6Jzu8Y+5nMxvcT7wHfCaAPq7hyx5XLrIWEAm8l
L/AGev+8wiwRSfZm/eJT+y8pBKb9Q9gei+2iZ+X3fBJyfRYNotCViXmnEYzBiiNa
NxWvd0jVDbOJTZ/ebftVaSq2QkMTIX1ZBfLY96ztuunADDuJNBNj91bF1RJQB+bF
e642vjOv1L2T75+NAzG1tqCi4sowNkwmiy6J5iDg4Wqekvh9GAsxkiG/ZRcovO3o
UPMzF+hH8l2qc7ap2pagbosTidm0xg2nYLdEWhmIlKPgbwEnyLimhGwEWvhJ6WVg
TTu7/A5+j0serxS+9cG8RC2/7p6Beaj4bzClJH+cN2y6cfpVObGpehLwtU/TmLz7
tBDmUHCtS1cghhdZk/hNoFo6IF4xE8/xZk6zgQ/6+RqOcwOWAND2q61qscljIx67
BtoOon7X/1B30sCuLQR4XM4B2XoK9SoMyOW3ILDjgL7OMnDO4IhGGAECcrXTgwcR
PpAX140D3+oY97P25QyRv1GxHU1+Im3c38NTrTEYJMPuwSzJh9FJUsxABqqXCgwk
G+n8jAo8bwpBlR59+LBeIf68vtYK6xg5OqygFrwn+ZpFaMwyrWaKTQNMZlZRKgh9
T34xjAiMKrNgTVYaajmoCCR1823vwvBtfWOPqHZJI7pZ3O4XcfuN22KTJ9QDKD2o
z7aBnl0SB2sazsr8Qi5ysmPTO1Y/C+1i6sL8OYXFXfz92CaF88MRGSMLwgpnBi+m
I+F3uq/w0V8ENLRVsFKXPS1tDgcT5cOkwBywZDeKTRgmqQnjBsIHdlR8LavAVKEk
1fWlSOqnfh1SkWPcz7JF5yyltz6Y5hVCORScSAa1n7DZky6sVGFvf4HigEW14Vfl
Lz4VEAJhOy2uI/OYOahJTa6Bl7ea/L6wNrw0RU1sewcg2qQht+40GLtex1VvwxOU
UiEVAjGcGT+mO5q1+uibkDSIzrxuIAk/w3jkzz6D2YLFycbcAwWr33ROQUYFg68b
IKvEwQqfMbp7kdsP5hOMJaSNib6HPnuo1Wz9GD/pga8GovgL0osgqzcyyGxCNZU4
S1HbVkmB7AOnbKy7uAenwha9ngj/hgHR2Hh/89uv5txbPoSp23EgQoCcRelYdDT2
sqHYsTdettAYZ8f+utupo5Se3WkloQrczyEYZqkWeBWNc2kFXNygWNnb7rE0RAFs
aSJZt6CgA4bq6V550kCYsNMDpzWHgaO0RU7Tyf6ohLYq1KnuB34LhCMG5zGAoO9F
sKoxRjRR1WV+6cbxj+ZJU0qw5vjF6RjBYlKRpjeTdVSiV5TONpL7ihQh2KMJ6tzk
TSzpt2oNcS/YEv8FezuUj58ube3NPi/7NyrPt6uekIJBZbHoo5+hdatH61gCS8vy
Gd+dr0JIADGNXEeMNY9joC/0b22JBrTjl5smCj/M2nrnUnRrSBw/RPwgcHYYthcs
mWPWWtkRvBnxNajVhaNwl57hmzDduRgkwVdfnGHVhjwr742KBwtIc7rRfC/SoxbT
G7EaflPYEHXZ/VPiZZHsANV57+3NbcNabWXhJzJIX5m5bgVIjV5C4S8/436ZcQYA
SFBkjarVWceejN1syxVUCKQeLwmbpcewc5hJ0VTY8/YrNSV3RQrWUSv0qhP8+dZO
hkIPSbQV6LVHWx44cYDcDTCHtaiLfH2OAs1N2N0EtMtCjCSPGMoK/t4SvsPoL94t
Gcxkp/xBOm44v4BYAcfnz5xPM07+XrZ5AFY2akBBI4ZPXZ5Da1Qhj00LQ4C7MBMl
CadmfpeSwdn+NPwgaPJoo0lRMiNjdQbtFy9/wlS3OWivmF/JUWNGDt1R41ew6b6/
M/ZtX6s11ILuKTZATR4Q1EDD4bZ/b4r0MuV4/2XMwSCyWBs45MSJ5cimQ0R+kfIG
O9TlKMX+QwVtfTKkZU5dx6wM41pBmzGpEJLf3CMoKQSp4worDJ/n2e/sLaWAHVyx
nmIk1nMcA5/miYUkui/KlmcfoiVRORZSLw+rpqfvkLvFhYWDkxU5rm9ARg2uHA+N
UHIXcXoJgWpPRTk/j11HVLX2faYvhdMKXY1ecoSPin6CkJRG3NAtvbVEWnerEM6o
nkTZ1jdVMsaKXVrJEPZh14vJF9/g7GIKDp1OIDO7fCeDF2FInyFyL5Gyu/Y7cK2L
S+vpr1KVMxw1phUaIFcyJqV5mRVdP4eyFeARDmI4ner1S/S1Ip0K7kjRSiJUl57E
glxO/aeU2NHLlixmjsKgmCK4aU0aMXXFuoU2PMTo9JDNOFeWn4Q9Ju/N1A4IbRyo
wP2RoFak7PjJmoRQ+bloxmQJUKIaKncaSofxa4k2hDW2pXOrOzQkL7LCbvbCBs0O
H4nLsMGvLFzStgRHDWoiJjcnYzX08gpxvfYsgbVVR3FTYqqZgUtMRdE5a4l041So
25uqT30pYPgMdWmf3DfR8T41T0o6f4yr/BPA4LvWwDWAkW8Bs3w5Z2uPOyRTMEo7
zVoqpq1JAKMr9htZ3X65WdkjW+RwmFmE/Dn0ncRxjTHmRI/LuJPuzcPwNN8mFu03
L0zqh8TAYz/tca5NNMV1z5tMVWg/GiB53WRHD2SqfsSw1DWC3ZdYS1zm1qjnFxlm
kI5mFGoAK8Z/yxVs5SqcwLkmKmAS9XBF1Ll/6iYgyL3yEWBoBpXjy0PbcVEucYU4
iy2MDWnqJkzpvgqS14Nr2edUHpsfQxhFTulJJGKgg8TF8J4oj5dalpX00Gk01Y+a
liNWn8jNSyPw74er8bbznC28Jmm30a7JRFZOrH4QSS/BaLzKs7OOfl6z0BEEaVwy
MqK3AEVxjyYlaSm1i5ek2PYeGGRzW6DpUMGpaab4LsjR4TPRsKDE/7x9rCquu4bD
H0/ySpgRyy3VJc5g+Mi6dJl1zpsiXlzk7HuS+XGy4hSJbSoFyNDK/sruHzBOGAMu
PT4ffrGNXoJgUA6ykY3UR9Eud65ECudQrZ2vCsnZPSJpfn/yF5TpC6rCEKX2GTNt
NYbpDPbAm+E2+9PeZfY041qilyHzFjfhDNsgnDP3x1vbcZdPQitqrjRNbLO4dK08
q0ZXI5mmou+xz/ebwfjcAdza7gvhGvsnNPgzBViZgNuT501j5Y/I6RHjzJ8fPyC/
Bkct+biMLzlcuLR90COertyKbrO8/Q0PaPanfK3VR1nB8eVMKXMLMtM36XOfxM47
Y3ToVBjqz6btVxP+qhmeIWTK/2owHQ0Ay75M60b6VjFScYGC4AdHz15vCT6VyA5k
PGDaYsiSbbm9a31fvrWWnqUoq1Q1lkhlwcZ1Uzyzgl1H0nomQQZATp32CulltVNV
+iLas5RuVCZZID2IB2MNnLjCfBu6wJzi+z25VU1BVG1uDUE8uH/IvGpXbkcdhfy/
J4/FP4yUJtztVGiVsB7WG7kFljCWRVMLNwmNBv/+P0nIB8caJZBh9d9VIsmcCqRf
2dREEjPEPFJBQ2MVHrMMaMDnnjH35bbxxtlE9Ce+/nM+Ytf01yHVJjnfvlq8Q3Re
9npbk9FaTM/biH+4TKUpdVz/D84zdZ99YWiFn2yloFsPHdE2Mq0taLpfBuiUBnZ9
uuxxhhbAAj+KEoJcdGcWkzn7f/uBxr522g6kE2fN/89k6/1CCBfFgr7ZLV+WqlL7
nbR84BY9iAqkX7KOtTMZJpemWh4bVdDTZSZnbMUSMlX/q3Nt53KQOBRWXTW+ulHR
O0Gq2FK+ogeSf6de7x9sjsfpibgacg/CbWCFAdERie8yCv8aSi/LRCisc5SNpbac
xH1H0yekKMJ1MdTx6GsPaWcGFmMpn2J+8R/P6+90Xz0arkAKPYFWFMOZTKb4AMos
y5YDbY2qVqhgY7VIZ5jrFVock3d0kRbml9sCWYkoa8+vmEYSrxlC/Ce9VehRlHHe
0vP3Mv3gvVqzPc+FI/oXFBb9lmK07VzEb3zLvQBBHl9mg+hQpJIzVdbICdNHtpR4
D2B/Zuw+DFQcJbjfCJGdirH5iFAY+No5SIEtSOcpeSeD1hEFkJJdlr3Lib/VEANR
4tYxd5KCChrGkbUKNZ9G38dxiekMpTqe3rNT2ppnogo+iCNGfyWEG3c/8qxeRXbp
Wzbu5zRrW4+y3sLJT5Sk7tdJWMMHJQViS4bxRlB0bxp9ZsOluQ7YmbLBf3Y5BKOi
Ks9qT9/ZZh3Epr1rDL0zImvx5QVLTSYiF91AzFfPt9dJ9I8hFtIgDlSjaFLKIklO
5X9uiqA1fZfEQtqE+Qqcp5NXyRvxIrMFt1XVas+C3J3yZ2FnUJMLnVa2lA+7zUSO
dMjRt1dU6PSqYNg1TkvRql8AOoBU6ZFm6M7ERfM1v9EQ82GGHqdTeirgXbWVeWm0
Ad1XGrs8Xpe+1HEoygrT8XM2WBoc9wxR0EbbyLbfqaRJl7Y8F+ik1GyiR4SYH9Hb
bulk5i0aCXl1/zVPu8SUracYkNkzkdPMiBt8mg/zG7mYAxSZSU4fl3N1mYStD0wC
j4ewKVzJl+5bb53ql8j8i1WbJRIAg7jSRIRo07CL3C3mCLUiDlR0mkU/FnsJTb3J
++fPH7AaT6TluEHTAvrCDVxpWyBUGyZrJUwWrL2//gGEbOv75E9SUsPILe13JMPJ
IV+RKe3mhJaqMb1shC/+lMc2AXJcOh/x6a63vbXC6E3GO0Yh/xx/DOnHYUNdPKQU
G+yKKXV2VJ7owdi7WEJAAQ+vhLYyQPCSnCqx+iijsHxDSd2MaitpKuU4eiXaJzdG
BXj0dSAl6kq5lSrDXtOxUQ1uY6ahEA79MhEeS/DOWe1GfnsNvtPMjcHOpRUcNCsl
wUniub9R44fQ/EUtdI4xnKY9zCCVbsB8TEUhv8YgYQtWSizj5wTepwhfG1qrjrYL
GtCPXg346X1lnz6qe3YPExLHTIE6Hn0MOTi04XtBZe25kEHcDZQ9C/FsHmXLWDG7
8vyTgaMxquRS8v+CFZpQnDH4mYtXxt1GF+0lAPrpRE5G61vzvOWoU3UVPvBfCxFa
DMiBLbyJTn3AJhZa5Ikofgy7Qxj1kXa+yx50zT9vmhMmHdiBHUDu6rQPG/1D5xxm
e+PvAk3hvPBEqRpJU6WsxibLv//tT8kxV1T6kSyIAotuvI+S0piNUrVOqg3cIlyX
Lt4k0lhSfwi2Dqw2zxpnSSB6H/mtNicl/GiD4NMuDFHNH+xIm7TBjkGlKin0C1nc
C6EPRr/njWsfLMI2Ch1FxpJohK49euThLyhNAl7LcIZ/S4K7P21CEVob7n8u/6H3
YsSqDdRU++/wVDSj7RC+SwnvLa8mFfML5nXxAbDl0BXw1Btwhy/BHFi5dwZFVDXC
JcTUMlOSilU02J7B8ey/mBj60EvRlAFUXfU21L7l8mSjQ2l6cxDLtwMiEg/csl7l
A01pJbeguAqPGqOzQ0BVLBjbCfciP3XbYXfTVsnr1OXbkJtF6NoL5PvBiWSie6Ly
HVAaUjhDAhp7ad4YwRGtips/xWXGn5fPKMaaUuc3bc4O9r1ITpgzdZnDkuhq0Q+l
krYarA6J4zpiTXeAJh2BRQJt2YbKSgSDlQELH3RGixoxZ+p0/nxi9wJkaD00hy91
lAUXcaFALRZpvA/K//bh/sNNqYs7DbsJY6y391b62CkjH3a9uJgms7wQMV/W52g5
Bg1vnKuSGg7AMYxUxXHIOh/trMkenVOWsIAk9dBs4ceBVcqUhz+CaOzJkxEFqUNq
pYQeB2cjspW2mWa6LBvEPlRexkdWN/6R/6HJlYVEGNjLdFKJqq23rB1LfvRErrVL
K0neeSQASQ+QjaiSGfjaY8nssqeFGlmf5kZn4vnQg4PjcC25prjSGAKtH/1MQBFU
8bq/SIqGgV8d6Joqh/v8iliOf8s2SOQaI3Bim0rrdbEOpszTqY2Qk0b8sOA4w4IF
7wcscUW4BbMUhw6E4DM08oiTZhKgG0qVHW2yH8BpSWzEA/DmqDJKikU5ZXe6nlH6
6eSm0ReK+MP+JXv65vAYYfXsU7D/ej/2H+4u+kzEH+iZnky+EduoPVap8wuR9HyY
T47v/1NiW4p/RFYOBOXU/6kVPIBNRqpyazzzBHqxKAHf9TsWBISlOvyaBOwMKU36
jH3lWIL3llvWtbh1OfsCTPhEeHxwhkTV/fP+H6dGnsEGljXYDmi4krpMtF/9XK2j
0gBDO9dWhLrm+O8htC0OriEkIFwA1Pcuxut7N6WLYiSpP6S9lB6HsGhFeWq7eSm8
S8lYrwvobm5uMlLBJhltbnz8wiUcZrEl0LSXZ+fE50a41dThLCMMmWcUpcnD7odu
5zcOzJOgLt7g2aGRxOuKiG0fXe2/OTbmb+ssbXobFl3ZR3O2rk4eMEsPA30TpwMl
xpX40l46yS2iYJr2+OljGupM88tcd8r222ZSEYj7+KgAc9WoItwIgv0B9Y5sTQHC
KauAaX9wq3VcoNlUOtpEnBfy1bs1jjYSddEsiMzbd+THdWxfn8wP4T5WvhSUbCGu
+hYQat+AVgIVzQCnXG3nF++KjxbYwzaVs1JZann/Bz+KoZm03ZX746z2YC2IOmRV
LMihv/2vhsZSqjRWR6skAYXymHTH8CV5q+vBMNEk8i5ebZEnBG4nW9F0hmREcX+6
TKX4ZNgLrHeMJbH2etLJseeCzCp83sdVN/NqqKTLr1qTzmJr/83auZen7fz7MZ5A
B/5R19s1/nN5CSd07QVKPqcZvn/NGiF9O/AWJkltUxJAtpfq24e+ubPZ/OQA63Mk
fWktoF13LTJxMD68CxHne18Q54+FP3jA4vldMnIabslHYX58wJlZ0QEpLxFLmYrJ
scCub5dQb3XpipQPoGJkZB4h3VtyNofx6wnhLCKWpvtvI9bc4xT9E6r9uqduHeek
04U7m6LsBM/CmXUToWlHQyTOHVELTo9Cxmsvp5nMU7s5X2/iLD6HLsh3NH92OI9u
j/qy0mQmCc2KSCFKXzT2dWqU+xaiu0VLysm6GUIptnuzap7SeemplDDw5N+Q/lWv
rm+t32P6tdmp9SAU2nbK2dCC4ChYBC2wLN5SvMv4GZvM3LksHN46q0/DAcpt+WyH
tma1yKuDomY78wfoYcaIlYnUp4lrNlxgDxzzwZZSbYzmFpK74oTuuV8FZwYbQeZA
mhaNAG5v+vDKdmsEVz2vOBblbpYb2DIkLYKtxmH4mx6kVMiQPLX6pgFCEpSan+PH
BQAfKZ1Kmqy4MquSf+LjGdOwGSbEK+MDlFEef/RVv+W6jI+heEw83+m1aSWfxkJ2
SSDIs3TJFwm9hGjDqK3wxxYos/U0vmDWu+y2IbDsjDFB+qUzdhBLNAbJyfuZSE6U
RCdkdXRKvZdmU9RJKFTphBEmo9K3ZWEkP8TeplaucQrAeoNRsU8ijTU+AFfuq/Lw
tnzlicXrPMBrQj2u52T0WcjKSOivMcZdIjdUkCIDbhZhWesitzAG0iBohrotUIMc
wC6UXQNd1MDm1E0VDEu3T8eENuvx9TuzFLE2jYGbniLny+M0Q3WQGzO859WSs+xi
jSAM3aszzNMyKPhQSWI5YUVX+litFk6GytpFWm0fuM1N3V/6xZlnuDu9V3nqZvUR
rOkbU8nzwgKeqT+mm/8r2lQEisgoNvCtze99lwFo8OPrEaEvAQJ1FXryXzF8h8He
Z/s4s+zJqmuAvUGXjHuIbrw0bnFuPZPB0byxE2p4mvFG3fLxlmASmJO6RdTICivN
sPEP4yNPvOLxHMLjufV5EkmiD4nawgX38pT+xI+Iwq7VQjLdMvYnp6Ptri4+uYc1
6qSazPpcpLMaA4I9NXP9Hwr7Wj8CHZnFqIOf9lzvoFeCdejwAIPUR6YI0lkbKw42
Rnkqj62pY6VhfuyjiM3eZnYUgsbuQ+3b0sTfSIUHD+vWkvGzcDllwm7Leg9WKefs
Q8g9H8rQlxG9G2FZFrb3opOs9+KQqpaxf9uSzTu/MzF3FdVuoDmTIGUjufsTBHhy
OoAX52+SsA1dVZ4A35EnysGWwdPPhzFFRsYU5g9ww9EJnVXs61wCGESYuh8DqrNW
NYb0ndgBOgppPoMgv8YEmvik7d2PK9AHjBgrM1VdZgRe5OJ6qGXe/iGrdGA1/1jH
kPBA4Qh3nX4PjYcL3xSL5BLIHsBUXC2qzAyJfkRb9E3ssTGCI+V8Tdzo0uuoerF9
2sPCHCylnMZD+ryJpR+K3K2PhsyrwXkerCmpn6OZmR3TYISKWL382NBWNQDrjfKs
aXeCX4tCPrnaR7TwPhtKw40F/FPkogdqmly6tg6BtR3R3DA0TfQDb8Qr5eMHop3N
+UBcaIQ+aKb2emtQ5OUHCcSgahOJRvML16ckcgsXA9jsD2pajL6USGs5RSJDKI58
xXxwdVCQTE+nV514i8hqMro4BfTQrC1hdfIz9LgBV3A5pAssB4urKY+wH4HEHIBb
QxFsDS6NXkyKnn3XmxTEl2TNAuPHiTkFbKxWjbiSRoQly1Z0afWFQdvX2i0pv6DR
zg6u4uEE6FWihSOVqrY4hvtOPx/SLs8e6xlglAQoh/4BnqUzfZLoc9l2f8KCoYNW
6HfksVUAtnJXLwpcYEhk2jfxYVqszPtimovM3pKOvAO9qcqXHYrU4y6YRaTnAtC4
hzlPk9M6KSBt/HWwpkheHaBS+AQXgTutLeu0U64TNJU6QAypaesk47vwILXe1o08
4+xEe3LxQX6a00MrC3zBB98wCso3Hd4VvPAX95G/NNqKfbi359zXVFP9oIFEtwmP
dzLgwyNjT6r9KqSrSgBR0paAax/hF0yTzxWdc6SAmchE2MD0oGZEURrft9CU/mQg
5yYaKYA9ydJAxvP5/VfvWT1sN2jVrGn8Y373nadhswxwMkSc96cOxABZEGkcEtrk
Ol+oKcNL/bm+iCvHmc2D1CjePfqXHx8YZery0FqE6sNIYn2hcwBuCmfNPsESxPEG
B13994GxFQXfUDjQHY0oSfGFbHogOR9bE7TdXH9/9amyq5R4K7h75x1AKqpAbWLZ
Oj2nNqEOVqeyTEOcGzhBY/Nvpwp16vj3mkNCtU3kZdhx6jwNxfbXXrYddZXtVaXX
AzjLlkfJ1qhEbXtgWiG+Xo/PVh0h2BIUl/MNWHBVytgUH6ub3VLxYixsnKmPNE1n
vHW+aS8R+OXHZwSKQtaQkAtic7OSSqf4QhEZGPEuYWglZt52RVyFUrVeRQj2vV+V
VNobwKHtYEyl0IuUeCTRpAbchvvjx4mhOtDLgRWh0KHepMpjhJdaU2NXdzcmDG9/
IahpolAoF+nCIScFoWB0FnA8an6FoRSg/EfGY+R3x0Y8fyN9Nidre1ro856/D8sF
gVu/rnTMHbkWqVG166G1eh5PHEim4cRGw+amJrMTgA2TumILLi60ZRBx46tG8SUt
AScIRaziROfEisMavM1yEXFlclg/34e/q5OdVAq7Y6BGWTosJq8311d3+GXkVBVs
hG1dmm42vHjchTJVvkGJ6Wbhyl4hzwEDAKHsqeDKGmtjp6aQ2q1Mi8itcksZdbq0
mVxAT1kbdBtmw+CqjvIy9G3pKXzOB0nuYRsH5Or2ERLt/QhdYhe844jYZ8gtqAFn
jUhLGfhkmWyl0ENgUKC78S39c4rkA9X6Mc8qsZ4+Whw5woqMXns4wZCm+qsTrdpg
qB1Vs9KFB2CdoCdHahrOLoHB9S1+5K/ftI9kf7BCih8uUa93aVh14NrO9tzgBLhu
TjRI7z+eKHznjZlfUmuHQs5j2Jx3Yg/J/1W+nE8eTCxh8CajbJzBKXUqmoV06OZI
YuPfplaDc0nM9JOmc7eayO7uOgNJ6usmDDcBAA+3r3IPa16EdAI2e9cXfjDmuL0T
uANm9LS3/NBsTgjjLuPZYX9te+3HoGhZJDBZj9wNdyY52kUx2Dyu0KVa1B2ZQvbl
LSPgPHtMl28mpYsENvQjDtAmFLqf+OGsWybi8Seap5teSdVDlcaJv5xxpHxvMDS4
YUkC12i0Ry5h7IT3d7NGQ17u1+YIrbEmRNWpOvSCg1rpfZL+WFa31eYRW4yjijJJ
dQo5EYaGccZ+ddhYnqEGLUga5qnmq03711CRPNa9vr1wSmtcdo5j/tgNFtBx5UOi
u8zbgJsqjj6eCUOOU+8l271AkfrWKLRp4Wo70kqCGkQfQ5/+d/OXKnbXKaGsc9QQ
nXI/dnBEEPRp2GtgnsQRks2YB/0syx7Hw52X/C4W75VN9DFrpeHbvsW27pPCVroP
mJbTTwUihwU92EIEqV66iUGd+8NTFNrQFx7lSgO5gjFVe71rBZ5JnPJiTWQ17jXB
bcyeyNsFkVgAFzxZT424FdjKEAN+Jhp/g/MvQd4mogAHep4VypDRrcCGoR4UQkww
F13Dx5EcYoJJjwnrbk6NFFomUJdrcE2xrtfEmxGVC4DB6x72ZPmA8rPjVE6jjYFv
oo6WbwYtVMz2ggKDI2IvQvaaSj+vD04jvQp7QailmCV5TFVjbfvM5dlvEW4T6Gm9
rnlBV2bSmF6TYuBZbJXJQaRUES6L22BuflVDGvQ09GwDtnW+483xBf7tbn5zqy9f
tZ7RlNhAnyglkNBiTB6BmvMIBb+Fe7+pLqK78sMAo19vmexWokykNb+8G33kI/ix
LctpDvCJm1sQudz9jpIQYmBCZBsz9KFfCE84BEapabdOPyosESPtm3bcekwBfqAQ
L0CAZQzXhas3cv4QGErKKFxdc8wFJXT9hB9lnESV/kfKtH7gBuioIWzK+CpM1GYM
lQh2vpzblY9GqJjdoLfy+mnOCXQTmrOGsP384NtQ0qnqom0nhQLBBWDrsxmJ10L1
lGjvoHJpuOOGKRvph3tPxAUZhKGVYEG/0wiOp6vUjcQsAhLZ6Rqa1IFiZivcQL/c
evyMby+bsXWJZnJc6OKkA5gEx+2GREdQoMrQF4LzF+oJ0W4KvfDv8koiFrL3l2I4
Yc4MA1QuNcUi/LySg7W1OV3KL1CTCEM9ptbCLMeayDPA1P9EDMZhse9DigFzYmM8
w8foDDtPN1UNRfCFgShar+TDU7QtRoN2HQaE1tkg06YrRqtf6B72izRVe2CH0rKc
5XDU8SIo5NlI+ah/LGU20v8BqmHTDp6kYFDFF4ijlS3O+8PjZPWXQ8T8R0zoU/ml
lbMS45QMGbjxNUtmOS8lnWjIHSvqWfJzVymBxNQfQAsfMUfxIgHVz6w1FYK/cKb3
jIjNPan51GHNbV92rszvIzId/w5s/JYflUSXqhtoAqXNPtPFP8bVDZp0EkqpoAsO
4aVW75kFkhWPieyU2Xpy7TgkkWS3OmTTx9qQXc2VazgvJhSSjXwxkfbhk2UN5yFT
h5gErqXS8FRY9uUl3Dse/zksUcWNJXPOjG5IxMLYTRyOfuQs0b62+HUMi6zGf74X
IUY1hIXMm/dCnJZoRwLLQWh4sd3GZtN7KASgaVSY9lzotCw7smW88G3H8Ine36Tp
fkX16AXa8lJafz2kABTguxZAGho4RqxIB2xj4jheObtL8vRDQeLnsuyiKOFaOMrs
skMgextOgXilXGQA0U+D627n8o1vZ3w2pW71NjHWZ2FaevRJYL46BCadaNZNZIQV
18oaRoY1DXxH6s1frYzCowSpvfPqs22j9KbkavtpdJJRFeZ2um0uxRlzerH2eAbE
qvsYRCWipsj1blzvWZcRIe0JT87qQZOGuuRsAcvELWcI5bg1eBSn8VEcfJb0KGA1
5m8kDOTDUDM2eLzkfktivzCkPILFxzzMWS7Atg8apWutrOzI6Jquo6BQYWvvQhHe
C8BrYzRtMYKqpqyr6v93MyKEvzrPJbsYkr9ZSYxkTnQIT18/qnh/0RAojuCC/Du+
QBar8afRT27/AERhVPlT4Kf8znldKre0xZNq8cNJ2Py6pRePDmEIcuLwZOiJWYkK
DEXl94p/son8QTV0zjeq+t8OcxTI2kuxtzvflm/tqvIZg0XF8u0+CPyBLi5Ha/Rr
OmkUxTZsgklIoUsojASlZGqOnzsgEBto7zt4VaJa6rB9+RUHdmXcFAFcv/KxeSn4
ZfBJLNjkaNu3Jh0qB6ZZ+/Wp5CyLg+qYYKhGAYMdtZ3bVN2w86uGGM0ow17IiNFD
LhiykKVkQ5TGsHRze8Kj00yAhCWCPltj6prVnVTOzHA46TJp3GeLBuYlW0+hXs/4
WYYqKmsAJUvHC1wD32XgeJUElKWubVb0TFB6eKSNIFvaRefs2hCRM7S6W0K8BHlR
CX3i1nYjObInUExTRorpFeP97LTFmBHpuN+qcMWqWDs3SVJuEbWsxVPVn0LmMS6O
8SiVGhxNUud3MgRwgEPxWaU9YdZXm/cIVGtJsrUSo03EPXD1lE/MMozPUvd843W/
dES2PucnzYRRSlCd3KPIKRGr9aBcTeGTUp1m/LaTnaZYUzAaSTu4ZfHkOK7Cu/XD
p1EUmRMCnbYiz+MpHcRfj8FjXouUUtyS3CvVflOe44FvdflnWzyDYFAbVZwifEdq
J8LFn5QHkkQywH336YjvxNbe7tNrK5fezx8aTqdDRqX6cfNDwoMRPYIX3woawDAe
awoLQQqBqLLfi05TeJh7ubvMnqUleqmNQlXoup+3quynRM4rTiCMgr+AYjzrCaNb
oMnzdVEzBU9iQCbh42qw7zbAAJj6+1bgZo9y7NnlERYiRwShs+R6Jdxw5KtDX96Q
/hHZK5rPAtv0RaVQQnf2ckSgcToW3Ze0u1OotJ/JLw3qOEp2UMA0Ji9yvtg35Vkz
p8Y3DpMUAP1x2Dt0R0Yq2uPLPcaGU+hXBZoMr9S+3PyN+PL/7SgwFX1OceNfMTnl
WYVgMMPilUipF/+WQZwAc5YeMxMJU5o17ymJsRlY9pde2dgWPC5kwKefs82auA7x
h4ndq6KBeLuJblbzeTNabSF9rhwAHC/UMZvi8RLd+gFcZxgURE/kWMRueS/ecWjO
ezZYyVvJPbCcKz4gXwxq5dimDJbQBPDskxL+/fUR9aRlJcAan5ix3PtQW4PR2nGc
NFdIXXVWmneNR4cbeycRBJysTwNKr0Loamn+WuS+riL0umMWWRXo4wsvuz9txwqY
LEhPXesyc4J2OV1D+rEmXj1G2AHO2B3drbJhhBZ7derREtFJbuuB5L4LRTjq/S7E
IFAENOOvUisLXnqBbHwch/2uGVzqFbsLN+8G7Df4maucvb7e8MHpVALC2Jr2LLOB
b9BiOUldqrcp/9W8gFnaKWoZ7Bzp7TsuG+u4GSNFokWWIalmqWfDC7nPwGZ2GUgg
4MJhm4OrGGynIBq+2Zbee4vZIWtR1vAi7YXk8HPQe/aJyXl/HOE9yX3ufqFwU2T1
Wd27ztKzxjAXf6m1h3oKaAswUBcj+DQOZEyrtqD+8TuDCDrk5FPwBwvl07mlo+9r
WD6lymEBf/1/9THPEs4iBzgZaqwYZGdRfFlT3AOTRi7ZmZCzUETShQE5/LKJ3Pyh
nEShvyB662XLY4llEvSh+5xNvQ7/eiLAoHb78XNw+Om1BczImzTMlqvOPD9R+hUp
r9hKC03eJ6ckpm8M3GsQiZF+Uz9Sa8/jFENTPxDGPJICv1DT/n83AoRamswmd2IG
1a1nYkilvPNeeY/3I4UeoZNCyQpkIvb68I2W6NNO/W1VTBb3LL0VXsT+b6DgkqMu
Mc7QgdPpGAIn1gGtZYMwoGfdSiatjV9bBFM5VY/yhsr5f6BSWbLk2IdflSK7BTam
SNb2kLzPrLVdTICnfn598OAY/ybYVb9t86hZ8fKaP5MeNlQYO2OiccTBBbUlhZYD
wUoLmhM36HERB2Uu+Lwxthc+GJTpV487rYTnuyASBQjt/ut7Aq9UGUUoyeI4gnY5
Lz8kGdXBLsl9gxZo0dyNIqZiSTtywztXgNNxjeJyC3KW0xNyvNpgy7/Pu8RYueZJ
bqk90ylGmyAbvxjINwmdNoF59pbr2CKx9bHHwOEq96wu+N1ZXU/KGFic5A4WF2kc
6YcfzoNRPLSY6HcOdAerN5Swcf9qsgdW3y4CnIXeZCYRzRM1K93TZjJKXq4ZZCtL
wdpEvso2ijT23GC6Nkox9oiZzVfzDG3BuF6Uq5dKkgkrwx/m/tGytUuZXE2KPyIA
HkxU2m+nBd7NyaHOC2ziSgZwJkDK6A4hcy7rsi42axvF8YJGTqOawvleKpZf3R9H
JNOn7E1yEE/nSij2yhL8homsRqfaXfToqx6iVtG5rAobXbvAxVic/FAI+GQyjfMg
EWX2W3ATK54xPjnT4BDB4ErxK/SqK9cXy7lf0AWdKwKLLbNjYAmVfnek/k0Rum08
SrNDJEDyKUJiVa6nR9B3Ml9xOG/0kijsvabYefD0RKb78o2SEd3EhxWPo4DqEQcU
yktQy/Zg+AiFq3v+9iw7fTqdrlpfQ7VA/doPNkjwIk2IbVMkix31d3oTIEQUYwL4
WWN35386UjwnoUF41b+88ZwMnSMUIOgLzkgeoE1z5rPObG+Cg7JJCzuhP9JMJ+OE
eZxRRB7z6Hgy7pLyJ8FwmhUFE3Ra0RlbUWVH+SoeZMH1Wj9iSdAKv8VXCpisSDpb
8/5yaaSEWzrnGx2K6K/FeuiR48UdLjH35ZtoW5BCO39LQZpgKibCPzWaK7kWcMW/
hGQhf+MT0Tq3rfAAJOr+gt3juAuX5zGLqfNyZsq5nrPZ1S58V9aTNvGFsBZbVXGP
5MD8h0LQcCvKvDhKpFaFKWxGjjTU3MdLuQZQwIzhyynppys+wbAu9GvyabqOF2Hn
J5GNnadqW2pgOWMgmzrI6BI/5BGuemt9CEPs1NIIu9tyfoNA2Tl2Abdslf26+wNC
u1p6QMV3lxFceNjF7QQaHgHzM5jTH5dQe0kyoGIaBQ7mABZlibJDuzyaVArhfMIP
AR1CNTPu3yqcG1N+vXSO4KJyO96+IohuBeSYisk3ogeV4Vwh55exlylbwAR5G7An
LZvjTqHWQ3hUEqESeYJ0SubpzEH+O/MAN33u8NXCbdwImwW6rLAZMa3jqdcEWL2o
S8t6mEOkGejLamfpyEKTwE0LR0tujapMDjgK3His9KwjkaBzeCIe5DqrH2F4FA5t
tSyxrZROLfyyy8GOFz9fYg79sFO29VtnZX4KaoJzUbXbAsjNkvSoHPIqB/iqQuHq
FC0QxL0B7ItIuiV0B/9pZkQN6vwVyEpMuxIXU7i7KjE9HpqT+ziKCWRqOpNI0gw2
8UZXPOkRjhNCMNr493ImoL3uH+mZtAyquhoM7HBUJjnwqFGCjMfh7GMkSEzufizr
nReBun5CPp49RfUFBz7OSGzBANncWizt8ThUFv1YYO79v6sGBiwV6bn39GXo3Ms0
nCpON6jF+pAOP0IY0bb4xHD1VhO6HU/An5KcAgnwBmFsN6vUqBSFwE1kXSQBGd5S
x1qnc+G4uFn7ASko2EbjKLC65uLbT3N+X8EKNl11EURN7NurhEgrR2s6Zz0va65Q
2qg5BBg7XMMT7WOl9fcRPXVBofpsRXA48NA0C6XFAsMftoTJmvOikHB+8fNIDsb2
j+AQmrGLbHtr5f9qOKnRsMESI+jKJEeZaitwGvEavCWcIHhP9Wm7TO+fY2+1y4xD
mIn20/8LqXfyXLMPdyVKWrddZsx3dmMyQg7u/Hj9A7JTGOLXaUJJJ0a4YSHZTXiO
FdEa+ij88AO+NxRORNZ+j4KJpJtrOuhuZW8/lnxoq+mTEkdhOOCChKCugY2C8ngV
jVw/d3DBRd2xYiFudHBrJCAVwwA9DEu2fIFwRy2k/R+0vW9LN6RXTaO52gph0L9X
C572slwoTF0LUIiSbBxzKDAhw6nZVIFpT9h381DJX31WwdDmlVgkWsxeJepZdRq3
8WtlHUVp4d6HTQp5WFhsWjLMsnced36saa+z0TtZsGPzYAs2ykD3X+lGva8Ogbl8
LRNzcFBRD9w0QaYUalzUhbYgN6BiqMOc/AfLeTJYrrXZbELX9j7VOq5pW+6H05v/
H/BYMVVykkBTY4Nf/NO50oygXz5JDbMWwjE+EgJUehd78SnJ2+P18anxCwUsS5Ew
H8Ws8vRL+i/0KiaU2dZ840Sr25Odzng1ssg7v4WlQqgxz1rhyNaeHcG6lqdEHRls
/ltIMIRyMZ9CtxlXiSNVeakdI6ufdoH00RgonG2Mv5mUUWlT9gi7+JpqEbtkUKJ2
VIL80jJRYsfhjwfuuGXBlGWvHcLygQclIjbUDr5fDaoq01C3WJt6SUy9lP/gxoRp
KhZyW3lrGJiPETlKDvdXuLWUcdgaw9YX2P+5q505WPOVreqo1fYYz9v6yj8KYtuT
KtmAHK4A0KOAfAZE0mKfz+aBTG6gKp94XZL18px83QtGw3g62pEg6es5TxvHKVGH
eV4bsNbp3GBYd8b4BJTw4ua9XxTbJCSsKWmE27dsN76ezPFSm4FIiNQ90xzIX6kX
YeE1yUCCffmmBCEeOhGc2XXTvCDW3ayf6e19O09ewitNFeTVrAvFvp4vend8x/b9
Ca1hh99Xez5zs3BXKooVDzWxHS/5o/hTSsgR2lHqO7mdnXBUqciwAEmeaoKxpSlL
tUtOMmOirNqfc5vNCKTvNv+iEMevLh1Q0L2y/mVrRnkcIfKGWUDgVcK2j/ZqSEs3
il/WAfUsRuRQIl2fYk6y+BThHKEXSTsjRJsSftsSJNCfLNDx5pTPl31tR19a5ZPu
5X38QwLvU7pjbpkhjppXAdZtaf0T4joVP5ky6NKNP7G+nTWFbYhPEVdWqdD78mKh
Ab/bT6bEuJzprGd7lWkdppzFoEpKUnUXxMnsHPXBF469fCd/NjS/vfPHHGWAAyl9
r/Wo959tkNZ5hj/QCoYDGEaBxUFoX9p0MAIBhUFcR+8vfn+DXxVGkdxq9TSoq2vU
HiqCEBIxIrDtaPv88KV9DyEbGll+K4Fv7krq7K/vau7j+wLCpmy7dVUhf9nXDJyu
/BQn0SZPUNCtHAtdUpFoR/MomO0TwP+ZjGsnyxgGzPBY7G7aKEPEyNudAmWhnU87
lNJk/BiXrbuj4PDeKiRYK1lLNAN+BUR1GlMOaEninYtHz/KTZfcp1gGqExRBhbxp
9C9lNXvMA7hSFeZ2A5c6kVsDtm52oZIEKLp0nzIo4JOe6VMAF4Z7Udiuz2Gf/ZWh
rlmXdJ9KgZ20j0xUO9jiw6s2dHpFr3NVrRpfLkNEC8Aff1ZJ2k4JRXROI8LbrS4k
NzVwgTyWdk6gPJsnUS+FrLcmzuxf6V/Htjd6X7JAA7EMgdxw8af69EbUcdHC7j/l
wscKCwN9BAn9rqvFkgx5lWjxd2spP+DEOO+tfoC0uJyhWck9LWzM+F9qTfqPLpMv
2Jj84chFAdCewMbzwdN6zN0O2m5gIwM9LRqmNXdWzOZoQqJU8zH45x7PaEvum2Y/
5wqqxyShyEAQRhMk6+vfotFu5ZbVEy4j9dmU1FC7nvr/glQha3DV9a3dn4GNdIaS
yH4Jq9ZS0tIHGgCLdf/9qNxswwLaU2b8PL/657sbt27WgLy6lReXmGjHQl+k8yiT
BO5lDPZTpazmSTkqjRlveI/hkVF5yM2z/20OLOEpXC71Vb1pNoJrDR27SrBCgcFx
T+t+83IZvwdEqLTVCFqcW5pBcBklWVGFYITljCZlx8Ysxe/+UUADBib8mwPwV3Na
VtkMLuAy4jA+N6PkDIoAMGJZscxet8oK4C5H4TcbeGjSU6b7EL5VXLmbia2zz6xv
qPYnRnZVNY4khCxBvmA1+1oZB+doz1FeMmf2o5Anb1SnLMBfTvGr2UTNzjB1WJXd
SKBY0/SHY28UQgRBXAxAwUhgkie8LuCjvUMFAyGTVhAFluKaFA+dNtalYs+bUasf
FV9+EBai0JxTulaW4wLpSM83L3izeYO8MHDLnYcBy6AIBgvYrh+nTBle11BX8+6b
7p1Sxkb0a4fO8jdxTiyHZmZlAyMgBkG8fNNHr3kReofI0Tkpt3RftY0+LBhmnUqr
NVkWtV4AINq6+Du1/WX9aItF4WtZctgho5iqVQFOpzcj7lEcdmQKPvtt8Wc7A7zf
LspDNnkryHhcyKPtHzpD99YZ3yxBHeOaGGnScCVeUtt4cGzrcIGE9inaxlcYKYfD
T5gTtk/4gMfPe6FwlBxIlTqMFKZmORay94tvNgL0G0lWY424+1rFAgYYKviI8R4F
xRxSuJLcugTXcdRbT6XLvfuZYj8imcuuCrABhkjVtah7t2UEMlOT5BM/MjCs9jcW
1v60J9ID8uXePnH+tDuHfxeM7XVxr3Yu7gojR/sRGetfAapCZJzZA3LcHl/RyGrQ
7apa/qUvPEKOJNjspxez4IQ28NBuLNe+tkUDqTNGlmoAdKhoVJvt72Mta+BdXQYE
9jivK3NdCLQoQ5alnJMTRhHJ45RWnq5J5fhMDPUOQ5H7McC3qxnS3gTJrou0qA0e
ji3/19t+0bXj8myG4mTLlsfFKWqqZSG6c6aWDSf3oELnaw3tgKOY0S0W4dsoIjaL
LA1o8EmOqiiQ9j604Q6deutEm1T6xq2R/hlUxpnDtmNgS89sYv6miZrAA1lWfrQw
/jmjszS8TVEIl8Wb782aeeTygOzqJEL24ud7OVWD8HKDouk7+0E0u1M0MYSwLOdD
5uz4kBPECa/PmDQRc9MNpWSd3UFDz1Ort2qois6X/Ui4pbf5+PRZ+uupafHB0rXI
a8ys/RioOclPw0KpHPQ3uwNbgBFOYb+9l1sqDYl0j/ETf7IV6XhA7YYRe7QKocJI
ZengPrdW68I60fF68Ca11A3ik+cmcoJYelT0fNghWpjFpaWBfbZAHPB9h5CcamCn
5GubAtoQLpVsjyhc8r4CYMFbwni8JAoozvc/v0tAiWkL1sEFpU5T2RC4BLr8kp4u
yUAk6Ap6RPP1PG6gZpe9UIGPNi8IdJkd3+8ZpIL1U3Z2qY7ZsyLb8HwHvVhhxdPO
XiIbZFe7ItZgsuTBRSA9uqetIUDsnZlfIucJujysx2lJKGyCFIGoKwLPKBgnRBHd
AZELyulvg7DjCpZlKplLvEluaWElc6AcwTAHl4D1GKdSr0ZU0M659UyPsruuxf9l
w6M2EryMPxes1qccM4IkxVtn8W7MOqusUZMC/VZB7kJgEKwcCxK/tjuerV+tRAQq
7474f0T3MbH4y3b1qoAFXdSRvGbvwhjTwL6+xIeJsqfGIQ4kr80IeeUfOmAuIfTl
SyzhZ+vhYX3yDFIJWPB9+CsaGrYOy0up0yu3x7l3G4i7oHr5z7Cy7NjLanTSNQ7u
IeIt8QGyUzpXiKZ37WDrhYimHOWdEomqMGchBMWhfhEnrGJpDfMQfmTtdYbvvd69
s/b1tZcTGGzcxRU7BTVH8PP9r371sHLcwRuLlD5MLfiyhvtwXEd8qzQajukju1OB
ayENFjM8HsuFAQTTj1xON6zn6eg6rtF25D/BqQk+hR2OFPCIQfamlsXLK7dpi2iX
cG8+WNvabcfAKTmdOhZg5mLx3xCIf6kOyTYA/nH8JTVUL8J8uKlAOJvDuEjJiZ1q
W/9Gni8YeMvBMdFBKdM1m94XkaOuQcyioUokC6ru4BX9zzqtjd6zvfeZi99YRVmO
KJUODc6jR3jWqTlxgFhH5T+o0u8UwYQsSvgC1mbEDuFpnyTvUVo8InmVTBPaQZAK
+ReoterB1LUYVRD474FtLEqF6GAc+HCLIi9nHDxbKLIjW01YeGR73A3H3dg5w5R4
Fx0JT/qfqL7v4plpoLHUJeaBNU7AcDKI/PQNjEgB5q7Q1zqOokHTd0/lIbXY2PC3
r3TtV5fDtAlJxFaGpMAp/Kqax699SjAE6XRWHCpCFlnelMTdGhsaoLml67zS9rzG
aPwCuvnvGAM3tzsOYrfQKAVsyOP4/x2DcNG1aGzCEC6sBSafSdRH9DRamohpLa9+
0tzmNfnWOKKOLB2QbGqoopC6yRTI1olYW0ukgZyWMgQ8V2BRx/5rZwaggn0Pl1X4
b6HL8fcHqs0TEMNDT9qqa+VKXSPdw6SEb/VRHcn7d+ASjeqWzzTkqhos1mP7Mcgz
ZEJb3cXZU4PnCEOLloll/vas5RkKWS3UOD2xNMhgiD8W+0yzrCCh81FAHgbO5TGF
1AQBW76cuApAU4bNtR2t+NqvasAbDVAMjdo/DJ8SZIeERWqqBKkBd5ij6pkRIxQf
88skSOKC9WxhQBm4WMk6SjywUl0YLVP4zV/WrOo5Olgm4IPqNekH6xl3PoJ940pj
wfCrPHEQB7Mv/Y7vsTjD6sJYt8ZcQVAtgq9HeR+RBdxjMs4tNuJLoZYz+JDD5vgK
xz1f4UHx5yiRzn9+jMLMPBB1YBqguW3r8CFMviNj9ydOirfISJK0O9PTK0Po0l+M
G0l4AduJi+CFNw9ke2Kysr7AiLBTHBe4aYHCqCWy8UwZF5Cg/aMyYXbAWV82OHFb
DeEcdnd/NAcZWC9qrPkE2gksgJ1YE8QxF9pwExFlI/MlXzBbMjJOdfq0AWg0Mv6A
N3xnrj4LtE35Z7qUP6VNu4h1PR9YfctQxsBViPQeZ7LvL1IomwQrJ91gLTk+zece
+qvOGGTQjsccVK2ZmsNw3BTrGHIuhnNlLyQqFdr0xJB0t2EFcSbtFIzmKCXAZanY
v62rtfHpC3XKVL5KQtY7Ut6B2w89fMzqHGtX2OaV1UvRfzxFwIcsUn4cSjOT9eB5
aURrkjnMX9wYQ0jieuIpzT1GYziOfn9ijVcjkU/PLMo1rgKAcT/Ati/XbnYEQscu
QNtVI7Fwc1IshrF7LKmiGRylkQlDc78qi1LvsD8VkWG6lcrnt0hWfUa8BAdyaz/b
JfquiIC9RPyyGMTuT2RgV47w7qjWEC3S3QH4Rmbh+MdhYRfTe0hHhiR7LXyJ3jnS
x1UfkJ+KhgASYM1/SzZLnxit4qrBaBK2MnGWP55Ek5jEVaG4RYxK3x8i0pv2vBy2
dCri6UIglK2h7ivIgQXKBjEQCBn0Io9K4/MGrgp3Tr31BSrO2ThCfnsCcfsiPRAT
PNLuvhptJmpuk9rZOOZ5bZnegOsL6asjEJY7MCQ6lyw78C5otnet//apOKj6mgB8
iCDHMorwUv3/fE1115ln1kHGavCCKbBkW2MQhDSTe1+CklzgQ8TVhznalnyI1DqP
L11SeFMf9k7GwDObVsKs1LV4XITYuJaeWgQUQsxNub3V8rshYyVsFtehuGy7IAkF
JxscWxY+8QqBuDw3bxZh6TGcHLTA/gk3vt8tEeL561BTwo4N9/8qqxm5Uego2QlK
D2corzREcTnELHbbVHuA+fBZKgiHGH6pH414xnhtKUX1y+Wke2mgG4p1BdV4+htl
3nktsqAJ0zYyBhB1xf+B72fIe22RxUx8AZBAtK3NIp122isWXZLZqwba21A5MXnS
riPzNroo8u+Z10SnWSP5Ip15Xh84uiXjTtaY7LQi4Zyk8dqrRVoPTBTeMtilUNey
iRK1dl1Enkz/cl4B88f0Gd4tVIpYfws4AUC7gbjJL2yNjgA4hCatU2xwiOcxWBVa
9ckbYg+QiG6Li8q4qQDLDTXv3F6ptanckY2EuaDKZmT6o+OCug5oUidHfr2AOa2Y
odtoYBrlo1sbOXenRTf7bKo7/NK3CtvExeVvdlMKVR2NOPFer9SUTbSEZKp3DN/c
VKizhNzEiErJrASDAy+FpNSEotw4l6B3v41uBD6ZYmTvjRQXNtuKbHTkNoE3LTcY
j4yt+A39TmirU5c4us9Db1MZ2JEg1v/nSWq7WITKWsAJsAV+5fPnTRC7+DmGXD+r
1gxPFRTLvvTWh1STlASssw2z3gQvMdIaFcvZm09/Gt4YvdUMzDDlxeAd7s4pOwbz
aFYiv4e5gYKFujenj8PxzlYVxuEF1h0B/fIExjduxfBP0JR61IokzmpMpX9RJl0y
jqLpNxkh0e8KXJp7IffD6H2pp8y5+iNYSrGj3bvRHh2+Ok5LPVZ+3xql51BOWBIk
9vhTKd6+6mHjAzU1hNepvjMHSrpgoQDOl1aHKptz1ctT/pNYACngGOhB/auQaGyY
ZNlvfhgelFKHHvhFiDc6hiHj2e6purFZlDAzc0M/QwItj7MraqcLbvt+CITHqMx2
xDXYGtoSUA52vqpHylKT3wNYszdyXEiwXIUVElWctfIqkEVhtyMBQqOH+fQXLVCz
W7YzEYCJ9nBZIh+ZJP+QEeFhHT9v+NWwmoQF/AJ4U0OGzluIuukNq8u0bp0NHgoO
zhSSVPmXhWbOC9l9MO+n1M+q4+yss04MXTkKnRmStqxgQv7Ujz/ZAtnuKswzmGdp
55GxbIZAt/bfisLbsRfQ1a+adepKIKgtQ4SNhHwhSngBNIiVTM5pX6vhYSux2aOT
+GEIVxN9vrGqEwRvwdeuSt7NTQDC5a2mPPYXP2rF+HxliLNpUyUzTXPzmei3voQO
dpSfavfBzS5w4j+kykw5grN90hw1FnaqS8wTYG41N3em/8Em0fBkmJNe9rGG8+mv
xojc47ZIHGPcXo1QeDj6TWoq91JUzcCEkVK110DArDmoE9xpwwP/J5kNjs9iQJ27
aWvOxU1RaccaR1FM+H3I8RGUCWPvLKeAsWhh3UxyaabQbYA9OF//vK7x3Vgt6lPS
S6wsTsVRhPq2edW+pt4W+TKrIONoNHeroXs+cndUPAZrYoK0y7CCWBXAUspDQqGM
YenslJQcO0pbjSGznnpSS709/ksVTn5Cab+VgTLLU/eGPjqdUlg7wVwwLAWVZwC4
pXr/KL8kaaTF1tkamFnMNswIyUo88FLcymS0mKyHldSkaZrjDj2tx4gGBaaFfcKl
cICgeV8dPZpgSybRVo186y2Avw34nTxV4TSAefxkcse2Zg8J/hYcENoyj44G8hhh
bFaE87e73TYOhItnlGYCd/d6YBaBOr9ci3U+a1Nl4HcByk20p7JGIbENM2hXZqo0
nt1Wf0S6MM/AyMZUEmDDd4qqcBDpLLDqfCKb67XkHR2h4oBTFTdQ1+eFLXUyDgA9
ZJXXgYMCg8BLfg99+xUvjrH8SWjri+ttt/hn4wpeSXxZIlxL6Cw+mETu/jwlohR3
BlJifSKLU7XbiI7Tf5zpWgeAwtuu432OUsYVagML30HBVVqs0ebhLCqLFvrLXvMo
jG2MAtS6jAKospMb6cuJclqVSpUewx4R+GEvYKBd/XmlgWgR4+wB2PUe5Qd72Soc
FwGb9CNuPtd6QuB24TTMi3HLkgkznOCTfZAdZ1qZvnQSKt+l3+BzPmvioTXgvZ1E
u5FkEO5IspPwj6udFqQ8YPpVxrQsBlt9PsEKimbBSEoH/IlPeEVndlfkLb78WDaI
4inj/ShKEk4ZEBOnuGgiHQTtqV6VqMAl5phqcls0GqEr4oaRs6vB/2XElZpu8rbE
Di3S1X0YTUlyB7557TRqAm0PnGdFCyfjbfBtg+Wt6ZviwYK4c2mWWcUpR2f89LSt
DlCsUtSKKGH11/Opb2ZxulrDKMm9Nsgoa8Ykhni8noWQyo7bPYhTXva5uy4GRDnQ
gnFgA7M/kf/BlIoD8JCVMydhRs1daHDrbKbnfOtmw9jv1RM7T+LACzvsFzp4wp1n
lVjiZIJpUzO6TTZATzkLJIbcdww4Lh63CQx2kPvaBdrh1JLFZYOBp1Rtu2FuBI4Q
jZJ/xLCj3XZHfDKiRlxAgU3ppmryiaj7Ae1+C4/0rISzmgcNiIhzcdzOxQaqb69g
GlvL9IFljk/PM1Z16SWjeCRmqxUF+XIAlAlGkiXvWADojbn27DeDab7l2rRoyYLH
gO8FqB6rsBQuGyf+UIXPua4hobRJJqUGmv9Bih+bWImwahDHDB9Layt+t5Vs4pHS
YoIwGndB4x5fnwQ6tTw9tugSZ3WLaPi3Yc+DIVxIRGNesAfxCRCHVQpd3gDxNFsy
W/9DUtrNwJwqEb7spUkqB3iMdoRjKnKPdeQ34urRDGCS5DMnl5RVvvMsf12LFuGl
aXBiP6cVpAG9Et/dh0gS2jG9GfjrV+s86XBaumqT7LMqBfz8VtgG0325dVQxdJ4L
SOCHbaRMO4Rv8gnGtNT44VqEU5UrZGB3/X8CIZSj8x3dxbp45vYP2KZTxwK6fc9z
lRpp847H/4oUEyUE+uPfJTebileJfWkXsTUcOYbNlFNRXb52u1UmKxXvyv/kQSRj
M4w6xTTByPlKzHKWgaKY9kSvNq8L3stHIL9EKMPiZc1/2lgBUuILSHgTfcO30Jfk
9vI7sMXBoU9UmXtyu89eOfYD2GRshdiSMBDUYIc1yWsu97Eha59el78csVgy6ubF
UBGLxuZWi/sjEhjMWiWfNd2K2Lz4wB+mFO3GiM1P6gPOugqUPl9gzIfQAFmMn8T5
QTE1kmA4x3NOKw0+Is85bFZuNT+l9aQ/i5xGZo6H9JhrLRDNtJP+j7pFvfwXVqt4
x+LHsR+PjxoKkGMcqwq7K1YsDkjW4u3Updbmtm4UodZ1Vh2rxyt4phn7s3MTq9tX
RTdtX5PDDIhN7DuJEHP2aSwRVsywaCH2nrG4lX+xCj8P/xx8bpJnkUUp3TAsQF3s
8AuOtDpPmI64Hk9j12sjDNtXI1AnRvq61/GZU0tQ/EwZ2fxSLHg8N3neh1KWJzDr
bFSC7GDKd6iaRnNhyb1zz1948Dg4ct7Zz8jw5sIY+XtJxOxlaxIE4DVbnWkxd4aI
kMFbyfVsa5ufZmckrr7A/YBg9r6eDOpAAeMRL6jaFHgQnu4SzFRl93xjuMULkJIb
E6tdObfCM39DezNl1pUXPDUfsZw/euWUOmaMFBG2vBvHuGsDqH5FzLVXoBpsBa6p
SYB4oV7xi64GUYaJrr5BmLJ4jmw2FxedJFmvhdQFhDIh4kYEzuA0YLU5/TqsFVxC
/QetkYtxB/ipTxA7RzXBMYewTvNJ/yt+HsdQMq+186tVq8gpCIYXM7SvexX54lfN
yDj7yMLaDs49qwGI8PXaOTcX6SCYoHf+TcwxrfF8BBQdrfY2XsDUjiawEND9X+BC
fJadTAJ3HOQto9XFzlYEIzJSeveuza0SLtE36wjgjHZlGlevqGcde/tldEtsAImA
Nx+uxsAAu/7gCpy6JuBETs/gkr3pDJsi5otDvd+NQWLAla+NI5SO+bIQ1t/+ecCx
twxdY1vtKr2hTnhezOSLo/6o4/oAmtX1SShevewT6SSqk6Wgs69HWpka2GbCcJAq
clhWE1CTvNnql4lmgEYhH7Zxc451cCyVB6pMhmbFo+a5x19ISabBNQcz2qQ2THqj
cEEX5d9Oq9AGwLKDZWIV2DfjeQA3foHbWa1yhfWlya2Rr2yKrnbBCIrvMtj4ysqH
w/kHHiUf3+ME+r0EN3B37UcaikG0tmF1eE3BLAmEwS8+fSma1ahhLaxvvCqZdUsj
v0yURhyKLTtSkZBbrQL+cg72MBeAIlTbUi0sheUanMUprKRCuRdn0jAzf6VMnug0
L3I2x+CE+UnvbwMOdEF9eEDbAtlBAf0GO7NqEMlUUjh4X1Q6Gm5vTvfPV93ZgCG6
6IbR471IkRWhr3vEM59X6B2Ent8NIVchHDpqCDYJn9z4RMgBEa9sQoZ/t4CinQ4H
OtKacTkC8LP83FshKg9oL6sO2vvsT/QAJewUQQLKyPceS5z8RbOF4Xo86EyO+jyp
5dhONpfzsJHQPzAzVNvOX00aubBG3VBylhvlQGbq1roD3BkIXPERmhL/zHKQaygd
FrHzkMiY7jAuPFdb/q+Qd8Ibf88n/XzoKQOw4OoJXEF3b61mBDrS0SZXRcVdlLMb
/cfd3YaDc8Yka+mwQffd1hB9L21lPO+TdNpRYWs1QDjYC64jk1MfQ9OTBu1zBmdd
8o/0tXhZxW4pKfg4xkan7kuP4Nd6DTY8y/HP1Rq+821HTmh6eUdm/p1mB4U0SJ6i
+XGz53HydKIRz8uPsKPrEykYYxuG6PvEAD2RH0WMOU8in1SkZsxhi6qSSyd887AX
9dffG5ibabZPr98ahyFqT6ORyxa1ZIuhZVu/AHWLsvY3S/hMu0C4Ud5IxTkZ/Jxh
nVPU0rukcUSkwsYnLKCcT+f3vHgn/0e+9ru/88JGVyS+KWHGlaGs/ZBzWhaK3x1S
YtG8C4HUQhqSRrnGOYcPCiMy+/xW0S8+B2Xh27m8mnSr1mMx3x2P+u/lwl3Dp5SI
dDde91AGzs00AzniGlTcJqkLknwwR12mU4ca3LOb+en0eHRPcpJPWt09OwmOkdvb
vEoHSyTh0QsqbIOhvOjItBdCCI2qYwiNvzRt3kYY7ptpzJ1wTyLbpUZcrORFXUu8
LYkGTK5X6mVQL/Qij1TNnrYh0YkN1bd4Tat7thb/+GC4+aVH4+Qn3C3YEU2eKMmL
iNkbT2Wg2HUMI9pxEuofS/6lgMvfvFdbM3skXW35MbX26Jr5HfJ4xjkwKkHYBsn0
lI0HIp5j2H94CkDJtm0gBMEN+KOv5uZK/F5I94uMnoAMRepffb6jeElYkOtoTmVF
29H9xVzLTid6qd1VHvSY2ceHnkOu2GhtWstTszf1VUulzScKPqTBCHaISZXI+LQ8
MNgamFYEDd0IO7NCOxb/0VdDK+ZIPMKxPVM0X5E8ouTPi2JsSGojQRSruWfizb7w
R/rWRgjqy2c5RkdD6hJGDvt1VNyuwP7bSczimoGx29JmYYJHq2u9K+qzqFUIY9Lf
UfPzqLgEHAyVGIZ1UxLqWBDYdX3Tiz52VnzJ02LGfx3/PaOb4NJIRB0mET6IefiG
dCRkF2xGTarG7YhkrfeL4ALoBlTMs6DIsdASX+VFRMnIgo+NaGugxn1VcGJGW2ax
cJT08pCgblZMAe5XlICZLqJQfe0wAVaFsF1NAxHxLJSRhuK0RDqoheu/g2rHCUdt
qBp2g7E1ekhNC8nNrITCmqV0gNEBDrLVNI+T1mouFB982hlibitltAPWK5xLw2gH
FEDuderxhd0afl2maBbuYtuP3nkoZS+OP2VzKhpoRVBJn7jn6LU241k6IWBuaWoo
ay0ElZMl7xYN8FxP7+8Qn30kfS89imPPOQGnVR4xS7l3/GrhXedQc+ZGM+I9Z506
QliQrWVFkJ6RnJdXdQ0fqQx0ylJeoDF5TEzlxRWBoYOCBCSL09uQa1VXyop4mjTG
FroHS52yLGNOlvUP5VFRGqxP9O7PLLTJAk5HfcAHeiQQh52jHxNTtQitJf5T5COL
F7K/QSOFsBwiG0OsYkSROfs4OiCbBgLdIP+nAeX1lpRbo2AATVkWbLc4hWqXAcmH
+ZAJVEX8/8K9e8+InTqdf3lTQJFwKOmXvg64eHVxeaRiR19sNvwHc5b63k6q2CVj
JEs4nguasRsfNhBOq6j5q7ezdH0zbNr5I0CEKy0qSn307BVmUEaQ7JkYI2jeCaRw
ACSXYaAxJRN1xWt9cJE9tBWNefwYCye2mo/qOvlY2HCN70DYQ2fRjVPeZnth2Pcm
WWBSBMvTn+D5B5lyZloVCb/hYDcmc3LMVtzmvplWwdHJLudMpdHUAiIN8jNlESV2
LFhVOYG6OQEazjhFcxaRKTp/HbO8nbXWBAEx2xH+A8RnQ76789zgyTTubsuEPBeR
91f4m2zppMQmZ5ZWG+SqNtWTx6wm44qP79mj4/fKljIk4C01N2ua9Ef5+3Myj4o3
cQX+3Al47ysQBNZe9bWqhCQCnLFKQY+rZOfDY2TESDKaukGnt+0BNEQ1gKFQqWiu
EA6/vJlZH7Ym7Clz1gcXZ2t6MLAhQbFoULtSIP0A/Ff7gQsEBTabRQX0s3dX/I2O
W1v/UUjdAo4/JO5mB3JeLb5KliHPFCXubBbqivIpd4Oj52vF+pYnpaCVAcQsQGup
o7F39YUJMs4MoSdVqnj+mkVX5DhFFinssvPlgVc/fnmsh79BNdfeSv6MamP6phf1
NPGUilF0eaPTcTsCy7v8PmdEysYjj2OMQUpRGh/mLDv4lQiaUE71iYk0cjFT6n59
fL7/eaxZIv+zGSBI0/drSI+m7WgtUjiI4oV1GQJP+ESiubIHhYo1RlBKqwuCvJ7y
bt+5F0PiFbHLdKUikE8mZmWALn6DGHr8yIzThn7NA1Xt3lBTyOfqneWg2VOJnxU/
GqoBtGS+sT8vZ/mjYxBZJn+bkoI4kY9NtpuL11myXliZ2RClijrRjeu7Bcwkf07n
/xVkZ1Y8o1R3bZKyFL8chlF8Si5oIjo8Hiocf3o1kUDuvOyRHYUhA3O5UEJyBCm3
VB/5H0RxMpKyqzUz/i/8TuNLWHmGalmRzvmzKuZ5s1jShMoKjHRQxqQvJJ+KHIwm
W01YgL4IV7o0eR5w4EUc3DHv/EtRiLzh4bEoXHfce9FFTvbi+lDa1njN9DHaE32E
F69RJCFMEgwaVD4YU8lX9bxSs0u7zAL+WrdJXqXgUmfdO9VWJpifEkhqXeJ62nuA
kolBTw4zQIE4AKTDyQE2ZapUGBg5xjSjEtb1imv6ZVu0X4BdvbT8zuzvGhO/DnAB
spgbYz0X/BxMdjg4bCNeyZhVHqfCoMI8vZguySxAatFe/eJSi94BxSRe3lxMWq6/
M3x0p62YzzV7d9JhA8FsmZRI7pNoFiNsKbSRNbewkdbYHlo98i9QcAZUVx/Dptxv
dpLM7L/X0ht8zV8sIf2MX1I4ZmP0fvSG4EPZSfwiar7Wua7SsESd3tSFjBycANPy
8MsPebkRMTXEEm2l20g4nwWxCxxqoLgaRUsGM8pBAZDnpkuT3SwprQ+HHS+pa9hA
0fn+I0AARIy6tV90EAx9o2L040vqxr/5ZBAhlhNuUFSXe0+lhhYeYK2m5NEkV9IZ
YF/50sZrkb3ocjse2uUICH1uK4FTl7B8I2AeMFL6HwOtOShELc9pET89ZJp4P9lF
zKOxD2DWPYd2F8Lgsz3jisOXcQfjbdvyTr3LXxC7oKTbrIsahuexw83RIyk9FQtY
Gn0VP4Str2/c2+lHBI4r/ev59rkHlx/1FaASU0jX+qWqbMF2l+YgoG6g5xpqTNRI
lBEmxG1TrWSeiOl3ZeQKZLXFLRMfhQWqhEC7qjo4ZS8YMrvPpUHmWC4jHvH7eF27
CEHrKdKjkyXwVojlILu0K5iNsbxg3NffiZB4eHFa7+5EhocYqtuTCsCDHGp2jBU+
fqY36hdxfNC0+EpCkJNyZcO8HaD62D9qRtKvp5NVLyilyfqqcP3bLSsatmO8xjUG
CpTZOn0cFRtqMSuqzNZWUeo8QvSnZJBLMSXWfNsBe8vUf7/cAV6B1elWK1HpW/NS
2CQbrF2fBqhgVKuiXeyEN7ydQE2k40XZOWp07MruKLWx4qjUmG9v0SUgL+XO3RBG
81sLfA4BsbmLM9P8Nd5wXMnqul/xZo+8+2YbqmiQDE0tABWQU1Kx6iqHpb1To2Aq
d1WVrre4W3dXYO3D8aOeXTA/Za9eTDxhNnJSSnIvjx3hBl4UtL9gf6FEPjMiR4mF
U+H2Vlk+Cn3XaI2zykg5EhswF3zEhJ1toK1HK9E5RCTrqkfd1M0ZyqJ8LYRQvet9
EIe7S4hCia/140DFIEuvHUzoMt1bVTFqetQaP5sT2DMDcc3Yo6p8DwNoelGh6gpO
m+cv99qOfb+louTzdtcHwyycsWtUzbuu3/vdrkNwNm5acDiuM+zuWYTMPfuz3FB0
Nug7mKOfeV5ZrpofdYruUC6ZQoulj8vFI17AXdFWqfA9KoUOn8rzL2ttbgpxYeWe
GP4+bI5fZPrKyvRScX6aBn+Fpt6zyQuQm1EStxwrnrjdlvT9AQOEDWIUSZaNc+Yp
G6NcbT50u1XlyxdT0ugGXggAO2nc/i58wAEKaA/n5aqrjJyBf8p5W6u5lvpUqvkm
t8YOi10i0hcrSBJ9hWQezTVNgBmpnK4dEX1rJvL/JffltQ9JWT7Lyj1juZDKiNDD
ZXV5SUzmscl01lme0zV0vQB+knM9FKtedSvYrK6P2ByBhtTEEARKS9ode4SFRG7v
Q3aJ1/LJmXUwHKjv35rX01Dh6OLjJDJLkkRWiSEOqxy1KzHwsHhLdRXPE5hm6D95
P3xYVxiCfW3li6aXtGx2QsaqHflH9sPql9rCirKiroLUlhGJRyCWI2q/vFSVp34D
qjg4XfGSwZ26k8nnGglee/2GmBX362RNgYX1WgFVexgKj7ehlk9U/W2NZNJJ6Xw0
QQB5ITC28C3h+ID9M0vyGL/WRAc7AJtlKbKmx3Hzw+OXr4p4sQ23FMJ9Y3P/ya0R
LaxdfeNheehO8wX9lTD6QwDq0xuq0jejJyHGKnpj5zSWIarTNGsz+VF2qgxejhO8
OEfuNksbjxR2K15+HZmmZFEOwtqTB3x7Xr8e7+nfYczOS/vrBRj0dMld1gagCI+4
6vdBdcM9xv9T56sSVuWDyYwL767hB41nEdqUHAU3Uq5LnNnbTBUjFguxObcblhQ7
FcBHeqzWOEegCdFn5QqI0B2FODkaCSCgwCNTijh181YV7h+gyz7atXMsy/CsI7P/
RTh8gjITTUd1ZtifjnR9DJ7kC51UEPCYBt5Q+WvxJVbusQFSmxlL9FKS0oz0Nm4z
hFiGtUQO6TkG1eGAvE3lO/E+0u6Ngc+YnMvYC/kJv9NylBjcFuJIQhpVDjobXcKh
jiNA2ErnycbD6+46faL3nYAWm5bakB/Ju9cOjBFjFTgRpEjacgfE5TKUXWBvXGvx
oql8RRyg5W78/7giE2azhMpHXZ1zl3BAfbXBaYKetjQqriIYQlqxKxYI+G/TTgiP
EQzp1QpYSiQ8/ITOI3ccrAxtFx64NFJPKFBQIH6pY51ulsujil8ZzbBCJxtyvmTq
AMgRLYxdv8/p1XAqSbLzT37komMKQMb9n/lq3obDp4wgDVgmh8C1juUJoFWxS8Yb
PGHWwIFkwRZADgxEp+NN3QQLFTzkFbjIkyt3aPi4dhl4kNk2j3rqLNY86hLOF/S1
oWix9tPZ9NK28agSM0p9+0Xzevj71G+bRxv9QEhg1ksweh0cuamj155+eQSTA0Lq
J8XVfrGzcYk9eETrLh8IiGThsfu3yUpH1WLnYTL7zJHkfBWNXtnWrOL7aApUMhRA
MZmd4KHScVkpsBnMNtUbzLrUhhTlx20sbTVWRskm8MY39D2CarEqoRZRdXp3LhTS
2DI3vtBc5ShaPNWyqEFCAgcuNMyNOTFUCfYkVOM5XnZD8cKXjCf64cumdD542VP9
uTXfkcZztQtzBkFISENOyayBtrN9ejmVUixpW72LlGk5lUSB4eFgF4a79HmU4JCg
QjCq3Wat1v+ytIJmy22MtUapCMmvNS7UeMthCgA894dwK3EmIuwhjsamJNTbRAeo
dabahFBD/Yx06FIbeYRw0kEOtwQVoU8wPN7Au+l8MjxSTTt37p81uni1Xl6HzRBL
oiQZ/Jeyfu5C6ppq63eZkBQQMwacbkgL9FBncREXXcWJmvxxizKMMSoOEwWv/e72
5+bkSFOuwDgKQTQ9tSAQ5s3bQNlQNFjGElbFNQGFP+6un9WVBTmcVT/e7sUmfkYr
b+cADe4S8llWtLLljQ+FOSMI91jXo/cnLrFIgv/JJZ+CP5Dq0lnSIePGMAIW6mLJ
8hYl6C74vC47vmf2BXZc9crbFeMRonqH3aMgIoEzyoq6i1hW1ION8Ig6YQXLVn/x
eKE7kvu1kB9RhEfvV7CrHIqr+AQfNKxO/AB61L/f8Vzjd8cw6hlB2sZQzd165QsS
YCcrs69U4BiQPgYPoyur1AkbFKpSUAaASo7wGw8Hl64FlIDc3ibBU4pxuy0o7Bwo
k+9wGjixzJ8Mrng3spaAR7ZcCd9KnnJKR7cWp2+w3EbF33lLqg0mUn3ufS7ICnqg
p7MuCxqEskbxSOOrhl7rny+00iy7Zl7ER5LoBk5qI4fCX0FgR1QYyF1WeIhZZo0o
PyK7fjDJ6SkiAbUPnR1lJl5b7L+vGwWRurVfF7M3J0jYjsTsW08hsRFF+ejur1aS
AzeWx87RPZgMcsQ9PQc7wRtLd70Tkm4r0ubFscZcCpKKTqDQnVpWMxACWVN/a5WT
tIX3AYjkJZCon+7NYK28sCeWLB5Go4aLruwg0eZTkJ3lLgJt9gXYamcshlrtGk7Z
g0P1lmJ3FtcP4YL3j3X7KeGRXZBxWblcWpGi+ZZRXMpTY4ewo7w1yNR0o37LCfZL
mO5EsqNT1vk+bwlglIwr+EVSbrQDByFIOUaV+IqTWFHlb5TBFDES2tDUjxR/M6B2
LL1BrY4CgAll884qsxx0M5C7pG7/hLsJ+DqATZWXNmsPNWCoTu8xHdxn1UlpVdL5
zqHEBpiYwFQzXZTdkEzuNrwM4pnFCoU9+qMiLKHImm7M7LzSyF2PePtSW6VSZiWx
xdU8r31w8zW6b5E8YFNjMTfGqcsFxIEmn/xPWl1WVmbFhlwHb7hqY0G9g3q/6dOq
YckGhspxfdP+XAfM9aHCMyR0wiD5uzz2VYc89I4/LtkZ9huIgCfJoF5JtB03fjLI
Xxp17/cwYi7f7YvFYlY/0o68zBB/HoFeeRZ80DhAoDJ3GFFUsbRz1MCYKYRNhbZ0
8nlQ9WkTl7lLu2F+lyPuqM5z4KcmXXxLOemIYQJgZvDaL0o2WACHi3V3DV7fIS0o
riIOmqRcx0qpdv9HbTCjQgi7QJzUI4+foAVft1P99zOWF2z+Y5qu11w63fIXTdDk
rbsuoqGnvPvXjfEBI0fKJqr8Lx+FnQnquqJ13c9iRZAF+WuQF/ri4m0WtGKW3/mM
GEHda9x9lkLsVUg/RI1vtYIY+iePkvQ9NyEM1w3unx9I8kMLT1nnK2LHx597H0Qw
ypkPiKvAkHAznDPDkIux+Z6BUdw4Zkicm0H42cpSj7lpk8UeCuafEndYvrY/SUo1
umTxDZ36jSnCzG8ibQw6bJqbjyrUiNUF6OLGls1WVPwjGfTNbxMOtoBqnh3Kdc19
3Cz1JAV7lpSy3ZSvqFLcks+qFSj8sPR63tKMLBKvA2i3JmtALX6QjFRT7dY8J8pj
HuHYx3byNCQq03jGMocDdOG3uc41ND5DSr6SXoORbztGlnG5CQoxqmDRwdAF4Cwq
eJzTF6dM22ETDGkK7rcUM3l6WEitu5YGmAwrIhjChrNBdLV068+8Fd3EzCxyIMhw
0BzUK9/FVXF37NakMIOzSFF3A0T2aQJAc9P9udmiSU4lHmwQkevJaxIfXw52hCH+
+EeA1mT9OejEo0lh13OPqla41VibEiCtbbh3MOg+xO0KrW0FTVs2Ixh53nNusor9
TyKYd8SZxuGhFLU7vrdAQYIUiGx/7oDPDl4ECNmXt6tJG6dh8/D2TAiKnpCG34tk
tr95Ez6AtzuXXzpdqOPe3nXlJ5sWXe0JCsaqImV6CMJGw6yLiD6XQ5Sjiqgx8jgj
zKU9KDmBWZiOIqjeWuQOI/kxzWZXvSh2moIIe3tA1sd5lE/AS4UfwFptsanXq+Kt
27WclzKAD97/vMgBetFbDGzsmSOuKvWUdNwN2X5q2ifQzYi7KXPdwC4fmKkIPNWi
ihPnHFsDHCVWWQ7ufAjg16lXYx3RE22hblzBWrHoOOTKbuE28nzY6KzYo29u3CgJ
A/bJmI64TRESnbNli/J7LeL82DRdVINqtKe0gFiNYA87YMuZcJUenk3Xq+DsldHK
FifOxJ6lO8I/F5GUrxjkAnL4OPeQ0DneFqkd3/nux9L95CzgXxGppclB6UZh3ZR7
YIJokaZaX012UZW6YHpdWIrtDDkhKH4Fc9D6gCyEbGTKkEHsax7zjQU5KMrfaLZb
sZordrNcn5cAXdD7wKMOoQioHsiss/LSQuFXO2exU49j9VEl0cS6a3KLkwgwBHW1
RJqjOG0L8GMF4aae24kCWe4Em74eg7yNBkHdZFseBdnQYecm0wDWxQLOlFcVrpjY
eDum7OZ49WJAoZ1OK7Gs/NXRVyTeeUG2nuoQ4ujTh+qs8CmKJ2/pI3o2le52KgFU
yLt9tCrD+Mcwc/ifVIpgUD91lC/1mhpBx3BLILOeThfit14AIpKPiHfS/m1PQo3m
V/UhuH3+aH7FX6oEAiwXMWGtF9dkrYt4NBQTZouCQBmlqOgMVb5vnjc6aF+72ZSX
9Bsf265xltXuT2EMRuD1i4gymCYtR+LznHO9gMwAEaLVY972UN7wbOg41T/Cso1V
6stCudwfVGuCvthOSjCKt3IYux7Ea1+LraWtmh1f7tdedsvwkAeNYJsPwgD8quYh
2ZmyWBFvx2/4nwV/7cTAsJnN2MRyaBBL+dPv0+0EfgD6j+6hN9wW2oDubH1sTbD6
JWoHkB+H+FIkeDPAnzhnT9A0Jmi1kxCRCyJ2IDH7b5ar781xUHgh6r/ZMUfX6lQ6
pQuCWUf8eoUmzgTikuB2ydvq/DNiO/SGgZUcdogp2ifpp42ac8o+iDlF+2Gk2bZ8
VU68Km5JCSmU4iD+vBzb8LDLM2YgV1ZhH0Qkf9bIgOBAw0qVLbkw0Ls8d5bMHj76
697QluLNQjFx5dJ0f/173pe8axw84TMefc7fShN5weI4XM9LNcMbvIXulxaaZqKs
4ribHtQrVoHmcjsVsN6iIffh3rsk/pAat3n2obH9tG5HS3GWh6nMp+DOA0Zw5Mn2
VUb3YreLuzjBuWnPOd5UeVFw3WN31Ho+cO+v+/6mrdaGYs6E2Tr4bBZ5U+/UeIt0
fAYipIXIw3DX96GWjtxcfRHAymxgm6ZhI6R7zRHYMZLrn/BIf/Ocvg2bSk+v3Ezf
G19UdhG0dCQ5XuztCd7ZwVDRbk6r5LWY4pU54By99EdsIIY8WqmyMA25R9xwEjfe
Te3BavFO82AY9M4BVF/6+aAZzKKF/deDY8UlLuOI50r0OhUoaPa/EOyBwZvj9wWB
qe5rsIispHWpxjRIzN9uwU/hjknGGgoh5r7kdkHgtUJFPXcWREVu/J9sOv0lXk/t
gF07RMVt5zZXM5qhNJyIp7/zSFNMi7Ps6fY/7sYTurZk080OUFRfwanLjUj3JzzQ
S7//sB7VnvpFqIdMsKZMurR2WkUHeOfZadkEQ4VPnZGHvU3o1XUOpRcokcdXLAlp
wH/71N9uy6D4hnotL7ohP2+vwV3oboOk/wC0BQfL8GumrXycLrtQ1dBIdr713NI6
++uKP4kBkCRhsZr35nT2Fi13je3YTnCnzsqRI64ySvRwvoUSr4XO5Hu+t2cmOCqh
XOaCi9BaKKlDWNYVBb1MG5WsPPKnCuZObvEsqAdLW/0K63vy44ukojSnzDgqpHSF
UkAebOsBpXTl/nEawc2UbRjZFh7IOQ8ZbttMlrmBeeE8tu4CRPoHS5/2tSp5SGdE
z0ei6Ej74nzucOkrasNK4dIm0ngAnCcF05kW4m0ESSaDtGHQMXeXJVr+3z5XToik
JLdoPh6+yf8gcAKowtPWNLtnGJCnqKYOOJvqfAnLjgYnX+0vDZij/HDz4XA/l/2k
LwHAexBt4zo2XYHxgtzHEM5kXT8lmLNj8mOBplJNUWyqo0zN5OddMgnLMfOgKBw6
YnA+FK7X4rHgRHQLa07ta+j2JfsiUABdBd26Ijus+GTw0UHobqhoRcuibJi9NsB7
GMKdXQSRSTcr8U1H6ZBr3+U1C05a0PNyWmWiKdqBPB9U65FbEFrq1Po5MO2HtkIX
RkqUj6o/02mGyQn549U+5uLLwP+iUIT9cEAU1Cyr6sTg5c7/PJJeHVL/kuSa4Elv
WSLJ8J0Na6tRg8XlIDpi4WWxAZjyrvaJk+ssrR3ZspcdfcxA6NIBPLNsyyLG3b+4
w+r/kOgDmJIq/0bneCYr5jOfA5GV1fh3yzXbkSNxbeBrWd/JHCfpbVQBNzhPHdLU
oKPKpY6BSNX33+tXm9TLqHZLfwOQRXP49JCinlrFgtqKcrH/HZhE72a1ixt14t26
fLBWKMSzAl+EM62JuDa5IcRYj56PU8ncuimSYb9zP8ex0C/Pv+nf/hsEgBNTQaQx
z7m6tUcoO36c8n+nhp2u1nFlN7tj984inFvO/YWxRspD3Ly3jjJt0IRDcIlYnc2u
IkCDpdU7+jy37cG1j/qOSGGju9hED2gBMJDOE+Scsn8lZPCT9+Jab5CdSzMFfQgI
77WVGMLx8KMTmalQPzpYO0Zgkob/Nha4jr2nDrV5SLcpVRYAX1QxADAhXApkSiKt
l5KZv3MceFdhmg0PZsYSiv5egHdaoMtnUEwnW4Qs4RPSTX8ZiqVxjxdw1rrmCwlT
eC6LqaenKWSl73abehNCSkaWHrK0JT/DCQs/V4xfAZ5jtQOMUFli5uHAvRJB39Dq
ypAyIawrzx67zETj4HiBGMBHjIrqhes2+sYHUHv+i9Hys0qzffpn2XZJgb41qmcb
T4tzZkErpyuDf7wcY8hIl+b3t04gL5zslNfBPyBYptdVssd5IwvWibuayGnawWBu
bGt4HTRnERqs/2ETd2wGNP6jSW4+xnJKkh6xn0k+hYf6zxpVINgjjVwBnp4/lmTz
m5t9nJDhH/8wZoS0NYO0g8VW5vDElCUmnP1pBtLXZ6dnnZkT8KJq1fQS5Nnc36sI
ZqY9VdiQS/aNyzgGHiu1QLD5/hSVUooBR7UVVvPD9UOVIPnRoBr2u3mfys+1ZZ8u
kltqNJgpWccI+6ZPD9o5VoCZqzmAf1Cq5HOlRpjRIjH1/ckScIwr3rSm2aPy2INm
s6uxLeCm6NwOvqgzmiGcan53yp1d2l/qdTuvSVKBdBLG/qFO0j0l/9ZtErcNZDiS
hiod+/guVTfKZ5YR0E10qrD0i28utavZTnJHI+5yoRSLeAHL/7k2UQMDX8mPeQMG
UYiJp0rgAq1B1lNMFeUbhoNbUQIZY6ZWMHgfNre7ftueq3jU1611LC2gYRmre9oA
dTRLPpFIKZmthZJRBfD29jm8JDjTbOvk3PzCqs/77+NehXau0ZyyngCFBT5Hf6Un
q0DDN2AFYljr5M0hgiKqtbWNyJtD5Xiult0nst9dnvVqNRrRDcfO/DjBP3aH/ePC
s0tqhLKi8f4B88vf+CQspFxCxHxl2FLy4zcncFaR5hY=
`protect END_PROTECTED