-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
FOIJnAcmVH14kip5FivkTme/qle+OFqBU2PZqsyB2AAKTGWQfay0R1X4Uv+tLKUr
WuOKGWvFjpdTn7V+21exrgjQyShJA+yWPgpjwVFrynV+I2I1Uo9oNYu956yVqg2q
nIxBXuxp7KLk45p9xoixo3X+YeUTxZGVlhrv123sq9I=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 18291)

`protect DATA_BLOCK
Z5fq+Dtf1b+h/JZjkABke4z2UzFeZNxR4Y9rA9ucy9rjdZY6rlSERKew6oGsX/iv
R8MbIbNbk+8Dzs+5MdLbFYE/QbnoQXFHaVWpsmMK2kPWKgF4r2ettxRM73AtASST
4n1eYyfku4tHpCSmYFFc6EZvfBcMxwdupqHTJfQQGQqUOgnFQjpOvFl/MD+7dgLi
4vUwma0TiFvgeVMLrH3FsveaAi1MnAX4T+v+JuFjOTyoV7A2FVuim1tJyYsHQWSV
qAuu5vF5c1yt1WOLzEpvAW3NSJD5aUeO/sECyuiu4CYcblJIbvmONV0R8Jyi3dnT
xsdVgbQtPaneNcO9Onh3dpdQGnv8/NxeaCGLMGwgvvYwfpgQZNJK38J92+wDXuSt
+6vp4cgONWRbc/OpYIu5BZSwfJ1Ucx45i4vmGMiQdWj+g8+C6D3RiCsQzeElipzo
PoAnLj0zTX4cQGPAlYZR3yetauAG5eH6DtvoxPU4OUELtTdtVKl1RGWM7XnjdnJO
jkse3W+ae5R/07ae54k6EHTJ7XY4gSl458DAMdcLrXn3GExqahAKnNIEPNcQoR6p
4obsE+fxUITURvCpuyOIsXkHqmYoeoTB/XvMvrRWdf/RKfoUwJGVqw5B6NcwRiGQ
BoVotUDXa9B7DyVSAFLnTRSA4VYT2dKWmhw23zrkcIy7yAfhbO1XoCSIqD6ikXE+
3vzkctJ1pR9uc+hT4tvCSdh8JQuNA02yWhuX8Ph6ElEyuxj5o+CJag5tuLz52UAQ
hlX9ip/vg0iC+o1Xd58nkTkUPUgX0kywgRpOpQHdsPDRL2LIXTEwVUqOWc8zdUJy
lGmPsRpZWReuIpff+cjGEZZAnqRIUAC154iAFsfEOoTrIHk8hocLjhXc9x41idGo
ElWL2wgh8wfVppnKWwuU9LcJOJhLs5nzHCRqbUsZwMBG/1Jc8ia9ULWCymJck2mJ
zQMhvUaRxrVvDHiGp7iLYPvRqe+ADRPNd1aNhQUxVwdH/LXtji67vRFOd+SSqlyk
TnzxXah2DQUFYJnTpq7Z3/CHF3P2kDSt3fIiKuEv5T5cvzZlvc3pdjhw3jy45VbQ
LiKD9uzbnFlcO325WVDo43O9krrvLH/xdHMJqs6qe9HbANgeUUDpwHzItXnmbnRO
PZDrnknhietvIAhHBhbVQPcme9DZK+2CIAc/tS6a62JYnrKDXEb62CFtgGbnKUVK
2blYmgO4vQ023nx9mQTWzY9yVI4h1nDLfEiOPHU1ovVH3TSuBmGsfRPUp+osW3x6
0P7rID5CaVgpkpSf24Aoum+KqEmZtSJtuLbosHXitzx8vMKKefRDHmPzhQQTJ1Ab
mCmFm9tu9xDj/Ye3vI3cQMGsglO50r5ev36FpWFrjqPNg/K01na6CR6ZqDFYYfaF
lL7fG4Kz8SdIjcErUYwG0ea5VbLL1BLo8JOVkGEQ+fAqx1WKrz6p05kc3KL+iw+Q
AXsLsVy+iBdkILKQOkI8Dp+OVMluAqX1DhUTDFfSVKVXJjDUqgunbzwO9HxoV8Qg
opyROgQ5WoS9sfcr3aYmJNXsAVkVrTdW6cOIT+7RyBMN0Wg4DG+1L+LZVKUprIa7
Aigd9WSFTYnmpoR8/wqNsaY5aZFwbgGk9ybggsX8/7imLOTd5n77QaZ0ReATREXP
JbojudwgLRBUxUFQmL5Bj4KjopkauScS8k4WxBH/APTv60DuT/SGeIQjkfWps2mj
ZT6bENgcPep7aqRElcIDYujXFj0ei+FtSX4s6LO0OL6+VUxfv8wwBVVWv4DOZrRi
BSQ3WhoSVayZAqtMU1P8Q5zm+ediWkReGUjOroj/l6kLRhq/N1jEnoWv6PI5nm0Q
b2eiZ1sLNHmgxXRgIbDq6C1bQqFFH79tjnzBoHD/UF34UTaCNAn0zcy0UnTPkIAW
nnTuW5hFu5c2D+Yp3xfDLXJ8+bbWcJhMgLtFPHF+uvQhWmku7SSoST1unyOBlSAN
Wb96LQBuQaNzdH8LuNAAtvpYQSJQCBlqX0xrLiBnKqaW6fzJzgppKixyt/Rv4J5m
i8ANRNrijdem4yxmHOwYT7k/sW7l5h5JT7HaKcMouUeOrLa57e6TIefvqraSPxB4
sx5+FHaFuibP+mECBkFUCeGAACL8kOgTtJop02S8AxsvYbRHTxdbiOvbIufnkRfD
cdDAsWkf5nXygbVyNd1mqgG1B2dyidMEKkkEJixMsuvg1Q3MH9ZBARdWMwbClZBd
L6RUbtWjt3Id8b8QXElie48No2+qWBLmIULQfUrzMQh4Wf1/8a6z+Ezh83yBbf+8
7vHsB5q9MAZRCQTXv0jLewiNAhw8tlGzdvmuYWtmmW7+Ecva2m4n9BeKOSnz82mz
IUxPe2MH/djMh4zvwPJlkpi3RKdcLMS+dN7FoVwk7J1C9BIormFTIacge0NIvRpR
nJFlFIaw32mBorKXlEqQSeseojNo1PRYIRXjGF1Ov/8OqyvT8enGoFP5GDlfhu/V
r+URpQju9N2rZ5aEyQAJgJeMZOIdXXyU89yW5irW3px1fSp/qWLL4E2e+KFDffTn
c7cRWSRmpuBKPQKWAqEFQl+K17dgJAX3p8EzL00S6LYfXLV7jg6L0B//G3eHVxJs
rH3k9+zbvFbyzEFg3KsdI5QwhEuYA6hOTcxz52nXYJ7Yjt1D4ItIJNstZDP8ppJg
56wYpED6V+3k2x6gCi0HU8VKgsGyj0WjQ8IIKHwgy/69/x6x0GSFA9FEn0AQVuBV
FLkgi20im+eqv1zennx5rwQAvGCDHQCzKev5c5ojPgNRRJeA0z4A5tYfDurAskZ7
V8cjadktLrTXxY7FoxHKHKa6Fv11rnOYyYW/MAD8fs0vpN7QGkqcEd6fIi2nAQz9
lw3G/9L2PkVkAskjOUseQYa3JvS6G57TP4JjHFHq7gIxBBCVEM2s1YzChg7j0RX7
dEvZcLMGF050uC0v8nQIZA9rgrZ3CtitdhwzbBvZUHgtUekigO7hvv5RqTcd4oU6
BOckXFCajg9rnc1arDTajTWEz02MXzOI6pcgUJlCz2jRwlXQTLNzqfNdOe0wxyQR
/b9RNePjNmMdcYlgmLY/2WrFX73UG3o3A2v6NttZc4XpFJ25JCAIFJEDHro4EXuM
Vmg6r1knsc4lbwVFhcYH3JTDRBCfN/3RbclIEX2dg6mYAzRaSJg4yAWa+LDi5ULs
e76BRjl2v5KuimSNEDpSwd47xSsCbDK1wrjONGOul3q083ej10ha14YWhNVcnX9s
5cJ6SYGNgOBDNzyGgutmXi5MszL86Fa+hgomZodhR1xmEtSl7qptpaMpC+Zba3ln
Uo8QpMofNEfiv7P6Tuj0epqU1HiD9iVHlF3Ut7diwdsSR5h72rYyGCQ12x3TgEZv
gtmnQ7w1w7h1vayBjWfjZ00UzKYsYKq5k14jUg1Rnb34Jmv1IGy6lppodc+HhF+w
vAS3EGc56ey9VhLT6aojphmF5FMfz97IxvnQJCFTC0mLvKsp6RQAg4mkaEmSQj6b
wvWjsyBCR6vwq/W+906JrDRM3wOeNR9t3NEUAWNilJtSCI9i8UrCt1+2Y4yZWLuv
tPuB3EOYJZjtWdMPLocAXxbuuu6vYkAdwqSj8AvLjAe/atn/oOdnWj16kEVi2eyU
9vNHhbtsiI9BtidyF6xKBOENbQm686EPyDoNbzrQwxJLJwhb9Cew9yPzc+oYp1a0
Oky7V15Ur7MDVSjCFMEWjthrnc2DXHspAJGGmUr8mxKBN/7qe70QYr+osnyLUk+v
YwkaPlpogQkLE1Onab0ohIoMHY9Ts0Mc83CLeEGMh8peBm5pqHpmSM70FBAAHFIT
rQ6SjGBDVvTYDF9MGHoCjNRmHoUs1hca555aMRnM7vCb6NuNlYG5DNodZj3C0/Rr
AwaNxP88YGANpK00Do6NpGYBi/DK5SE/KYyqgtzF7jR8arcgD3eCPgsPLBCO3MOF
dheYnDqyk1rAkfRrFAfPKxVMLwS3fBSmG6S/nr5poZyfVRcsU0Cbi5EtGBIQErxI
BZczs5o9j3iorPfReD1nUNMHP053V/etyJuREfYG8LoIGp9Mgu5nL/W+xFjVuSmC
pZzBti/i1KIbpVLBD2fDf5kPFMH5cHIGn1i2SMs6b2mBExYjdbnhhrWQL04Ba8/W
zX7o9gbkybdjBSO3Rid0EOP7IkodLRmCIhxQoDShiA4vhyV23sSrv3FUK8zyEjAK
wlhIuhRpQEsDV5Sfcb/Sd8CY5koEwp4TzT3TU6roh/9tcqOCb4C+MuIICt6ntjSl
f3UWh/VxVIv24A3nTjjrp8uhST+hb9IxCCwdDaYJ/GckoxSN79LKLxh1tErYGz7r
rtXy3318fakR6lgCYuzf6bR9F2xzSjuBstdu3QPwGZ2PcNT9yEPCnBUWfDKTpN7N
iIbWZgw4Mk/esMQKLOfLe0xvno37DfPt579tkOvkgXXWaX9g5K57W+ChlWdoR5EX
UjndiZ7TgItFUewnrNNl3YOq+84jEw+2ZZibc/VCwy1Puf+SvljE4cGd6KV4U10d
MBxMzDTtY8ONpSPzasL8H9UBRnAA/PLAQlzRH3XAEsUQF3uBZpaZLIZ/Eq7k9RCf
JSimo7BQ3RKpLG1EgIYb+I0xT5EdJ28ErINGuO53NiMC70WOfclkDOvabjyGJzL8
qRjQpj0836V8fvme0LzoWszAlQJwPNZwVQErguW4RXWjadwkBfC4ijC06UCHMNNl
GsPyGPEsjnfM2Pf5fCBlZkOJlTnf9+++BtcOM3K6KrQHZLfCMeeBIwFDkrdn/aSE
Q/zVO6qlpPzxF/5h64i1KFYwQdgZTEvwo7wMa0zhuErKobyfBdPqoPnMFxdI1eCU
06BAnDm2Y4iiDWkkwhYX2HDu9YEuRqA6K1QyVC205Rr5X4Q8PXOsffBrOFtPxKNC
UAjV2hbDat91h9eID/wcJjnlmtq/MpKz0yOAW2T3LjFLHzZr6hCeO19MWp4kFLap
f/npAAIIv2HFI5WAZ1uHdmToLuvOySCCKujnkoYiKiyGI25goxgepz4ivk94iXRN
qayZ9BuuswMUDQ5K4vayuJSYxc/HHfjGYqR9MQsAl8JX8sO8lc2oFWAscuZteLcD
sER7bb7J593UC5mwAOw6OuXY51dBCosYm5IIoagsYzuq4KVP1f5LeBmP1Z5EDFIj
3WHuEvobMYXb43LPSRVnNngpB7SpmvMO1dxRNILejs0ULSWWxXd3JWt4AXZBglsX
tayFd3lfCimB06a/VjgbnSZcGV+7o0dOSM5dcKenqqJ5nujfJyIWBnGZQFbm5Om+
El0VrGFXw2+2dV9NfYXnchCatUdb29YZ6mI5GJM1EUgpjw7eYJdaQHsFXEMi2S40
8pNZPV10Zes3V2+q+1glEstLCd03RiAo1DAzL6NmusFeabOKflQv9dvRkbs91/a8
d6w8RfwmHntmt+10VNrk2LR2mAYjxspSkIE4xLNVmRaTRi/cQSeAkaAL5ZcfSi19
wIbrWAmvI/VlKUYyh3LpWP5eoDQzu2sMmIXXbTxt7Qm7jyQM22r815ikL2wqnVUW
eVskUd3ZUMFC3OX20HHEC6U5hGh3PTYiWTNBMfihGA8a4hxhsKd/qttQwFbsn/m8
oj1swKwxL9UAZbUXkREsIRKEwXD32DuUi1kydbLR+Vr+YJeLF6mz8TWiLOtJrDtH
o1TodvEXbFX8mRUILU16O0exVNSiuMgSGpUDgeLjz5BFoR9LScyz74jBsDqBrkfx
US3sjjSo6M4A1TDXGgrE9BW7fD40EFSKfVKayWGHOJz+mpTe9nWf81hfZd2vBvjQ
cvHmXao7jxSa0tEOQ+5CMZdyDWBfqBNHB6/bsDX45OnoFQsR6LfroivbiA9UBx/g
48zqO8zJwKSL8uxt8OMZo6UK/H0ku7Me0bH2xHjrdpUsmy4SNISt6Z611vH0bAsY
qG9AdXqF5RA8xWCm7oaE8ivi/47w1NwORnz18O2htCgF5FMtacWhONR9jvrSNK31
r4/6Rn3FSp1LkwVbdpeI/MRIpviNqsWOEoYAQzYAH3Y0NeyZJeXR1swHZKNGJ6cZ
uFJsOiQSwC/7WVElSziBzpF1v32GngIQVqJu+jy3y+A6JBP04Tp2vl4Z972AlRFo
fexXyl5zF4turzgubZR7EsxOulTlOkJE52NR5lOd8Mal76KLrzSg7InZc/IXE1rw
jEMVMwmAl9IxSCEDu3WSlB+G6dZfLFfGaqKvIuBUFhgNk5SlB9YejJYvvJNqT8V/
66Iu5CZmNY61dQdeqQr7Ethp6TyE1NguTWhs49ZpKQ8r9S+nd/O2Gy+6CPz5vHir
NZXo6fo0eOGocbO6wCqru7se53NKBQosl0B488nPPmrvpEheRj+emoSA6xF0RX5l
ypYcNy7tiKpcGxJVtS6HWTGZV3DfrVvb7YzzhunNa02/jCI3Op1GND/KfZUSf0fC
/J+LZyJZKCM3rVYkNdpbpIDt/xfZwRR6MvlAe3UyzpWNurgDsH1sDypUr6SNo2Hk
bOheu47xKM24xsbOSk65OiVjoObKBUu2+2Q0f1hQNRvU6SEuYIIH7zDnVX66/LXN
IwHgHYZ6WcX0AXVzE/BwFLU1Kmwc1leZEOk7C/DwljBcYphG2mPk/eMfW1Je5iRy
5wqBQXTRJ+0oKDB8p/B8FN76B0QpCHWU0toCtUqUNI8arf+MPmz6KHz4MmLgLCa1
OSbjFoxiHCmYHZaMByH4yv/1otndt9HISzOEyqxdCRBSS5IkUi+JVSvnN90Ke1B4
A5ZJU9ESTUdbN8ie9jbruBqr0hpjefwnUJ9YA2unngib2TkR4Zi69KigBHTIMZlm
t16Xw/+OyEMwEJhAzq1TERCvE93JxfbX41mojkkuLC9OtXynZ9969huaaidfnqrH
AbeY6Pq1qxMSqrKeCkdn5K9ixc9v+0uSzB5Pc+CGfM47/3Vxwfn1mqRSfSckrRLD
64iSYyPqqBfLsaH0drdf7/IsH48gvXp7TZvJi4gznMqx/w3yBwTXzY+m38cHGBDz
hDTYybSCCZK4dSSKBdDTOw+8KbFPUBi4eyuN8ir3GdgYh956oNP5HJFTpQF9Uq5G
+cVKWw6iuqdMyl/KGS3kvo1rnFV5Fnl3GmHLC1lRr+v2R5I8WtHI9E1utya8KEM2
gyedkHUpSjwKvgdBJ5YLi3yYiAA0xP9iUmMoE2NRgTlonm5Sr51kDag/4CKczMK/
lGEr4moaZZFJ0HSj+MndwOFjHwNHNailQnYD6FXcpxW/17ut8d2WWXHAkuaS2jlJ
+mu3TjxYUHzNpKuRipNNpzHrxbQIBjIkyE4StbTsZtb5inVqn1MO12wkP0J09DRh
yMps8vnK+HOkXw5SxNAinRBV3YEHGHAwdArjgH8RRb5/S7VmuMKVXQ2/ynmrCW2H
Hrc5G2hYPwvwQwSmkyhUbhF4G5h6UD3JWzuiBuQZj+88tXpL5bf/XmUCMtmHeR6P
8F+MAH9Ic5S6kpsGu0kbaE1a20WUv6eDgakLD77IYcob8ILB2UjgAx5jv9wQIbT0
BwhyHmIzz1XbNm8KqofXic1aCnW7sCLAJ1E/DXht94hvbGTv6SZCqH3kGlKC4YS5
ndgaQE3wOQdCE6w8AJn1+ZvEIuiKb6Etc0TUQyIBFYC4XiwPeAE8MxF3QF4pTcnk
cZ1VNMr/FiJUMwibeQPumjBrf+3Y1ku3wvHNS030PFTFkjtMRgy+ox4GyC0M5pPM
P0ZU7rdPFXbCmVkOxPUsS1ENdNO143IudVZc4i1F/G6pXneSJH/ag2o7Kmo/ObDK
49whPI6QPYA9i9qMIAMcSvqrvoXWg0yv/biMIWu1Dcob34mjy9IHaRKcIssdZD17
nvvambACRm4CKlodCSMsxMjQG+qG6MXLKAAxYd1LunW/aD14v6mD8JOaav/rTZ+I
Q850f8T15/3VnBCVG5i3OhAiFxRllQcbv6HtdRT69r4/cG9rf78HK48lOtpJwA1i
okKsVxsGYZbcfH5UwnFk41V0+K9cVmzFCuJZRQ1KByNuZK/S9sNxYBghZ41YUTDE
KwGPAmwKTHFyeWpzrKPFkPELSXBeKZdrKvAJeFxH7YZ5QbCPGD9c/yr/QWFgyB7C
e6rtnk6RR0qQqbvPWwQoHrvolsv0KJLrpuVou94JIjx3zdwsWnxqKiIlw7sFHee8
M7ZTyWlgdz7AjKYiknrZK7qdZ/N9dYrOZkrO4FpjIGaaO88n4++uzhP1mSco+vo/
kJCfmwg0GXhmB45WlgDpQ3J8rRZZ31O4/6wMBniUqljcySbvWcXb3VR6MVySYij/
Jp7PD4PlVH0OEnXyhrNB6ocKyXfYS1rwFQcdgrIYIq71KvWVBwFlNqXeA/h8Xj9i
TBAf8kb7dO6GTiScyoRDFdjI6yiL8RMnj2f9SfaeDUaUqXL8TLSj8KsF6hHUqcIX
NA3dU7gUf5fmtqaYERiur1v4efG+SrdQd3/Cx1MKM+ojOK3emi+mhZt2kjEAmZHO
AA+z1bKpMqXYx/L2vjJ9EwIZ+0XMp/Hz2fDEl4PqwF40pci2zPYmtckU08kqZHFH
/nbq7opFJ3GLICohRHyNH8pBS1fEHHVv6TGZn5xsqOHTeGaTDN/t8h3kBOkeAWI+
u+gP5v+94XAi/jgCQXXuWbU8XujPrJybdBDJWck4qJlvUGrwTFNiFF9ZaXyZMRI0
UfOOI+dU6Bwu4HGxn5uBWSoXPny5ihfSQVD8uhK6LVf0oIEwvWp/25HPTmcbqi9G
e47MvLLSR+Q7UP6YIduyGnY9MthxBJsFoUyF7Jg2A2pqvCW7qie8/0aiaRSZP7jK
ylKv6seIfYcGlSGoVpZCERuBoHh7mGnRPdUp5qvHjMkcpPnhUmxpmLydz2P8CRiJ
FmpqYo94yVf/OuWJcABxb/uQJ88RrQeYxsM1yC9ZLtpK8QmKWgTB6tHpzZbw8vUm
cGFX2pNsUcBk5aeVdckYT0lg4dp2aXn6mlUgm22M4jKKF2kvUN62OOTXwdDbpO85
BVz/3CjxkgxXDlNPK5tA5I/Bx/CRMs9PPcq1FJwWMHkqu4Xz+E0H4KH8IsJy+vJo
fEW8ak/o7tZlD0OUFj+sgICUbmVRsB6w37RoaBMZxitMGqBY/bCGf2lmRFIDv+t+
MR5npnR5UqX4YS5JBy9BRi2FhXULCkFK38qeGcsmJjtEWWmta+sVTY+UQWjbXOED
FANS7j9XHAt7OhRenFInKEVPbavCV6DBvGTUEBqpb7UuVdNVqn5G5lgvAr6ZipO5
KQobgLOhtHraqdj3Vy0X7oE9KNl10zZalpWzNTRyG1r+Ih0qFgV26B5ok+AmewQ9
L5CBNVEEEY7yskPuSj6TO2jyW7fRXBPzY2/3JJRzB4v5qQzLVkLCcqVL3TXYLGGm
gbfg5iLTsKnG++W5Ht7TUozo0KbrxE3SfzctIK8oIvzwCrS48/6E1lUhFp8Pp05d
qRf0HC9+xCg8Gx5ON3PNn1hwHoAvHafI1vVqeyORZeFKg/Qu2fiq4D5Nm3ydc9dU
XOZGWOdrZo9Zs7BBVhj17RAWzuz1UaXN6x03FJ/R/QB3qOFt/EMbQGBkSA6t/kO8
BWrKRFIbdhOmKg6kOe4zlC4ztY5hQkT8D+a9aQwTlypwMQe5kYUwhN51vqqB0jVm
UmVTqXzDG9XBTxLLbYTvU0UiR4Da4j0Z2nK4m2wxmtQzttli8C7ilK/DrZWPd/nT
Osaduo7PApdGZaicfnIwTa6jbHlbJnCESzZtLu3vlpC4J0Nlb0esA4tkrng0lzLl
Dwy6wKaueymuEYxYMDPMzxKZdwYprg3zPsLVGeHgxgLV4RBnKPDO2iSgDoZ7adLU
mNi7iGPqTNtP00ozDPVNfOI8wayUpdGGwXX3OoXaruk9WutO2nA63pRzqeeBaIfZ
NGv0iJ9cE0fePSCLsfjCy9q0EUhvbcmlyFcnDP/SlqPu4RCwLwMc+q0yLLBzRBI7
wH2IlKvaMRqEWSV/KUFwxUeYnfbjt+TS3dkRtL8A4Z6IO+t7wMMzu7Oz2zHPVL0N
ZNhkuCI/Qffrqme5xjdBsQfmLV16ryefKcz6UDiycPPfWLikWb3R7UpexlJL4qur
+UdxHM9oRY9rw/a5KXQSFXgYiwStF6Y2Men4zxSNSzUMGmYuOH1nwYeU0/JldKyx
TiI69X+/vDyHfvda0icUoGm+OuDi8JS5rg8qcU71RgViiLNBbhzVkPMtMo8q10iq
UaUIqrXhvxNC/Cb07RE4GdQ/8OOJMK8ribmueKCs3R0rEzF3q8HW3KAfQ6HwpT9p
KGGsN4Y848QmxyFtgP3c0sgQp2eM3lh/mbvAAgZzFgqnZBLf5be3z+zFEJBHsnCB
qRFS+UYLJbJTW9BmffddjwswsOZ5zUyeycGV3zbxQODevtgeX7DhUF2jdz5/dRdj
ZGpGuWy1afUsQdGlqNTmZoIJwf7LkQwq7LLQxYUCaYQ4L7mH08hs4SC84MO8fd+o
f18lKWPfBKexmuqXAR0nhCBXm3dWVkW38aOvxef5BC5ZYs1+TXOMLvCr3va5W6OY
1X+DPDCtds/P3l6BVnsec8dLzbYD40g0cIsSi7vnUdwtoEJIzUgHxJfoIbggPPPu
+g+mmKhQ1wchryXhtuml6EDM9Adh+S1CVcRUPHmGJXmBk8jATRMI4ohAd43tCpXy
0VUigf06LRZ/fAkwWYi0wY/jscQdtY1wzVMO91HTho71louPQcGSEXnm9cgXBHsd
KSytN99+ifJ4ue84jwTiiAK5K1N30kluL01wOOVNVLQg9+x5aWQ/dUNq/npEV7lq
CnS3v+NN9SLUPQEj0VTdNVs9kXDUuyBTHPJ2pJNWSKHGYdNWRNXK2Pi1jzD8251e
6PbyMdv6YZtulzYYMtap23+9lu1z3qVzTGCkGQ7kR22shRroM32G9oyGKOuy06Qx
qhrzn5CU5HljdnwQwzTVhJGoQLaxyhokHQ6XQge0KnT4AHj8PsUU0q18/cv8+qlD
xHrw9PgU1ojLwT49QnCHkZX32aZX0jEzEoHjsra30eSwzUbKN2u77MsHraPRHjuI
s6aPfXMb0JMrkg71Iwv2Zkce5UFK28o8IKotGw4JTaoyHXrrBws+1FBKo/Um0I5B
66l3wS/eEl9WJJqzBiRWWvRQ4TI/HYs+AnadNt6kMnley/lF5R3SbHtEDKZ4pN7o
WjkaS8+GK+4Ix3CzCERJnquoqd6oENjTr/5lDDa+5trOO7EpIv67Y+h/4ff1/dTi
MZNHL4MeCqva2Qqp1qs7XQoPg1skf2keYDlf6/Ze5pvyq3xpuukeyREhM0OKbS8E
CmppJGN6t1Fy/n6GNx1cqw3zW/y3RfO93Tpr7LITZRkRU/+rqaYtcbh+AJDeW1Gm
3CZthqFqFFH7Rl8y3sWcbJCrS7ItvnGOkru+4kczgp50GQ0XgTKKlERYXBFhc/Me
+1Y8+AH9F0VIqzUpFhtHFRPHv8EiVhvQt56Xmy3T7t+ZSOfzEZigMUrD7doZJTCz
knbBOXzp1Hct7ItQlRDvlcKMcku5+0JpF9puTJGaXiV7npDq5HFInUl8BTAkLN2Z
6Diw4AksQrzDO/wtT9G/PwCpK1tY131Mi40Pt6VtyXFNhUtuUzfu6hzuc8SV3P5V
UnTCthdOckAcOddMhT/m+HcKFMhSGRP23MBuylHu+iSbofI+LSlA+rIYxD60DTjF
9QkLSXZKpzQhxW2ea3vgMj3poI1iF1U+F9WGSKPFoUPsHPAd5Js8ivKdVn1uVo2d
gRFr2vkU3iaYqZfcpcXbgov2zDcmBhKB6pWRYqOnKqhZugRWJf6mIoX31H05GhPs
AgRVY4uMnHZpAwdcamUDUqnDXRwX7UlnCyEFNahJ9NeM0nASkRSks6QWpeo5WzqF
mB8J+UJRHFhs574f4XPmSuYR1quF13K6rPrVuRu/T3nYD1SziEurEDiHaTJuWQ68
nTVwJlvHm6k3fcYKmnjM4MddWioz9w4GC01f2RnbgOSFznl0OGwGirupRbmutclG
oIjHElg3ONRHkgTU53YO4JL8sTq4u4uJ4NLJKN52/rPf1pcqZbAfd8Lyvw2prLYK
wAO2cgWK6B2x4PrEUcaFH+dC/mQDsTJ0M3O9obJ6DUTm2nIT6vCpWGluiAMpJ+mh
kxt4mP94qzQemfpMhzrxTGeAagOYi+4QgyjNHGelsKpMVBjMiMwp9y+e510Y+g8b
fnqt6+FB39A/aEtZ0YJoFExZUyBNEh+/LanmGF9v8G3nPTRmmD7FNqeS0d/TCkF+
tEB26ckU4Mqiw6SYQ4uEpIWsvij/ZwaUKCMmP5nIbrf7S7qi17ehr9ZFN1w0VzLL
EFbzcWdr146y4+yJ8YB/TdGV4wEJpMFkxZs0IOdgamZrWhvIzNkWqQ/R0d+9igvk
96mvVAa2QckvDyTduCKysDTCE1P/EhzcqYT4bxqtS37uLmOAgjaPHQChIpPcQXbG
v2lfdmG3v8ctU5bWZUct4kC2G1O8HV+Cq0iczt6cZU+yVbevfnOS/jcsJsv30g8F
okeTthx9UVwzdi3MHasfMtJdk+GaGZbvTcVyFUpAFsS4QtC0Oo7OwxLrbhgZ005q
Ht4rrxKFG55tPG3S4/GcXnEKNTL1n2lQMpX6kbK+90DmK4DpOhf+VDwBT3qHznc+
kvPKRtgXvvcobH6D3CtL3Zsxs1Tz9yVbaMUgizi0dq8se905KBpwIGrW+KItiTsT
gY1mMB3Vv3G51HSAETBlBC0UVewGRf5qa95vNCJ5EHKHYB28HtctshI7MBnJGsjP
kw3jcB3SLqjB7J1YRcieIVG0AJR4znVbK1uT4S1vHe0OSFZ3aMAbZ1aVDHXPOsa/
wQ42QZAQJ/2cUZnyTMp2gyq8T8cTCiPOoKsLUbfogQOqUJlgVinz7A0ZJzuM4adl
a/FdwXCIhda3AxugwVif1saljU0pXV6UcprUbpIB+u9eGojEmvuGxIwwLb60STV7
vVoW2BLVLDLeC/fn/jqyYrIIHzUqLKmVITBnXqP47hDh97L0axnmNvIB8hXv9GYO
SaCUpTS52NCVv+Gjnl7v3yqQvb+K5ba5oR/6TpLVPpfLHsWUZhOOpV89RsFGHROt
mtEvcUzTOs7ysqN04wuhTPKTAjs06pBpas6BqYeqJxBQ3JcPiT5A5htGShRbxE5f
rFlpnXiZvboINdsC+7x0pKPnx1AoV5wQ15RR9c0nsg2yQ2TkF+3/GUjcZ7bH/7T6
3HoGziQf0k7GpBTz9rDgXJkesbYAW7Dvni8M0Eom1eDr+/dNCzG/kY3+06RkA5Ty
FP7UHMfAUVqfOiFIdVvKUoQICe0G4HQDzYafBy7eMso0Dqchy9MHg/kyrEL5uXDo
FlWNHkfMjGe0s4XhMqywvRvUGkRihPkXqsGkKpWJ3G5r6AXUG4rSazLJrf2uXR8N
HLtW4VKmdU0iBX7nlS2wBsCLfKAQNvoEHrelgZwS4v81kMoYW0ybDkHzhY0dtlOq
+HKI4IzZYM6W7AX22OSf8Ps+epXe7WNAECIgkQNghReq/Wu0q7sHxuO+zk6TutHB
qh0C0So3TIDbst/6/61QpcHZCNoVXPynPej1ZyVowsQHtAh+0kYkv2ajX4XBrYQ6
S3ZNo5o4tHejAGIPg1I8Hzt9L1OuBfsvYJO1zJGfn1IPl96cLB10XOAMgxldB23w
UUXlJKavHrIkxteA23b4sIpSZIJKcouehZKIYw9POjMjbVvvDmcshYZny1dxpgPS
rZ2SKBWfZ7OyyqfwS2npe4fnyMdHAst+H/H7FRxGmAat9XuPXXxW94Fx/b9JNrgc
fEWt3n3QuvUtFYtLVpMZtpCTq4OTjn6aDsUCSpmZ74bU6CVWKgEZxdXUNQtAa0Ff
9GlXCkdwBTLmzMQS7i3BOVB4dHrIHCootB8KabtWeB+U3xAzssAHvyqKgafnRfc5
10T64N3c4RWkdg/zTVQhKMpghlUNuVJeEHMefoJL/QLatoXHDV6WrjSlGjMwGAST
BLwfx1FYwj9RqimnEuK6OAYl3JDD1ZVhAzvgeeq2W6tYvcRYzJMoCu+c0+/2eMo9
5BD2K2xpgzjDEvgAqjtqmrPkFtyyAl3MUVt2c1kJtc/Oc6PAHlc1nIwsYajxYn5t
CaFkwpuCgF/2EW77cfO+N/aLdGwXF/tr7DCSQcqn4FSFmhLa0xw14/LRIyy8evt4
SaMb/usDNfwtUHqGGY7Pll4zbOoKeEOG015wTRzsKFTdo4ZyV8+Q51KZEHxYyoUu
+SzSJzzHKWMS0cM/sAFLd9q8JVBhdQ26g7khD80KOAfmDmzSc5OwpReQjxSsIW8B
R9NIYimVVSzcVg5jFcBjA9JuInsrnf9x1aRmPO79OxNPjAsjvidx60oF9rxAycVW
po3VOkyqes7SiDqjmH9cbEk+qolCxi6I/L7P7Ge8JAZKXUR5yZ7AFDhWPqs2N2p3
+T83VQC3lm/Uam5Ec2g2dn7AYx0PSJlljOArl0sPg7C/do/C8FKZoKCb4hKTHcPN
OWpAI1PAxdJ2XEUtuSbZDfTIVXkxWMSPzYAsD8ovBt1b05vv3wCiJTyo8yJUDhdG
e1/U7y/2oJ8qz71tthuvSsYkKE5Hzn2xcVOKsZz9gtsJpTW1G2W6295UULWIEohU
tXtaFEitE1v6y7qYg2zB1l6wbm1XCtqFzAKvjuo6z/UezqQMnuiqY7iF5+Lnkldg
1tVV3rE6nymW4QsBO075ecVAQG4wPMbdbeCoa9Fnn/XSTwlhkmVKZP6cYMztli8p
baoNvGJbBjQHYoO3szrUiG6y8/l3H48jrQ6UCWp//V8lARDe5TOqNqWw0k0fSvFA
loUD8E5vkanMSi4OtY23lDLmWrRYZtklSorMG6QnwU7DSBFfnVQgfABYjFIyxoT/
WrHD8glae9a/VhFIwchy+XJmm82dIwTa286miC8zRhz8yRV6+lzPrKjm+bc0iMPo
mgxN1K7/oNqk0CbmT8/QdEnwk7gb5sYV81nNSAb+ZJHA2zQ9SoqeAT7+esUG41lN
H3gLYXqLBaToZ7628u6+3Yewss95J/zBX1JwBZVlKxkxvKq5xbV4d6tt2yFuSf4E
zxPY+9mZl4GSoj7vz/ZTgm+0E48l+pvMz5xSwTA2+/dZs4y0oL+Zbh/ftZuhdhMM
6vlYeLtQN+3hkyjr0Z3CvPaMM9YtY7O2rlIv5DXe6QaIdiQ6t3VQ5EHfB5e2sS2b
ENMPXKPVVmLSUNgQR/Ax0EIZ6SVOJCEv9cfYt982yL9WfeT9jxJaKepzaAwfcQN/
qTGf2Ho3u+oooFe8Lmc1ErfYDGNmQifhanQngybhpxwuIOoqUaHI85uu9AoJcs8b
gXRMjRxXT/h8JrjlU/d03iO7YiEMSrzaiFMTf+ilfbJEnV0h+IwLsV+wt92D6ncj
5+1rA+oH7+ItarGqXu8FTbAtmY8sdles5REvSVwE8q3w87q5gK/SR3LTv7DGzCKz
8Twpv2R2fRy9pu/VhuP/DO3sTHcV7lZqZP79G23vME3WIfIyjF8jAtcI/YNGtuj5
RpyYYQ5rJ8rNU3Z7UYYDbzXiAR0ENZiVU2Jo/RbIsTNgMXCSFFACwEHrx3peanFy
iQImA7u7tLhVNY1uHz48mRr4fDcoYNmH9YaFbCMRA6BsBVyqwYrryfloxsuOBDoN
U7RRwgdq1sxp0TPCQXOYF+bdlAnr6SSb8X6RIU5vLoRWtM9N5wyxo1/E+q7L354M
jDnNa5mIx8IPo7v+qwzfUqYZGo7Hd9EDee1GF/wOY0LwFhMV6A4sEYYYUBRwtKBk
80DRCAfePlcuWxWOT7+GSQdFRsaqH5ju6dIMXezPyaqMcm5AJASjklTlrxCrmhWC
Qx8ddhnHm8Bn9Ggyf3qwOyvPk8Aq8j+qsCsG7NjnxzxGhUc6rTOK0PqDdW/r5W6O
rxtUZZGvjl+GI48FklgLExmYQM6TpWZnX32s4zHkAP+Atge/Zpgr1NcIxZRB8Lq5
xwpPGIKgk4OBR4Bubw25dVfDKDlQQhGH5biaBQPsgzp89v2VTre3IzRbKGhuYvbI
IeNHMpmN6oSIQJkHlGQVoVYcRMe+nUNTA0LT++zZHzTlJFDBVTjahSYtMmh/8Ifm
H6N2D+7cqYaDo8X78wTRZ83wUTUQ4dwIc5K5RQVBwsk5/ZaJzUbml6b8htjPdW7G
aMywQ1e+1SACdhBJL8Y1EuMa4NtZsX7lPZA0HKGujZGpQmKZCIMv3I1C+MsnLVTb
OTShHh/FDyRab4HCcXFyt4l7Y0DTa2qjcqmNZQnm2ONtQ+m9bNguvAj+ztWFCJwp
mMxY6n3KmLbd03C0/ydK1+hqVGEYOGcJ0o+UD9loOi8DxSES3JKkOvfGX244Vqdn
CfKhZUsZurO2ztTtMX+0IT0p1xZ52CCia8M//8KVtSYzUGB9UEoaQUjyGUHy+iAc
BYuAGoRAVNWfGApjQdTy1lh2xItPnIAX3iSl/PuBha8jkbHFw8KJXS+jam9L6H1h
Fu0s0caCPXMO8HmFxFqs/TpMreMxOFSaaDn9uTvTVL8KD+ckQQIvF4SPLr8lDCnM
vGOYYqZU9Uzl+OzjjGZXIZ1dEzydF1NlVNdHumyA1y0e0T0pXV6Nel5/rn/VzjhZ
XrTeoLXCF63TXZ4L4TQXbtpT8qpFBdwZWE0Kq5PhHjlfMoEzIsnBu6lTMWAGDIvb
ewciKQte0PDCBRwJ4mPiUuU6Rqxry3lHAzPti+2BZvSw4YKx5J/f6hvI1dDEq1jb
vJ4N5BaLdHEaeTTacaxoXjYXuh4Ae0DxAAGf9eWYpe1Z/iyMDYvJeL/wuC1hY/Gp
4R+/ofCdP/NyXRfCZR40g75FDvh0u1q0gZaooXGKaDYoI8tB9BTawCfXlMRQxAJP
noiV6+limXtoVYxiDZau5eUpc9ggqjcqH7rV1HLQGmF/U5wrd5TswxlczLknwCOM
7bn1bbO1cvlOouAgqaPTR+ZaPgPZBFVAo/OJd7tC7SqBCDK4ESX1Sr/EiJp0B0k5
0Snb9qCJKn/IMV5HqMyFJIVDj5xFRbGy0gDwYYbW+GIy8VYHqL+iaIDOeSXJ8+Kv
+NOcrumK98ClaSgMXxlumAsJpTcMiRtJ/C0pdQFxYjzg8k9kkvybUWs63eHMfpWe
yhKqXvMmOGYUHcFmePq4sB0NI1IkM9SFEYrZ3WjHxNoeBmYOPLveTXQ4AM8GIsEu
NWuEG0L3ZhgoaGxRdxjYOphdr5xQo15FAf1Z8MOKGav+7ffcoEOtpNrEKBM0fyyR
mfRzQ9hmuCNOBXCpSNFCvvr8quOFdktGXDl90FvIm7kC9sKnLdqW+zxo2v+CHUbO
PblpxyKUlsKUx7Jh3lEAfqaA4rKNTYY97az6yzb6OeyVJ7t07Jyep0Z33KYKoGdG
Y2VR7N9dgVyX2DNgAZ+SGQlk572NQbvxtW/cnAYDLISRjt7G7cwZ+dGsH3HXKDst
TCpsX00g3UO7hSobNPDSIHOOp3lktn+uLRblmlrxSw9ZxzXqoXdcP+IT8NIIyBG/
ZcrpFlMIIBTjG7lFcJ/b+eR6HY8EIbU3sWNB2TJvEJGRkY8uLfBt1tiR/Q1+n6mF
BgJpuHkXE84VOsT3znvmslhYvfb1YmlDdN4UmIifCQmPEiAnym2NA1KaMYeUj1K+
4j/SDGcHD95mfYe8modsclHtCexQxymVcam2mF4O5gYDoxRb8kraNnfNBTJGllRm
/zlSs5Jh3ewLNTLk74RNgC5arzYphsWwvHo2QfSZ6mBKBkWsCT3H2ye8lVPdL/e8
NGD4wXvIbNopukJYLn5n5Yy+hGl4hNLQoUWMQ/otH6EoPs01xhuRZUo4WJ6oaxge
mc/7KG+lQbsKU9SnMfcvzN8vXx+kVSN1VPJW7cBVZzyPIM/kqds/nXkqSUhamOuy
QlrDfSn5/A+WAsmw2ozoVjcl5dkvVgk9zfzIfyHf5s8ZDjLdWFSE6vHaP0bmavYe
ddSdbSwkruRKdOgZHoMHulLvLgbutZHuV9QlQv5kJKBD25sQ9GLhwZjKIi0uhZ1r
CKl3kbv0f+0YHSNheAGlx33U/TgtGoLlo8ICMKTC4pczfLf22uyUepQetZ1iwxks
pANSVxoeiuucGBaibNGYOYuWpm6SLVsm7eRnaAkewAZG0WdhPR8Ff3Swz/iRPGyV
kgrnWfGPYr25zOb9AwQ7JI9xVnjrnDjJzc5xYVIpoA5aCs70jS7CaTTR1PonftN+
0Xc+0U5k/VZji28SocmI8Xp0GuPB5MjYdQtMweZRi0DVu6I0BOLNfDDsCqnLSw2E
m11dGLYSYVIgt0UOD/zl/xeaIGXebc82auONVFNMnJfCiclxYhvtohY/d9Apx2Er
JQYeWiVAvSud3l+Cl8vSFvuVezHbEtBmDvJLdZiyYqgHgYSzBMPQXsP9NChNs5lk
X9oc6FLBMxW4/bxsr7yVSU8mT3YnVB3S/9gO5qejHWETZ8u7Awcx/4rC+wMBIjm0
5N2EFA5jIj5FlDLnKnF/v8Lumu0IjnwUWEyX9c8hn5mOek8sAO7cyUzscUHRcaTC
0//idsw+sDCFTSZksJTQnXVUHFCi+Sg8mSi8vHkwSPeefbo/a/nZTWJMO01NTapw
J6XEaeUoXuRf+jIEGeFyY3Watu5kc7sXheQZNtRbrIEYRgMjhT3kxQjuZIjYE7mM
lgodZivzOS/OdlIPblYF4cqiINU2S1NZNI9WLBsmICkqP9F72PpApIY4YLFVy118
N0UYAqllTv0H1TCXKxaFvWxhlvvAzixqM0z03MFmL+0WpLw3csCYw/NJrNx6U5HV
XcY5GkiLlEhciZ9kgUhHOGjW1derux5kc6DMjOG9cUtU4Qq3AL6iFZ2iw9faZUxa
U+57858HLbe8lmqHsm7iMjmSU/zasys24aWUOd7AtHHq7HaBdFXkuNeif9YrOE5B
Gjc/xvv2sxlONU8vnsrhWfuD9bv+54jJzpNyz0lg869M1dmK+MtFurPqPwRUVbsr
hth0UYay0HwZqsMkKnIfkgA0FNmHh6v2Oqwo1BUvsdqjI6eiWGVD636DukFGuSFg
8IehJTIAozGMUhsogJwbMwkrVq35P+x329PiVkOD5KhKtgsOu1AP16pR9qHYGW4C
rHn5IEIg/ZhyHXPF/LeM782gvSLwJaKDuFux6yAviA+uthN7Vu1V8U6D/9C9IkXO
25shx2x5TZgTWRP3dxFTWrEIGgiwEflifmiSSE8NAZuaHZhX6bqDqcSoZ852MfGG
+ge0Z7Q41XBzfkbSTgWnxU4kPC7vsQsQPSMvFdG63z3rJfaN7uhdNMUcvc2hVlqA
55Zxy0GykYBJOhASUxHh35cskvUkUYByHF5C0pBoCDCChug0gSk8rHAuvhYJgATV
wGqXF0ARkjumJYGB7muiHl+rGcJr2JSiYhisTJO9inlUY//bywiEuvG4vBGo4r/f
x3nt8gC3u/YnWm/EexbG9ywLONpXqhln2jsmCdHYO3nVA67WqklvfrIaedD2LbOt
/Kpbz2DIGAXk10l18egInvUKeMOokYJ7B3v9cyjg2Vqg77fide3KJFbqrNtLQVzo
Lrw7LyepV9cT+8e42xrIwDRJjOaNHoyHRg5BKVReOxthzB6QE6YRWaTdwH+3b+jR
m/4ZLswTAyve7HnOseF6dfCxmHvZ12Xx4PFZL8BAwKNpTu3OY9t3w27UoKfr8xnV
bIRlN0TlXiDNX6V8BJ70YANKNM5usvQwacc/8TaW6XNB26cnSv+FnISOM3LtUXCK
HjeZP496FM3vk5v7aGu6INnkwSIh+Dsqabw4UJCtBAioOZ5Mouo8GcSF0C4FSVBj
syvIEtcCM+F1Jdy/yhdxDsuoaKmjL7JknlBsd/x7O9CgxKFmqUnxPEvxQETgtKK1
yvIxEIusGWnI6WTcFgHqbc5RV3Y99tZIx1vYXGRRhgEkOoK1BoEaoEd6SrqOf8AM
eWjBrAaPDdO9VpD7MOUS3dGvUMLWG2s+byWf/iL1tF7ySwn6BnRbEBbjzeZEcbB4
A3LbIIZR+M6VrWLttBEy1hk/459X53Z7Dz61SarIf63pvfhT/z0Tb1gkOd/ukDkN
YzuUwLYtgfAfSr0FM9QP5UO3TR3aap65fD9vQGf2xClNl38hKuNsS6OW9kcskyG/
LcltApMx0C7XnPJttHo9rDT4F3Dlk3gXYYNOXwP3L3VhKx4q+apx/S2K6W17eeX0
92h6+iR9JyegzLCXxBYcSNp4a8c/50zLNywBspLvWH2nSUduB2V0/J+i29kWmF1E
2HoLZiQK45FxPRRnmaV6FHDH4dd8vVGSs/MLc1qwPyJLHg0mh+nlgoJC5VUNZS3p
g7lVfsWKmL90v0WHwgJ7jyYFSPt4N5uYonThRTcU+O1AAHmd2lUdjOUqCUEA9NkD
JzSM9plpLc/AMKe3+E4TfX0YVSzG+LyKzjrWXE+9hhe3RIPy+jKS1tmJInIOW8I4
f3yYE7UdRxRyM5aP3+PVyeciMfIneyvAwWl8abRl5lHkt8eZcsuzcEjhCNq6xr9e
XtGXcOmFheE0bq5QZkDz67ZZ0S14vp4vciB1sGgk3YaRAzUVGdK3BT+tH1VkIxEG
WiUgr4vKLXVo4d6VNQ4s1f9j2mAuGqUgunI5XdUF/f8kJBFMw58E7iSa0deXd7M9
62Hyi/cLSMGGul/gNHGGCAU0N17HF3RrOG8CdREsQTODzAkmHx9IP06WznldeYU4
Q67RP6CbC6fWlhgnhnFEgGO0P9Hl2h5cjG6vgyFePrl20oS4Xb1URglfUWFObpTY
TFQ34t0/5/JQi3SOUBvlRSSuQw89IN5yQlDVdYEp1+Gch11WWQIysiYSzk6W0rmW
4HcU9oHDm+/gy+xTKPTfgoRPGGJl/LM7UD1hguP5of74eSz1QH/0dEKQJBa4L+pH
p0WzQojBZovhM0pQ5CZ+IoqDds7EpiuaR0a/Su3DOpSwJLd9sdHo6SsgkxmnHDIC
i8P7ND/dw2FGTZkG8yiM5g2zfB9HjGThOhO/QGOdvWp887h9HWRqn6KJ/jO0Myqj
zaTn9qDkYjQbi6KWeXlw4lFEAhWCVBFVPPql+4rKpH21aV6YZE5kv3x1oEEWxaGr
rG2zm4IdeCInbv4rzU9awUuh3qAyml0zU93rmyp62/atXPm4BwrWZ94t9Fccz0op
JeH9/oix2I/NLwLgYjeFoBV2orzBfdlOaQ6CbV6h1L9qI8irmSiDJCG9NTui0iP3
kebMik7ucvPCc0IjeU629Cb+FVV5XBNouxgABNy+9/DkoHR3/CqqY+O/IX2ClEN4
02iZQ7tl+g52a5p2YedpDz+1aLZQOPAk+jYrOJpZHIAMQ/TdwGRFdfz5WzEhw60i
+wF8JjGC2qZpc66YvHsT1yWqgGIDDuIJQq7xbPcofR6fY0rjSof0yBzAENg2QyDk
DVegwPcHZnRZSqorwFPH5XPHTIwFQgd/ARHUCpkCQgP9yHd1Lr/1rb5qdfJ5V+/K
OtGlRs+UZjToxLum/fIUyzVcCbRvXUu5W+/aaJjddrPlX8r4LvoVqwBMi1K7S9GZ
ghNwvhyaLTvQUyxoCzgJRnMfam3ssuvwAvrxuDGr1uldkZ5L1YXUgNo6eY7D1AR+
OACH5DlpPTjC+TYUqhWEBhE5BvGjnDIhD0xCTy9toe8YD8pZvgjkFbzvkZJTtWQx
+Xsv0blYFrTvM06irvqYj0r7cMP2j2XSdaL/vpiAxwjE9jwA7xc/AUDjurVUD9lh
CoGYSvXcICidbcoe8vLUm9BrjEi+92WE6CQdKI6SEfefuetNB1PmYv2SiEUXrYp8
sVhHgh0v/YAnjcvsEbVPfUqvcPj5Z/pT6DWxukhxStUghLVjnmz54qg9S/CSPCHo
NOZRyaGeDccKjt/AWBYtx74xG86PtkgMO9to19zTEGGMEQxk0480jWvU36+wJ4sV
jw6dKQ4fJQjGzMD8LHSOyHqNDRQMzNwQxZv1pCbojgR4fIOGPmdd/zKiH1sRwDxs
jNkAxVqzdcnJZSjmpNgNbrVHCvTYAyR1MqwKSdZV9CV3V6D5hXRIbmXIgB1DFuQ8
AeUp/PFySKHgGAb/0g3hsIPGWslqq1vhoe3j2J9mtmTpdip+2M01vwXwtogXP0zv
xzSyN4Pqp/NGA0mkTEPYjBlDj2asS9dRxm0qosuCCy004rwjgasUAMXizHQlT3Pc
Edk+adsEsdmYeFvYuwg7fu5rnM/e5sltZaR3arm/+EuK9WPbP6NAHQSQMo8XxnPv
/r9LGk7LdgRvUyN7EOT5zOlNpD2ZOh57oAgN40vZXwEk49gRBgRS1F3nAATAVq2u
c7GQT7dRXQrN5w2rO7/bmSH94SotEa8eoxKxbysEbRjjQjguljhm+ryRLUWVOd+d
O2fzgWlBfz7QhQiHfnMxpKnMape0us9SzhYDPOD+U6OosMqYrQJUDpyEYeeNsDsE
9cB7TeJAexh9JPXRWt3qOZROcEMVsLckDgJok5uLAW3u3R/kl1oQFRRHgteoGKlG
novt2wk/ZP5QbAYeiBOpdMI6bB6lds0+yVgI5xkpLXeWUyD8NjXJqagge2mIuCBx
N5jkDdVizdHpEERWzk3ZZSxmPKLZcs1XZByoAkdHEUxsObn3VpRj9oF86ZV0UPsg
ATdY/IZqmfeuBCI/ZroN8HQ6lyLBLpTWKk2FzZJJWiV8eZsO21iEYN14U7tmgkgF
1MKwA7wA3+AaLQlYY6tWFJcYn4opBBOKghdWn3jNkxV6JNcl9xuUhI0c9b2wbdVM
47/k6ErT1R5EQwmLEbTeGEe6CO8dTA/3z/rUM3rmaOMsE7Lup6H/XsPGPK9Hr1lj
iNL1CtZVULpfcYAjG44RxLm7RkzUZTKX7oYrEUGbZzWa5GeN05vdy9us5nye+XAk
mGCEJhMpZQ4kj6pCiwrh7M1mPE4RRfHzo7hlDg7XQVyCDmkzARzYLpeNKi7hEV36
+coIxohgLIFMfgW9xnbucA87v0Nlk6aShmiEQKRMahOAUMHIU7lhwsZFBwNqH14d
u1+0Bcr/Jv0Vpdk9KYAyHurmIO/IY6WYdHZRgrGCZEh6ZS6JzGrwqrf+2MxTqyBB
eeWOZ7cf82QRcKzab5nVUt78UWGByABOZfKciTh7urYevpP/y8YEM13g4AT3g9Fi
Q58m+FVpEfIZtSq7iriHDPH71IElwQ+g7kat4vA+vAlgc56WQz0sViyQZwtzZ2De
UZzvnhcEDpfIjN6iaYmNb8U2bPxsSpby+7nD7pjS94Yl8MA15nvZVyUS/thT09nE
QzBEwlken6cvbVCXGDc3g0dPHKwS9y0uxPFyexnZlxISEalokzt83OYINJsRzDqs
t8JaxO9SrLljCkYNo/MkSTI+/AalcVI/MrMQ0GWqgxKfXcBvGU0uUDlE1L40YaMY
F0ve9SbkEdXhPCYATBNTYYytm/c4ZpH8k1LyBALoo66pPvps/kpxKmMw3Ag5lX5h
XPLP50zJJhbt3Nie+dQGH/s+oNO+hNfqzpuKt8YJJe+oZ61wo9oEpwGFnkDrnSl4
MPp/+x6w0al5ppgD+03kudmB41Zi9KiA+n7glHvdGt5qimAMCjQgl1/I7AfdOqTD
wHCmq44WDog0pDEGErx/4dIIEDYtr3TyAexg3B3vGUCY2pFbH5+fKLO8dUnb2nPD
f8Lph5ZWYFZA3TzUc5Vz1LiVT4idX4qQJhmimuN5lhnK4xp5sM4pSYx9TUtwZ5oR
mFWG6m3fNxpRAHqThbvSs18Kwy5qg2FT5U2oVFQbjrhG3FCNvAEeuJ/5aWDDx0aT
nDi0CY/qkMNMSTM3vWoXqZbveacAavNcB+BOIn6Y+ezT7uQDwlqUofbcKI6/EN1s
eHrNAkqYMwTO9YIdG9KqCAFNHf2zXdr7s+syy/D9u/hzA6bj3MmBpsQzL9BpgCRr
3Gxcec0Vi0rAoT3Y+NrO4/vp7CHfznoULnduYzOY1P2Sm/0Lh6jdBl17Lj2yIrqK
c5CLxnfsA0STLaH6Fb7TM3yGku2V3qSmPUAzznSRus1E7vaxhqdxqqY2kOlaiM/C
8TPVoAWn2CF2jDegxWsfTM6Lwek+faf3fCBKuC17m1mOg2nr8NIMqtgDjGZDu435
j3pRiojtUXFhB9QdCitOLisCm18jTj3ZjCyJCE0pQkLMYIXk9mPGQbDmn38lwqyI
IEYaNngddTZ3VFXHdITmbt14mJC1zz4qBLJN5iXi35MmSg8TRB7lFp7G/7Pep+0N
XfpwSfBbJiD8SaXaoeWsOInxiNkVgVx9fC2z8Ut4hsY5af9llg8PMqUOW7fJTSs1
37x/+yqQbJcysTGBYB3odPTCoMoAh4RKvm1PH55wQCKlS2NO8Ncd1JkvPSmeaOnA
oaVTXSdL0mp85kxw+kNj0DBT5GcrZhxo4GzUeCC6Exg=
`protect END_PROTECTED