��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���d�v����0�i�=\��A��?��� (��1_B�f�	�Ѻ+|n��y��Q4�]�aY�����*2�y%����>��������K������ �
�D��z�z��C�y�B����
_�U��hkF<�~x�ܕ�c��P��OK��F��/�v�<j�}.[�6�Ć��6 �������t'���5��(n&�4��ҪX��Zr����r36k%ѾW0U&��:t�)�s��C-Uz�#T84�^$:t�(�}�N ����&U���� !��3���>|�{��z�qZOb!�$Z�h5�}�A�7$���D�x{��>8�t��> �$��o��?�͵�O�`n"*;�L7��TS~?5�#�H�|��<,uS���TJ���4�����4��g�@�Lt���uSV�_�������LՇHbE)�*TdlJ��T���y�Np��!�м/��Pk/��;1"�7SM�kZ��|9L�L�j7���ҽ�p���԰)0G�O�b{I�2m|�,�.��(s(Z������ta ���%�7����P
4B0�O�߂N�_�̜Y�KhF�#�Y3�$�=w����f�ך�?��&o�doPI;xi�W��$h-ш��^6�����1��/�	��h_H!�I�)�&���s�A8�_V�|6u�q�����]��I��ԍ]+����1~�V���÷o[��MH�qUh&�¼i�5LC�=MXq�$d�*�[EWԛr>x� +���O��_���o)|/��i�̓�A�o1G!K���\�к�twgJ[�Y�.;*w�Ftac^�i/t8�@.�� uJ��%��4$y��p�\m��;�.�zg����e4R�^�4=�����.�)G;Ir�"@� ����b��=�"00���� TG�4�I0?
[2��(:�Xu�8�h�)�:1xeļ�oF
[���7*���ꋵ��c�Y~ъ��T����{�z{lj��jK��,/�E�7���(���h����[X��4	%Ѹw�S\$�BM_�.�9bY�������}�� O�'��ѯ7��1���E��b�����+	���B<-��(}�|�`��	U,�1ע���a���Ү�+@�g#�<[D�U��/�7D���L�,���^���Zk�6���������=�W��tQV��fC���;f��Z*˲��u����;�V;�Ћ}k������W���w� �K��6ʻٛ~����>o�����Ώ�9n5\�7$I!����F�!��5��&j��`��g'9���F	�~������+�ms�\>�e��qM,$z ��L�K`�ܞ	���7ĩ%�oΔD��(0CL^E\����r�'dm4߳C`oA�+���.r�Ϳ�?;7��F��K	�|�����i�8}��y�Mz�>�����O��ƓvW�2k��9��w<`���N� ��O| !f��;Z�}�T�V$�������D,<��;Ǟ��2Ӥ V�'5Q$�g�� V��M�{9��f0�]�J B���D�꙲�%�\��)X�ӹ��R-�<ri�vCI�`�����R��:�{Y�yؐP��$D�����R������p�,	�1h��9QX�?NJ�6ť��u+\�b�/կ�0!��0XH�`�ӈD��)�3҆93|ԕ �{poq�q�v]Nt�]�~���p��s�~]�qo�Gjc�逳��[#.�c���n�v��艸��F�J>�3�Y,Z��,�C�t�Z"Lyu=c?�')<3	_��!3�I�A�%�8O=����˲|dܱ���]�n��-����=PsN
��T��?+,&����������j_���ς�<���^g��$�ѐ6o�+!DzP�te��.����Ҹ�ц���JOլp{����wq'�d�"��lt�Fu����O�O�T�R��Bo��Xm����}L��fb^Ą�-�$6a���[O��S�2l��Ы�
��=6�t+�K� u|}�c�����&F��Ɖچg�Z�yWi�^Tvk�2~�oc\?��]Q���g}JUn�Ɓ���x<�SJ8�xLh� �|�[!�x}�I�<��Z4MT�w���g������)y�rp\�G�>AT�>���}�)����K���T�=���ۗȳ��OaN����sN��e=(���Ͼ�e8y��'�i�Ԇ�&��`���#�� s�009�_#�p��b�t��G�}����;��,��.};��/��"7Bg5~��.��CU�A7����zҁ5b�:�'GkđVe�6,�+����:D�R)ԋ�����k�&6J3�D�j}���z�t�X�cm ����s���v5�{0���_���C�װ����t�eX�#�VN�8Ԉ�lf�!�����z�j?�	��ë���1<�Sk�+I���{��$�o�D'����p��ص��#Z=֙�*��P�[	����8|A$�z����9	RٿȷG$�(���_��ҏ���[��g�0#��������N&/���2|Q��? �^�MpS3r�y�n�+C[d��=�C��0�}5���X����t\��8�	��$sP���]GK
��lc����:�3UގM�cSQ��rlm�Ќ�OR��Q��'٢�S��mI<�<��y����Q[#��9��:�qCB��E���b��y�TՑ0b���7ؐ��!�����<��A��=�|:�?�}��E �"����+�=h��T���礇-_�V��{9�����x~�A�A��� v���JYZh���=��(�����]����ΖN�r,��/3o�m���˽5��_���&ZA7��&��D�u��l����4�ł_Ĵ��<��Y�M��d4��w@0�'W��p��p!'o���Sn��:Pӽ��دY�i���Fo�\Fz����_%��13%@�\]BR��K�c�`Re�'`)�"4��G���[p	/ �CW���{�ѓ�Y����![9#^��K�bR��r��욶��X�!s�K��+n�����Ѐ��{`��ma:�����\O���T4e]� �>4!�<Ƹ�L�2J�-5�?�(^����J9�t��F-ҹ����Z��n�ud���sxi|Z?���[9����9�&�KLg@�����/������%�1k�i��u�%C~�&ӥ��Cn��	��n�����}Ůd=���������+P����tZ����.O��7 �̗?s���ׂ��#�1}��a��2v���LGM!�l���s�n�5w�(�] ��@[5�-BK	M�0�fZ���(�x�*�">Y��m�j��J���cDFZ���c�W0���z�.�@����� e���� �^�l0�]$:}ǩ
�������[)�΁��q��!3O�rw�&gt:��cơ�	1<��U#����V=>L���v�-"��E���/���_���S�;�w�Y^k��z��я��9�+�jm���<���	���t����~Q{몥��f��E�8��ÿ`�b�!���|���1l�P�|G|=��|�9q�R���&'ktt�3�o\�bW~bG�;�Eԏ����6��C�(G��7��k���}<� �'?
!F'e:q�>�t��)��q�����do����K2z�K��4��\#Q�̔$,4��	��oO�<�8��n�[_�� �	����k���P��>�{��L)Ӷ�&���H�(Q�@���oqVu�gRT�9.�.����b�F�Tr�_O��}�{�.���W�###���X���X؞rs��I<���C���p�AL,e�Wj��&�����?Ȍ+��{}W��5���b��Mr��;�<�w��5O��i�-co�N��������'	���}h�Ůc4�"�M��z��x����jx8	�����Ar����@��(u�*Fh��қ~ȘK��5*l�`}��L�M�~�����ЇR+yE�V8���;����.��6Bc��O���K���jɐ�i�|�-&jH��b�?+��ф��"|�
���I=Y�����p�'���R>�<yB��a:8��ZyQ��6ɏ���;�U����i��r%v�??'@����e�r����	Z��.~`��\+F��{t�F��;(��B�l$�U�[�\C�Ɯ�P���	W��>�q������I��`�1 �ˍF����:h�3��3jl��ٙ��m1i5u��8iO���L�`+�K��R���%k1r�؋���!���Z#V�|�<������8�9K�� ��\	+o�G|$'u�1M�Z�u���*}�R����NР���O�d�Ow�B�d��x];>%��	ϒ"�X|h+�����f	��Ë�|��m���b��D;jD����P_n�����]K���Û�3�������Q!�A�Bl;i܊��K�۱9�63C����	��5��UB:��m����'T�����<=ú,]��8�%l���yͤ�O�ёO��8��uGw>Ǧ�@�Z���+��M�����lrwL���� W�Q��=P�!�Wn�{c�8��s�(�&��I�B�6k
��l��i��!6ZU���d"^4�2�5��+�,AJ 7���$#mgٖ��Bh�+����D6\M���a�d��n��3��Q�pX��-4�J���Ys��`q��E۝�2kH����;�۩��l��,P%k*��>;�d���4���}_����&`xF߇��s�4�vi;6�V�0����[��b{�S�gx<#q�����7c��3�'z����7i�DlAƭQ�-*�2r1WNM�+V��8��o.\�~'<�~��d����4D�&�Mj����'��z�Q��d�.��ፑ�W�#Z`X���� ��^�z�5�5��)4XAs/�i,�9�蔭�];GESHn��L�R�����k�bz$"�u�9�%�la��E����ʋ?J/�P�0t�>��ǩQ 1:	�ҕ��Ck���=��,��˼��Y�L�2x�u�W�|D�m���0]�B�jc��db�ޯ�v�B�pE���U�5��X�XF�yHupY��������S�
��E�v-����	7���D׺���^�^YH]Ҷz]�5Jr�;Yk���؅�BI�; E��N�n���@4���ԟ�x��7\�ʔ�s��ү��x�{�T������^�M���H0�LV�\�t�3~*oDq��3r���ښh��B�}�hx<��$�s��?~��M�7_��V����CZ��PP���&�:�B��ܕ_��c���~��)ae��c$�|�V�_q��A �:ɖ~����Wҗ�<,�m�Y /x(��	2G�OnF�(���g��.��`6q�@�!T��.�+�Ku���ҹz����*}v�]\HHb�M#/����M^u?�ď��r���VX�J%��~�#��<=��2L�^@�A	�/M\i�P�] ȧ?bZ�l�Ê�*N��׀�&��S�eO� ����=�nt�3������iY��b���杖�G�-B��}��~y�-�*^� ���kS�D�	�#�?( /���K2��G�񄧂�VN+���onr�al�����=qי\}��X�x����D���&?�����e�d3�&ovj>����\���3�6���m�!��'�7�p��:��n`^07��y��Գ�qA��Kd�"Zt|�E�Qz�冟�$2!!v/`��D�
�&=�$�I�t��oS�#	!��.\�mTZ���Jd��ݢ����!E�6�ni1�ʆ�U+���wEV���=�I�e_�S���]R�U"�����y�H�%����+! �ş�U�zw������u�ҕj��%�cH�v�E��r��|
4�c��:%(w�����P��W��r�#���P��nv9,s��Ըm
�g����K_�c�g��*���uI*�G6�J���	(
S/b��1��l�Kܴm�48�R�㐦'��c�r(��X��wf��p���:T�p->LR���k�+ҳ�](f�lO܁��$��>gJ��-Բ7N�c �+�s����p{%mc˿L���Ͳgt�8�e+8��k6Er
���'�pb=S�i��W��GX߇��FzhcX�[�0�R����d��p<l�a�*ﱠ�䖣IVGx�?:-���A!a}��`X�vh�X#�ɁU��6�π�WET1x�q�>|���˕��d����j�o~+d����l�
o��Bڐ�����l�^��`M���%@��
�B,'�OE������t��`�2�l��q~.�!W��Rᰈ��C��|�}C�~D\�F�&J�����1��,��Zڏ=Q��/:>s����3B9Сu1z~�K��W to�)Ǥ�m�=�~���U7ചO�!�2V���U��۹�A�	����,����7琄/���j��d�u������b�ŕ�D~T?@��E��@��0�N����P�*�?}�l��ی�D8R��8y)�G��V��4ؘ �� �0�`���"غ))L�"X��s��#dO��l{6�6��E���䍲�2�d�պ�,�6��7��H�a`-�����i�wè!`�.[.�`X�ן�{WN�Ӟ����5��hј~B�¸�����X�s����2(�� �"��u�{�e�I��F �	|�9}�Q~q���j�t�`�:�C����Ӑ��(���S���k�%/���m�'T�k�d�i�t��:�s{�?�,XpM;ve�ٴb�A��x�u�ɪ��i����J����d�WP������u�N�&�S�C�����J�&�=E_�8�4�0��	�����K����V�%���!��V0�O�g�=U;�%�\{ ��9}�v�8Aeϴ��+��_�#N� �
3��˅Y�A 쟏'��@.B+G��4��#��QX��l�4�
gz�藒�r�������u�*Ji��V�z��JlW�I�gvW>�Е�M���%�!��Å>C]䳂%�..�KU^}*xlhg�
g>@�s�.Θ��b4Ht8��[�Iv.�*�6h����LW��n��|�I�!��3�`���0�N2��;��l�A k
����f����}��%ŧ�uz'�e�4��Z�\���{��j:�(��:K�/�~��W㢓L{t�)��|� �*�H|g]�+���^�������C%�	g2�UV���M���Y��(̉�)T�`�q��M���0��W��l���L'L`���h��9�������6��Ù�JRב��59J W1F���BT-&�.U�l�B�nBD׃4Mk�k�V����,L|���bV��O�����=(�{��P�8E}�4�s4�64]�?v�5k�����h��kj�&l�2l�o�����<�Ƞy��ͫ�J��}q�� ���%����e4��%�ƬT�	���İ�,/��@��$Z��s�5��WJ�#�0 �1����������z����!it/gN����h[�S��ܽ������`�SSw�1�e������h��F�FϜ�Em��),����Hq:�Ը��
��Ƽ��F����'Yt�+*^�6R�QQS
3��2����%��(!��#�-�P�0:Uo�nб��]D'�i:��k�$b�@Ás��Fi
�]8ن����@��V��:�� #_�,L��h��%8�z{���2rX$��yJ6P��g����)��9�6M0q1��׬�p78e��b�?Yn;2��I�nZ�7طtr'�H(�{\�%H�H'�g�X6���'��`�V+~T�dwQCm;.]�Ƽ�~��H�m��Jq�6�LQQּl�9�y�uZ����8'��a��������Zт���O+_B�Nlݓ6�.1�Q�L�S������G=3���8���2&���������V|-M���I��<'��i���EO�w��8�3S�	��jS�w��(Q]a~q�X�gd�5a�+�D�Y|�l؏^"��ן�q��-k��t��-At7��煀�$�F ��n��Y3@iL^QT�*o
���+)rEv{���;���|���͗![����&���O���[?�.g�!4�F� �_R�#����j�F���t��:��Ձ5a�&0�+ ��.�+fˬ(�0���@2BH������PW(��4e\�����tjcn�߽P+�&Z̨��R��5�hA)�(y�W�R�V6���o���/Q��[����N����o�lQ��K�?�r��.+�q�}s�m�����iyR/���oh����������qV:ż�<2K��T?�o�;V��گ�k
CQ-b]�{?A�{����F������7��Dd��� zHrv��v1�S���I�v�k��'[q{>m��;��H+�ꉕ�W*H�k���j���]��?=F���pp��<C���M5�'DIy���'X����EWX�>Z�ӯ���ul�xY|w��U��M�(�f8���Xe�����`��/�A�1��hs`��Β9kj��
۩�WD�RZo�k�0S���p�i��$���� � ��ɒ���jfڶ���E������  �y�yJ�p�m�`��<¥�fa��&�_�/v�ё37����L���C5���Z�6#�x����a`lP��6�E�v�&'ɯ�c�x���.�cIv�K͸
g��ur�ט��U&nzgnZ��M������ �OR�A����+y�+Aŀ8��l���1��=��X���^����E��8IV~|V"k�&� �.��Rkd~�d��;��g/E;e�-}��O1�_g+z%�||]�.^&T�˩�Q�P�+ ��,w�:;�V^���Pq)�&�u�
x��9����b��ϑ�*����N�.�x�0��p����5=�9�XUµ��1ʂT�;m�-�-�y���+)�H�P�z�9F��C����A�^�;�~���0�"��>��15dO͍i,=r��[�c���w����
ٿ0-Ƙx,�=�O������T�c6� I�p5�V���{0���4�<x���U}V�� e����VY�����X���qש�0$촷�u2����P~�)�V���;vF6f��Rm)!ɜ��b�GaQZ:W�Q=�V�V :��h����y�֮;�+����+�1��=�89��E�v�R#b_@Rm�[�d.�S��i5_�ܢhg�s	��@���	^z�g�Az��bo�ވ��;�����z�^��E�Y���]�UrR
t;�s�̔�{{��%�3<iMc}��t3,W} v5r�,�Vؾx�G�F��M1o֜08"#ug�!�t����
����5���o�Y�É�T�Җ����hTB1v]r=�gha��ۦc�MZMg��S�����.�E�T:�����'����G���H�ţ�)
�U���pPY�4�e��i׀
v�>Y���K�*�U�鑂�XΣ�T�m��E�2p#kɜF4�d�K�N�к�8��(�NY�7�V��nS�`�8	�U�wKFG��;s��P~��bQ��V��^�a"g(�D��l�tè�%E�4����v1�<`q�
0q�\�� 9\�n4��!�f����l{s�q�ڕ���Y
4��傽�a43�Z4Ե2��^ؼ9Cy�+�g0\�9a�Z)��^4ޕ��1��A{rf���17o��
E=E(g�H~k��$&�\��n� �ۈ���i "qF�y����?��Q*�J�����`+^?"P��c����Yp.d�
5Γ�����^�l�^S�]����ˬ7A���ŷ�v���Q��K�}����QpxB����5J1p3��w�R��l�Ә�Tc���7"�C)zB���*rv�A/=��fG;�����$�R��
GΪU��Go�R�xzt�ۛ��dVViQl`H���DC]o�A�z�4"�/���E�bX�EdO��������U/q]j�����RM����.	�&W�,���:vC�X:�qA[�7�ӝ��(�
6@ c�ěK%@'������q/=%4�P%��a�匎�4^}I6�w���6\)Q�X�L��ձn��u���zҝ�0����i�]�~���րv��V1lk�1����A<���p!�Ӱ�a$Wr���.vv�Ϧ��1*uǧ,�U�!gle��y�ڵ���}[�`�Ϯ:��$�w��9M9�����U{9��;)h�6O���ٜM���&�3����G�\��Fб�x����U �G;�V&�������Y��Ӹ\����d|�!���Vz���&�,��F���.�=��>&��$�~J�Uz	���?�����A���/�#U>�JI��{��-�HSr���|�ƹ�I-� �#,"	�En�Ҥ��G��m��;�V@�F�`O��O�DPS$m$~ )Yv�C;��؟}�`��̔�:'e*�9��mOҵN�=sC"5/�<?�G,�~D5�^*����E���/�=<b�,cRdr���/��	M�9��U��أK|�Uq��(�U��]�¦<��ʹҡ�/V-%
7<)vt��&���>����j�	���U���>Wu��!��P�)5�h������ �������8�)бpaD����l�\����R��;"�i��H�!�!�"�3�QS.���/�9kw�{�;Y�d��w��T{�}+C�9�VA�p���]�:�J�,�ao]�P$�p7�T.L'*��5�\���� j�cM{�������T0��K}�>c�u.�x���Js.H��~�>�I>#��:KFq �tQQ�_>�hP<M��K�i��;moW�X�$V��.HG�$Oj� �� o�G��ޓ�P��|s��V	�B�/^�RJ�P��5��j�`UoI���A������^M'��+ފq��/���O�f��:���%z�#b����HH7��5�H*z@��~�&>7(��<��E���r���'C�ok��|�Jx�RZ�W;�Um��7֦�7K:�h�묱�)��vMa,��U�B�"�V��r�H: +�
��jB����h�k��9��b�o���D�G���BN�����\��j�N5%/*���2�7��U�?�����=�V6$~#����'��yoG"�q=��G�S�E|!Cq�U��J�W>|f2#��gm����ɝr歙�n����9Ǜp��Rj�&���1+$b�i�;?�Wy��VH-祣Q��/��{�@��rI� ͸3�3��D [�o��1�߳_������n�}�$��.��R`�)Eh���e�Ou���,����T�Q�^mV��W�J��*�7<MRW)
�=Ф*C��5�ͣV���R�P�7+�e~��YGו��ol��A��F9M"�'ڐ�ɾ����(��fAq�§\.mHam\�>,�
.���%�����V�e�7�7���qPx#_�S��޽��^� �A��;����f���������]�+]Q*0�Y�����z/ڃ�ј�o�Z�{۰R�;��w��"��	Tp��0�FÀ�1e����1�S�pǺv6|ͽ�M��2#4y[������Q�"�SA�����%@��l�Xct@DnXj3<?RκԌ {�(�SmKJD|�_�n��ӹ��B���G�<(�:B�9��PM�$'Et�/��䐍�(ZM��lPcc
�	���N��*��ǘ@���(@�J'��x"��^����:%��d�I�Y�$���*��r��M8�/ �����K�4[���{�*�Oe,I�wk�ۺ���ۡfE+ߣ�wN�ǫM tw��
&n BR�N�~�4��V�M
���)��~�.��n�~�V���1c��M��P��H_#%[�A���Ưu��� ��	��ua	i�-��l� ������]�D�Ӿ(���ϛ��H�rZ���i��3 zro�cl<��Y�tY�|MB�>;-����dÄ)1�:{�2�G��.�Q�c��g��z������Q�6��[fҫ*�$���s��:�D�:/�I���Kj��`P�yoՏm��ԯe�eW���핾�JT��}�o% ��Q%4�_XI�Vs��&~��Vp�Il�����j�;`�MU�>�z�y�_Ad����{��ө26J��0R}e�����z���������M�����g<*-D" ���K� �SBP�0�Q�ne�qx��RS&+Un�-�}�B!vb�a��%G1�[h{�wp�q��|��|_��\��7�	��WDBvn����Ο�����jY��]��|���	+)�	Z@;(��������kDZ�P��N}Lk����w�',�we���ɆD��@Yj$�'����f���e��(��5�^h)Z}�>���B���:��N�Fǈ��|q-���C:^����;XJ�~+�%u��u���Ѿ�����&����=AH!��]޲� �1�A)r�0�1	n�,�u�ݶ'n�sY�jӱI|�{-��`"v��CK*d����p!!�-P�r7_<�o*0&8�%p?QUBۮ�]e_���rp��QmU��m4#MN`S�Tary*��b�r)tU]F4�۞<���2�$���N����:z�s�ጻ��	#�d�	�AŢ(=Z/7��`�`���d"J6vy�@��2߀$�%�|�8f�b�p~����6S�TUDj;4�:�4r���dj?00Z&��-�%�py�!͛�/��d��,囻W<�qhyߞ����2F�6`�_������y�m�)�H#q%�p�G�we��u9|�P����="��Z�
|񕜌�\i0�<���u��#�[z�0`/،�q1cV���e����ؕ���ݏ�������b���AJ�%_����7��6P�pu�i�=T��|֔Yĉ����NQG���A��s�������n6'�S�)t�Iΰ���t����]Ѩ��φ-�y4s��PO���K�l�.����7�J���p%i
9:AVx��'՘�7��f)���i�����p���{�.��͠`z��GdL����˞�kǚf�����D�f��h�,<3���3��O;��ޙq�ׄ�u���DH(+��N5Rf͋��q=�,I;;�ڤ��e0��Yn�j�P��y��(V�m���ԃ�UˮW�y�B"��D�������*>�N �]0��	 ����楪+Z��v1��p|��Vj����	?%�q Tn�{`�����mE�����na@b��� �b{Z��SE05�0H�=��#�0��)U�J�h�~_g�_�֣���F:���,V��I˪<����-8�}VtC��s�����͠�X�"gʊ9�)޵�e�7��ɍ2}��	L�$a�W(}<��+�1����#zu
��>�����n�'z�f�Q��ɇ��;�7�K�h����c��x�,|�b�m$8���`�F���4�ɵ�q��?>��w8�&r�v$�w�t��h�o���۴ݫ|�S��	&���9�fm�i���R� 7�O]?��sds�b�9 H���.ލ�;f5#%zk\��K�n�s����5ƻ�8U�Iڈ�Xƌ	\�ъ��?,o�&D����	�b3��}�#��D����Q�1t.��<>�W{j�m��Q�����)�	��~��^Je�Gx���l���M��yW8*��4qH�� ����ƌ�;nfK	�^��o�ޚp^ 燇�[	:�X���&��1�"�$��N<h��=>� �q}߂6e��qs�+�
�i c�!��d�n�ԯm�B�_�B�]�V�df�:qq>4eu��UDC�ڛ�XYT�k`2�_HP�4Gᡂ�]���|#-��5�� �$,b�X���H~���R�I��c]�W�˄pD:D�Fp����g��>O�K��g.�V�^� �󘗀�x(�?�sL�Çq1�e�c*���C�u4�q�+뙼'����I�ʍ�ǥ6&Q��8�CU��1����v��ֲ�����!�C^�I�\YXWM�imq>Z&��ג�b������R���F�|�t\���N�	,�)X/P8@��?��B�1BH�,z64��E�&�e�k�\�j����/�����X��ᕼ���-0TA+h�q�T�f#l����9Za3�sy�/w���fxbc9}*.�Bh������؍t�������'�#�
���I�W�JC�O�(ل�v
Qa��<A~ocIP�Lvg�&:𤞗v�l��K'	D�L�p���-��@�HAsj�E	5��zϿ��?���X�z'V�yF��qs�����t�����QV��t�Vk��ufu�eN/��^��fڊ�%$�fR{���X�!MG�,Dz/�̗*,%qG���k/⿀џ��SF�A��z�%�7I�WqF ��AL]$��ecD���;5���.'F�R��tC�W�˼JݾC�1H����9��������69�06{����Г�wR�x���-����gZ<T�EX6
���/t({M�咈(*�/T� ��r��2��	��L���@���!A@����;Cڼ���X��-�� .K\ts��/��Ur���kw��͍�C o �:�&���L��l`.X0>	��0aM��	�M�aRU��AB�����&ZT4�\j\��&���c�s�pсH�����e=g��ZV�a&�
i7 �1�����"�D��,0���$���h�6�3᫺f�"|7!�����\�#ĥ��?h�K���z5���B�p���y�Д�ݱJ���������Y��eA=('p�Ŏ��4kp%�����(����E�8��')͵��&����I{Q+�d�K�P��v4���_����� 2� n=�<QubZ�O�o���!�o3�
����m�k L�m�?�EE�������f :�;�ѕ��>{�qr�¯l��C?C��R;EE�{A�vGI��Ы��=���^V^.��ʻ!gU�9"F_��x�UO�'����%$�:4��
�`���C|pj��
��R�e�����)�m��d�?j�W��F^��VMU����ŗ�B>"�Ѝ�'I�"An9��m����u9��/ �`��ȋ�	���Ӿ6i���}�����V��"� !E����h��$f�\7A)98I�h�S:�:�E!h���)��)7}�b%�/������05z���`�ͱ�<�ƛ��.E������������_�WL�ǐ��'�j��X};yklU��L
��0#|M��~��t���ナՓbU�)��5�B)��p�zV�|@�v��I��۱����^>�G �j૱:%���|�}+$W�����k�q�uPݘq/e�L�L�0[j��g��3S�\�K��rb�k��R�ȶ��'��t1�O�E�����tN}T��,���7wp��lO�$<\H=�����?ӡ�5Q������1��遮���3���ҁ�VZ��s�s�i�;��ik��eo�DU1�ϱ�S�Yx/����eԓGH��i���j6f��l� �f+Cf��G�IB�m3E�708�I$�W����:r���#Ѫ4v��.���A�'�ay�tL^�
Ǉ�?QF�"�dNʈ�`$VD.��3p7���	I�!��	�d�B����f�3ht��EJkaܖ�J�'S�8=�d���sO8Ch@R��8��9�f�,�L��t�<��f��;�5@Λ>Uu��6�u�-��u-�{{#��KvY�OYr?��T=X3{��y��f�"َjߓ�T�Xf�}I�W�`쀴Xe����:q�ܪ�e�ݒ�u�vʟ�xz۞ &`4)h �yi�G���k��GR��[����%��}M~'�<������dR偙�5�c/��)$�
;�c@�/,���&o$Wp��o��߮�_.�"�@�C�5����"��ٜ5�={&o@��\=s��8�������Y�:O�te�I�q9�W��g!_����*��9�z�K��<-P-�L��n��$�`���Tx��,*[�i��f�X`�:����p%����:�ǶdU����#�����D���=�/�r4�/�9aǙR/�U^�D8�]�ی��&z̵Ǆ;���x�p���h}7�(	�:|���:����պ��E,�,���~����3�4�"��H��5�t�^?	�J`KSbc=�;8XH��������U��m�l�	,G3�˛:�{ -�|�]�uZ-k�M�SmGlP'��3s��>�lެ�e��'���T.�'`�yK�&2�1TK�e0`N0�� y;s�V��9�iz��!�j�*)�iy�[��{�\�mb��%^�A�#������fn^	�s�O�^����O��d���R���&��N�i,ZBNW�k�2�)Z��l>�.�Ǝf�U�l��CL�U)T�6K#AJ���yd}T�t���ւV���#̒E8�{M����6�3�sbz�O�}{��,�>�p�4H���YU���������)��J�Ww	���T�Ed~��>]4�ڞ��l�����NwDz݂��q��g�~����)^IK�w�Q��s��S��>�f&݉� dqٞ
�^G��̯5,Ej����������g�E"M�([�Y� [.i7CxV	*�~��H�`��Y;�_�6�����:(� \�^�Ƅ"7��ؠZ�Ê���dU�7���e[��;�"�B��.��\c\�F^gf%@��ݛ��]f�^Ki6�1o��0��a[��[T���N�f�7���k��fK��nq���OjBGj����s�lr�4N�6���Map�q	���[����t�r��>�Pf>�툡?�l�S�캻9�a�@
��F�W�Q��%طxώU%�����r����{����LU����P�w��msАƭ�2�S�6)*N��&��xo���*դ���^\�!0
(�d@��
?���b}		g��q?�y5"�}����H�6i9��+W(�3%�h���Da�K*�ZX�\�����s�Մ�[���-�f��M�,]�[�R��h� �O���8#3)�U"ʘ���G�d�i�#�{nr��p`��G��Ј����H"A�՟��������L�# Z<���V�{�Ar���������#x,�{b��H�'#��+���K�4I�ƨ�i���LӋM�Oݾ��:k��)�fp�0�(�`�X�z������O'Y�^S�u}r/;��8>e��zf8U�(�T�a	��"�� �p�'���^�n(��z�����kt�V{g���(P_)����)K%�Н�T�����O̺��OEn'�����ѫ�Un�}�����6�N��߼h�o�Y�Ev���N"�^Y$�]x08�ѷ�}Z��|M����������\)��+��]^F�5�U^ċ%�:�'��,C!���A\�K�q�d��Q�ai���7��2?�LE�%+�vdE���{�����+�<�2?O�/��w��
@p�e{��	2S�9�)�)��X��}",���H6�p�� l�'}"�pnE&� �~v��Ǿ����~1�Q�	\f����C�S�����!�e�7<'�t�K��s4ō��/�� ����
��ݷ�r���0F�A�m12'��H:""�H�J�.
HIb��+j�E����0;�ZNH����PZ�3𴇾��Ip���Y�s�%C1L��81g��5�*�C�>����	Y��+1��0<����Ҷ:8��\��jQl�}����9�h^��6��t�F�olX��%��͆6/r��t��k�)W(m/h?4ԋOhTzhm���G�Ѽ�a:kp�L�S `���u|p�ȬU��"�v ��Y������Uz_ 	"x�j��2SBE�����Ij���>��4�Yտ�2�?�hm}�e�{�b	czV��c��j]��THO@T�P�
5�
A*�����qhdL�xM�}�Ɗ�]��2+g�(�zh�������U��E�t��'��
Q')n��0�L�hw�����"����8#T⾋�)kG�}����H%��3 /�f?�KY����&p���ؘ� ��}@���y����&�-l��-���K���Fs{O��o�~��5^˥3r�I(���g��'I��9Y��c���I�tb���~�����5�#��hU�'���?2޵���Y��n�y�%��s<�@�
7��b����(R�9����`�~>�/ت=!�m�VA�w��dYd�,�����������G�%���г�ĳ'�r��Ȭ�~ ${���Ɠ����2���=h� -E����1a�P�������k� _���Ga�$��V�ed��#����p�ۯ��)a��z�l��2�L;�;2���Cs��d��f�prl}	O���nZy1�W��2¶���hyYo��g���.��I�)�L3]�_B#���==u�����A����E҄��9�&��:��u1!��,1NWGu�����p��Z*е��W��h���1�F�F�ݹe=py��6q��1{&��+p�*Ty'�4`�YڋZ1'k���<P��tq#M�5���2�'�{冊e0Y��̴�g_6h�1Go�V�ݰ��B�����ǔ�,�-\�
��s .��,���q󰬲��`��PP?��qq�^��C�D�C�(��?L��6�Z@�*�;ّcx�4�R�5W���`�H���}���a��������^Q��Z�X��X|ְI����_:W2E��=��{��F�'����7����E����7��^/�Y�Q�v'�t�6��Nt�����R_4����r7RXwZ�K�({OXw;��z{ԮП���<Qsr��CxЀ����"t��s0�n�@\tkZ�t�.\�8vIB���c��
��e_Ja-CV24�,�0p�0��Ԏ X4��g��������D?��y�le��\��Sܕ�WYĿ`�b�>��0(g6�~���J`_.�8��eO���W��V3�9`���{�mY��^�Ɯp�|�?������1e�|�LX�����|P7��c�f�N}E_2Cx/���!��;GS�H�AZ�	�����`���XC#
�C��l�C���e(T~�B�.���[�U��&)�Z�0��>��<j4��GO��bv�1��˻�!�9<��9��/J>�؝ҮL�3,5U&j,�;���/'�g�7���*~�"��g��4�I�E�-�c7�[����t�g�,%<3z0�ڔZ��\Y\h��_��*L��I�@�#)�ڀw��z�C��������J/����E�=K�b��Wx�h�ĢRS�������i�^�0[�5ˋ�E��־��S��gp�*7]\)I�꿜�+@°,�6�/�@����R�$���m2�:�%�Y�w	�%�ru(�ƝK��"�sr�<���Ϥ�xj�����}_�W$��-����ũ��A�,봪�Z��%������N	d�{<��dtV��6%��I��"�.�F�ׯ��l��t����X���mmbv����sm!�!`�E/�uP��}�0��{:�`�����TH����'�כF��Y_��H�'��}������s�Z�1; WеY��R)�6ɛ���SFP$��~�vt���`�$@�=��<�Ҏﯜ�Z�c-?eY�!�Ġ��hǝ�q�;��*�fA)�\8�^�CKnKz`~o��z	���]��^�0m?hg�b���0y|ޢ� �@,]���Xw�a����@�g�+�;�>S��]\ti��L�l)�*v�]M` �m��G7���E��ĽP�8 �:�Rl��/=�ۙXN;������p�%
o7i����[s�hf�+�L�ci�/�4
�>m�Z�3�SV(�/j贮���V���c��G�"��X17�?�6���¶���!`PK�� ���|��R�N�Ǔ�''���� ��a��j�ރzz�>9O��l�h2ݰ�o�������O@�d�^��$	�$�r�����D��.G)��me8⾴,��n�%��g��߶�;���g�aL�g5�ip\����)�u����Oh��k��/��d���P�����[�3����R���m����	�oE����X��+�k��j���2/=����P����G���oH'~f�J�qDQ����H��T�^"�Ŀj�Ք�(��^2�����?;��2��w�'t�����ȶ����I=�����,��6�0�����������i�q0���v�i��� �u/X�2�TI�|B.����Ĉz��1���Yiq�S<c�,F޶��m�2���
Џ�P���!$��s��Ϻ������U�6^Qck�t��[h����j�2���QfR.@������u��2|J98�7/�:+��c��x��*�*�����]�%36#���2Oۆd����>���윘��;c�FRB��ߧ*�|��H�@s�0 ��,��n�PE�����K�h�;�e��6��щa=����|��=��bt #���(��oz�	c�� [�7gHo��Qﻸ�KI���K�PQx�9�{7�����<���S�b,�"�#j���X��q��77q[�J�ܟ�����@:���b
g�5�@ّF�%���t8���§�"�9r��w���ء=�Ř��s�/���˚��l/���o�j�������t�.V��4|�}�mh�Թe���c�� ��>���~nJ��y?���o �iJ3��1Ӟ*�7��c��v�7^c���?�7�Jx��'�(f�"��~2����NA�$��N�j��WP�-�!A7��;]���Btl<�U+��gu���5��1��]5�q��i�5�{�����3�����ilM+"�nW`S@t�����{�<"<���+�����iOג[A&��W霊��$J
]��Z�Ze7+{9K��"��8���o�/-�B���_6�'���9��"�f+:]�&�NW�6��W����s{5��Ew��_����a���k�Ď��C=+�N�T��G־�S������:"������]�:�P�������ܱL*���F��NEt�����u:`��)�/��S�4��F��YϾ���>�d�6�g�Q�����88_ٺ犘�>����h�m~��&l��;��f*��$�yX��?ǵ�t��2�[�~�'Kc͌}��n��"���ꂣjb-l��k���k�4�1���f,3���rUx��m>��'!�2T�F��A>V
�::��ۀ?���fIk@(G���V�#��v��H��R�� �G���ŋ=|F>V�Vjs�������0��#�;��]�й�G�IwՆ��z-Z��r������7�_���:�*��N��G����q�u�8�l�\>V9���Q�pZ�v'Ļ�
Pz���f!5&Xf�~m��H���}�W�㲲>� ���^&fe��I��y��+���,�ÍF����>�KVPÐ��mFf�i��pgW�}�����[cQ(���
�h-
�Kb���s��^��n��^�d2��Se��%�Y�KFCdl����:��K#vO�B�ː�u� �#8�{����S�*��׆�i�R7�A�F
i�����*�`ǽ�{À3��Tp#���-�?3Q-eaЃ�t�%~�6�a���"Wµ���(gO��U�����q?��hHx�6~+�o�%��C�9_�7HPj�/N����S&�QM�y�f�)����AT
�� [|R���六���4`r������E�v$DNM��?xH�.����Ƭ�}���^��y��xx��0������*oc�fƴ�d:����ab��)[�gO�\�<nd��el�v�N���!���G�)�Y�n�{�67���.�u%�������O�M5l�x�V|SA\K�wZW�2�.`m�WJ�����>�w�[���nr
�ۯ�L����~b@24���O�P]�,S�_Oh�ʙ_���8hb����b+Z�s�lו�>�<�ْ3�.��M�X�6��]G����
�3�M�j�7�[��ְ_���?�q�7I�a���ӳr����\M����� Y��_�o�	��U���Zg1�'8)�P�+#%��Oh�C'��-�Nۘlȩa���eei���1֌nOn3G*͒L6K ������E�T�z�g���x�F@����E
�(y��S� 1u�~���o�qrI־e����֧�b����J5[��[k��U[0���Ҳ)@�H%Z�A��[xwnD'v�i��,�+?kp���bv���RQ���uyl�m�wlku������|�vm���˛ uVb�[�q��OS�:�U;i.���j�[� q���@�no`ا��4��P��?���~��1)1I�F���	M��$Eފ�k+��C����
���g��L���o�E��5<�l���D��������������ꛫ�1�gs�dG�G�g_��`k���M�q��b��n�O�=ȼ\$���p2�%����UjH�(�� }w_�r��yF�4Ąa��p&ulк�g��%g��p'$p2鼉�դg����C5������=G2S��o��9�`�hé+��OL���g��!�y�Pj�b�~X�8M���˘�b���]�}Zv�7'��v
�M:�Qo�u��>���'�4sԔ����K������1|m�M�`~6�@�g�����C��ٷX��hH��C�&�~��C4�<MrQ�6kg�����v�U���X�$���:֝�1�e�c�5�U#���\bM�`U�
�.�e��Sv��n
vm�������v<FT�z�4}�/��v�\�r���קU�"l�����~��
}��~���R��ǜ��
��@j�#��ƞG��*���٥�&ګLo���Z/���= h�����Ԃ��9w*l��Q�)���q͙�Ƅ-8'��I�=4�@(����[��V-oūiF��V��������Pު��ti:�$�i���]:�9 �}p�
��R��F�D��	
̓jx_���]��7&����<�nd��%X[�����<�|�d��o��&~9DB�[r٤B�l�e8L�t�����������xR��l�(x/�R�m�c*NS�y�U?ι�LL�����֕`�������z2z��˻�2��s �Y���'l�'��(�$Ш��=l�e���A8�+ށS���9]��`�#��-�î�9�~��Z� ���L3�T��Ӥ?/ِ3򜃡�3����=oᬲ��]�a8HSc���ٕ���4�58̤TR�)Z�h@�C[���cQ�g�>v��v?����D�9"t�W�Usw��|�bP�D���L��?��BC �W��>��,�]�WQ:�	c2�t�������)�)��N�8h�2��@?�7�q:���2^ךG�iY������#[?}������?C�	���\�B-�؅<�U���Z��Ҧ��Gk��oYG��WwZU÷�(���|���mUTJF�B�o|<�[����r����˓����S��XK��FZ��S�j����m-4��ވOqظ?����C��Zp�}�֜�u�rw�8�/�SP���ҩ��i�(��7��F�g��ѻ�	v�����5�L�V��xg�oF}�fqb#���
����F�Ffk���V��.���
:�'�"$�* �Խ8?M,"���Y���Z�$w��v�B���z7lK�q��
I�8�(�%��USi���n�7�j�H�1�WP(k�uL�i���pV-GA�1ȸ$�[�鈒uA�0̃�i���������e�ӏ��j`�_R���m���散j����=�K�X7�~*@2%��?k�Z�'�ho�5%e�
��:�����mP�w�^�Lc+��� �v�1��$b�BC��~��G��<Շ+�����R`����� #Ϗ(����F��=ϩ��3��h����í�%O^�+y~�	��cv�� ?�� L��v��#4M����s��L:�wz1^��R�oi_�+7��{�>�Ob��G9>�2��K>�ܻ�C�����6���H��2���Ʈ��	�<�?P�"��>�U�G^A�~e`H�Y�p-U/��La�D�tRs�� &`Z ��A��=��|[�Db����3�ov�O*("Xm�X�ᙯmm��Uv_g��`��h[����Nڅ4iˉi :GBz^�Xx݈�Da|�fo��ճ+G�L�g��*��3��4�«�+4T����0v�(J��L �#. ��R���ԚE?zX"1�e[����%c���N{�9}�Po������3�C5�3�S��l��fL�������j��bc�26��Q�.[UJ���ĭ(�,-�Ǔ2>�z6c0z�p}'�v�RŰڻ��A}�/�6�5�H�z���=�D޵3�/��F������Xܯ��\E���>�"<[��eL�]Ʃ�M�� hh�����-f�T
�_ͅ�FȊw����37d��d������50��~��'��XX�j&�Աٞ��=4͙R�r�������"���wvJ����;�Иd�4dZQWx���C���j#���I�� +�u��%�������/��J��;�;1��N�VNL�8]�r�vw�Fdyߊ��?}_a��Y�G��$��yP��,���Q��QIn�L�]�K�#MEO��y,�d�?b	Sx4��0#��K�L��_�8�M��*I��1Lѩ�C����}����n���Y�^g2֯V��ʄ��jG��f�i�z�D	W�=*��k���4�W/��I�Z�:��M�P��|�o����ˀ��A�k���|�I�-p��;>�n��pH
�d������+ ���:��l�-C�QZ�@ap������; � F �]�T��-�1�䁰3��ն�&W��ؗ��E�Vם�hgR�;ўΆW�+��z˳m�tc6����E������s%�F�o��*r9S<��+��]9j�d;�;e&}��p���Ӎҵ~G�/�F�*S ���
��W��i�ѹ�A*��:���ޘ;U�zpC� �ɖ�kg�vٟ�Ҝ
���-9up��ѻ+y��Z+f4)̕�
�1��:B�E���4�iz@E�;���GI�$.��\�C��R����/?@���\��Z	S��F�ߗ�7 �.J%��@��=�lJU{|e\�i�}��_�S#)U�p��y&r�u����� ��A���G��.cΚ�6h��֡A�F��y�de�b[)s!x��`Z���;����Ly9�������>$	sl�F��4V�����|bQD�(�،/��	PΗ}3ڮi�8�@�0{��I�L WD�[]��_f�rv�"L�@�ǥ�%�zC��BPV�_��߽��j����Ӵ��l^�w���/�����H�6An��l$^�3��1.Br�c�$�'
���j�e��α�S�`h\DP��+�\�íª�)�A*��a>���؂!����x= �7�E�* ���@;|�@5,��F(7��f�Y���L���'@{��YJpёZ┺�H�P��H�D�>�C�L���J�ZO�w��FA���?�����Qj�|#�B���"��?��!���VR`b|ŤJ��'W�X�CU5��(��H�,���B��,����㫒yM�_%���M��4%�jŶHO�����8�m~8�>�my�%�R�ۓ�����0&�@��V£qW��@��|�~dE^���H�V$���g�m��c/��n��'j���C���`����Y�C���a�Ƿ.$��n�Y�TJך��KC�����m��?[���C}��Q��7R)02��쪸"J�Jh�~����������"U�G)"��*�oaʔ�'�=����$�Dg|���_#��O�2T���ީ9��Y�1Ϥ���Ƴ�b�XR���3S���f_ล&J��n`H\�X�Q�0e����������s��R�����q�a6����(�t��Nc����C/^��Γ��p�P�;����Q u��1Q�G��P$#�0�����䳷D6G^N�D?B]�^t0+��=�?�,�!�������EHW�>[\<�!��_kx�H�eQ��4�_e���Wa�ě�؆����+���,o���:ϼ�\M�}E��d�0���� ;#(�O<�g.��Z�p�4%Q�*���[Ǩt�^�0d�G�����<0��iԊ�o̮wԥ=�6W$e%���L�JrO/T5Twr뢉�u� �q��UӾ�=�UR�@���.7ݠ2��ᘂ5��v�Zڍ�����yy�DG�9��奟�7�t��ȃ�X�7�VӤƂ��aM�T{\�U�	�_
b٦1�̢�����~y��P�����*��#�Cm����ph�H|�
L�j�h��4�