-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
p6s8KYO8CUttdvUk0H3l2GHJALfONKrr0z3gH3fbDNJ0sfe+ojmeElLhCcNNAyzW0mrTyNfrQGfU
uRsQxRPffllDPyrE35qIKZvWUk2EJQov5Rt+9sP2w/+gv3dlypBhANVJUwC/5qhForOIJRJHcOXP
x428fc9kRpq7W7qprixF+K6tipeMtSRYWRT7Ha1hZbAs7pI6DrBxv40BSuNvO+urM/VgAKaw6ieA
+855I5u2es/ZUzIVa85yrzQEnVj/ThLDDZ7dhuMXVt4a+jDzx+jH+Bq/z8tKCZIG3AXmdWwQNTAl
t+b9v7wg3IGDbtav8PQuh5A8pRShHKnt7Ab9OA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 24080)
`protect data_block
ila3ZmsN9C7lF5HVpfdFgNmbigxNI/L0w58xUmxOS+gxgt8/n4m9c8CphUr9J3eyKoRyQzz0v+M3
mPJeOwjiajyfhHte+DXinSxHGU0Gge9DE/5KLqxmER8mRyuizHrSG0g1chM9h16co1IMfX1DBXVi
1IIuhDgzduWpsOA6mJEwhYJuOai2G+QVKw5xhF4r3HFPfCWb2RBHeIPsd8lqlH25SniUjs7BYDhd
scKz8h0JJq/6xiS2LvOWuOFUVkKCmbZesUDVeCzowIer57MPQcPy/7kth0Ahu/ISEA7qaggvgOue
0WvHUuhrWBdQHP8xjBQJHtg2qN64s6+BBAmU2WXcEflWJsO1GwHZ4mhQBRfwPDdF2uzJZQL/rqKs
C5nvwA/7bFVezm7fdq98oVT8ekksnZDTIqEKse+vaaU/Sf4nal7lc3SHnp/8r9b8o4H9EPom2N0o
8/ANYcW6zZ/XUWxAtMdXrsku5HgVJ3UnZ0lVEyiUJqeg81uemukaXKh/9/M4+OS83TEec+Z8FMrW
9ku9pQBMT34glK0IZ3nM0NVz6L8sWgmETyG8UtkcYWMbcjHIoT9rwiVjMa8W4mkyPg5DBke5MZ6+
Wu0Gmv+fEKZ3s649Ia5jkTrhh3K8qmbqAzA3avrT9h3scjcWG3yduyXYrUowkmGAZz9070S4+G4l
jYtmSTf8uEsNVQLiJIvjhfz9uK9Ew/ZTXIK+aUWrXSFdH22rJeesISFR4GZbq3slrbOxYrWnrE1Y
0HtaNEWV4Wu/v/KefYPKxJmiuWiJJ59WG3j3wUR5w2ySTCh8JjHrH9bI46hLAZtS8vXcFSKtMTvH
fvUNW57UzoFZ1aeG4Ab/TpEPVCpX7XHVEeFPyD1GA3pU+08gbd0uOQNN5NiuYkYOd46K0wIs0859
B/WwhAJW+HahJymHcJOdua0mLTJAMDZJ07QSYFO06xyDkNBleF7zIy+arUKqpAquvU/ltKpemA6+
MahaDZj2puA9rpFZ6B3MKaRZ4ZnnsM9MgRXrfsvmqmSAzPu6BXKKZ8yi50maSrSTVQxXBAZ6AsEI
axKjAAcJLaooKKc1nAA474w0hDJnC6R6D1jR/MiOvbE5QybBzQmFR+ZalnJDaSlauVy5qSY8QFj6
cfvg1VRyrdC7uVeU1l0ekFkOGXjnvxZ1TGKZNlhjtagkaOeidLiQpGY1/vZ2w8HratWz9D3n7l9y
OlwA87z7Up05mtwozYeXQRIiYScqBjaD27Cxxjp6mdwgP+DOnHFnUodMOs7+tMtDWOX2Os57idwh
CqGeVOlmG8r7TvOrAYU0fBYP7uxYyNrMcV3qtygfqj0Ru7XJxR5ZxDDR9BJTRhHpV76Z5qoXiVhY
dimNMi0TXLYe9T9qzm6ZIbgzdIjZDyuO6jcqt3u5hkIrfNqR2JzV6HlTWKFMvU62bnA6gjdEugPH
1meID48AptEMldp6rydLpOVQJqTjGOsJhwM80Au9/5nTBekaOZNIBh4kAnqj6R54OHVXz+zKheOe
w9sKohh4ds/lvpFWVqchpjZChO8qBh5sMMwVXQebquLWapM0X/wkEXcfeF2XT94Gpxe8rVgEmnKk
1+lx72BIEe/b8fwkWDq6Q1Q+QuFMQhWEQwdefR1Wo/LhDuF3hskoY/V/grUyaYA4nUQj2EY0wpTX
ec2jpFXWGuvIHLNH0sJtDjJo5ZYQZOSSgW6Ah0x32YKzRO56NIxcVwUEfOp45UxOaMGO6n5r/Uoz
z+RgudMf6XZa4KZlultSU7mOVIJRr3Wz5zy9Nv+uVjoLEduTBXuDqBueqC/hPbctkCh+LsWZw3Qd
q2N624dwMvex98edfqHXgcwB91tMcSJ2kK8koX6IAv7XQnY30Qe2mbcBofhbvdNwlHkeJ6HFIE9Q
lWraKLK3iXXXex7iXRnSbvgc8dot6u53WrD+VBYfiGSYRdZwsY0TyOBxIjPQeeULDAHSDDixp5qp
A3pxUeDt1xNqn/YLOxqCrVk4ZC23CzlAcvsZSWLcXKMsHnZlpp2qINIZHdPQND594g9LzLByS98c
Vc4t5bRg/NfiaLRLSep6m5GE0+mn8F7guc4qLyAtaJAQKfNx1w8g6GPaWhzBDmcPb/El72X10qg5
BOZTdBSVPhYqs5cQIhE/iXPUWMab4uiCMXz8XRitLGwCZ/78Os3EyK4pr1I6ygRnmwdmubmA7OdQ
BPCwPA4BR+hQbyJP7B6eIF5xAV80r403PRaxjLmj85Dneh9SWNLAKcg91ceChjbOKBFCCoRZR9yP
CeuAmceRFWHdXw3AyOuRJ40Lbilq4FFUj4qEFbYHgUt3k3PHEBtGBN1xUJmQWjQqY/9s9TvfIwbl
twPcna8dnRQPQ9fsDCQmVxiJkSqIK7aaFr9+tMzkMm3+S5mDpGy8UPMnq8A/D2v8XGvQC+X5Dlx8
IuoaWB4YChMUIlEFRxg4OchKYKoNtNth6Zig6iSQxPoPgGk9b2LM+/y89kycDWVFgRk3WiCRmosk
a2zBbpFEHYRsqOaJ5FkBYkrofOrEllgoP46fTevaonVhDB1wdF2oUS+ZV3HkgMX+PFToay1MdS/m
Okl7Zvz7/I0VRLHrcPmjm47hjYmj0EZvnM4etbOX9oekh5aEFeCRY7/sOjHnzpNIwZ/FISrPB+Mb
jS6zhyljUNweSrNbC1vtUjl3THEHRdN9tSOYRLEU2l8LNfJi7+pAuEyzBJFBhQvNkRmPzoAuUY/7
4zOzHUeZKoqiVZfBnaC0YL6+UR/OaoWxtp1BsWXRPgjxqBcKQZhPkniRy9+ndNDZkgspXPA4aK/o
vta7souXxQhUMjr+XQ84kKvqn+uUNYXT6yDiXX3zejAWNb66oqg7G23m9AEVAr6pWelyOc1VsMxI
+gnzzK4VWPwxSnIkcl4C/HrKTXaM1opfohM/zXm/dBTWVwIPUi7J0f8k708bnDxtzRsdtgBz2Nru
mFRNsosXyXFasmT+yuAhTWQH+IVHVJvctzfaAvR66VCh2kXh7/ylgA9IJ4VlxB1UultedGROpMfV
wUZ8LRe7jUXshEvXWjaN6t8RUwUEu20oYg3FiA4qAvV9QupnYn87eW3b6awyRPxLcL0gFDVQ86gu
UKjYxf7dWmutM2FbMgEmSrtC4nxcz2TAZH6GozEupUIeFA4Ltxp9uooYySlSs+du+4koqpKLQwMV
ObzTKoB+du/3Uz4MVDEEcJPQclN4xtDxc+6KkfkqjLOJMk86Harc/JQM0JB5qN9zO+T8DZlnZw/h
MDgcN0K+OI42ULinvwhNhh6n2axkB8QO4+okdKcy0ZrldJbNKktdI820O7zMA8QZcmSCFCzw+R1e
hwHB/NALxOEHsz3hs1iwvlcPOKn7Zpw2PD8D8zKbN8bchiYhWFo5FPfs/V73Hlk9xUrf0F0HYDix
Pwt95ZVzYMJ9SjxIX9xXUjcywuCvloggDB/MTPye0ZkzUP2c5a5XTrFcAIHNr9CX3DAZ/drAvHgu
Aof1a2X81uolH/YolYygdMI6F5U+wyfgnzSePn0nLF9HZYdMrCqr22/oj/EzXvRo8P0kEfuOPSfU
vzU4fX5kFilJ52U+M7pH/4tAzvIk5uHnmAFtBA7F6X0BOv+C6PxG1qu3gzVmgY1TmImpWIUb1yLE
IB3OsCSsGFVFfVEauayTSIuy3nABBpedGG26z5YU/jTCr5cW0SycC1oWsoPl2PYUS0duIbRanQLH
9oqn2F+U0e7/udStiHyTWk1obL52r051EPB5nUnnJXAnxFqLNvV6Qgw2eyUCOafIPW5NlQXxE/sU
b7ZuJAXimvwA0UvdYjA6PBOROo1P1GbAZBUCfjmt/WIhYifAmhlP6On5/vW+FtZK9ydGcUX+n6YA
3ZaLWWkcWB2cg8/JZ0EOLfDmVkqfI5Z97Vi8GcZcrDb4bN97LgkIvSQ9NpEbfNxmX8VQ3ueDIWZM
AferdZTYbXiuM/lOg36M1WuCx/VR+OPfjJgdzhOuFzwLTa4qF5aBc/WpnEMnc3lGlxb0JfXT/J4V
RerLyRIFBh/LE6yj307Gevor+MBHwxH9MhJ9LrxGycwpQvYzzTl1uITyc7iFiKtBzOk4nx+/JIBb
Pc09f4+L4fKP0mWrr7XHP7EJlvuDumRV1cYx7i0aBIf6ojdWmHuGAL+joFJEK8ueHRG6ISJp9dkz
pKZ7iz+eaLWehPY58DVMHc/VJW74JWGn3wHihS0KHOHMP+vfYCx8N299a6yurTHJFOWuKCcewbdC
HmlPnCV4d35cHcT3gpnRDuA0VKa+0KAjmkw8P72JtYV1FD2hay61mM0sPPsyZNwpYxjgyyjuH6sG
c1vSaR8nuD2ESCFs3rFUSmtOTtiU/adwCr7goVHjmrK2e9lxEpOvC2VzJSD31vft9KTEp1t8WQVg
AL+T9Op8ieg1mmm2HAh7Uhr1zlXPYBb6iCvrEGBOKkA9e1bcCiT8E70/8UTgQkDmn7WnPUbpBrJY
XU3BD2HFEUAAwa6gPzthytXmxITQU41jmeY4j6HO+NqB7ds7YT4xmJARalz5rwQ9QRH3zRREJ9QG
f6IHY2K7oXeHIIX6lcSbD/iGovQtD0YyoAMKlg3OwBzPF4KezxqKUKPT/ws7IN/fNjxYKh61P6ZW
gmSpagtj8WFE+GnAQOlNRBTl3UB1VvNJNz3jGBpZA7nyFHvEzLMT9WYWCvmad8RyhULrX4OdevJD
ejSpr4asE33LxDAxGqpYcjdHBrGi9JisN+c46GRhERGD7L5MiEWwq+fEdRDf3coxrQ/Cxg2akrlG
GDBk11DrhWZ6JgRokl68skTX1rVRg8lmVwC1fwc2s5ymK/seLDGJmVGeNZBQITjgK9V5Xtlhw5nf
rCW02CW/sGZKc6YTXDMfKmP/Pz4rlC4ddnjVRZqlb/p1mP8/JKYXzL7jQ1+//9U7RF+oGJcurDJM
5ssfsWn5E8bCqCkDrrCGINqiXcUi37l2tUFhsXqSVBKQvdQtfWckhKiF01C+8mAetSW5o9SgsMT3
uNneNpRcYFOehiVQG9H+kH2CDjonUFi6V2WZvbw0rFq0FVlh5QOp46YuFR3ziYA42Y/nVGJACG+Z
ULUjhSzWqJNTDdSmt/eOFKWvkxFYmeAmbYxWXzDfMYBOn9LCeal9H1jP/8w05ZJ3ecIcSR8ODj56
Gp7noqsJ02ivITWulpNr1cc533uSvTgKWL6a4MrUOf43QgbtFLBnceHhBAB+E9INurA/JDmF42gb
pA6OnVja8A/uuR/o8/RIgVUCQBD5MywH4Wijoj3fQg5HzoGhabLHz1VIAEKKKRDs+3ha7gFucCjq
zMg5/XR1zw8Vv7yXeFjwkOg8AG59Vp7unxltKlri+r91+xwOY3MCveqK8D/sCUlF8/e9Hk89JMsu
hxYWixk8ROUkBvEZ6Ns4blySZtTfGE7Myt+aiCsXtIxONYhyy1yndwajm8ZY/wteM/b5w3FIT6rR
B00qZ0fxAiGpqnWh8hUiJICMlpoB7zCkMHD3oNCbUC8hODJrQvUWAg5sFGE7IpvES02VZrmT/vDU
aUd1MWmhXmwScGGIYSXQBTujTDSZ70P8xVpT0+lScOGUMwY8zNd8rtbsZvoHOffXy2fvfY7CL6rg
oxH7NW8q9D0XerGX/IxKjtWzjS93/vU649vvUMyHLUlkQ3tOV8nb41bmAcCwfJtxpZU1fAMZd4rU
tfUGUjsJZo95DfxNXbcr/Os/uJT4szLObJIpTjMTe44iemnQNW/PWOKJw7GJj4ctexmkjm6UytNG
l+9vqs0hKDMFRERwex2HJWRp8wW3lpYVYDjGq3j2W8TDGtqc3rNupiWfAhyk/t4mv4jWQWOt1ZPm
MMTnIwYcqVKsXNUkNFf6hbl+ZwSdHzSQmRazYYKulF2GpIounT0yuKHkh9VdmgA9iqNArBB2xaWA
Uo3ntzUhGNBWgBVWy1ZH/KennB+2NyF8zOw3/PHGsM143cptk4erQ8LVRAh83qeFxUJdCo9dag5S
KWMd/toizGlX2BIl443+yMEnio3USt7Ywcbp1y4eqTuIDJgOUc7Qxp5ua+jfyPhOrS1ODNxz8qDa
rsycLo/l24dllaTouAPGqBWSQkWxd82ywfjFKsHJ3E+T9B/P1pyYnUlq25eJ5WCbYY46SSLjhBql
rjfPjoXPmNzbaSlZvMkhXCeZxMRBLzGsANjjytgJ4QhRWKdr75z1pOcbc8fkT9nbucT7sWqQyjsI
gy6WSHFsvbfwmMUqgsuj29f091CPYIIz20pjY+9PL5grYGz8d5eUNYOMKU8r6xIx9XT+uWqW/mv+
OEIpS+3j30iprSKu9vZHL6F4dkzYU/QJcPX/oy/TSjNiH4j8EfNHM/QV/yPDnqr3Frois4z5xtX1
xIbbEHad6iCGalw1inuhs6uHSA7qJWwsnZ+MEORH1x2RyMOORtK3+jnHnXDdDsgh36RR4jC5orw5
8Nc4OS+GG5pymwKxPG4oq7Yv9M5r7MJxMIwAxMTMII6V3VESjGmxUm2nN6I+e9FDGP1G3Zn8ssL8
YPj9G/Wb4V/iM4bZFdbFo28mxKCA9mn2cwrwBZB9N9NXmGe6nhbhKlcIT9uDpqMvUxidv11S6Gm7
f+1lMyS93TBUiKyVzgvx6kVBHkRHIkeBo0SffxBK6W2+oTqObwKwN214Wabety58vF7Ux4jtHX69
cOKZsjBxWKzZkagtq94SPokck32HqAL6xtmEaJqTdWEPx/VgAExP/foxNylKa2AqtkYK9ZK8zkMP
/6KcXkJ8tLsVeX1AsmUXlqyiaHzDMu7AlEGms2baZxskLOT/ulUxg+wONG0e0YxWzEoyVlKfozlx
eMHiux/krMAAIfteveftmmAhh/6QxDkXZDLVg6N+FC2PuSXNsrhDfdDGDjhffABCNyc75rVc5mlZ
YXGN1SJE5mqCnvTvaN9WDBY98o1x2c5OqL/fOcWZiC9Vfb7A7GQkVUHr4YHwXEvsOE1EfxW2dxcP
oFVzBOXc+f3MIP8oL6nMyezLE0j6OZioYuUP/wgD3Yu+rufXf3Mec9l3+LdmGlOLjE2DZ6SgM+6A
rumPaML8zJ40j2iLzEfjZxRYj6HTubbeU2ca7cMC5uOuOO3hHgGRwplvFuhp2V7DuU53tcClc/gt
oVXdpcQQDbId8pksuClHWBhrg8t4EsRAaUXGT+k9a2BrKmOiafQ1gCYfqbTE8hVTL9mu0+VQZJaO
2k+tdABUydpd5XJsyH1lbYzhTzCJVc32yIjejnXW60QkMQmRM1drmLJ5NvPqjNBeKy9xNKPkP6ro
NQMy6BgXRJcPEc1dzFU4l42MsxY/vjDv5zTjunMnmulFvjEFAKfHlQbszbejdsSpkIJKpEa+LKbP
5pXJC+SKP93khP9UA0PRklKSwLDehT9k9nvozsiZvtAYGrXxPCQU4lAlaWj9PDCiZ2gqQyBTOWDV
eJtwbUvTqtj2ncs6p6n2R+zNei010qY88Ge2cGxpF7oHjVEg0GAVLD7ODLGs3G1JvhNZbAay+nPW
7SRNkN5dtY110OY4bDUNaikzCVFdzCEy6nUt9M62g6mOhzOPK23UHwZlCcx8v2dhs3n/DJBkNE7O
QB2jJAM8DC4NRO9u0pUW7tx28Gkmg7W0XICbQMCoCd0XbRFS0Kr8bvlYtOZysMD6cGSmvxxQ0VzT
F2q9WubsLeC6N86cw3tD07b7kXcprhOLg89NfcgNjirm6NUNO4d44/5lmOGFR8is07sreHEbzdRr
p/HqjQhltzQW83sRxoDYpHmcX5LtkUGWUvX8Y5GBNMepE23BxhHf7N+tCBC824ByXoz8RuIGeGlM
pi5IVf5wpgtGA+ZLGKanHKOB9UH0ZNW6Qvr4IIJQGwe+9+y9lGNmUFev3l6R8qsDVDttPPbzdZRY
2UXjDBHQByP+J2Z/Phvl9j2Y6EMmo7LDPICFhq85mng0NISgusOVi8zOmMmYwvpg/af+NVL12XBO
AHyl1yLpaUYnWLHN4C5gYQfd0xXgMRiCGdCNQ1ed/8MO1WRIxb6te7geJvx05kZZgKm0PY00M5mM
aCOBEvMzY0Fkn6/C8QGFEImirGCNg2mhDpn0z7ontL43jdPS6YK2Qyr3T4KK3CswE7EqK9UhsZHx
eHRJ5p0v8d7Aw1/saCGjYe5C36oyk5jnwcYzUAxVaykV5ABOuJQUtmNq4dZNyxfc+j775yt7nbOE
ap1z0B7IjuDWHftoxUG5PPiArqoaOfGqyjoOBCqklLcumSn6y4yeTKQSDc0CAJFjCZVJAI4gOK6p
5IHp40VIwQZ9FKKURbgDg9QLz1Tsu4x5Te/fsMF59Hbea6S6LfoSJXbEwA371F8iuaZZnWG0Ea7W
9kClf2iaPRi+txqjyH6vXPKsobBpmDOJrvAfYrd2saKhceeqsMdX71B/fWD27YkIWjxXgifCUh3E
rzpH0EZ9ojJQXSplHYUCkKDHL95iO0jEkfzO+EDXEsQDWbO1AcmaRwMeOwENZDKN6r1v8EVf/RI2
9Y/YOZ77Sg1ZNHb75VOr9FXjxBceKcEl68PRF0wSTMvs6Wq5rCB4scGNn7CVrgJTFnUtALPLExYl
KFZLYnLtjIa/SbExJ9nwukvNP04kJB4kV2VJ9zHqHXLc2Hy2vnNF/CBlOJ8J4URGquipOg+W7fkI
QWnOfXKN271VDJuvwbUOT9zYfBbpXvF9yjA1K/3TwOlYA8zMj9anwpGzS5ezl1RcjFqAVXBWRaWR
wE/N+PrnBBd5Xyl1o1Icf7WJ+fp8kL5OerhaTRp7/CavfHycH8dkn/VVRZ08bIzs5ZMZIu438Sww
7cHSWDuuRhDDrFp/Zdlwnk5mcLtOQplyiof/m2tVBJoWPIbfIzT63swsv+Jv2WSY9aMxDxFTJwyJ
jCpYnhVAoiz4rLyceV+tgk4Zi8FZTKY/EvR7KS17zvh+dw983r8Q3R4j7sqHZ6kKq94fZPUeDDL6
AzDvxQz3i8Ln5Xg7SE+imux76aaJO2o3Z5IsjAP3ZdZE240L6TZ8YBmTWWUn6wKhVsNHWIvui8UX
jkAucpcWwbT93OjGs8MWNyvheB29SHsWn8Yb6cgDP0tDK8fi+Mmc3XTwdcghIyTf0gjIyhVbMdbC
Ft7PJlgH00ezKzJFoTFUdnthEVOArWkxaVXnCwJ50yUVQ5cXQTEKgaLmFa0LMPOiSvbh4YJZwLEo
FD2NzL4ed15jOL88I5Gf/IJfje3i0r4STAFOoTNGRRnjpiuORYMzVSe2xkw0nw6ZX65Mxbfmit53
wiPzzfdqpnPKzrn7kTYVfxMx3dHVhREoAR9Z3UEqazMn5447xmPo6W5pJHU+IYnnWVfpgwnArGpz
Q8McEAEIqOXjFQaAddJekxZKtLG4Xxi7BBDJgmnpZAVjYY3wA+fYssmX4VnwOugROkwzda8Ybltw
V6k3i8USUCGM+TecjJR6/lQX4Vv73sUo8ZOBAtBFB+umH3OBITh9lwUjY8e06aqR7DbpIfbUFtzy
91l7TJnI0xp9uf/QVNIztuiEcb0WVKpDEYCYTkIiS4uLlo7XL+3tcgvQZUG9Nkd1slOSANJE2j/i
f/iv5QVJ8glTDjUdyQTmIZxnS0zKsxDgy1zurkoM7wZ0Sw6m50Cut1Ud/0SZi/gPCLTYa0DW9CNO
0Dj0l8P2BaIR5lwGKy8b90UXzOvTGQf681Vr+TuQ54bRc5PbtKZ9qnFXLujhN67J2zHudw5u1VC8
WGd6Htc0zGksRR/Kb0MPFvL+2v1I4boh9MQJUZ4siHzwXxSvbWBm5QBd0hH4iRcpV5wYZXwirlPO
81rBLvJSwt0aftUMzAzYlMZhLNiwecCCzzBPC/rwU7t9TN1bSTUNvM+IguW4Hyq31p5MTminkrRO
UZ6x3YjRVtYeht9qduQGFXRBdKWdwpgF44lIu/gy7QTX9coeNtWZKDSp4N5rIla9sjt/8v8BbL9o
cavnDd3O/s3t/xzOLhZkmFkbkYvS9bBOrMiZOWyBzKV5PjWdrOQ2+aSdjLVVJUitjRRY5HXhcaCB
d8nIt1DLTp2s/DNoTlr4jD+MJgTKwhOTpBVer800huMU9HdCgT3b3x92B4MUw02iwGYrxjC9GpS3
L6AuR9VXRAnF+RtfsSJY4BLhSxPTB2PLTIIdaR65zT1yPrAMgBenoQ8G9Cn7vBBskJNYIQgjdLhr
/liiCKyM2fwhnurzTRMwH8bjPbLdeopvkegHbXdnYdB0/zAD2QbHjLUoKFiUWWW88BuVMs0kMssR
nJzzqiVVeYkgwVrEbG80BYGWw45BTwyhXwgMeqFe5FyuVII2M4wrgPc8cCILoX6CgA79vAz2/qfc
D77gKEyS4OXhiUGgdfI7MLFGim1h5TsdBJzyV9NC+MC9lRtz4FKTGajloU5kyPrSHOedBHwhZvOg
oGoFQUjgZUXXLaGfkDbusviHLUfP1uqNFnUFZnzb+AAxbzqXbcxAOUR20U0e+eXRu/LH2bsT8yEA
doG8tWKjUXHiZFdAHhcVajk8wUCaRu6bWPaWC/ODcmkkPvlkIktVEq9Q8daZlYDYTrw/6i/asfsk
xmorisLCJPH/rbcNcTUoSfD3fbopcFk+BkzKSEsdlYXmiiWFgYDT7AhBzJr+316EvdZbFT+XTIEi
fuS6KdJBqwRe+dP2fVrIAsrOWZmlNGXTWi/W/X4rN8UhixHgRflDuRzFQgiPl5ovfqiPi1q4c/7j
PW0eZAudeTQEZJ3j7yru5TT09wI0Jk8Qnuf2xl9d49M5NKpRFeMi93baalDniYu/TypcoB2TSnfT
qBBxppG+pA+s5Zghcu3AXNOAl7z7MfoDk/0yNoN6ZZwI0JWZ6bhI8CPdLTTmi6oFlrx5u9nApcng
7ms5JYCybOyVd38wmSAnM6lm9SJYDuSL9HDKbK9/6iWq7ZuJAcVcmJ+6c2KKlWAVVPaHNiE+wU24
ovwG2KUdimqfr4ZC4r7hWP0FHBrndnl1ljfEQjTLMSkhnEjXmvFOXmqw10q8uHx/+UG5xff6+DJs
hdJAQic4RmGFCI3/dSP2/3DH0K7i//ZdwxObEqoUbTbGQ+w1EpwVQV/c8jeCZcSNUqyxEEdfPMyb
LghbdGQxaYn5URfSn+UL6yEaWe/CgwzBuF2RNUcVpLe85sz5wo6zr6aa6A43cAPmbamq9Wc4+Q2/
gyzCVeNEsTKU06aCguxlVPR536egEcsFIbuvgMkW2Z4PAiKKwN1KbGbgslyKbKAr3zgA6ps8hOW3
Gut3UPVLvpODoDCPQZVc0tC+UBnFYgYbLYL1UW60WpY/5WXFWSubdqtJwygnMGo4qEGGT24mNd+O
edid852D0yPShL1jE878L8MAdQFtnmkf7EplNQC3gOsgZl/Vj+njcleHHIX2fQEG6owIdY9ldFvF
jZLn77NjCQ8/K2oZI/g/OSD+0oY8RCoWI/M04+VRa62MUwDqCSeE/ZKQgdY4DhpQiG6PGJWTJWq0
DbpGYya/64V6NQm6b+PslO6FzG6L66Ol8933DOBUFbRwB+XXW1lrcChxmzQZXJ51R5Saef7oD7pM
FeEUylDahNqg/iTx4YUZQgc5aLrKTjYLAMI6kzjKxwEFHooDaYRSZbXakzyBXGZJn73SjMkFr3o5
rEQSTSCSbj1nPHnly1j6JKuEf10DhgS64Uv7Ptai+0FRKob5stqAaaEep3rVZuI/aIJgKd3bd87N
t91zlYDSTmIuymII05P0EskAp+j6jqyRnrBuM1iD0/e2VknEJDlpcFo/wUGunBvaoCO5IAWsyBqg
00hdnsqwllqwmbWtWvgak3txHG/xUj6hBfIXyGYluL2kT9UddZsn084Nds0VWF5Zxpb+WWfsnBYq
RZNfjFkI7T9xV+LoCH5QRxWiPeLAIG7SFLXlLdpJCJ94AXllyEt2cowoZvVqoIB+1ZuMpOXYmU9C
gV7LF61yivbK50t5xcrwUB7gjys7rFOLUng920p5aO/zMknnC0zE/IcbydreOURwkCXOkElQyQgC
vA5jKyPleaHgNUEhwBCLGGKNAWvj4eTM+lpVWz11/wztVEGDYYepdip+W836FTKIG3gG6T3n/mq9
3yiB2n77pWDmg6f1qaMzfqUmcArZq0jsxtEeVqiiP+cjBxfRBXQimJAbnKpQnMkChIyhLaGIpVRF
teAI2Rqd4It0GIAV7gSDtvAYSkUR0O8pauawmigLub5gmNTHZWT2gHxN4Bg00xuebq5ptrdMBQOZ
fy5KZZaSQQE70IoCdryAbWFntm7eLFAqHFciS525FAx+9vtczaj238mdeid1CRanUd969cyY0UGb
AwwrnK+JslDMzLEdF2teuwVEqq4Wj70gRkSljKF7EUUfnUdmPdD0wlYmHSdsS3HbvfeK2ng3F23Y
eyjWWjRb2fcv8b0zt/8h0+hHloxHmtzb9NoKTkhWi/T4CY6+5gXY3ZGBHmiclLfP7jCQTEEKpBPV
azP2+nBQN/c1zStS7GMLmCNxLlgDOsGYhuUf9q5vlQEFOZTUqgY9/ZjUQoYTzdr9M9NPzImRWoka
Vtwg9mx3FXNQ2yK77VjHEPzqoGVuLHekYqhoqa9fKRBDZXhkAI89nXyqJF01jyJa43jSuBGEaI7/
pSFuX96RYcIw0l+H7WigL/lyHbXurqVjduEBjiWswchuwvHiFaw5ecWYneLopUnGKawxMMiMeQdN
Q1hCCcgVzXqGxPVnKtiWDW/BMRk9bRwRFJJgC8Lm+UtsBSV44AEizKLnEEbVEXR3fx71bVeEmnqw
jSAsvgWr/EUsbSZ2HmuflVax1YRLY+lD6e8Xhv7mTyrUy5Uaal2QI76sE1IUDksMG+k4NtJ/cvd4
AG6GuQHStYv5T/BQx2+mcBUrYa1zokvFGvNfGWgnBRbM9COnE+vgDoUDy/ogWsMT76ajun80ILPv
pKsQVpgpatsbZOme5YzbTn2/RACEk60BjB5Wpj11r+tcrNcnRcXoWoJw5mnxP3/bv4zYJQK1/sP3
tlzgFR3XreNMamidpRz0/eJ0dr3T9Tu6XagC3T2hvk/5oJL7dgY59NPAmzDRIEQ1GUJQDeHGyV5l
ttRmwv3CsZxzuucX286vk3RjlvCQg93j5MBHk3MjoYrXEXJ5GTG5Hbc5Xo3zfkzRMrMLIpkCA5JR
/d4rsgyCypHdzVTLISD2gh66dnfH0IlVK9yoeF5g87jFixrZRHSZl0XxcnziIAkRCrr7yqVLoQN9
MOLbL8Ra6XysnXZeArXBRIox/hGysKLS2skh334/qoJrFGaDG4STNr2Bpbhe1eVDQQBo+4vmlJgf
C1l/rIDOL08oBw985whJ3mdF0P73lILSDypF+dJvtyXhT6VdoKga3lio0IC1snqsUP7k7G8BrKRp
hXZ1wrKwLbtFIpafBnmCTMVYAGZGryfMGvcCoc70i/HVikbJQkLgYApFQ3Zkgbk6zD60X4MgXEvY
qH4Od7uOie55su9lRJvL0kuhOQuy3Aq6my4DFLF4bO2sYlO+1yzODrCLWQwdEAjkebPiMgvnt4e0
4lhVQ8bkZRQBQls2yEmdRm3+mR3zDT0zXRzH38jlM4ulOMbG/tJKIoLtUPj0NhMOPEqsv44wwLqH
ePIMil4HlAWcK34Or4+XWPSp5pIrNI08cAOCCnNlzUd2Ul9IeuNH53noReEr1gm8ZxjD0d20+iqy
RAUDNB5O6J9kkrPbBYcpDh4aEmuVXeVERHiyKDZ0brRCh+eryEjl+YtL8I+k0EGoKWH3EAFzDkyj
ZQOIfNJZ5gsZCqDJnY+Ee/wHLd2mJkan6fkNiwZ6kLzmjfSa41uVU7ZoWzG2fC0+al6RKgKOmmE/
wuOH28N+nGFlz+RQBJWmlrz5yBQfzhuXnhLCfCK41yEGzfv7GDcUVa9FuWBRURMTry/ZdK7aeXHh
qN3iaD4nkJ05rFdWKh3xV4MoiI0gDD5+TXRmU7cFlrBAjNxY4SsVI5xw3tj4bAfcF3M/tf+m/ikn
lb3s8Marl/1b6JpwmD43nin8p1VQHm4cRA3ioMJRHpR6ZXkQmMas5wKY7qWYVI1SMUqScl2sdPyz
fON5dfLzPBJ1q8iOs03UEMKoe2gSafFf8YeqyrCW1L0IpwEK/bUAbLCggjetK2fqqmEjnmRGq8hF
M72EbNOBtLwkApOXnT4lRIEJuBOh89B1TKModlJ7hgeqEapCOECDgFF/zer7QjsCYpCNiMxEYDh5
gdl6MXdpF32BJeNITV5H/7cP91hPjLzYFqZm6iChOXYg+HsiDDAkEDaaXP3gp5gDS+Ld5F2F939B
Ikq8oSsWrfl1kKTJvvncZDKBAPnyknjUN1AxahHR1TjsrzLE8cfgHpC9w3WMhElVKTY2Vj4X+8sG
qWc93iY+tUW3iRc2LQPONbsYcR0UlCW5nm/fUPtBii9PsrF6n1iZQ4JVP7ghC1nAM3+xf45+bYYL
i3q8bdeW0JCHqSagiVLv01Hi+KgQChSumvFFHrKwnD9ANJMrw1Q7Aeqbaq4+rQ92XtxrBxWFe6pJ
nqs+ZjxlDMCJvbHQ55vW4uJJQXl1CnJ7ZGay5uz8Lc0d6XMypVsEOHT8xlhMwlX8u11E/EXvWrGZ
4J7VSwvdppCqHZIFPV5hCJm+Rp/ZVX1D2LuRYPERoxqu3Lzq2UR6UlgCNemrjERsBaBpRYCs0YA4
yD6Lxpg33RUjP7iWPZfAC+2HJpg5yZwtyqVfodn/VGrzdjQ4hJd883hz3tzBbMDgsV4CFdErtzIA
7QmyCpX0gn5hJLmosDdj3cOzjzESYU9RRk685YRHIJnH5Ei4ZK8KBoByOXrS9xGKEAkYR3mIGdbL
7HQunlU+1BD+CeGbOom8JgaGZwFdsAMNkBoyxk+RGc+8sgbNLKjJxI8hohWRu86ZmuavpipcTnBd
BxkUz+uh7i1zoL+LZeS2rFgqjy2/3PScgJ2WV2kb5kxK5qq51YOWCsAIb3HXKAFeOtwdBgGnzery
/pPai2OHm06gdR0EyBTsRxhgKCoIgNDTKHFJ4isg6/dReBQnHwLNBiDGMnM7rzV/tNX8BH5RLmaJ
gzuqbVKyfyFVJO056a4QM4tW+ee74cRDaVMKswvgtTqPBP7Lieng4VTcWsI4QRbnIb1o5Bv34Tbv
8RnoRA/N/Jrc9Z4ZSuE46ys1BIRQugfSBDKQROsHTpjHvC1pp18PbNJ84IpsWcoMCPzODbdgFC0/
hh8f9XOjzbeWqOmGeUhYQN2WQK8q+zMDYc/L10DHJDbhnh3eFOX3QKNvOLUfPV31FPg7wZhd7bpO
eZYGxSmOQcb+mvWzcGArxbYtGpegOTuWt3piNiXpyRAj/G0xLxzuS4B1x8FJ6EfXSTfIpZ5dORRs
bBZLR0fnt6eSrtT5hMG5Esi/ulI8AUtq7azzsNSZKKfbrzW6M7b8ge+Dx1WXuMTl70TMvq48Aw66
ayHjW8bpXnrJ64kFudrLqp4PdE0uIchA6Go7LsFRxQ+KSWiAegZNFo63zZfaDstV6nC1GGydAjJs
heXN4/UHMJFpQ8RTw5RboRjIj016VbTizJH9XY18idEFn/bmJotNWXveaf034AK7x2QeJ5JsKquv
3gDnLVw2+rm9/u8Fvl8xcEWwqXytBOfHD+Ck1QuJ5k2YiePmB7mno04W0gfVMppO21RWrMT2Bb5D
4VTlStDaaRsofxhWb1ZqAfm/4OGcRlrz38An+/D9VpOEuvdWnRlREfBc2QNYgXBxdbB1Vuf7hU2c
f1kHMD4qBETEGogzYC8BPgmfwgZb2HKJM7AW+VdthzU8bW3/pALXpMZ2BLm+4dEU9DlF/DzAOwKl
bOfyfzQm81PpeUlShKZcJrr0kWA+VsP2nZw751piwSjM8h65KIXaLODAY/rZGjSXIScE3GpOGdMV
sZj1DLwJYwdnnvnqEp/fFBsNeRPt6VqzraWPFA4KkAVyTUypu1lqQxNjqBmidkQ6ldLQzgudstWC
4RYL7+JXy+WDy90oX+5lED4lJcRAExXar6dud+SjUbxUkk10lrZNG+mTUWHkkdoUX24wY43UWnnd
kLvh/txWwyvAJO1edKfg9iMDN08EhL4GXyXgqAjoPdZPB9hm5G5cEryWlG5CiS2Dgl3K3LD8kC7i
etyBACoaddt3fYQqGLEBMJaR6/IKf8R00VgW1ZRo69ey41bMMTCJc9Tt81fHermyGA46bjs5XN6u
UTd52KL4Od482YLONyXoCAgwGbYPviwigpeThEPUZHnds2ZN+pHSVXqbVdHIPmoPLsgCxuFbrBDb
aXPxISlHS+PSmfIQxQZNr33Xwf9KbLW0ywJVIdP6Gt4SZcpjmesHjZkKJ0zCRx0vOTJNKkFxgRgP
YHQkNJ7V0lRjj5WYaXgpyDhtAdG0vf852kNIsW5lgRQzWBvnTx/SLb1xp8Eduw5+y5UzNEH/occS
RUbxGNhglAKwZVGGVvfJMaIkPP9MXsVY6CmP+4KRmCNWxMd2uLSshKvAUWgNSpIxUrQ+HDTQ86c/
BspgXWSOx52WTv3kMK47GaUUlw0ui+0S8/N0cqxUzQGmSCe8lkreW/0axxovfVo45BDlElsH1wgL
xDUpFmzurNzZVIh4v2low6b2cwRLpX5kWLM0wKYedviBDA/H/f/q5SQGGLPHMvgH4FadSIYEnAQX
G47Em0uOk3mnQQmZP5s4mbwPpREc947TzlUfbvJxDp1AA3x2iy/DYxIUE5bVyeIkNd6Pg9cxZSIg
6FS+P56BXyIYm4lva3XjekxR/UtgKeDRBqGbTVmyZKHP1wxjXRWyk5i6rYqDctIFYKKzE7dZ+q/O
yUe9S+B+mCZD/i9Uy68PrvZuSkohnxYCrxZVyDKkzsWdXOalXw6mbkkipQ2MNPuY6O5M7u87Qzfn
1+9O0e7gAJMtcJQkrGh6cliaa8Ga0+W2SKcX8FRoHA+1q+8nJFPs3WwD6SaugEwor/849eyL9d4e
1Yt9mk0UidgMwmkRl3txHjsVt19nN9UXxOZW8xYoKSpNgshh7yqIcyXaPnk74mMJ2mFwKYiHHwPh
KgSiA/RBJR1o2Z1USCymu109ZWRUSuNM+zniO8cJSOv55IwFiUKGvH2xBUi7+6ps55dJIGLsB2VF
ZaSSoPQBzOrP/1HxHcadaN8409pXEMRyERDZBJK57vJxJ4nQaJEkZ7OBLr65S6Gb4MvyV3pgVr9t
z7tMBuuJ6txyHUbNWif14sjZAeCkYqlxBQoVaeuzROSFIdYL/0QOWLfUxXevQ1UXkJHodOUmL3D9
ZYRw760N9Q3UexFYREyHRSqN46cEmRKNRaOoHthzDikW/G4WePC6kzEnB4esNblO+NrIJ5ibePXH
NjTJzC2IePN7HwLF+Cm+uPINMKTm8vmU5E6ZLIkLMUm6258OOgXDX1g/P2YXsoVEP0aPKTDf32a1
TUaGNL86mTAYa9NeTjTq142JdbtBHIruDI+CkGBh6b3bpOeUIl4AwThwUsg6kxHua0gOIrKHV0hK
krZ4IkYZXhTu8Ln9XYj15hW5QYMZhMRgJS44JFdekgd+8bMA2AIskeSYV2a4WOloD85nW+vw6kml
jWcH2/rwj6Ch3wEXVY38jMJPULDcdF1KQtl+twUZKSCzc01tKBGbR/VNGr4Yh+inqJurRbVuvwb+
aLC/rqpJowiWQSzYD+zMloRFZ8M1+whn0Xp03iT01O9zPpBoR4A7A37aYdVlKqwNq4kjdX1cCAcu
Vey45dqx73kDPS6z3vLnyywd2KhJGt3sKeYLi8Ltxq3cRrWR+sBkWay1FYdClJXrSaBJYgeZmYc3
Gzz2IwnWw5Oi8SETE5ihAMzQeGrIKWYM92Uzs4mAzvAl100/PE+DOKwvo+MC1DaYaVtZ+FSoszCP
jtC7kdRfCPJGNo4qni/6KnJ1rVTvX1gXmXCVnXmrI16buBOtPeY43+GGntcjREUKHl7jXIYtWp+I
F7jRvb68Gyuf+mFjdVY2Rnis9mHw50UCtjrF1k0+67gQHcExh/vwEsL2OpqzTMBnvbuzlMZnJXKe
ncnDwYWu384cCram8O32pgZWjxtqme/vZHL4lSKPw2pSrUQCo9QmWHavOYOOB8043u6Eh+BF5w1v
fA7GCCKrD6mhBYqFocZk2qhH4b2LyPlZ4ALklaZ8zZLZ1xzyzHmmwmreP7OuOMGVd604DNly4lbg
RO992agVJiurcoED5dx1ZCfBvGuEpESE3IxQgC0J8b4MdNViGhD16pTLI0gBmOsViO8o4L9KV+OJ
YUxuHe3Q/jlwxLXKMtFeJEc/yfgjgrvDoUadjKHt0zFb2sNvJZNu5jeR7s6A6aVHORy1tvzU8uRs
ppW/W3NUJoFlrrBbYe5WtkAaKoNfY+GVMmDnlawc998hF//8TR3ptHLFGhF9Fxl8J1z942hJgmAm
/hPRHlfCfyDFl7OrQSTEkcyK3trLWapi5QEeu3Id9g7vR9aKk3uaei9oWH8VukgrbvcejHYoCnzf
P4WDC3RduleRz37xNK7io42z/DtyF/vwK2MUqpeGCbtH1c1204gpHuhTBNs+PdqrKVAmYxzKpa/R
Yz/TdcnZYo0Iu4djdZETGS+r/8zIVa9WzWyABVUwvtgH9tE848tJFcA0+OSLKhJeQimWOZwtvreS
CcYq1WndkN3tufQkoQa/BwH54JDG1r/KdiSjG8eYn/enMxpVIKqvYeDMnsiCE63QoPzlu6ZIYilm
dmmvm56RRjacC2s1a8Xcqpaqy9qXBjGREpeCb8IKFpoWW5oBFIfRppsXKXjcT0AJjT8WvW3+ThLh
1npBubRXuqvRMjtFDUJGsNPj7rsO2VVDbU5wH3P3Wk0y2nZgj1kFA++eqg+1JHJHAltdIUunJesO
aQaH1KkqWv2zSU912rDL4R6TbeCAjPAcK4aHhlQ5rXOiZjHOQAWVdNTiM0ESJRebveYvXW5WF/RJ
seNq03YlhgGhpTluda5nIHgz9wYZK/4XPcGAcld1b17CXvggsr+Kmr/BHjP3p2afJfj3Y3UDVrjY
QXYbgFJ46SiTckz6QBOylb+f9Oqyc0bOqf2CIfedBdPIjMnFEP8XCVxmPwe4MokrVCcnHJWU8RCR
bBV+tSDS8jIHT4WwiKYZ3+XCi/l5LwRLy+z8NP6OUiaydWB8GqlgUms9irfxNNmxjiqP+wYKrqL2
3nwfZcC2ioQ5+QtAtyuVC06s0UqCkxbZODNZhRPYyWQnagVmEgvaL7Bb98PbStveZwjecGGtOPA9
e0z1qlvadtNDCGMGD6YdGs7KbiAzL4aOYZrDKLuIGej2SPvhDt83Wrkkfxcf+1fxOj08q1OIzcRa
hOc2EhhETWJOsG1kQRJqybtsUw3CuXL0GflzhGGT0zd11wCw4GQGqKyr+Pjqpl7d7mgwsFP4XXcJ
iDnItiJrQQ3jv6J/3Ya9rwPXh2pZiJYenTksuE4RdKRIW50y/d24poeBWUeg+ghdJ+j7naUbL/Cg
zPpqJxxYzgNnaVHNx46MWnlQ53CPYddSEPJoO1c3axrGkhy7XZ6tLMXUYZvdDT57wvWa8S+KFCxu
VXU61LGWRxM16yEXtj083t9OtWW7oIsUgQuWZBQfgjt3LxmQMQrd1VQEXNEzvaK41748Miyat4Mk
rdL/YK5QnO8ivVOqzhtg/LnuxJJSgonrsfzgukk8vjcUuameGklS5B40D89mqAo8bp7fNcMT3soS
lJ+T47sHxjQRTOBS4+4sjK030AjUJMsXj7NoyZ3YMB+3zQuwwdkMHrBsDYxADbflZPMFMJXwFjSi
GQii2oTQGe+hkFebREjEUtSEl+XXXjRX5mDgzcep13yG94FiuVX+7QxtZn3HSiWJTtffgJDE8wNt
7hUJnE2o/bRQzcpTwv9Qasb3VAmjopB+AniZhOIDdHIA/iXlTVPzeLEqWxf5wqfAp8JCJKBLLQ82
CoLom8Ufm0AQiwKW2823ye/Gcw9nxE1XKzPfiQs+r9J/EJMfpkm9dfl8EAf2oCZ1LWFQUNYtLhCC
8CWS3UQ2S9oW6cvMEjsLo2LQaC6r8HWW3L5TCdweLs8eAYnKLjhZd0/uI5G97djX9lk9jjDNIQhc
5tJt/osGZTManACefSC7dQAQKH7pfEZXvwYyZS0UUgHVg1LFjQ/Ijs71Ye9jZfMzCfDI5rfx3i/J
vHdpV1Qh3Ed6ZKL/6CTDmJ/AHqIyU1a9E36k0MoX3YsNePiJm+VdQlJ3FZm+D2FMXEHCQ4FahwHa
o7BGXRv6hB8X744ilwQxocty7DSjZE3FuVhp2iTKJ/8d+H5GHU/YS3AiHbDQ6CMAZmbn/1NUjUNl
QHrpm3HHurO4zviOURi9NwBc/f2Gm1cklUquC/mz5mVHDhJvkRGulvexl3UaPHXJxSOxDvQzplIp
GuSh7KRGjzQcc4MzCns7DDtdGS3/Bd7c0O92cL/ISDptnhMtlYV2ZO+qLJJlNga90w/MK0UE/0QT
nmpsexefyh1A+HRcD4edy8OJnu5sy9PPHg2IWQALgxlC3mg216mGqbAf8ezuziX8OFzwzBFdKE4x
3YhNuDfNOqGz+Rj9Rgo9F8u5j1ugyM11im7SkSAisymCaN1AfPTsznI+5V1Mqxa5OWOsu16XJ7vg
Fv3q3d0bLd2nOwBToaI3hsoMGDDiFgBdV5C/0syQQmbWcwRr/zB2gu57k8195fawct0Az62f4Yhg
rGNoWNLIP7QoOUpRU/cYlar+s5mtCgWeN5mhqMCrW2ZU4ZypMaVYBem3/XRxl4TMJJk4hRSNvYD1
yE0w8t7R6llzLpqU7/ioTPlnoT+D2WpEb0vcN6RhKRY7gHN95uTN4Di3dsbxBXnvlhb/47TeNh+I
Koj7P+K8ORSbiYQDR7o9m5DBR0KSw240LecYSMDWa8C/ShqnThdUqlouZ2R9ZVgJKE2fFhHch/iq
j1gutFEsZKw3Ie68k8bm3goLq5MhwHKS7O+teqwQa/8eef85YpXqS34cv+mQUeYO5rj+1fIU3FoV
LYkf9N97UbQmjZXlTriWfGXZbp2s3CmLCjxZ4pHfM+wkLJYZA695TIE01X3LPXEVLxQYqz+nRV1g
Lo/AeKW6AdspMERkD6CfEU3lk3C99oMvubyd0d1VVGgbnbZzTH3/N1nAPHGiobQW63xi7h87/yQf
WcMl12tAwo4jbqjdjXq+GaUNsLsYA2bNSRPXJoKgUD21rST8WQILgItVKBzE0A9/9WJiEiLnc05w
PCGq/9GMVsuL9TfClg/OTjnyfEyC6RRZnhyC9AxqhBOEZEQ2Baw1fnXM/pfCHzETU7j9y7JwokTk
EC+Xwc4Guzo1DXadmKRSMUcnvRkRBJF8PUgBOo8yofjfujtjpXqeKcyA6xbrTxd4GQLAkSht/Q9k
eTmro39+bDOBEEKNFEhhj+WdjH+qryCPQ30vuntOi1lLyw4VXstbHw6FPpxxNelKQafAuxwgwOV/
Pk4eONimDDPmUS195Cz4xT0SYsMqjmiSnmVon/6LRyJPp+Nj6JYrmaqjAIzquMzy/PGYQ1VzaaOX
vqI8GWFsbRC72iCtedmuwU7IQZ5vrD2HjqOEXogDOXUyyMvYquGO0xjuW9dV6fKilclbwjSLY8zr
V04jd4L3RIoeQGUX2MNhYoWzW3NHZG8Iw+5AHj8SJzLC+7IzLRJc1H1LltSL6Q5HBaJQHRLOuUGO
FpLRMiFyTT+Fb0HX2uaoIb8pm7wsBSZ+zr4vUEwpckFoFcUieo7nONcLcXR3MSwQjBdtCL111C80
8LGJmD+H7/gHtJXs6wC2v2F7JlO+AsOelmO6ZSVdys14t1RzLd2CDA97gMKpmS+9nqtekfCGnjyN
3/X3h+96AKJY+UxUYNsSznDq1ZXmQXCOJr86IN9DpiyA3gFq/iqBsC48HSF1DPSP9vVqKP4E8BEH
FLFJH1k50AwYO73LUtiolytuyK/7N6rO1xX9vqU/zyqquuwUeuylr0sBAQszf2amhbtOQVUrMUGM
zpeElub3nrsisiVzJqt55MV7QG6UGUaQCBKbQyjP8WA4A0Li43MGYNa3nuBVEKjbdKi10uxD6bTx
CXRR4TmL24HyP4mPYf7Ac9Jfi4BTshBLV8bJT7aSm5X8s53AKXJeg9hsV4jO4tUFpoDXug+L8Q9r
Wdmu8AxzZRlSCxusipHkEMqA9tJtem0hk8mpqF8PAY8uw0VimJHDZ2dRvLnyb7jAYRxeALQqz/Zy
tK2xu+Nb+mTxFKU9cDa1n1SqFQvzTQfyB+2GyQTdRliV05fnzWavvWAchpU/veP6Ut6Xub88QVci
K5GAO4kBReoJlvl6Asn2Y1e9WaB1RSqGRHNTivJ7rKkFDarcsJVRqCi50jWUaDGIich4btkVimIZ
V4EKPPMfFa0e6zCPNN/zvgs+98D1fccfiG+iqlI4X/prAa/JDFFbGH+djKXf/TmhmOAawUoINt4I
l6AQHr7w9nhPYL9N5GzwXeHpQcIeaqoskRcQ2dkFlPD+k4JVyrUkP2uDLrajCXsyafejxtSYD1ex
LYVgxy/zMChWDSEOU117YQUinK5FNAo1Bu6pdbNF/nYH7qLAplu17heX/UctJGTB13kAGDTSCFZQ
1E/MxbHwsUpzm+fHuhDEe2PuJaK7mQaxCdcBAUQmkWkEhP6s64HcsrEBB+sSI2vM5wWWDb49EyDo
T8j/D2FFmvzrj2g+oy018lCLlCqzAo1hNJ1X5fnhufcpIhPUwaAeQ9osGPeY2bxsNt7Cagruccci
R8pX7zQuzZGPMCrfi98Dy3UwjAU9kjXF/7Wd1yUBuK27rXPnRJ3wQN8+5JfgdKlAP8nIF+fV21ET
6v8qbit6KLGKq06B6/M8D0ahr1pqaA8yLDjgKE78w3QGYxntL0tU8/9QKYr+y4eERFnVKvTjCvYD
GhTTtIut4Paj1Cf+w29vdr7aNnL4qCTLEop1eI5Cb2vIjKqw4fUcmO7N8Dobp4kHFNEVoOHPRCoO
K6yNvZ6Eu8YcLIeHzlidiU2pTbmFVsDd7gGSUYkjBszhA3GL8GiNyRP0vKrJIzZg2gBC4kpB5vr3
N0wFJCPt3pTq9lL6BwyGOCLRzhkCBgVL7Ee9W0obDGvTUm8JI2alh8hbutBGb2e22YXEq/V5nmjb
6Zj71CIydQ99+ChyzQ44c6f+ges1OxcQ8HVB6dQPG+7z3pHhn3lvbSS2hTAYBXQ2BmKw1XtfGPKk
xsxXRYtUf6ghTeujkYUbebiHd6hCoRInTcTTbamdzlAo+HNOSfqX4Th84PQgXBXOUEoCrgRFTgAn
s4PSs7aeblz06UZy47kMkc3poIv76C682/rE8tzWv2amv9VkCoKjbGMvh2KIQHoXHxMFT9Rl9Ptg
50HQPGU15fcyXGYrQPmVkh+kmnxgXKVViXyzrY4mSkLt/4kUndOzVyskukeGdTBA21ydg63dl/zd
pTNtWKp2H66BzPRdqFXPZFCyMKaIBTySjDJKl/2nuc5pfGg9LIJb91S2pt65WRM/fEWQXG+HpxLd
42Gr1QDndORdB1nmYRFd8j98gpmQJv5zJxKIZz37wmhNJXApvq0OB/ygHAGekHiJmzdH4ZZiIzVh
UvI+zUqatxVRn0rlTl6C7bPMvn0ptcT02FeEIT+r6BaUPqKF/SD+nH1KF+gLN3FzlPrSxHeB02VG
AzhFZZ8RR+pUczpFCgJ10z/uYskGzOXN9jY5VRU+iffKz5URt4GKYvZXgD+cPLl3DKnbSfrq0Cif
l2ehs75gC8+JRB68I1ak//NZEgxspsRfdbUaWYKrOYEKGZYRzUk2mXvWK3NwygFb+lYXwfatqEFH
1uVEjBMEap6mZsd3PvDKOHp390vUIk+KzBSgVqmGfzG8VyRDGUddYM0patN7p6jrOOl7S2KWtiNG
6LNJgHER8jvEKVMV2mLReBGcoeutEaw7HIMPBY1AC55IyhTACSrsvCdFg1F3stg4Fr8reOx87SAg
dD3XKiKV2P7Tx1bVu6hQvxIJnRZ2v/msrnWIyHeU2OXl1aa7TRbCbi61rES3K7s/2qEm1dc5f47N
AUwsnXDUVm4G1lUQSNBx96ubx36hqLxYc44sYffPFXWFa0CvHUL3bOTUMUmYXGDa1ZpPIlvvlfNE
dgbqP230bOlcWFYOt0N5JGp9Jt1fFa/HKtpCv1Bb2j5B3aGZQnjzHmeqrDcxuTp17ipVSvHufHfB
7lGBBZ/6fOamsrDDcTjIJ1Li1d5g9UCojm/BuG12zynKZNIypYvkVoIAOehsSsPlNjIwEPLjUjRS
hgSqb5noDe0dTd3SxO3MtTQIgyat+ERDWu/mjvBb2m+ooZ3bcKUjkj/7FCLxxjhxBkZYXr1YmaGH
MWAabypnS4/keY6jd2VKqldeieXLl2XZkQGm3WmX51vqUsmNtfeaVtdLy+G4W21s3s8EgFmy+quF
EOrgtzhZ+kxtnfpP3TvQ1IqHnVcRy91666LiHQE3L8mjhBHQSrpyIHAFh1TRI1bQ1lc6aCuQ4Fdd
Y9a17CnmI0PJi60KdcwtzeAiLXwUhkeUI7gBB9NVM2eIVBP71m5heZnk3yxcINUGXRh83aI3HDbq
dbaYX+RZgzb5pIathgs9PYMh6WjQhgRNA40EYtN45ZQYeohHPSRZkqQlvtgerxz2U1csoMjltCOO
NfPXFWJLTb1NGlIv8pMuV5gTD0rqvoNJR/9hq6sIhFVWYPHZJdRbjVLAhKkVgrDMYrfH84sD+2xF
B7piJn/u6EUDJZ8wsCMpzxYHn6PrGODTHwCakYH94kCxqf9avS9PPJh1+gL5Xbo5jSFOA+Ir7BfK
jZZChMWXggU1I05pStEb8zMzqJLfqeSQRYsYOpMhksk5Bvw7OYle/QzCyPaZL8g5UDJ8NIrTzbdM
O0oM63Z7Jbsa6CpxOnV30yQYY9uDBODBvDwyUy1wMFv/bxqNXgXEYDZiawWjpFOMckSP/Qwn5lwx
aMl0tiNZgADyY/lQbV1fbimSJhrFNTdn8Zl6oQa5uFCPJz8hA0q/G9IHUqic2zip+dLYpExS65gs
QpwcLHhG1H9oYNCzaWE0aQc/pp5o9OpEZ4rDnM/hvqpgqsQ3M4IVRV//LNWRY5sp5Scf0USYWYKj
NQwjXL2QFEBAsphrDyXRCcMWfSwbsgQCPn4GNktH5pi0+pUSLftc8LAyKpxKVXTmrnTtt+PK4GV+
6moKCKWsZ/XM7KR1/kbDTtWMtAQHcZIpu0PVuykB3ki+AjWBREUnDP/4y/XC1V5wwxoz1uK+zwUO
jiOPoQdDQwafO/gvhVq069iDm9/U0+56gWOuewkzGF3Klzzbb9192bBesNmzS8H05df+mHzEbJsC
YWGWc2Ogm8Stys3EqC5odM+xnfiu10wCoo4D10KgGZaJKLt59afRZmu5wyVDsa9Pvn9yAQ9FV2+a
R+/RdsnYpFIyR/obyp2Eug4iGSAfZlwDGGFUSshi39DpKWkhKH1TxSkuDo8KpFfXNKWFrHYsgzfX
/ljNVwYj7KBm3kXfGGwqH19KNBz6AjCMj3Gwk25vRD7TcuQ4CNQbiGLXcunbzv2IoToGHhPMDlnT
vaFtGr0YiTXL1lHHrgLo05vpte0GtUvOSGZ7umvu1zv03NKVvFpoXIFUJ2gs37jYuTp7r7wMKkSy
MRsFuKJ0KKcz4ZxxhpxgjO3ds72COz0oFLl8BTdjHman/Ufp6vcMTqMd5Qxnx7AoN3PPveIAtqOY
9c5B1O6jdXBoujzI4mIbUxOiMT+UPcvaCk90ap0HBtq4qQsbop7TFj8dnWKpBX8X4cigOWpFHf2W
tS5IFbsSRdtkqhsO5WXP/lSm7FgxLi/exkQDKarvXo37o7BlBABsw6DcjIbuUoLd7j/+Ks76rzwg
EiB5GAXvzyO8Vu+GoawjAMtlwXb2QIkDC692B178DpIdwk7OcbcMjVEl56amHPiatZTRZwx5HsfQ
V92EMPaghECw8UsuM9lMqKTucCfFffJZy3EFAtixyAj/NXYisIb0v5uSxcSsSms/+iKVK9/YsJUs
kboGYonOUo9OWJZazXztb8DoBW84BaitMpMp39nT9AEW6Az6S+qANq0r4lJ7far/14KKQe7Bqz76
ouBi8P8jGhEGlMtUaYGnKdDxcKGIOATkImzDbkFG5F86rw68KOpBDgF8JwAGWneSulsGb/C/3wst
4CyHf5yH2R5W20ojSThCKStbw71ZoGPE6oUew58O8Jvb3stWSzr5R6XEQzGg7CivttX2aM0IFjDL
jLOsLl7dtsC1mQCXYADKOSvGN7eX1qTR5HnwDozs4zd5iB1TScgMyeeoHLIXYoG53vumNTbu9GLy
Tbfeum+lb7oAr9oPkY1KMhDy92Qn/9/X5QYux4Kn8HtY7yGmnr5ABqJvlImqPu/rq2o31B2KY5NC
GZ3KQEKGzx75R2J0+Y/apTC8o0SeUajPUvvainbV27ADDofoFS7Oye9jyAPNxO2LgNGX9x4wnBy/
YTJB+Ei/JogkCMuwiHWakPSdn8UzhT7bGhzEKlVTp2GNn4rnIN+2cKf0J5DHOFYLVJLpFaPaCHq2
a9zDDwA+Z5AEr+J3wRX5sJiZWVU6gioF/j9G0JqZtFKRdmUzzu6KsOesOt4JJFbaDOuNqUCF4DS4
vuiF7kvdl8khvbe8VjbufhBkRTAvFeRGsvGB82xIH6+MybylablaJ0/LJkGOvXlRSlyb8+PSDQye
caLxvL1c5H+se8ykhyApRpx4ldu5Cn05l517x+knf37WxXAz6HK/NCbFbx/08m2bXJjpX2951OkC
hXqW0IeHcbIr3+bQdDdGwYCkHkNwEm//LhLps4TUYvo/BTKx8aKU7/PbABIFY0vRBYi9HzcWf1YU
pxQBL2HaPQHN7XM+g0aTqoJutoHjgFujfbdgfQuXsGz78JcsLx6jmpEqw8ljrCQ7iAofywEjHN/8
Ik/5Myp1UhhqF0c4fkve8vwJGUDFIRJGvo5R2CZr3eCBbqvI1CZTNzgCfzhjW4HJbnVfYnW2qSlt
TRO57wCuabReamU4frvfMXN5/6bGHDo0ejm9MR5igF+zcEMvAta8F+rrx5UQaO2PIQesLhQDAeyP
Vzxhcb1zTZHSgRog28gRWIcZvQZbv8oVLHNr5c3Ggy85Wyp9yMnkWHOw1c5NJlBnG+kjBu3Lf3/f
HqMi58kPtxouSEvaOtlprOXiJVViWSMNtmZL/HT+P6dOWjLjL5LD/3LNNJrXU3Ps83FAaCuV2czG
P9XyBSIXbn4ZY1uGND90p4R5sdFpY23Ebm2UcIjiAS5bMuI6LC2EE9NypBPenoOFJ069zXBA1bPj
7InvVWmMgmi7ZC2g4AfihhRN0xZJcrKKXF0QkgMbmYBszDaoMnVb6hK0DNRuiyidMoJ0VynVKQbm
Y0cT7Hv91RRmUQdU2dDA2iKipaeUdzfJcqo8w3MN46LiQnyhfrncILPUgPqlFhnkB5v8tlXX9J+F
3f9iOLf6qzOxoHNBfUk4uWl+87WRLmTXfh0TUTLkMv1mJMxvVIzCrum+TiuIcipDPenX/AQqtaYX
1vySqbJdqLRvGbu5As7iYbqL5JL5rhxlRtzLD3mJgkq6ftoU5nfnThbk3KjIs/mos3n3qTx6t7L0
+NndbjPPl9xamh61ChD3qibTb9R6j3mqwwxN3LoAe2v3yRGYN4OVltdsA8C7CNN+FVBVXP0nNPuX
RCOOQ/YmqawD5ZqPgPWi/xbt21OvJpy+Z8Mm/fSUayziXc1XGLkoyj3C9tD/5Mt6mOdhP1TWjIcJ
q3LwqYn/XDIlAitTZp9AK13fRQcXK7D4wS+6sTbjPgVipxE34XC/WDjk0ynk4Z9jyU7QVOYaHmvh
DY79/7AGBYIZP7o6sr0JvDcqp8ktC4KSLsmJK+UZ1Wmd+HGO7dxLCRFTfipPv7Z5OWXDG5FfBtu7
TWfOvpgqwLuh6lSbp+7Et4re4nRxKn8SmTf8quluR/NlquspxF3qiLV9fduzUG+B0qhhcyHLCy2g
Sf9vFQVxFU6g/0Mo4iUEqXuDKKS1uBOx21B4QVhjIDXLU37989VBE+ypCRcvCO/4INzth/keKojq
ZGVgqzJWiK6IyUYJtsipE3gpUAOE1ILXRs6FOsgSOOnGvao0IA6YZ6uDwcy+mQ1MmB71Wgkq56EA
mGevB9Zj+L+184WlX6EYmf21Ivkd4Z/sKX5WPJuZ9sjwadjSbPkjkR0boIW/NPpNJjMQiXvZTRLf
nQB9j4y2ygZkS6/dXKQPI1OhARvNnlPQDjGrQKncbzYPjCn1TuM5P5usKTz5FB7mwY4tRhVJomFF
mpkNdz5FZb3fRHVpPNIZqZF9p1gUZNZ9p87tmZP0cww+ujqFxuGn4zVksWbRaOikYLTYRs7QO34+
5NhQStzvR2VWQLXPAaYi6807Yd2Q267RjLSwNz6eQQy5JhIBMW15N7Kt/+1EBcJaq8KxBd1B9CyU
9WCwTLAXWKyc9rmWlY4GHP5noltUoPB48pitLzlIYVsTbJhUWgtpdVd5A+nGyRJpzs0e+sl4yEL2
mcu2FyUDKHnuV4c4aQjD+OjXPCF2CliUiesamsZ9eQJOvIGw1fu/2jECfnT3WdsX+w5ozex/5aBt
N9g5tNu+qjAegzkIQeHSalQfyHIAgwzAx22K9ZnprdVzS28IO7uUTRRveH9bbZCUMX5PFNSuD3TN
613kNTxup3wPFamugsQttPezaH/wZ5YL+vEAatdyyXCC0TGrx/w4Fu3COJjmE8EWT3fil5+fqEKf
4igkP/0XpIoupWanzgQa8vBXmV08CG8yEwQospRUnQun6xUWbQ83UZ3XEprjVnNhkbZqHUZEXcMO
mfOnom/g1eKvzjfdXbPl3Uhfc6QSzMhXONaS+7s/mW6OPgEw65miA3xQRhcYSGKBYu29HJX91M5P
mMxqKU74QMejvj9KgSqiYPVysLECfqC4xjoUPzYA7Pbm1eqdNDL/N8AY3ZHzMg6JnwHe/IKNhcAS
1tMhVUtz6A9d7u+STE5kmWue6r5k9SrI4k7LNiGIaA1KSWQB0326PodSZdYPHtC0+i31BndX5eAk
IyzvZ+Z1isizdnH2+hH9RRyGuvjKz2lBNHszINeX2TdN8EO2kWGbJdgsIf+iXGODyqZ0vuuhLCYU
9izVHMaJhAfN/n5DNCS9YlJq6QN5Hp0f+qwHOOXBnaEs/41zQJy53cI3D8XTyP6jxnvEFvImDr0E
lCwhlUggzpdHWwApZhtKNCo0fD3EZNlYbJvOJhT+wkqge33u1dpb5nEkfZO7gLB4tMWEuBJzF35P
rAAkVTR0LHFjIkolf5UG9BQ+qAzY9G7+mhZa9DTOSUbGPWqk8H4s3/u+LKDb45+IjabKobEvJef1
QHrHhSpGkoGH8PSVdVfBTmMCRQL+RpN2gsWBZPAXnnohX8HlLbAF0e/gjFxM+/qaFOYtiBIqXIC/
WKQe8B202bTkaQ/PkKDR5cH8EcRgrPU8D1g89O9+fk6RcCWFv/VA3DjWGwqNqV6zCkxlDxU2ULfC
cEQQ9G4J8CnkLnHKV7SRF4VSSlawruJVzo8MI2VHJm1FfKB0U4hoc5Z7wB5Xgne6WAWq1w/xVNJC
VyKxkGnZd0kyLzCl9eY2loRwVFjpivYpLTEfFRSLteBdH6HHa7waO2YKV87Ws7TpRRbKN4vqcB75
P2qJtGqPg/Hd8FWJ5Znjj4c0B+V3ZZX6nn4I/meKN8th/GINl2sPnm3odUAISY/B9GxHSiXBlPE6
3jVPSs6NgHkE7PBD8M1YaRtafvdDxMhbll3/UHYS8A1GqrH4Uj8AjAqPbiuAxuNIo0Srpl24ip9E
pZ+JDJonOuRILqcvhJo86AncFz31jwEamZzC0qyNYO1WsjN1mVOSyTD+N+2ujGNrk/AFVy3v5hJY
PJHiRG2YzE4+zlhkzcDxVlX5ckVFkIsGzZ5GUT9GgrRQl06NB9dRvvqO9NQFYGvbU7QI/asXBO2o
2j/IRx9p6UaoFz/02bNRWQS6BYm3olIlNQMiRkIYIaI5eSvNd/+j+n0vsVMRciYc0HHheBp1xg4a
+pSnd6CkWGpY4Jey07NUX1n9WZRIa3dWePm2APiRXBQmZ3vKzBQrIKFzSf3FwONGq6Jw/QCpOyAF
HluSpo+y1BEuWxruL8DxBs2fM+CADDx3YOKUD2QvxiOp17U2n8U0cFstH2K90WJf8i+A5GTlnyCL
VSq3FHzzvHi7/9N3kcNqicl29z0wj4DgB9tDXPwzJKDJ8J/Zw2qOnPHwOBiTFGuwu6KoibEQBsX7
UWYcS08bKR+aN5i9Xt2CO6taQb0f3wrUBZ5W2BpkQzomHlHJrkR8w7qMBtj2irt0pAh8jbcS7MRg
SZ+RWUCEgHBI7Te9ym/aIrD7V9PkPAeG1XpWgBn1WXYU+i6DewFzeX6cqHxt3GEuqkKJLCM4wroe
1Zim8c/RgliUHuX8+XAKI6bL2ZXurwm6Djpzdz6WM2khsqKbWpRNc0FImRFs/ifVUtnQsnWXz1QJ
smZc3OKwZtfUIuoTqlJWmdEpukiIy4pHjWwNKYOg0QTO2URvPif5gi+pNExrI9uOGmU/d/dEVd+U
ld10Q4aCtMqAMalV8FwDtgGm1kI3WvvSfuF3kKYQBb3kTCD0sBUAu1Tc6jjXbMfxJGOyw4kOhBQU
5xNr57N/t7iU7+HBFw4NP4B5Sz30awaCMr1DDrvcd0RyZG9wSnP3jPU6HNEzGflPDkuq5ZSYKhJu
StZRkO4RVYTJtK1o0PSVfBp47aPkvvaYw/Q/3DNxbyXj0BPHmC/DymoeWV1EwkOJTxnKC9rwsDPU
caTMkVpdI9ckpbMZHc3sH5gIaFoqHWTOPdC+8k+qZuQuwcfxrv0zb9xnggEaqy97/rEbOwW4F6R9
QZojV4q9ODE0dZy1J7by/KX49vKKi7BlTPAfL4FcZtyB/GpfzwDn41DikFUqVYNyaQ1hpJI9M+gf
dsuzAW0DHfhQO4nD02sub1PgHcjPPItXL4ge9dy0J09WR2GXORUElau6s+FJSF+s0OepDqzruCf7
iH1cT/p9FbNIImx/RAv10pscfBTc3RR4WsR4Q546zk7ST+wHPz0qi9GGFZ2aFepPJVYdTQnOjVaE
WJ+ZpBLqAB+bW63WSedfTD9DMEh6SczPTAKLu3kYW051xL6hRGhuc4n7whI2tOokMZ1/IUZS9/LK
X8Os9gv2MXbBR0M1FKrQw/k3HfTJTCKkABYTpaj3eWonVRGzHoURGfEL778hAe00sIn54rauDZ9T
vKqSzqYW401E0J4LCKGrg/q4AXiXH3QhLx/m8ngUXCz1+Hh+JJgvCz56RofQ7+3ZxNOxUB0/vKhQ
U0VhWEQXepnIICV1jya/qcL9bwdWEYOABze++0Is9zeMzxJ252JTLu8eHS5vFwKIpacHcWu/gY4m
P4xYeHGyoYBi0TkyCwE8tKI8dSAHEsaD/E3m4SCLQpy43VihIZYMwUuTc5JDbSd+WwD4gIJsJz2R
boyVbgF/c83QhG7xrfN0YAKa4dCwF/AGyE5VUGQGdzGpF3nE8Vr0/yzbqTWB/EX+n41S4Ylpvp3/
hlTML5EGH5+6ss32Tyc2mMbeLJS5L5rUEUEvBdwer+EMACe/0GBtl7Ce7v5jmyFpGMnAXBCLcwv8
CztktxSF7zsw3GYZRN9cWSaWdUB3wz+sqWkOK+Ua6D/nBs5xMkDc5PAS0l4w2LMRZm9uhcdwxAU1
4ClpXq8tSwD5SbRecdHoYbG68M1pNdN2TnZKoR4k5biG9kSHVaBF4eT9JDQxe99X9mYeGOrBdhj1
yNHNpLVUPy4p4/hYbJBzl3c0UTbMA8gyZDEY9PeyqZhmTWqao+hjhMFe+rUmhB1VmteBiun7Xqmm
F3PVjAO5cn7fSawR4H+Gt5hTJDkClnY+Vjk1dgjvkTyZPiAlzhbcpA1qiWxaG6TWdWwVDP1Hb1yb
wbPrfiGfPvi/gHp7vxrPnWVbp+oNQWRyQhhgoLfVtzHVzglmwLgs34anx8oInfVAUQIPlNB55YTX
y05YOU05gV2a7CezWE1IACvNq3HMmu1GRFKkoTtGABESiLZI6qLi3v85wI8/TsQ9rXhyGSV7QvHG
fyb97m+8DOmkJJuN8h7+7txLBCHGcmzWeOU=
`protect end_protected
