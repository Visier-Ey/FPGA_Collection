��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���J�l����9���0?��l�ȝ6f
*�
�7��;�5�I��E��������&aB�Btkiԣ�xyx�/�L߁�#�(�Ʌy�f��vp�É�5�"�*�v*�ْ�f���k�f����h�L=�`5h��"�����U_��n`��l�-]9�����Ϋ���/z?���l�J8@׆\�h�,��3G��,�O	�"0e��)�1�$u�&h�a��'w�� ꄭ�����٪��O���lWљ$Zr}��e��u��hm��8
_�O�6�0|*����Q����8îv�׼ɋ�ъp��|F5j7'�M�Lc6��/9Sv�\L���K�&����I�td��OhfEA��M��g�A�ŗ��l}�-��Jv������)W	ż+�J����d���	�rd����5>Q��65u��m���[|��5��P���%�'Wet �(��	�5����N���D�0���ْ�
����Т~�~"�T��� 4������^eh�'Q4(Ȇ�m�N�[>��y��皓Ē�%�7`	�j`��3dD�e�SfP���ۗ�;�fS@���x0�
O�(�T3!�c��k���32��au��t�Txh����D�I�*F�D;X���=���'K�	0w}[|\�����Xf+�>��*�ͱ� �΀�".!ݯ�����XV�(q=�oAZF���] �_-�)d��ݲ��tle�|��	�'3�j��Y�)�9$;S"&'qV'X�kS��,)��L�D	�R�#��(;<�fr�Ym_�Y!�i��M����I�3gҖC�����71�iOV�~ED��[e@g{!2���U0�1�2���L(^�����-Q���=���^������](q�h���	N;�]�`3�s͒�+#�3��!�<�yA[�%�tJw���͞�}�3.����R��@���G��M�@�)/��RՍ����yc�,D���&���V���u,��.��:e�?�L9ۇ��|�5{�7鋣��'�}t^�%'� G.�{��g�A>�_4`z	�A��S)h��g�SH..|���_�y ��>9Nɾf!�{%?>-���
���Y�H�E=��}-�h�w��@�#��}�BM"�m}�/�lԆO������ �8Ǒ,�ONRa���^:�,C�*�4���]���������{=�L_BY�#��1����>ɄWA��ͽ��33�еE��m}��##��9�%���4�W��9;�G�^'���E�O1U�]�E!� N=`�2<RvxO^i�u
R�?���^+�=�y�$��-��!%g�Ԍ�d�e��AXQ������^>����:�>o@R��h����i��vXf@��db����"�tr��|"���/+�`�q�ݕ	t� ��d�@`�^}�wde5��B�RK�e�xvw1)2�Y$��ǂ�BV�1�:K��J6Ɔ1-:~��dR�(��������u��C��h܈K�4L8<E�@�4�K}�AO�"0^U�Pb@+5�է�T"��8�;� � @x>��et�}x�"�Ӿln�\��*��k#��į�ѮQj�����`��/N����7�׵E
,ۛF���j�������I��+O�K�r��t'O����AHz�fȗ=>�3�� MN[2��I�#r
�s��qp����~�K��Y(��r��4�;��DR%ǾQ��֎s8wz��_p����b��j9�֮�J���+!���jv��jR'�I�F�`�U�tP6<4a1��>L_q���:�>�5?�{�_���?ʃ
����3�����{���V��Ă3�.�Hh��>v:���CF�Qw�������"�(��^�J���y�v��h�/�̢d�Ӝ�Dm\Т�ѷ�N�,�J�$T���*�Isk1<����!ӏ���L�jt��2��N�_�^0T�Đ+u&�b"l�*0��~��I�B�#�L#�{��"�'��]���=���[ͣw3�5z��0���I�U<P���橭y��S��)�2ZZ�aÉ���6kc�)u��ٕ��6g6���֣\Qf8:���GF�R.C'�ϙW-9�AT��ź\j;�&.s���v�)7c��4�@�H�Ȼy�D��<8�iY�P	�>�OPn�1�!j�+�E�T1�Jf����?�1�U�����qW��~s�|9���	�i�Z�݋0�'[����PŠVI}��@�l�4L�iPN8Ǝ����� #�vv��C�����2����ng�6��b��Ŋkb>���N���&;lI?\fl���
�^�Y'�7'[�~/�eh��M�S��]5*t����?�ˏL4m��\��S珔0dQ!�cU�\����=�2���4�C��8��_���]�:\zM����r�2*DÄ����DabZ��|LGA$;S5�5���'�#&JX�m�:rxǣ��V�QL؈�����{��.�`����IL|镴��v��d�R`l��kB̕��+�`�6x�d��d�ۼ3&���&����G=�< �ʾ� ݊���o�x�D�d9����g����"�wH�s�d^[�l'����ڧe�C�������rGm�M\��!!�yO��.C;j�ْ�B=��@��bH��H2��+���!:��iL�T��7{{����`�S���:�g�^/'�y�~F++Yl��O�#����ZN�fE`��JWU)��s���(*�N�˸'�k��\�h�󘡶��n�!.�$ǝ��H`���l��m��wl�f;��A=��#_CU�q�x�d�<���۪���$��RЀ5�§���!k��v�Y�u����)��Yۘm�����1[T������kOr����SI?��E����YYSnx�J�A��4��0D����wtw��߷QΜl=�@�Or�Y����)�UU� "q�q�gxHL��
����еO�f��_~vq4wfa�p��(?���`�MG�:KM	yPѭ���nl��͞�qk��"�X*���1�(Ԡ�c�]3��8X�>���p��l1Sf$�q}iM�{�ę�B���Jt�"��A�:�}�����tK����Wۼ����-�;�rʕ�x�͌�\4�h�D?h%�9m� 9�����%lA��b��@��78�����҃$�I0B^i�����xbSD�_Y�  6H|�i�LV+#g��xdn5����ۦs��+�s#|#� 63�J�$�J���^��e�3M�Ri)�B�K>w�p���|�c[���#!DM�l �����y�&��lV����f��n��ݭ�ב��P��>�:w<K#����ОP��7iO��F�v�ӂO�PZ&?��7���^��o�q��;��0���Z��+ĽB�t�'��bw��#� ��;5G�g9l��4��d��\3RcL4��3Vǋ:4��(�Gvt3Ig����h������ق�Ys�M�n�\�a�8���\n,�d�(�{��"�:�6t#�����2�)J��͗��UJ���_ԣ�M��өk����k����]������|x��Y[���fZ�W�5jz�v؁>̓XV�G+/?��t�F��ޞ3�����Q4����s�����8W@��7�)�7�1�����a��J��
�%RR]*x��Ŧ��Z؝�E��1��A�<������p��<�}���X�ꀵ�2�NB�c���B��*Mts������F�e\R�ƻ3����	�����Rz�.���*J�����W����a�
ߑb�$	j�Y��L��*1�f5؅5����K�!4&��N�6�X
�U�)�s>cuo��l�� �ޖuܪ��h�fڴS��[�`nr�z�==����a�F7���c��l��r�zh�Di�f��5����%�~�"�S�3�$���"Cc���3���i�Z�� �-fXB�ؙ�;�7`,���s��R��첈���;D�a'[x/3
��L˱�B�x�w\�L�-�=���b=81�+�}�4F��<?|�me��XH������<���t&��L�����k��D�"ވ:s�k�DM���o9-�Z�d���Yr]KHU�b��N`_?q��o�
�{��-�@���3b&�ֳ�zU�{�
�վ4�� E���z�(�B�P9EUɒ��5�j�`C{zĢ�gM��{]���(�x�����+�>w ,���?]p�
�aZ����u9ѢA�eH���B[
&�?{�Y�uH�h�F��4���-K}qK�d����B=H'j�|�b�Ma�����b~����XQ�S��*�9?bo�*uNC>���"Z�,a` ��K�H�|��x$;#���,z2h�wj���fz1f���G����%�Z-��a�Tb��2��xՖ)Sg����y:�����Ln�K����!GB�$�:��tc����^2|iZk��Ϧ�rG�-���eV�08���_�O�IR�0y�UBX��	��_$W�S����)M�FZz��@Q8���A��e.o�"C%�b�q�h\\^��h� }P��jk{����ш��ށ����PJ7���I�r�ʚ��^q;j'����+l1M�cI�o�6��\̑�
���~$�/�
y�˕��(��6��Zֵ8�~�jIFL�)3���'y�r׫;���-���ݚ�׶�ŧ��(��0�q�$5�6����1S�5�W���ȋ�% �}���55r���8	O��|�~��"��	�"���r���a�6_9-f�_+�+}G��F��!N�޿v0NI�1@`�~�8�b��`$K^�G��Qc$m}�سRCGy������
)��r �75qnꊆc�`��nc� M������I���}�Y	*��`������G����Q!�$��C�_�*�n���k9���i]����'F�5	�������VlO=�[M�2x�	���(�>]�A<��a�/�D&��%���{�sOl����->�L��-���#�h=�b�>�4x����;ϥS��-�a�I�w�ߘf�w�]�HѲ[җ�rƻ+V�<�$W~5�����8�(��p{qI���,�ŏpjȞ�0s���< �f����\>]:�U9CJM�|��S�kX[;JoO�V�T��Z�{�����}���ɚTY�tօ�X���Z�1���-Y��F��py�ܛ8�T<��&%��&#�V�`1�G��ݕdT��΍�7i�4�B:IN;+��2�t�Nˍ%�Aufy�A�äY�1�Y��"�x�F�,��L��=i��\`q����%�Yd�N%?ܑ�����X�."��Z���`C	B[n�U�#b8�2�8\��Pa�F�6�����113`Q�{9}�=�wS�֧��]�4^�6�8�B!�n��a��_�l�n���p�~!�Dl7�����{,��B"�	�Σ�r�c�!�I��6�)ɴM�"H;QD�|r�OLZQ�>Y^(��'Ҫuy�T�P�����1�3ϴ���(�k&���Bً$�h�T�5�ǘ�&N��io3b����t���Uvu.~��3`�]hf&��d�e�J�h�;])al���c]�� �NZ:��Ǽ�c��(@�ܥ( �����=w#���w���>�33�]��-�Q���)D���G��}'!6�9��4 �m�מS�b�b���
��c���?��.����Ƹ��	bî3�a~:D��v+���FrOۂ��p�a���'���o��ty�S����`�9���P#�W#2d��|:1^E���}�1��e�~:)�����o!d�nh����E�׾�/ᴪ�1S�y}��o.X�Hw6,�"�f��U:b ��F!��wm��B�bwt�N���)c����]��� 	dnu�H��H���f
�0����p�� �m�S>V`<z���)��
��ƀ_�6@�J�s�3ʠrE,
��P_Y4	��{�a�ԼT�m��ˣ�{��[,���^��U�0���������� �}-H�ϔ*�Ům�WQk�[X;l��%<���_9�[�����i?N�l�` �O�	�G'�~m� �<,*���M���]��P�$no�e�(���r��
|a�ei:�n���M��ȳ����q��.x�cQ��i7�<��L�J9F���5[&)`�ˣx��sC-qL�W�tl�w��7Ps��d�wG�Q��I��C�Vg=TK�C Y�Qv�r+pePBo�kUꚫ7?e9xÕ=��T^D��l���H�����i�e��{V��s{�5El��Ds����=�c=ڬ��w��'�� �	a��4:>��D#Tϯg���Pw}�95�|���bu�`K��z���>�s&� s�%��(�$�YX�Q!��PI�%�s��܈��B�l.V�tA/�n���I�qLp�0��6���-Ghw�;�S���4�|vʗ�9ym�����_�J�NgW����CM#}��Y��
�b�h�>t;/��d�v9
%a��B&�b��Dr���Ȭ�ګc��Y�aB����c:�ڔ̑�"��Gǉ��*���y^qsSF|n�槡�\ ��<�5G�V[��?)tT�!{�YI�6-���j'�/��q>��q�ᩢ(���g AG��ԭ�u�rEz#�b�L8=��Lo;o�n{�3]IJ�#a�|���tǡ]޻���w�5��ӫ��r�`�1���&�/��f��l�.�#fS].��w�Ǧb��c)��F(�O�W^�\���M��� �vA�0�P;Vu� LtZW.��A�4�W^&�u�L����.�_���Kâ����TSD}4	G����U7��|�ud��i�������g�s�Zx2�sgL���zh�¤�m%W@8��~�Aш�o�y�����+2l������h���}� ���8A�Ӊ�={,�W�V�=���M4��g���h�]���ޒ�,����[�e������\�ʛ*, Cm��c���=�����p�g��t�8�ULt;��#(:¾���?L��yQ�v�;�[�������ڥA>����a�Ȋ��&�p��8]��}~�ע:��ŝEJ�AyZlK��M��,`�`�e9g�CB��s7�{��b�P��q��W'L��g����|v<.�Qf�ɫI��	L�?c�ǼǠ��mڪ^����D���5`Ef���D:�rڤ��(u��렮��?ے��Tofd�"�Uн^W}P�<�f�=��"���WiB,M#�~۾V�*�o34_���k���>̬�P�4��Xө���H�s�\�75�J]_j�������͕��m�9������0:�̩�\�:�x�w��_f-HL�8iC|���߃(]D���c�|vM�27s�8�/��R-���Y �\�\�F�g����v���sD��� �M�,@?��`ƕ+{���ŎX�(ei!_7��Tԅ�Q�I{�kc7Ӯ:Z'@|t������g��v��.^�R��}�ҷ�~s[#ĝæ�<��XV���E�6X���!����7غ�>^.�Wr
	�R<�g�4�K��͠?��O��Ùѝ� �"cy�#�IF7���[�%̞��tW���ǰ&p"����U����Zv6��/� 
y��}/}`V�k�pW�t`fhS�i����p�I/��}S�5c�^�� mR��	4�<HH��i�͊^����̘���_��CT.��v��Y�Ϛ��:���#4���0��ſ��<x�EL�l�Z�D����j��Z͉oߵn��u�^\�k|z']�J�ٲZk��P��'����FH�}K�c�	\$S�у��j)��&��y�����,��]9�b6����c3H��1���P�κ�-T��(��?(�@�����[�6`��SSq�@�7�2��t%m�a�g.��o��I�.��*�m�<��1��9g@�ď�������;��`��d<�<��T�b�Ƃ�ּr���&�5�^:�;���:8�w+��]��,�G�����G�TD�����]��r3����\fS�k�b�)�7+���Bx�*w����{�by���Hٮd�D�$�'��(�}�=�9@$���ϋ-�I�Ck��y%s,�P�F��%����<��"`��_']�)T�<�|�^�wqr�`��*��@۔�bQ�`���QM�c�&��u=�_�t&^o����+D��MyD_=c��>��qo_���"������5�&���E룍C�s������b�Ֆ�U���E~�u����+_�ՁZ���s�ȿ�k6k�2�_G.���%AqPށ�������T�O��q����U�S凵��O����9����`�ڀmB�"�z5�O\	]6V�_L�~�=�IL�L!)������!=B�P��E�j#)��9C^�w��#��	y$e�
t�Z:��B�o����_!<KP4���A�V}5	��Rv\QO =E�:���|���I����y5L���V�h�p���5�Z?�a�qP��1�[��P4��,&J������#���lyB6��\v��FU���<Bb�WzӞ@�1��o�U1���XM��OpB�%u�`)�܇�S�:�!�x�l�IYv*�`*�%��!���r��?!�'�+ؓ�I�o*jK"�����$���kO'9~	�Lw)��r���sG�azu���م�,��5Jc��a_��J�����7��I��7�&\:v㟯�j����ÈD�ܮ���#wF�P�A�x����+hE:�P��Ȯ�
���y�5Taf���A�4��<����נ��e"EH�j��j^+^�m��p׆n��y��Ҋ�i��o�Yד�b�6�ΔJ����=3�wL���2V�ێ��$��a����M)�Yy\�̫�L*�r���ݩ�Ӂ,�;�2Tҧ��A^P���$cdq�C&��2$qz�'%�����)����x��`b���ag0W�e:��)0��=@��ۧxjX,~[��D5��V#!F�`�:��c9U�@�3�
�m<0F �58�tɹ-f\�.�>X����K��J��~9�'�0k��<p�����~ן�>'6j(I
;�.$H$�υ�m���#����Z�=�񍭓W|�'��]��Hp���|�Go ���n\d��ȹ%e,2�m�e�!,��QR�s�iy[���e����x���q�x 2@*��^C��WD�ܷ|*�oFNW��h�:��g x�U �<1k$�����70Cn�����r���?pN������dD����&+G���B5`}��8c��LV2�$�6�f��^�4��x����Lٴ���ZZ���%v΋S����(�~����b�=Tc@PHTò�FV3�Y����^�$�?v�-u�*De�^՚E�gB�9�5G��� �l��lPi���T��lKږs���rAs�uoj,��ݜ]ȚH�:���4���\�����7MY�Gr�8�R�OV��*	 �w)���[4�_�h��n��O����w�r�k�53Z�5��o{�N��t�����RW��d��`#���֩�t�á��S�xS�o��������\�f��t��3\�F���k���mOՄ1Ax�)���'ӈ��	cn�3�U�������h�E�٘f��p��.�A�s�$�z�+�y�&�j��AEN�"1�I�؞iof��\[��Ϲ�2`L�2���\����Y;e+%�c�q�	�K�y9�oA���5�H���^C��h�#3�`��v�JI\���Q�<�_��|����KL3c�� Ft8$⑃>q�08ON����:e�Z�c%�`>=4°�����������?�Ī{O��x��g�7FS�O7��Q#��=Q4�P.�7�p�����5%l�����]�N��V7V)�J�"����O�~�>��pH�<���ָC���h�18��T�x�F1T@�Ŋ$��G� F��.�F[�@��_=e�|�zE�w]6�m��3^�}��P��pG<`�~n.6���s�_�%�a@��m�ޤǪ�j�ͱ�8���~g�\�1�I99������)7��.�A�-�c4���y����ga)[� 6���9&����̃q��fRa�����cF�n ��c�������Q�'���S��%�����?)P��5����4͏ y܀brşn��%xl(�ȸBK����7'lE
�םc�*N����)J����{H��/��eZ��#�1W��Z�A����*�$E�'ݼ_�"a��xpjuKu�]U��w�i4����p��>,7��H6���Pa�?��h_=K�8�FV-��ݬ�*���ǁ���GG$��v��'������̬�9��+Ϣ!�	5I�zj�Uwa��_��Ķr��iz�����#��\��܄Pyj�k�V�/�ǻ��|q2�a+3�xtΙh�`&�_�1�+Y�<LI<I.0�"%x@SҪnX��@)��1�jy��$U����Q�>�YȦSz_�������6N�j��|��G�q�\bGծ$�w��
>�O[��}�iD��W@+�p¶J^��4%!A��A���=�l
N���q��P�#s�[{���x#t�]�e�xK~����B�.f�>L����\�X����鍆��,}�c���9�}�!"���?�R��Ѵo�p*X�E�
�����I&�_ �dñ�0�	l;�����T��F���N�U��?ɫϾ�`"-N��Lu?U�
e�2N�'��Gu�N��1�����b;�9[�cJF�R��:��Z�&��`�׷M�sC�B��>��P�3�e�!���5R
2N���'}=���3�#�� �]���.����-�=�)K7���ɢlsw"�f�l��≅~B��#a4��֔� kS� 3�-֗/kR�&y)�6���ָ�e��2uF��2�9�.��%�^�������E�H�u�Pb��@��^|���]��ϭ!�� �΅��"N}���V�~��^�|RkI6�GO�`!���� 2h��r���h4"��ꑏBVfnV�c����_�[���lw�L{���J��)�8�����%O�ty��hzP,����( ��}oJ����j	Aq-�kq��)�į��a}F�>%�� ���9Wu6�.f>��n'q�Kd�嵘��� ��	NT����מSf�[-�C&��c1�eC�B�X������	�Y��S)2�|$����h��vF�U���t�a����#�{�-�B4]dE�|��5�+�c-��G���C��X��N�E=R���1��G69S^�e���R��� /
SRG���|ֵ�Z.�����y�,�z/�Yۛ	1=��˚���D@զ���&J�*�|Țo�a'�WY ��ع�njAC�����`To����t�j�>xś�Vs�,�8��S����36�����Ә���㦎d�nOab;�.	�
�W�Q�B<��b.������/�(B_Z��3�q��E1<
�¦l=�.�Tσ�=^O٫E�'�S���g?k����V��T�T3c�WZ,���]P�}޹�}���M;�(ǚ�AZ,o�>f4�\ ��y���!R_ 7H�"��:�gO�L��6�ߧ&W���	j�}�������=�'��i[����2�m�F�3�O`�"<�ec�P{&�;�s����ZiR_����R�1��6��'AA.��@�ˠ<�����"�>�^����ыh�{��������ô��7+�e�]��oѢu,����)6���l��9
�7�fAyј�d��*�j/"Y�P0�%o���c���aN�K���x���!��k����� UI���8&i�^�[�&��#/���Ёy�	܀�}ɬ�i�`?��ЙR.�#ؽ �>����C�����~',I�Ƶ��PǶ�1Z0X�>�簯��`�O�~��
I��ꉻ������lc��{��%����Wi�E*ZƦ��Y7Z���ӱ3-cp��������ي�������+�И�P��!�4FgV`�Mf[�.|��D�
�D��^LxN;|<��5���b5u`a%�L��a�o�ƃk<��2'2_�`�0���,�`��_�x�M�O�$��k؟��~+\���ud���|.l������E�O����?<��#y�\��MD���7���K�L��	f	uQ�~}kh�u������XpЉ��_�9ȑ��"��|����L�=�k�I�����C(��(�;��k�!/ڲ;4H�S^�By�^��O��qf�+P+�?@����uRdd��u
���u�{M�8��<�t��񩦞S&"l��H����	�7�:�.�:��29m:��t�Uҥm}�7�([�K�.y����'�j׻'�N4�M�����g�y[��6M��+��hS��T�8���w��� >J� �h�g�bZ�����_ <EQ\�8!��@`����k6�Ӎ ��-�^�C0-,Z�p])��c*���1�DY�A	_�t�U���j��o�ȓ����1+L�צ�Ƅ�
_�7!+U���Ip��N'������gx��������(f=����ܷ�k\�@�ů��Q�u�s�aw�T�����Rɋ�`�����_�)Yl����ߗ��g��^�W��oq����⿪�DQ��4�O���q�V���R!��]Ôo���
귟Q��S�v|�p��;��%���['�ڻ�6|�q������etQ�s��s�U��do�9:Bǲ&�U�CY�sA4f����-�BH�s�2j�����^��IC���ӳG���i>Z�G4W�����o�4�ӽԱ(�C�Ɇ}I%���u	!7�5�<r��ח9Jh~U���i��R���H�#����[�,GWM� ���]QN|�����ܧ�X���B�V�<P6\ف��e3�>��#Ʊ	����k�I}�`!#���q���A{�(��&��rm�o^2gXK��*����9�b��a�C����h+R?�����p\�
,i|0T�{�6���>��9T�y�����������%��ڑ*�,��?��t��Dߔ���rbuj��vҟ�B���X�\=�;�(�W:�z,�M-�\�Ъ�������M}"a�ݼ��.�Lj��̆���WA�7\� �� 걮c�'3�f���28���y!��.	:�'FڄD�
�f�04�*��
亣z��	���'�9�+>�5�5�X4Nז����ȥ7�S����YJU���3f܈�ݠ���$�E����.�yE�"֐ܣz�"�o���8�N����5My�#�>B�"����`�����ժj+y�#���Hj, �,e����j$���R�}$�ĐK�=J�ݤ�ùz�11��װG8��A�o�0""�����8A;�_-AL}�f���u`��;kC'�FI�0x=�R���Ӡ;$UwP�k�[y�.����<^W�j奣;��V�Xrv�p���D;V������{��7?}Ǖ;�!=�i5i#lH�m��֟:��'����GH�o92�M' 1>B8[C����.�FI2�ڣ_:6��-,y6Վ$��i��*j��͕�C٩���}��Q{�K��+��4�
�帾��+���]U�)�:�; ��π� )^���.��0?7�W���j<5��0�>U� ���0^����w���Ȃe%y�x��G5�-�)}/B�� a�¯���&�+?�l���e��n=J__T@���[W\���XL���"tG8�����,����2��ΖB�u �b޷U�]��+�T=�շ�����$��,���+m6걙�~�da.���/=��'͛�
k�̆���"�D��}��U/Xrwί�U�:�������)v�ӵ���1��+gڠ3	��lЭ�(-Kf���9l�S��CO�Oa����ʷ���F�Ҽ=�j:?�Swa���	a�)��͢�k��>e�8��Ν�s!���X����~fc��_�lv��=���!�(/
��Ǐٺ}ozO8s*�l��ω��K"��i���򑆹�!ÿ>�?tnQ���a��T�̱X1�юy���Q����"�S=�ضt�[(.i:Ji�R��Z)��C+��7����r�
�[�h>+�����
`��h���p�SۯG���"��_�Ց�Nv�(�{�PU���`�Oi�_��p��ǽ��a���h���oFy��V}B0�|����,��~���q����g/�����]ݴoja�}�J��2ܡ��:��e����b3�"����>FsF���-���y�N]q����P�q�=M��u7���r���R�Ƭ����q
O�pV<��� 	�04M.���PP����Y�]c6R�;�I����$�f� Xr�DL�j-�o�d��#�k�(8��kY�d�%G�iy�8���)����7����'2��`�'�n;�aC@d�#�!�}�����c#I���C������u{m�t�Y�S�����;�I�zG��q�ms�Ʒ��zc��+JĿ���4������-p��>[��J)|��uS	�*��m���X��8Ҋ��<\ 
Ԉ����cN�z.l��
���fiN��-����l� ����>����e�KAv�
��'p6*	5ʫ
�q"�� �y��C��Sb���;�M���]����-�_Q�|i��JU��_�bSz����r����EGȽ��l��B�+��R��`�����\��(����AJ��6�E쓊!�c��(vD9e�*!d����?�$E'�����H��}�GAW�M��P���*�����`�$��*[�j,�o���&�;��!8��V����k�D� �����8yi׺o]�C��Xb���Z�M0P�!�w�����x�N����V�f�J�dD��t��W#Xl%��x�@������
M�݀�C���L"�+�9п��p�4�n�����Y)�9�K�wIt��2�̦�n�5;9�x���~����@�k]�͟\Z�:�R��*���$�*ͥ4؅~�1򰳛�Y���Tu�$NJ����p�=]O�_���˩>�O�Ӈ	�Q�|U���zM�$��i�鞺��>��P��>%�]mѦn�C�)Z�qe?ٛ}R��M��Ȟ%Y<��^��ug�4���h��^�ˏ���"��~)��H%\?��HI�H=t�r�ު�6 s����B7���4\O'���R��<�^��ޝ��hz�5�K�9$�<fc�KH�J��9����sP�:���|��g	I�������.�O�Qڗ���Q�!�ô���%E�h����C+�������yK�+��m��*���(ѿ��x�(��@�-3(�~z����k�Wk������J������pnβyA��њm�xn:/�JL���~��8��!Dp"(�����Ӌ_��,���s���K��So�Ci��aЮ,�(�	\!A����H�VQ+