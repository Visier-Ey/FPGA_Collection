-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
0X0P3XAOm/qD+JcQNGeNwSq1M/uiZB4WfgCuF7h0LrbZpW13Lx1FNFFDqLbE5Ff4t5+/Swv9/eUh
wk8dLZvd+hUBd2lwuTDuq//790F4i3af624JefLipHQPXB04S9AifeYiDkzPuZwha092bOby9d3/
G/kq0T3qFscholM01NVDlSRtJalvMCphxIYZyCO6ZoHFCQTHtDsBc/Ef8SlqNYEvXKTQWU8E4Jvg
60osWMRGJdvKX9UFNyTKULLOpQNFe2NQLPvHx6PSeo4skH/dk8MsE8D3TwClCB+DaO7HcEhcB9kH
vr27neZ99NJ/a+Dv2/KXwVtQpcFX5c9kf/mznA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 18320)
`protect data_block
7Cj5pbIr2cyEiYD+lzTEIGe5pcBkIBXiNfUfHGa46IpO0RYMQzGrbv7s/lfyw9bLQduleOaVsVON
eR/5vlsKEVUGyZ/qdszIyYk+EazfO9Dm69l5eKP41uAW/oi/wi+J/Tku5SWU1mNE9O0fbtJ5quZr
xYLDRrA70TGXJ4nE8PK1Tby2pkjwpa9xrQ6Xi9U6Uq/02jo6j70qjq5oBMAzL0mSMINs/t5YoIcJ
1cTSUP2FixZM2/nZLhtfcrH3QEaeTAfwRiq723X1lQ+PYJuvqMcN9Z7AfRTAaMl8S+9Q/1DHbU2l
P18quIui5kxHOOL0d+++X6rF40hBwDrQhwFmGWX7uFMiYDgXOkgTr43qzmMGz1ij1ntDZIfXWnyW
TMK3Qae/tFspEqhfv0qlCjQQrRcQUoiFVsQlWGRx6BOAvWYrMosZW5K/+tVCgXwEbOxjeJB8B70u
xqxPcocvxHj3ug53pSaAaIgZd3+ESxevaSAjACZqGooUYWbo0DCCzFc3wnuf76M6qJKCs6Btnbs9
cDmWAuuWoc40vvgaE9Ytl59eza/41jFWBoar6NiLWgrB3GKorQhmw6hk5NcepquLbM5+j1EGU05B
Cw2oNC3TWzYUOnjT/bj8CjIbw4s+rFBFJSjRgS8quPeScgnefip4Tg2x6mk+z54Vh6pc7b2RJtQi
sRnji5H7cm9CUMMAI46JxzsVwgt8iQ7REowgNpowMlIg1pmr1Y/TxmSh8yIKGNArr2z9NhlMSB99
+j3n+QiGSjIJdM2tQUr6BVp5UdD8MmxeCSL+M0w/ImsXT9RJEHnAFUh+SwK10Cv5+g2/wpv8JWOi
ROsM0kwkbLLid91mmJJXuQAqL0DO8LMmRPq3AG1UEsNFaZFvWGVlcCHqNEk/Yhfn21kPjtU0MXgX
+h1GLrEf84x6E0cLYBamcdOZYqZT2jokQvY5bzbnCR8ZYGs3SVG62x28ufPcaTxcZKFyvgfY/umV
LAYNJtz7vfVc/6Jbxv44budX1FwL0+Oa1LHMAJ6hL5HhFlqGpCiW6rgpGTgfN6wWwUsL6SnTNKq4
PkRTi/SE/y3THkJpuLL+XxtX/+4GcvVSCKuqnd2Eopr5IquzTU0jSkdkKRVCsgGdbVMXNmSD5oE8
gTCBjzv12ivqLbaqHl6zyShYO5Ht/ogE8AJx11KlLkZOwlNCWH7lmVzypD2TG9MUuxmUtdhkbJjO
bf56Pag5iV+iL/TBLwp15gmCr3x5ZCyFqMCHBWAMieBRKj/yGydkWSPYlXwtIFbtoy/7xqT/Ntc2
3mZY8oho0wKzGQirx0FRNVTwwlySFA23UjrPPBn1yV0cJI6gXSBj7REB0kjdY9mDTfsB1cbb+x68
jcbCUSQ6st3IYXj8KNkCzxH90hZJwQARttCb3DVrcz9KrWO/iQUz/S98VmwMzzOjh6SM0RnBt3/A
07dfwKw7Vz+BxTGEDIlMGWOnohXeIhuXPyp17fGtLibHh/ZLkWzdIgIfYeZBm/JD0RCocVx/c7EO
9+iiD/WD3StsPKdwXMRmPkp4Mqt03Rhx0AehBKFa5gCV3ukj7OKKd20GuqaE8LL07yHYH9QQiZQ3
TJp8FhFd5mWCWDKV8S+BIAq0KUdftNRwoKAyIV9wp0bQ2gpNwqShsxZjnjRfPT6eq7WRAYzbvHnl
ZDznKMJMnaDZjtB33dw3HxfiZ+ccgwcM0YStri3vgJN0m0oq8qwNPxRuKh2J/53bfQgkncuYbNq1
CbRtb36E6BzjUH25amXCpvseJ3BaYwRf3CYD7xOPwWvSRylqBTlHTFqX84q30JOO5Z+BfQ4ppIcn
xmnxWqCmy+OBPij6PGFnXdy2PrnJjqhoLH6nGkD5fOJj+JbxEATAqpcNW1VMUMDeal1yisqFScFr
yen8HOBjKlYpAtDmaFcaYUMOYoc7j5Mo4XI7ywLQX88GZlUSfatz7iQe5O/5L+4p61J/0+nEGwfh
o/Ew2YijY2fNbwYXisVlA24/1VgraraBziv5XIvPKPLI61YT4qtWd43GqQzr3TL55nOkjAN08M9w
yHn2Ao4mVE+axXZ9Zk8A66SMRpUSEmPUy/3EWwNHSRxQPB25oMpqyC4MeYdLLlW1ef4LERTskY/k
keuG3VaSFvR2V1tSleIctitrHVJuUqMk1DMqf876o7glRDcfd6EzkS2guXA0V4a0pZqeRSFOYNMk
bF7ARon5siUU4IEIu7fH//S9vxnMIBIwrQcQcv7v/i3AQVR4trv5vKJ4uWLTJAY3wWbDEPNFrVrH
Z2RqcnczlSQvFbnSuqvbmRz+4vN8tjugruSgZQGsUsg2GyRrV7G9TfCi/QOuWe5jeleS0kwRyvBr
wa+aQXHZMY6LNYgROFaUugVYke4ULxMf/VXJyGvTtkhjAYxTK6VFqoirgh5pM+6geyb3G2D1G4v8
ng5LwwNO9WzQTDS3fc9//X0+gUKkI6pHaLVsxnocOc88fvDyLFIhfcQyFOnROHa61xSMNOtjm+ai
jWMg7TSiKt1LPp5nqCcvZocUlHuw/xlFyGNUCSPnDXgciZVseqafGx96+qoVA3jHqLulknCnYRbQ
0S6oFsyq9A90TUntgOF+6t45SeH/5GtbdFzEpIWJ+/ARwQ/tqeyLy1wm6fQm0i2DBw0W5BkXHeMi
OgLyXoaj6D4dgo5AoSv258l4vINQvdByYlDgdSJnzcd0ad3TLx15DlP4T3bBh20ewlNXYGoEqoWv
+zXJ4K9Ugf5zz7g871+hlrQWBDd+1EDbP7Zi9L8TQ4IJV8SaQ4IXnqJ3G/ubwkn4E6433/QqMzcD
7J50gabbI/79rWvXUVxXDKWbKYD2zyOfvFLd/84oaNJNAguGr6nKCRYNxbIcqkxm1qwpbwSNRwEp
3kehzo9yov+cJ5NsNhAfgO+GA8H3Bo+ObXXbay9XNCgOw9br3DYZcbTemcjw21GLEjsVYTjAMv8T
0Kgn3RQBz8e+69nWpUV1KqLlPDGjAVAtb1Eu/Q6hcf9UQSzTOZwFv+QxTCMzE35yiI0H6VDEARHw
4cbq1tchmhiFK+80lMG4w37mnJz1WRfPu0YrfAOhtuvEgt+71Mm7+3l5r33rHA8e/Oq+qtv0zujX
2K9NDzqAlfX5zbt4ENGKOj4vkHy/3LaJPzYzDSoCASAZj+TcTZv9UUxd0h6Q1H/+hwl2Jx8Bzi4Y
P9Kkkr/TtNpa9NRmTIUK8jWUEvsAk+JIUmrDNQUUt9Qz6+o5VUPAaYw7ziK7u/4UPQwfXZU3y8gP
LS5zkrPQ8o/i2usdeN8rvh+wPM51GfHdn7XmqSTjGFfkYDvrjPcIOJVVLDb91O4gSZ7Pf/W3ah8e
KQZGjDrMS5/geFIvnSd8Wiq506ssdUVoxhFTaSXT+x5xb3RxlHFBcO+4nNRo23oIqhCzWKw2VQUo
PXi5nnV56I5N+vyAcstokuxj4cmTRz7bi85XfCR/Kwc8++hHXxIW4UAQ7d5cVslRseJni7PUF0by
LzyBjUCo7kingADoS6y4o/VS0X9c1WLJz1Gy7/WvFaUkenLtXBIb1eU8sfN2+NhhHtCFE5NJi0rb
VkQXUnLmOEyQure12rDHWuY0uFr0oM4MrfPvPgZpcRsKCFnFfZuDRlJ7ZeHLJX07g7i/MkTo42Xg
pWD2/t4LmUk9THaLSPXGdV/9idSDyG9v5sj9l6w6bvLC9t37sJPgCp9lsXWirOeRpMKUmYH4B8G+
Bbz02Yz6Oa7SnpaARtgMfZus3CLCppwEZfWUBMxytDG6YejObuVoC0sP9FdAq8Majc4Kbo+zsY8X
NTUwr2+v3g8n6fDK+ix2aISy6gP59wFv6VBxryA06UfrykWCdtthnwg1vxFyP0NMJkls1+tYQSQr
OKkzn96SiyubaELq+05Q5uQLT8KreWUxqDyrp4S+oCpX7UpMznQjxWGPScNiqHYmx0wUjR6SyPXI
kYnKYZ6ynsZT13XOgdOjn66jVuglXjY8k3Em2uhYockJbsvYkmjfjGAxQu4EY2X2J/O5U0Ilndm4
BtQIs0w2Js2fR0J+3t/+Omlq9VSevYNDO+voxgf0AyrhsMMThoDKM95y/j0qwlG8gDw4V+AUMHmq
nlUU13iqvAfUfRQhyZtVWHVSlE7VVSzDyhu9fyg67qhQNXa5SaiH8jGtUVwsznYo9wk5JtJpEHbf
R3TIzK0VCEmYZ0DrGevIezlkM9IivZ9QO45vJ+0i9v+jS1CZJNPFnmN/8OubvTzEYOm7a5HE87w7
nWYAzkUTr/ra34PwArRyeHFkBtDhuUZXGVn6nfqIabI5I7sYu/KR6gHK10J6s+zYquVQENxnGBeK
B4CaNDaFthWX8868tlj4xUxCv4INv4B55qqAodzhZrEqKyEVlIJJ/q0huWxwl3znyCY3OFy+v0E/
oNP/RidgIjbHQqJujsb3R19uVe059eeCCCIf57EcWPYU5CBf3E9rgXkEDPPcdNglbxjXSC91RaRz
lPq3fcwf1aervzyNmetV5VXsqYxZZfZsZ0+MUPiHjqVKaSsTO0VNxafCHVZifmnl8CW+GlW0O7Qk
5gzwXYGlvps8oLNG7iov/UOP9nDMpAXLuQpWlZ1LUmJ0h+lfCQL5bZMS02CeQ8ND91iwO8LRX2XC
N2U31c8PI0xIEyWDo8vHlaCHo/XKHM0B5ecksXUsARYFkADtFQKB4SOU2eGTHhOjKb2JW3ZkJJpa
hHd1tyPNUvcurWniXaAMILCahTx7t0DhuvtUjf+AMX88h6ksXflyxM02EGRulJ0XcaJWdA1Mwji7
QWEs0RL+ttlGWwquwo1DjOf0y4eW78yQTMfvG4PqVMEl3V40W7dHphpF5MjbnjcvDBv66fFppdqw
MhgWXE3y/aKJ0F+zBhl2qKe+qkcGHlid0UUR0SmTmzXm+pNzzPkaPABfqX6rqCWvZN9oiLtrYoqR
LcMfd9JVRUxbC26Z6jN6cQ2aasw68APOyzDAK533U6w+eUoKdRS0cRLwvdpl546HebydnUQvEQUJ
AfjPU4JlGyXbrOZ8bPF6yJBfzKAgxXO09to8ePoGQRy0L1xmRBckgi1g1wp7DwFqkWiSFdpgOyxI
ChkjDmaWxcfQ5mQruoo7IG3YTUhqR0Ewb3lhrdep3yewubHxOV5A1g1rNMo+jS/O/f/nVxhEvq6f
egUCD3vcdkpPSdi7/LEC7kfBUmAYLtDpOGxfAFq+3jzhIno8ZSdWKCRhGJdZ091iCpGqF2dIBOaI
R0BWBvSLEUWHcwvR1PW6KM88uC7jUkYKeDs/tFdvzUql2av7pho5NEAPqWvoirNSM7dk10SlppLK
YlkzPBPPvcVHSyXaHuOWUlSBUAYeWxphiTGRVjooI0QKo6gDZKDikV+AnkdGAk+tI63QuGXGahEE
uNSK+Qpe7+1F+kND8/A76c5YJCFBwja6pf8jGJZIjyswXjY2o+x4G9m2AplskrkwG0i+booxoYix
+hPA6oKfnGvT8TKeVX4+YS/kTE23I+AJVT8rV3A9BSJikvOmw6Se5jGFya7BaQF6z3LFF2hPM83C
SXniDIkoDP2hcHU3J8cpGeWcaaTm+C8V7OVZIzpMyEjTXQweuzb8Bjr5fblTZvOlU3trw23MI9u9
6fI6KkJYO9WLTa9D+akeareptQK9T9A7Xh13FH7Y05eps7T1SbgnNcgnn9a1TTpO7CIL5ZbQJSIS
yJvyl16Qusj71vFz3m3KhQvi/hQI5k44bmcVCv1fsgAGDABXaYuS8fulPD20N86Yo6fhz4M1HB6Z
EfcTfw4AGfFzgXuZtmZBI8VkJQhOiYnLCrrzZkp76XIv2nzKsu0pGHi/uj8uKapHguTNn13I054m
cWpP9gcWvhYMbCR+5PZviAnvbOZG43o5e/SjikpXMs1Oxu6zrQciYsMaPks6IhO6/46hOU5pIGVn
C/syrOOu7B0dJxVsRgUkJjyB0gig0pY4jxqt2UhCq9+5rBlOOHKsEDlRhhJYaMe6+yGq6mtaYEcn
2KdkzOxjdiVpFqfKFGOo5/WQdbayGs8Ju+upReX5DFwfFxPlr5E3MEj7HYQ+aeiniW5ZyPoAfve8
zZatz6jpW3acvjkQi33IBlf1FzgiW+IA604ms+lLA4pTUD9ev7CCfNlgB6g9j6a2wSNJDCw37rb3
EAnSV0Ir6cN9vtC5AivoPS4ugpvXGJnREfj3NTrrevI1czeP2Oza4j9GWVn9mDsW4S5BtI4/5h+d
wEj6kpxm5+hFbkXl5fxCnDaiPi9RDJhC+eECQtZKHzn8dD+3pK1OoPRBRQuFzhQqfC/yKEBI8N6x
yjcwz8JtmIPmpph8eK9awiU3a5eBqoDDbNjz80uaXaIHVgzesNyzzvZozd47FdC/R6e/F+K11PcI
eBx8td/hORm05Bz3Kb7W7cakWp3pwp03zJYUvTmVIIyFP0FCp7MsTXIdbG0TH030Cb+kHKGD/+Ii
EyWlOvFtvzTdXdl7mXyW66/MIj+9cXgkn0q964xRQuUI8sghoRwAxmTkZow/qVS/6SDMZ1stHB0B
FqFwfG7PZjsMUBZ1EFmi57U2C0OIKqRmqEPsEzu148uvSJSGFUYGl+kiq/HL4mSLsIlYcWR5/a8K
dkmxS8nmiHxiyUCTAnyZsuqNsyZXJ97rVt6jZqSjis2KWCyomP2PipuS6id7umbS/Cuf7+M+pqGh
/9jcLgsGB++WJiymHC71sKjJQg4N01it6CuUhY6H0FuaRiKNpBCGfPrg5VwJACheQsQ/VFftRf/0
e4gYE4v602UXY4TE4VvnLfPxm7H/TXAoP9b7y139CNmkdkTSCQEvvz7xA6J+qkUENE/9UOGX/Tym
u3wkDqGGVnv1WwrD70eAjRFanoxCzg+kjJZjfgAuqWBx7ZGXfk21xblz/kywxP8XhRFmpPBCBEX9
NyowIB6lVBcJ6Kp1jzsZMbxzajZnLm0XgptzdfSPlmV1NeB4sIcupy/VOgv7jRZ7b/aFTd5RdDJc
Fted9sU/DmkzvTDFhe8Kr960gJtgTFIInu/FL3Yb8uBGEYyRjlsrPVlrPKANHvwJH3CCUgqtcO99
GdX/DlAtFKMorDkVbFLxuwddwnkt7EcFr6ywVfTDqyrm0oHrO9wc5nhvTwHJriiCdSMmXBAiveCK
j8v7NC8fXJ/G7T7/BX9lmj+3481JCDVKNxkC9SwAXEy2WX43EzqyX6XQnEABmi3yfaqQgWxHXCdi
IbA9I8zGH1JDFpLdzmYjuyApm/OCqFHgMgB3a4jMWHWOg8zBkS0HfjaimfP3U4uHZtA1LnHL9xWi
5YDIB6UBmOx2zS/jLzk5Vg0c6qLV4JB2in/vuB5alqizXDajkhVyOOlUY2itQmAQ4CGN5t7amzvp
qLC6e+2eSdvm6V+BI9sbpcVVpJKVrO1cVDcyUqppE97kZz6tPlGuIG1A7+D78PeaM/c1lxvQhmNZ
u+svgyy09CnhYxtLx9eUlNln8jVrGVhG4baFteIRJntd1EpWvaJZJLP5rEvRIgr+gKTIBJ+Zdj8c
IWzu/JBggG6+285TcZ4YpWoozrNoR7G3xdhGKcq/5MVzO3LlEXEBjaaNFbOFRmlzdV42W56du+u7
Y9m56qG/7cRPXzk5J0HHxohS3CqMHyK2F3pFEIFpDwgfW9NdvHhM8c1c6ec6OeIhXcBkNAPmPDLs
GTTuL4+EVrVaCMkz/UiqgKWu3g+42UUgj6vEWZL1NE6zs7f3sM3hXQggX5+p+hPhcCejODTRHBfM
kErgVsuDFWiMoCLyaVv8av88n4NfL49AJFI+NgfjF1Y4he2iBKG4d4GVrVspFaD7sjcHfUuxooFJ
jjwZeStFcqbnM1Wy7TNOKgbUWec5QipbOysv3k0SWVwwWii7At9ZIM4V6hkwrnzvUeqqgpPpAHOR
wVog6VxE28jfLd+az8KIpcdhONz5icatQCJNikk2BkLZOzgtDBFTce6Z5B6RWye+vQpoMgF67ol7
BVjvMgpIAdC/Fah57oMWt45g457f6pqcJwrKiCFUBNcyBhwcnZCUSqMBNVRmsibpOD7VumPXzrp3
egKHB0R2MilyM3QUUuoClANdul2lBLAUDT1ZlX1aEZSqgr0pXEJsw72PA92gJvNbyQ8lkeqvNd2R
qehZ0pfr+KNn902s6cTE6Jw2xbufOHpajpD41mEXxpvwi48Q56RsBRpzYxX/lTClVEccfEOTj9IW
cSAY7GRvW0ZehkHCGbs5MboTj30lVDjHTEvzrH3TygyDDKma4PChSeMfCRsR3edCknv4gST0HR9C
0GuTaF9dugXoo09uB8btfB9cKkls/yvEG1HXiDH7Up9R6iwscoMdp3oqLVzD+sdv0Zg2CQQmFYkU
TGkaIlitzCh+cBEaRT1+u9u7WsB8tRQeU+00F9g8dXoN7yIm2M8StG1kemy0hLHE3sKDFPHkXSoq
HN+oHlrjb4IdzQfqpJu4jcGj6EjV4W8wfw68iBhY65xAOGzoAYxDUBx70A/d4lnSKFgDyHq6GL7b
oL077J8XMktPy7fbeZmWB3xrs0ictD17rQH8xeU/4kVWH98VTu18BHd9FxEgpuV/O/DwT2qu3OXV
nYjwpt2/HBMNGelFnYPyvdLSF6i750qweogXa/+9YNzzTcYeZKecgph5Xeb1QrEKTIw80CmvpqiE
PI3RKkOxWxvGxp6fKbR0+ZdXTu7lPLMiksUdMHisaF3WIo10XXHRn+NjitxsLax2p3qwUkgQupIs
5gwea6hCb/ikLRPTsR1j2hIjp9sd13YlodXev+0w8fF2XCMHj0gImzGga01b9tZj6L6DuCJpt7gb
v9utkGmTBOl07k1fFyP47/52Zj9vPcH+/VXfLCcTX6q7ztYjCSAodKNQ4sT1EoLT8CmjZc5unjb8
ttDBJ4gCxnPFy4736nIrAitxZtJNR6Sd1Eb7KcmS8GaTM8JirSK6p4FF8O242czdP2W/nYJG2SJi
Xci7k9q3mBnq1fl0/o6TQrF8jREcyDyIxW7BfRjcrxdaqs6FogVkSgwMBtwwbjIO0WcWqrv0V+uP
e9kc8YwS6YyTMAVOMqex+l4FHnn5X8IjK52J/oXowU50lZHm5KEratuHlbgrxwQGp79g6ZbPK/BH
xlsd9hCawitv2MV2TUwmxn8UGwb3Z5VIG5c03vCJxelXosux/dgww1YHka1sv760lG1MK2AORuxL
/riLA6cObNkGztStvUIAY4C5CGYm3xydDXMchLzAd96at4A4hwrbGw76L9CFDRaq2JaYciUOkI4A
mPad5M3MojXaVO+niGlvzSEBj4zVsEv+23dvaTFnxbxS14uOBpZmj9vs6DrBRqUTbkshqDNNe3ut
xgazN2jlNt9BqrcqFwaY/yI7fmdO8Gc1jmnCA8UEVchGCFTFUKU/1LgWtg4LWtOS6hNhbOcIXFEG
C1QJZUq5ZoI3E7uKbbGA57pQNoAqfIj2CWbpkPtrlXGz/mGu/Os/YkVOshAgC7leaVLp+2Trtql8
52m6sa8ig+240Nliv/R0hQuVyI1DYuhWmzxMN5QFXISLyNcAl7YG2O34xkMpJ5IEExv9PwIYOTRE
eG98XKpML3H34TWOJ6WdWI+azTB+Qz1QCxr9j607X9MbV4t4lBTzeJSL+cHeZbUaEUzeUCeGwwDP
Ac1pA8DOxgjlfo345sRUCmelj++b3zLMv4nwQ9PdR4hFVaf74qv+SL2t8uMijsRaMZu0dD+6Gntr
YjfkWWhWN/5GIx6gQVsTwroGOTd3Br3/Ss/ur9dq8v1rMXvmUGnzb+Emy5stfm+zAxMz21X+AhJf
RWFptYLoZSc+UTBaqvBrTMeK8RU3vqKcLa1kKVPnxwBJC0HRntPhW9V4ofL8wangYdBp20VNxgi0
kc+FL6zCinX2jg2D4DHiUprf34e7RCCEbZxK1r24HN0GoP06kw673W+EX84TPm/WamGamagUTkoE
yB742AhXDG220RECEsESFxDxR9xpemEhf3RspEFeu56VSIkYU5JKK9u0bFlhzcgZKJ8WsCD24wPv
VS4oKw//43Q4LHEC3kTvYiF9+CfianukzLtBVkZeRSjj3kKUMpPwh3Sh0KBIKtK33LiGRfoviNjR
F75+77h21UPOWnG+BIj+Ca/D4JLIfEdUhjjtIRC1tIn+UuTHcUKar5xzL+A9r4pYXQYDiUC+lPNk
YHF+xzP7XIZv1kNZAPcdzU6/v+njuGhquhw8DruKZ9C6E0Z8Cur0iolYYYAgVVxQ72boZeGJU4Ge
avZvUw4QvvVaUcos5NtjJjSQ5nAIUKl+NVMoQt035nZXaHLc45fnOhqC7E6cUzBpYIR6l2l2yUN9
aNssJvHJmB/BYsmuYzc7469/zmRreRScKRtBXKmuAeqp3/SUWwN73jzsy1kcYyOt9BFXzT8sEmfe
X58qOjDi3+WQw2IHaKl1hptw4nsgV/Oy/5UfarW8r39vhY9XHl19fiMhDAcgRjE2Zy5di4fek35j
HOIh78Zj7Q1MwJ1z+ay+TPzF5ZK4TYCqfIYl3oH8wmqFO6f7TGt/zKZPIPeDQdo69OhLEL2s4sew
DdPBBqozj8DQX03omVAh+HUc9b0EUgYE5x8rhL9Pp4AF2KU8DwFbtv6nrcuowqMqfP+gQBxiUOiL
jV3N4DlN0C9XQLlJLQTX2GaljUQHNxeWHjSZH7MGREGTboMBOl6GgMNqtFv/GIWb1Q+RYnH0G4TL
+8BXaZRlQceyBuEAyU6u+dHRK5g+04aJOdhFdQaY4qlRvVK9ay3mFV1HH/0F0sMIaI3QlQx3NaBh
6tSAybs1A+O4fsrdkMvg8ri5XUjK302Jp434q2Amqvupf4gmw6eZVAs/6YkkazRVNSxNBRDCeDp8
2SZ6iDqLw5fsp2Txijg59fgEoJkwE2Ge/OzriKI4BXkeoDh8KdpYvyskw9gAEYvdiYhBqSsTQCKI
qF1axw6m8ae0TpdEkvjtpVYijx8Vrqlp/lzhSqchHdZ409sEmPvgfPGcBiWbB8zT2dXDBbutPYtP
8wn1nbN5TySRwQ1L1kdYR3uv4bDFt0w65A7YDNcsYDvlB4c0iXZyffNKjI3v9WjNRIoe13kKbOc+
0M580l8oZKGI5zyUn0fUKNXzQyKYaRwdQdO++2wmRWFI8JLgmvrwskqD2eybvG7eSNbnET926MlG
WM7WjnN0IFrJIvpWhSbRbbM6D/reCpN6l1vV6E+4h6T9B7rgFTfJ8Aenozq0wcYIOIvLxLgkyxhz
unP7eB4+lcsQjyLK9BhASh3hNqm7mo3MsjEteyF8rUXAh9fgkLEC6RuY5d5duJI+p62qnR3+928z
UiSVOdHsLJ0WHbk3JHHzn/D8uGcR0RugmjqFwAIyE5nnDpO/UOEr0ebmwNXx/A7MqdfkSu0UkCOq
TZAcBnZbTA61eGVnjcqF89QPIYDDBcRGDD6AL1dl9NfQlAGGjRp+Meoy93Qr8pNa86RTSFI6hmrQ
lwckVWROpARSqklnGu899uT9RSfnC2LmXZhsBsrWJLTl8dbIhQtVF655InBg1gFAsRAhdvtZ4K+K
xRsePvXhGjG+uv7G2obt7jjVXeK4UJp47+j1/VApZeh47xGbOKuuJz9DEm4/1hMBAFRuyxnYJRrm
83iB9I1mNjtHLimMnMmIW954j+2MQiV4vCslo3U7MZDSzv1VUkPycMPmgO4/IEDHOVqIJqrBtpq2
rGe4fmouG7d/ibsNNV3fXPd5OmHZ2Hs39bMNySEsvsUhS2HBn3t7bj21UKu71h6uwCJLIjLr1KuS
/JamSdhnq3lByWrVkkEGrkTHbTkhOQWpEeUofNWJgbZGJc3Jz/PI2pdLSeTd2OFwhgdKNSutUr0R
RG6CD8pA+ddbOuJdEB8VNdqfYW9jbUMte7UnGytJTv6drv/7fxCW2TUlSb9H23yxUP0vwbXsrWb2
xLltirJDeCLq/a+JNGj7Wavg+srLiIpd616+gxotZ9i76Oz94aTgZf1NXIEJBlk5FjzFNMkxWU/c
A9isTe12PCyZ6bx5o0q+IzdKB5/EZal61arZCHBn14VHkXQB/aHPgOm9p7UwmiqBWYX+w093sWzk
iqaQTAZRuqO7XcVxK1+it5Ey8k38p1KO8pNDTAfKFz6Ax/ct02DX+kYj3pVZk5DN85g2Vz3ZMuzI
Es0203OEmeja14HXu3ACxalSiyddbRVaW+xUdt0HFvs75tfgrUzwS22kgQBULegDA0uvCgDdlmL4
xgQl6nCtNdvGb7ET++K9gfsUMcf6GyGGJp+EM9qb+iG3LYoukNKW4TC9b1wEwAe6cvDbnczxY9by
p5GDOKFt88Qq2Qf4fcZ5D+PUuuMXJC/XOGUsypm/XFwQeEyVlfWdQ9BDDL33EVV3qMvc5fkB1oWO
a0qzo8qHnJXGZhPLd3jsXneoFaOYhbDyIN/zDQ37kL2WT/czMnCrClK2MZPrszjq1mjNCodbaUPd
FFxqcpEIhHRrcH0T2gAoyiAJ71hKp8DTgCch6Im4jUX7H7rJVI64OE0oXDsgOO0/00AmSOaJsTJA
Dm6WymRjiwZGBu4PWnwEWcHV/C4bQVADMWMuuUb0mycCMkoIwTWGXfEDajPzCvbSvdTB9wEklMkj
8kExrKV6Au5FOt0Fq9uCUE6lvXMrpD8fbjUrISvSnAR5jtnIvlq7STRfqwF1ei0vi141LYkT12NB
Mp0QFO4kEydtnJHR2gE55MU6oosVsguTGURwMtx3cLaIUpqfN+XCr16kfCFqw4f9x4GWLp9Op8Et
ZccZmIR1m6mqkwZjiIw3gRf/I05lZgU46Lx54P67AKMyFWyAD0KUtby0gVAO12iDRNrIXgPfUmhl
58VfJPlNUz5GZlhMSgME3PwNX6ZFDmydTzeH2xJcF6eURUpO23ZJKaqIogqrv16KjLhbwn1nlSdo
8zaHzcJJ2BfIirdRNZtZN1yLeu/myHeipAPFGUACU5qIG1Su+36LIirhvVVtahTZcKkRq6XKbN2x
lE/QloY25Z0/4XIoudbh82Tr98UuOoi6EKOAhRP68yGJt4fTEEEJjNxlp/gfn20cuD8qE/PdLbqm
VrXcQhtk0LgMzEsWWmXMrJHfA3XcBbuecX8ilaoqtvZXij8l/7gg8kQHhSn9zbekp1VSIzkLGVeP
Am4KiFBNmFMGV2Y1vj5btG/PvIar0wHlqhlcJ/WQjafRKXBWS6yUIl03AtsQqyXPuFxsZRj9hnny
Zine7KGauKLrZkUKJ9SbW91AZlIXnyLg8EaLT+sZxPlPeBH+vpZaLFbAOCdEgd+FM0gOlGuZWUwF
cs9LUrMR1b42yToAXfOCMQ8eYF70kOQjCgNNw5Qeb2AHdd6rOlsnd83VBZo7KGp/NQkw1typvdh9
09ZUaEbuluoaCNIzISynns5st8Bh7a9hjmA1YmMfU7sgRR3gKgIRw3PbKEzulBFbw+9npTyTbZHh
OUhcsuv9ddZ3ZLWgaEyO45NF6EiymSNWtfhrcHAsTyhu36L1M9bg2L/n0WlSZIbJ8jVG+XbJf4/J
Sk3UfJWNjYsEtvzYQrvoIY6FEg0v34Mx/p70NCRwsCgXrlFIsWajXNFhhuAH25xSTL4iMPuDALAI
ME1O3yk2QGnEIYnDR0h5lFWPzCXMmdkJO7Q5saOht6gUXcgWUoNCfZGxrFM9Gcau8E61iss1QWHN
Ug07W3oC8RR4LgJ1gI4QSz0l4SnXZCGP7vnxBDGA+SlPSpz/USTscpMlg/Rh+7NSmquzPs8rkjqg
E+MGgoBeXkkYPEb0BRDfvw18eBO+Wz3QzdSekdRSV2wLEORusufmXMPVNb/llotCWmo7BuiFO+pu
qcRA9XMijfdGNMPiLzFymdOaIzZfhX7ocJByBWcVZ81h2LUgGutMlzogNyaVQvfD+sXFpK0iOryW
tapAmbz+jhGWwYJ09S2YhRDQ407mFQfLjAiKFLXlm6z6xuLX26L3EZx51MyHuvZ/9pZIm8QmWcYK
Po8FXE7kD1og7pMgtvNUso+k+ogXWwEq3q0j9v2NlostG80nRB3IeFNgjzUqDfq2df3HvdzWOU9n
VTGUvKmNr+wzOsjYqvhJbJJhZpjWizrEBkvWx44VbPmb8Oojj753JK2zEo3k/+V+o8r99VBF+lOP
h1u8LfvHgn+P9EafB0ynzgcwFrog/wbnsVV93RQin00oUQJ8dStBul9FlKWKJ8qP5OMGrX3w/yEH
7x2yLSdysZsnxtf0LiFZt6JgN1tQxM6ZzgLy1z2oyF10fA5TKGM+mF6ZNustf1FTwqrv5x3gHEcW
CBFSsx7TyyAnxiVUZFG1cImGiiOBLGLPaPgOGLmUe3BM8pWI/n0R5eF0EYfIfWKhAA4izc8s4QGL
Z3hP+ARFi0eGkDJBWkGmuR3siUntyLjOc6Kn61DiCKTQ0oVthrBhO8Esy1s7gX6gSy0C4pInY3p7
2KR5qmwj1HaeIY+BWTonr4uMxe5SCIVULP84ADSBA2G+htMIBt4xwu1+i1BTRP3TEfQmdVKksAZ2
DznxhjWS+f7T3fycI3eyKYEjA42UaIL8+u+j5H26xzQwpcPnbYCQ2s8kx6vDh7nxQCop5nSGrtXV
pPVexmDdZvL+Q4GacwiSQ0AwsP94yyg94gfhli36wvc25clcb3U3olBGAWZXUkwjeYc/1tXCO39E
7YcFaSm/h+0an0g4eoi1iHxYJvtJWYmbXJXNz69r1UP+rak5nVuD9/5yjbP9ok/awuKXEkZvfLCM
nu5n9roncadDjOX01gGSD05jmZPgYuCp50l1IEyKsTTHd6zByVqB/1nlLwXHCv+cvLcxU36NgQEC
1HTv/+CE7SputGeXnWQFpgl2deXjOJICDE8RsALLaO4AMkiPbiMiREbYlddfX6JaIlETFcpbD7Zt
cJbds//f+amIzhMrrxaW5V9plYutsv1TK5FLClNasuAMw1shcwHZjP2hfXZ7xBRszgO/uJGZIx5a
y7K/e8Zaom2aNFa4rtzrt+eAE+3VtkC1g/eAwF19XEYeF2dSDkSHItpVS2onpP7ty9qI8NKRVQ7T
RDtKgyGjdUlg/Xx/nRtP0ahz3StEhTuEu7n/sCinL+rWj732PM8fghLQR/8ysYL5B0Ui29kEJ+id
cPZjvVdhz+R4ImxOMT+HwetM00LcRA86d3MPjyOY53BszhLanlORMIfkx/+fSgi0PlZSbF60Z7X2
19PtqaNzdGIyeOLxy9lB/KEwXG1+tr/zCwm7HlsLFQnbJ6bXyt93QygwgBP6dVhUobmqb8FPKYOg
psWSHTQkKDWNlsFA8tX/8IJ8yajf1dnHakJJqPlP4wA+JBj2/IaoahNST17YPs7I601xJvgSHTFP
z2fBJf8N2ezuobmEb5GlgKDCfG7dytgSQ/PLfdP6jF7sN0dUzi4lIZI4z9GrJ45ZY4PE/I7mmQVo
X11jeOz94mMGhlINQeVkBrcd/4iC35tTet/wsZo3TRFLWLhlIdkwWUIPeBHGaXf01FIbDyOYeo5c
z8XbJSkhM4VBw3Oz63ysChulhPYpJDc/rijXh3+ACQWGszAt8RR40/yzStmWJEgniJaYlRmdNK/v
fWdC4R0aX6CvvbGfH1jA8FTRE8XAL2EH3IZmi0fNXPNqYpGI3KTZ7fzpSnOzPhLZpBdgBYj2qwx9
0Y75cnZejLvlCVwdPR5meN/UKq5asr0Q+JHzPlBEONkjoRz+EgRJrX2SZ14mofUxkycGowvL84pM
iNJU4bVEWrz7D16Ub2U5fZ+XB6AQnmO3Hm8gEWsuhIcfvOpU5ZJmQllkpJUT9WF1mLm2ZrKcYpXT
ELNMukcJbRbTxyx0fp/wKcmv7nDVAUgBZX26ed6uYPzAMeR4COzZYcJtQfAdM4V6MRs4RsNeFH2t
TLVHOD6FzW7gvRf1vMneKBUj/ru8JmeCWxGTlOCQ/1RA7Ij80BpM0fl3z7mA4br+e/Ei+6rFR/gh
NGi1mMKe7rkgNfoShSxPlqj5fg7aapWnrfHTggtNMHWzCfKlMpk5z+p1Kw0vRYigvoMNVQasccSo
DSdL2BwucKPKsYIyKZV7OH6IsS8dJ1YHfyTtmjaHRZQJqnsOgZUWClXg7rpdI6BcDmgrQE96TMs3
5PtA1AjXMR1fpWzk1pOfOmtDFNYBTSezF1quzKL0Vu1i09zXuzTo2s6rnsIRJj8TAwyUL3Y0GmO2
Ra+PnTph1wWeXPkh3qtDM9zPxoDY2g2kJGX3iCpUz/b0JXjX4+XmhM6zQsfVwiDZHhsMt8gn7QRw
qRe2lVo+q79AMNJHyi+a5TPV+fM3HHv8CngwxjKt+vR/BIgmvErcEujEnmRfTa70il9fgqDnnD1w
Vgr8sx42KCGmgbsJXCAmVs6AWkbihIQryqIM61+VgKSYWZ5J9MJ12/rxCyqu/CHH71OiA4vGoeoi
dPlgm9PBWzREogI5Luye2Kdv0DLA9qaoTqgsLnoXVcGspKUZJxkWLB5oGY7Lujn7KcRbgtCuSbzu
+5zOFHo/UL3DCB1MK6hV2II0Yo0C7LxJ2bJw3vUnCznhAeh/q39bABplH9YUz1DNP9N3k11o5td0
5duIgQRwF/wXDc1TsGcQtxIradKdb/TQtc1hTGkKb5ixBLqnfPePtfJ+0lETWlYJ2vuvj/Y+up4O
RXl5a9n+4w/i6UbG/e5vhpaqpXfClzL7R9GOGku8demdQ3raVpGEGVbjeFZKxzWbzRerE70XfsX1
NCCVJbfSRcA8WyjcoZ5a1xkqo3cqBCia2G1rhE9sL871aFOBR7Mf+tFhO+2qut+KY4jpZodPoky5
neTEZmD8Aw+5fx/3ZTbv/AndDdqopApcD12Vynulbby3S3F+cxWkDMA7ij9ef0d6iWAt6iu0jaPK
ikYc48DxLOYsIcrQsY/WtHa/uUW/dDSAfOXepHOJXOsHYAO6kt58Wzrix4jtO3F2MAbgjM8nl2ti
vACpoTl6iCwsXtb8HXHzVi8A4lPysul03I4zIQGE+8RUtSPaZOWQRUmN93KSzH0bjAoW5MJM2D5W
TUl36r/+dJv6d4+Q/MTjhorBG7urIq2zEmAfzy0jE98cLVJWXg5RZlvyzcpghaBMAqOkRYd6aqFC
jhWR0LRjc1h8iP4wyJQzOl0nkqB9fNpAPZN6vH74lP+shJtis3U3my7IyBIhDeMlYheWTMKiXcVo
cYzj3jINcRNw2aiemRL9/6YCKiDBsj5yhEf8Lb5tSbeAS3n0X5Lt8BxoFqmTazCIM50R8uhRe0hv
jlPg3yXOxKmIuKJtKRuHXlV07ZjwJ7PI5A4IHcF1ViwjvHb8jCzuGYzdX745optPaCduNZ2roJsK
k7cBhv6TEC9JYgxaz5gspWRSkLi0FBpAE5w3Gdn/CSOivTT1Clc5eKSYMUW5Ne0KivwDkZSrhFmN
cD/ncT7vqqcVkzMLWFZOuJGSKHGgmJ42Qj36hm3E+iWiyuE/NmaPtSlOQgfWwoLpaAZP8/6z9WMK
NyZfUH9sNYSlF2w6fESN4zbhVmJuQDszB+Q+5xTZRDzyBk1HrCAVVjuEJ57hVyT30hCIFGW6e8MJ
/UO/PWYlGFUMcRkiBJJk0MlZExWy1/m4GO6lhyuQubvlb9ypsBCXNpAbSpTcrfua7yb3fqGSw7Gq
AAIxB8DveCmnCPQw8bBXnn1amLcmYtfcWu5rMKIbqv6HnxvTLPKyVdlglZGvgqIMoxg+0SdM7z/W
EGA7PkDsKFVIbReYigO6+5lK6rQXW3sZNf+SbuFK6TQ/hRqtn1KgwmHw3o8egzn9kYd+aHYseg6/
x/2RAafBdYysA8+VWPES9vUBYDgBBKN/vrYkABDA4y6u7feVdk5jxXsW7Chj2iWIWW2pacPknZgc
viBXJJaPeIwEc48knMUcXUqPk4XpRQcBJrMNm8YuPKlqjCemBS6xOhSzxxjSy/lcUgg8OHX1cliX
xfIXq81A3gM3baZy+v+ATDsa+fUMHKLHGmAZU3iuqqpebzZbxGYXjIckPkGz2qLvLhZgSFTVnnaQ
srV1PKAhrO1FHacmT1uUk75Fb4rVnJfMwhDXaBvatz4m3cKcTGhXWgPNkn64yDULVGs6qafrd9ls
hoQz7g6JKkqMIEgj9RB44iaKHdoxr9irCSMiYembH7xEihi8V8TPNi49LfJAiIbALtDnMe+FhExD
Dt1/4V3Cg6xx5+bue0AJ+TOYhoNF8PwVT3lPMG9RJZQsUsFFvaueIn5ZyRaJH52SWwPBhqIcDZgQ
R8PpqyFKKUrVVhSbIKmHCc0dTRRe18vjE2UQB1bcWKgkRCKA0ErJQEkduXXH5hmJC8lazUkXgqN1
NIO69ThtvPynEfrO3QGasjWHC3QVjAJpswXTfrnJdYWZMt82xrSnGkkelg0v4zvNQuOuOQ4wxaz3
zC30TSqlYhxU+m8F/bDoTtHx5ZeQUftUWmhHPY9I8B8Psrnf1JImDq/0/SA7qZWfU8XkdGlQkG82
5T45GKy9Y4k2nXbTMgOgKu1W5kwC/U3OctRXUHPl8APhE5XNZQUuLWTVKF7rNHmrYb93qN9+z3Yq
QO+IRTJEY3QOoqEkyUIavKOcEgCHwwoCq8hFQ5wNu77siXS9WuaqFcLwzBlrlQEfl3zKdoralVRu
U5ptnG3iGBEIfBiXrmez4SjUgGFuEP7Z/IvmbFsc7clsMCFE4ga3kngz4X5MNwEQDwDJJvb3TAJa
dUy25129R3HGBIUox5RXQ45vVGUTMXg5t4nuIxEaTzUlfbB0DW88FPDKYYgkwBl3qvWZlBFaYGiW
ZF37P3ax+RiFmDz6qEhrenpTnva4Oi/HVTb24f4JdeKaZ1wclwbgSbYjiy7ASqfcHkLUXvNp46ud
26QsKyivN/RSB1KSlmG2/mrBtZnPCKy9ZJ+iYSRguRMxQieRsDYlOQPgQe/sovAr6pjCt6wOYC0C
IYzSxJN8Mo38G7zR01ntnwuOEc2RHHUvO4PrJrPDjHwlS7PDBtZ4A4X2KDcRjUGne87Wd5NsDvnZ
zKCh7TTh5EEVZOV09lWMnqnJp+1fU9fIUOp1gfu1XtMYG2P2vqE7/2+vn/sjery4w6FO7bjOWXVk
f3pm4Cg5TfMDzfwfiXQ4dI+noY/qixmsZC2CKT+3bNfDTsRaIwGbt1cWK6dZywbuMoM7WQaT5OPU
duX9PN7ypSL5N0qD8tE5J0RImB0E6gTlWl7m0t191rMOyRwQXxoQD/4K0SdmBsf/PVjX4plpLpwv
6/91z1P+k+lBNgkY5RJEVsrIff00j52Qf32A/v6+wy7K9DcohFeCaszK62JZiHtplj70Zlmb7dmB
geglviNp+58pDA+Bq+bZ5sWmdjPLKojbj+Z1O4WpL/ZGR7S0F03VSK04yyDnspbr8GHzYeRlC+pn
zjKqksZVelfP8jYyEdOPy3eZ4QmpprDhl9QT0WgQGe/RTgnjQMA9jHEjLZ/+YcPkCDg00VUU/+GO
H//kGvosYfWURJ55uT8CE5YjKbnKuU/kB2Sb73y3dYOtnVElX1meTIONWj1kDUXr+yOeyUM3zP+X
aNciO4F4tZrzCt2D6y7aWkr0YzABMd2c2RvP/WWfUy+xNuBFCjGltaorjEz9GdCLqVVQNLqUkKPy
PctN9TlYox7wIYWxP/98/E6A6x/pZbrb7NWL05INZiNHXpn6ljnoRKB7udQPTsdCrG3uUPhwjO1G
GeMrD/3kBqFgh2d5gJiVAL/cqpJZkO1fmanoXhBhEb9VO4VIIC7JfLzrj5gwBx2E+6ixglUKbmA6
2uGzaloyy6zF00CQYvB9pUTP+j3OLMoosNKA04MffggVxxfryGDWweXMWCTL8mS9VfaMBKI/Vdb8
wZ5KBwWcOnoQnpRIjouPHTLJFa6+p0DO27Y3GzmH51Qy57NaMr+prKIVCHE4Yc77BCxnMy7Kichq
5veC2Ioc/Z8IALdm8cPGW3vcBi00bYrErSm0fPeFcl0dkoD/I/sX+YGV0dZeFiwdPt/dY7QR8oo2
FsJt0EfN23yqrBdF3fy1Rf3xqd21+Wvdp0hwYDtqyvT3ttLNwKioX2PoLyPfPIuhUc1xODYU8OjP
g+CPDQ3L+yQh93Ae3o6Mzk9WeZhhsgHxOPyq/K5jKmYx4yBwIP00slCL4tzwB+lG01ih0KdJ7uG3
3Tngs3YNZcRVUZ5+OwhUu9lAx8u8nFOegWc99di+igDPeG+kYVyo/hMqVOCTyUwf4Na85C3Z4JKU
W7jQkJZMBwqKDm80Lo5+y96c+pYrLp+5V1Z8hd4Z8B9xYvmPHYxBW3X2iNffD0XClUAYS5Axegxe
MsZP13mg8cqzexgaNNAVtGjO2sc+DWZ1iH9fK/256wRzZrBVJAu7J8kvR+oVp/2dhDmrw2LWhABE
75L8og7igvV8duTt1p4D3pB+XYqyKyiKrnsP9q/NpspcTTCwna2BBNY2Hk+fZpVyJxyPYxSH9Nrd
QmTbV0F+KH1YRLVCtXPDARPnVT678a3kqyCZayZq012wL1sNhmTWTGV5KwR3F67cMFQ9NGisaZ2l
KwIUD+sZj2eYwvZnP7iYuz1rk5lIViWLWwhJluOtHnDrmJ2INAPnzYhWKNQz3cns3WXZwiMt4afh
scREjJkqKy5t+AxbImXDogTjo4v7wuVY60gn9BOgAkwFTjLJAVSKlPTOnHqbm7O/QDtGuKj4oyBg
W1tKiNN/FwB0xSp2b/1GAuHc7RzYiPJFAiqaTOqVSu4T9wdpOFWvV5BSrLiu+gseOKNknYIO8Fn/
PjXC7Bem260vSj6UXTdKTdaVmPphxAeFTGrPPFr5u3x/SVKZr6njsqyKJJhJt3pCgVlApnc1nwh5
CQwbmgiWABSIGBXq2kciqzEiPdvsLVwE+xXWh7cRjU8RykgokYPg3Hx1Dtc07BLN4tIh6YCBgTOH
wmyddMIrvntdmp2c1C1Dy/0vjw+UWNocr/RPDFrOHTZMmO7bMBFRMcAkTqqSwcgfcjOQs4fTwdKK
MtkCnwFI/YWXtM5kQq7DnxxUerr2QHjhYJ11/zNndolfh0STFmX54iJTZxUGGnagtHe0vDzA8ETX
z4qJg3/Ij0JpebuHKqeayhFnSvEC/YStPPEBRz41yo5S/jPYHI13LHOPM4U/9Q5wUbuBhZROtNKZ
xUE/LOEeoORhu/kKwCZIKTmJB7ulb6Ujizuj9JBJ5OGLHo3vX/gw94ckH9BzlQmkAinkr6xu4hXc
lYXwP8OcgR095067ldTQVwksd2dunIRKCtMgN08E5TiPuCii/JFYmhFCkY/H0QWjLa8UkezqpO8K
fxEZf7zewE7jB1LFjC1KxQd+nLTBA3XZCtcbP3ei/rM+tbMhuurIrXotsKZnE2fsx2MM4SjUn9NG
fjWTV67gXEvyy/IL1h+Nhwe/o8cC0kAWA3rHYRy5aGV6DPeYUGjZTTHZjdGUnYX2SNsv9w8X+9EO
Ss07BUWmZCiX/w9xJrC7tqx3JwcE7C30sTW/pROfxd/5uaa1zmFl7mFmgJ8TPXWqavC4mACZFukH
61tOv4bWrq/PrnvNY8EUGA9Rp23XnQ3eEggkD+7SMp8cjNBAGGQFE9oWl4fw/HseOEXgi1BqgLz8
C7CFvPwGw6Y6MNXcP1wGBWosSSoLkS+TXTw4Rnwpospch9p9VDwXU5YgcjLohv5NO7d+5pu3imPB
RHumFSou1F4pMYmDXMa6X7KwR7z8PBkZU8csCCgIGGrgI6fqemHKyAWobH40Ws2FlOhgvj/+s2ju
rM+a1uLrBKB3xKrA5nJjRfRS07Ljs6c6Y245zZ8rKLScJYQb0qYFgj/FirMHaOaU1l8joOkaCLRE
Uh1lSvAx4AEaFM6yAxhzkQmpkt6Yk4+CEDW3AWHZHMUzhZxjVWRvajvWPO9h5tEw/pt15Wn4hLx7
cD4MyymXYBKMvXu9xPPR+Z5uaUsiIW3HHDWj/4GdshBds71J+ManurIOsJDILxqwYwsw7exNIsnr
HpmwnUhcOs4O/6J8iLmJq4sFBzff+xTqMfH3ZaaVwGndSyFC6DaQRk9XaTy3thqZO0bKmXg0LDVF
W44z64ujwfB4zvIlxlgoB0jsJbiIKQfDxtO9OCQkEQ5kpWYaAhwBR+Lb3eAJ0XYSpMrevQo0hV4u
X6TrcSMcmvlWFMKxUWax7k32BUoLCeKp59H0QCcTszY1mHebwRde1NKMvhh4/O5nQRG2e1COPjJM
17SI601kdlKw5Ol1k8nalWUZjzLVMTVRXFlSS+moGuDtXT+WAHnE65K/NyFTbHEpK6C+WwiQScOT
SHPgIT3/jTliLb/6vaH8FtU25GaVT+uEAOlsLra0GSWdWZw5jdn+VhJpiAfLCyTDfWFqaA1xOXem
2CKYKDnWVJi0OsxN5Km7To/5Ni549JvtSZXLW4OFVcABs/aly7S6Ia/QiYo6/swUy3fB29HWnm4c
G/zB0aOE1a3ksjkdXmtCudYqmzQkfN7tecWGLwbNUAS6PAv/ys+F/rdKa3QOPT2jO8H2TTgHqctH
l0gc5K3XHAyTiNP9XzhH9asfJWZfR5D+XNz++r5IIgjLD94ibNwp3CXfK5vxwgHn9dYnaFvwvK1I
rVNfM5lr23D7mpEew+6hV+uOn4KS8HZdH7iritNbz017w9x1d3VExl/Wdsl+YFwnmghFxSLMKjga
ChoQI3iuG1p+r+WeILWzs1SaFr0IYRA9Zyw3EYMEUrugGuf5G8EjyPlTEXxpanhiwiQBJGqpiwrc
EXkcPyplh+/v0ufKo5YUGi2R3JAbiqkY1G+5x4IzYr9XznmiJSCv4e1bgO1zWkvjNFSrCgKma52q
Y/oe7y7+A62Qhq4Vh4IQmvjWYZuwCbYe/mXrg5xfrHXU3d78RoPY7zM5OBC/kdP6OO4J9dRYVtM1
3oQ6dCqxrNWyxwOqUlPqoxxhq34CmXe3BCgs8gtvU7LC1z3IVErr0JSepabz0OqclwzjtySxkmxD
Z6DbxjAGb070Va/yX9TR5pjsumZStSJCic1t1wWKO9zvv5wMmPT9y9vChm0ut/wPhXeJ7qUSrvaD
ggyl4cUAj9incPyKCtjLuF3bc1Xfeti/S/iermJ/JnMcxVtAHYlHOuCj2XFVZq6oIepqaag8JM4Q
hRFQbu4XTgJviguZH6DNRUdSejRfb+vcEUlaFeTiA2znTANcOW2mGfsGfDfEUfV7tjrGRQL2ZW8A
8DjNOmACTEGcjXy0wEgQVG6DTC4X1cL2QnUEo5UswMTYxJtTseYz9RURhoCStUV0R/vm2fIs7lSc
k9t2jio+xzifRQuTRw1NegLC93T9I57tblhgJIPQVfd+k9ngO3EIkinKP9p5+sFpweLWsh55U0lz
gMZywnPWn+QQvYpDJGHwyV3CrBnEDzXSBf0oj6bR4qFxL/u7PyqxkhrpRPv/DukodHNP3lGzMWsR
TqkzWDdv5sZcWgfNGOw67f1u81fx2RJA2kZzmw69cze97TdA1UcHtnlyghYva8nTw8oBdIR7qjYw
8T5+TYzRu6AqefJZQ/QNNwYY9GoXil1k3x94kG6PlAM1FetCUdm2gHtLWpZQaUQD0bysEPYi/VjS
72iMxeKGcU8vekXxlhNgjxSQGmM3Lkkl0eLI8PvIx2dAZQveSNL8ionC2z9wiaNnLUeB34MD/2DF
7Zuf1WNiRqa8Pni//W+iTkI0KOz6PJ7VPbSIjeH5Cej4LAPTpdvpdHWOGXUaOFlk0qDo9gHQKit5
P7Zp8+IpuVM8Sg7o8ZEWjSzfONr6EZRJjqZK+MNKS2Z8xZ8hThlr4Tldc4FoZgqP7iiKifPcr3tC
s9FpkRhgTfHaLT3FYW5fX9Kp/+8Kd8UYkz20ZFzXA7e4lhQAcTAcId1U7wz2LZEYY6WLTCJpqx3Q
bT0dnjvSjSPqkfqib+LQFVQKvXBTuj1BOObpkLnfdg2Aq6YWswo+Skq3SA2HjmjR800/ECW4sxA6
F4MYHGL1C+JU9W8lhRQdUUUznUccbVgT8GP9QpRkz3Ma4YMa/22QM3i/yM1JgxZuuWBq9ZyECJG6
q0gIvtmd7Ti63umkiL3Kaho9upFqvQ9Oud0ygaihk/eZ2eco6J59rlKWx5HykltEvAAIfkWsO3W2
804epfSTGCA90RgEKgpqKJONgC2Aw+GXHnF0OO644cNEhOSGeXM2xFTY2C7zTI1hBtXWstreLUy1
l8/ZLTBZ/12K8pHL1WBuyibTeoOkEwYumK4M0kfTTXuSXrJ+0vcbzMagChMqPIg03cHtuKNvQZmm
SGnTWQE05gweO7A+5ltAo4oJcnZMveKj7ita9sgsW26scGLwlDVEmOzp7s4rdKHQbIxMVqWozpVn
amhp0RAjQm9uGPz9CifR1QPj7J0aESTfrrSZXxn8V59UJhd2oZ7PTbtEY5fQiRwoKNnS17ksGdAG
+Wh3XC2fwaWqQlm7AuZ6OPJS6tPFOx0=
`protect end_protected
