-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
cUS+g78kdQGSP2IZhUYSV3lsMaetMvfRv+mqqmfetgd6grK3M8uKy1h3r1cKnI1q
JYsscjBvdGVFpbz73RsI0GI+2ySZmpQzOq5JSZBj3BoqW/gC2bT62MNwbBFc/0xN
+4AYBFsIzZK7m+CEXtebCE/YtF5NFdINrfhuwD447Ws=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 16508)

`protect DATA_BLOCK
H+qZ18Sb8qSYDbTs+2G0DV63lFEwp4a69cURGsGt93ZqFHST+/InyeRKmqZfhRkI
9Ixz3qCzIZBgFWa0PyAmYyFUmFQmBPwPlkO7d/ICGo5s7IJqYPZrpz688klMk7EL
OsYx8f8De5MkF3abUrfip5nFH3qDqrmlshPZ3+AJ0u6vUN1c5bPeI4AkSisHWgdk
dkxKQ8l4BDkV165F7VU93mxZFrzSzNQP7xMHuTwHzlol57SSS6Ed579nrzeoNsjM
31u5vFlaEue8u/zrjixBMXjB8AViivacojbi5+knC3YO2JrV6O3M29kxgvtl1adY
+HbJ8q0C90p4FchJEOnsrxaqVlZo4sBfSN9UBHysYZ3XHTLlp+RS0U3sdDV87t+l
w2ZZ/iy4lU38kWuozNTv6nb6qT7mT8wUsgCgrwz9LnubUy6GcU28aWIQ9njAsHT9
fXvYiws6MSA0xREt/SQCI07Zu7tzEXbH239OmsLEClcGspPwRbksdwxgBws/+P9D
VP1gof89WCquvde62dTTLIrQZ5T5RW2Dk5T/6TH1ATjn/WT05MPkV3iqdU+IrdXU
sCpjHnEVYw3AGwUHQ5fZnmPellzCEfQqjLj57v9tN2LJ1UHGUDkfd61yBb6NHOsk
8wyaEa8Bkfc4BMkvDI4UZ6eiwOEtM3GMlRidGsvlVh1KrIvLga0/5S61DSdzweLx
jcruwkc/DrBzOuHDK0J44jK9dZqKskIAOEa5Qm2Y2sc8DJjzPWjDczU1JKJb3zc9
F8TPj3mbgAGDY7csMr6Wo0ggooXEGZZWnf82/AzSH0rPWJgdw1d++2et8LHmoWj3
GzNQt9WQAipf+mdYvSIfMfmxt28DOSbtlfwciYGQqImYrseXUMEjo2FNGKfWMSzS
AnnVubpOfHoJMQWLF0uONY0yCGHwDiN9E1y4W5g87y8PuMZNjQzk/m98+ctQ+nbj
06HHSChU42JcABQ0RkflZQL3uYLnEwzQzx0VVOAu1wL+4WxV/4ZnwMlaDZzjWR7n
9vMn+cgq8JAnjEQFP0j326/QbkFacfqwBXVf8PS25HjWOoArIh17FXghLdOEu4F6
Wph1xq0Wkjsll8LSqGcV731yFtC+uDn9wk/oJwZWZ1/LK29ApOmIRgkflHHbreBp
dwpEf+aKeKpQ768eggtSTREGax64wekSd4aB8VhJFJYUcOJdpHRMpbaK3oZxNJXC
tsve4RMEaw01BkkulNa9fzQltCCbWRLko5l79+zRAviPoss64ZFYVSAY6grHIKls
YA9ZI91O8umx/sER+E7m9PFuWF5f3HEtf+F3++BcyZ8tQvmMc4esOqWCmXz0wliT
sDzdFQlwUC0wyEpcN2GQaORdtrTZ9FtNij9G4dSg5y4tUJW0qVt51cSbSvXecpIW
lPIX+x0ZX5vHYF0pTcmAeb9h7wRdPcsX1IkbFm1AidTq5wRlv+dsYiQ/hFjnfNZb
lOF1xCSr0L5AZsspoS5Vh2CEtCJ8J5JMNfDlOB9Ds/T/9RIVoYIMnCoKlSAgZFeR
JZYFO7uMH+l7I33o3tiK4EklRpwe/1/J+ovRPP5rqUdMIM9jLDVov6nU407fgp4Y
vdD5qN67I6qfs+sKQvHtNtY0T/1fkvUh9QDGrcNXkCpccO/1IU7G9v7bGVekvPnW
XtWhJu06ENRd4FFn25pCwcXilUABf61MaoxJhEK3P7d06aOOL6HcCE+CkAqxUm5i
fSB6h4zyXVvK1V4HGbBNkyftGytcm62ADc0w60WNF1w9juphp+VRY4WDqj2UAbcj
5Hd5tU3TMVgSeM78jSs2lO0s/GhXCz7YRlH/Bt9VvH01XurVFIRwgRShEZ66mnrW
m9ufZDMwG/3k6FjVf6aumx4USPswvdcpEdZe6/SFkE9Taly+jJHKagXLutHOHaQX
GXqfcWh9aB7nUF+g46mcjFt2uoSbFvyVXGCxoC7+edWCC2uRoccrtteuFQGtx0rH
bpi4zYrRAg2nOAAz1WVoUzye+iwJqVeHuo0q0ozO1+zol1qdl0867naTrWC2bd3x
z2xFQkguBa3OU5LHzoepkOvi/fbW7IDAsABgtEbomPcNEcoFApnOYfhpkt3oZt5P
s0Po271KtK2b44GNF5NFjLQmMVijV/zw32RDRXhc1nWM6MKy8CKH6yEQCSZnm7Kq
xEXTlbY2dc4QnAZQaPnfvN80UohsSviZ5e8fNzR6UQIkOrXJOGjQCntKHDK4EDaH
56rbhCpw/fUTaG820gf8hSilEPITl2GqFuhUrgWuVd1mb404viMf3abrWQOReu62
2Qo6dDmrRpo95vhcwYSylytWWW91+NOsZjye6o1zEYzjJjXbZs/7XX4FmWtRP3xw
6O69asiNp6XgT8ESeXOYz9jNHqCUWws9XjzarOrocOOZUWBySF+SC3r2UfEiPzpJ
LEnbCQDqO5z2pEZBIHWP3kePRgv3/HxyJz18HNDOijdZzTDa7PI4U4uAuNVQEEjM
Z+BVN9Y05ijn5Hn+MnbiPUS+tmeHB1Wx98YV03OZaSW5JG5/HnJErTgdLs86w/zh
ocwFz+c0iai2daGLU3MznuYkZZ3QdqAcm5pXYb7Vc6ZCJ+3rJcgmAUoI63oHVM9b
eS9EpOFAcShT21ArBd4v/ltlyhzWKnmHKiGc2Z71Js+XEl2uFaG8d4IPyOjmK2P3
XAF9IVM9+ok9HUu29JkVL4Kz/SzNqg1AMxcqGNsTLIxQp/m3U/prnUKJTi5COWhK
qoz6GocxfVQeiRa3/Kjh6tm67aZRICJlpBO0pa5wp39keJN9GT3XDtd7xM+OpVrQ
F20IpCTMo6KMKE8bgTZDuU3VKt8R9M8W8EJXYAezGtP4HTIXVhUOxUFUgsAFGHcB
9ZNobFlHdLDOfIPMqERt/HmMYDcYGaIjb5MRwI6TFjbU2BmdQwvk4Pd+KV6RSIqi
UnuGM2LmWNjYOWZQqnMb6/rIbTCou3kJ/ExAhoUAYfHuoQ7mrCvI2YFL4I6dOaAN
RrjfDixwZf6/dDxUcsfmn1OuSheyqtaQ7/ZKRNDK+/wMh+4BcEj7H4rdRBezziqq
jc4J5eWFdKmWAHCLIY6DA+O8YFi6DQY2SLsowRMWBGtZRulL1xaV9q1IcsfkhU7Z
FkBxxmQXRmgr+9yC0ulvhpgT6U1/CUiNjK83zkGJ6uMgEX+Gck/Zbg9Shpe6EcHT
QI28se1+0PbKJrZPmuCfmHAunLI6a6L5c6zecs7TcMwLljgGBf/zWxMDZFG+vz3d
xExTFZSI+/Xt83lkqa7x1ghK/0LmiVd4YcuxL9QmN3p4ABLfxzoX7tSlVoea7khO
OP+Q0wQFRRjAujzE/9rVHAxx/J6iX6RxBuKsBr8KecjdZfW7r5GhFC8IohEvo7pU
7eJPPUN7iznQ6GdV8rrBZZR/1POSG8Cu2rZ+am8Sk+gGaa0HP5e8JQALNVOg+Fqy
0mZYCSRyLeLFV1AIKlzFMCPLUgEG7uh2VS8eHz1Gn0rFQWUG1oEUElDKZPeK2B8z
AI5eA/U9MVmvNwLVZ/DbXjq265kPlzOPvSq2bop8Xh+jBJGyWLsfCDT+ANcr1Q1+
bQZLcU3w3cF4DXQgyht4PCn6VmtfN4MklAicy409s/q+fPeoiZUkbWIrxdf9A1+/
ObS28RmSXEPZivuJ6X1Qe6LR0szeokpgbIN98YZrdFFA3irl8503CWSNOTJg3DDz
JtlzWlJT0j/lJ+s9aw9PWFhwusLemlFwZni0ITxteySJmwdbT3rDis832aElRIHd
RHilQ/p1F07TJsBRg8pA/BRsIZOVs3qtPvvDuBSkl7x4qCdqGcNOATKtF/ejlmrL
EqtB3RMCU4cqQ3vw7akC7BezOWjU81kSxklZqH0tFSYSTtw0WQPvrPpCnPSUdLlZ
8TDFVozeIPBgXYCaqzmyphFiJXNrlTaKwZ+aD7dLT+yt8Vn0o2+SsZwL6YeW6eNP
x+LIAdw7h1AXxJMzj9r8U3lU0Td1QHKjnpWiVJkq+qbkulE9HqlVEXKW1QkMJ4fJ
ePDmMXQh/l2Wy2/SyUOzwa1QSKNg7+Q6TcHV6uBmWmzu3l/JiexaYcRV+WlB0euf
ZTlg/um2m3cpoKFOuOQiVVXbq8UCDmsGMjT1deN1G4QFcfHiPwgKcORKRZAK0UdF
SleQNtBxb7mInCsY1mETEATayy6USApUjnOT9NoNNpx3i6RxLuOCFYnD3YRHCu4z
dh3p8135uLx11RIlbrMyWY3mvOV66mgpguHGOlwIlsY/PMCEZqPdFULas6O3yddr
zmTnnerja0JJMp/EPJs16EtzL53xsbcmfjJcjO14fNBirAh5NWNFaGHvI6TGVD89
QoRMhEZGw26mGxG7OzaLgg3aU89CSGEulaww3W62yBTPZUMyTEe4MJyk2AAH8/Lc
Q6h89Es94FMJqWXKUpvfoIi5MbaDzXpw2PyEE4bKJ9JF5WfOnObdvrXp/bd5N/cK
cSenQJqmXSIfMpEfRFjIiNRtO1IINDbwEDMtdM9Q+olEEX6l3Jr+HIfEJ1W71CGC
ddnuS8ZmtLZqDyeuJSMrowmC3ZVUCZSBSx9665dQSPXhhta6iWAc214WL6Hfomvq
wrmoikNR10DHrC/linLA6LzYnQ5HyBPl1PuD54kB2Da7BnYnUyEWNh01bMgmeNnw
k2Gy3KCySr702M8ZY8kNNJoJrh1TUgZVgDDMDEvVWprMEZ+zMAys98TNtnuwvAAi
WmZvlTDKJ9hRpVGtkoxVjn3QJtGqwqbAOHTBAd8x8fi6cGt4T2ZIUmB0zD3swpZJ
oxgH7bMMey49QS9NuKW2tEtcrC7DhgzYFTlwAT7Bo+MRblNy2UJzP2bayxoDvhba
MtRsuxgZaI1R5j1VVXWmcosndDgQk6yqQUUxPMP3x39QgAlASOrH6pqjG1GjQSQj
H2m6J6skKhDXj4BNnEprPxkB8fRQnKFMl8NhpenSAQjeL1H+SuppIbj08tIQWxqx
Gkg2gziWCb7QMvPJqsHYe7rOe70MKApR4bD7rbyhA8cT5HmG1rGnbcI5kgpFepMj
qM1d7xQ6Z5BJLSvozkr0jxQojybOT1MYY1XXzQ/y7U+iULWSP/0ReTt1LKc68+Oy
Jcm0+WEu4uPZERJWGB+SAKWsts9GK6h9AUIDjrMImO3sqszTloDnD6SfbDM484l2
7LBQIC5MqwoMEZm1wz+9TGHiChM/GeuBO3ZPykQ7gae6qFK+PnRmYZx491UO+MUt
HPdn5ClHcJlFIYqGR1XTvw+SEKLCmtLuxeoLGqFgDsiHbfbuJY9mMh6svBvQxkJa
ADqWN62leUOtwTyjGbs/nWKNi/7PHRk6XkX4u+a0iunjUmtnsC/OKo19m9GBfdNg
BYvWfqyB0w4W8vuKrR9cnGLFowdzdbY/2lyKrXTKiGus7Rlxjnhl95sIzBYrJwdg
7mLB80XCv8TkCHLl747euyYVutAtAvx9BoocGQ9kV9BZiCtMpV4mX5Vm6nLfGm3C
8oddT7LPGe6M6qb4V0agZHg3jnErJCuoLdQvxPMyChDm8AoiAqoCu7bjkVIv2qLg
spfstviKtYIdj8kZeV3BDXeEx9DAnIukGjnWmhoH+UuHVlzwaYVp8sn9EkYjAXMC
8a5gQto5yvSvmsfcxDyvWG4jJjkTjf/Ho0fJJ2WcFrrUnNr/9NYr0feXiHcYkeiM
6rpHzF7QEpC7ZPruLk7Sru+CrpZY3+uzeyReqZ4L42TSnex0OdlVEBXG0H9KQrbE
l+YN8QhXomZA9Bql8W8fnGSEgtnEV593jcny9xzPXqwCnkkaFepXkvbd6PaE46T2
O2WMX0i3yDfBLdsPn8TRH9rpbg6+82Q9kuYjmO4qjlj0uBHPnEfbLpNNkF23s9KV
Ulg4pY/qTlRPFkrabdFmaSt9Iti2Er0G+f4kgoNGVu8i+/ekvHPmdwX53MNrS6JK
DmrP7+cE+2XhcyEIvt0DoO/ySiVSQsvX9uNRON9Nkn/5jJFA4+zi8qO78CUQyj9z
rZA9F0RkYLi4m7R58d76g2ylXgnkNPbrIzncgLaZpc9RY+N93pYSvMvqtGVq6ThC
ZGVOTJDiLTR1ZtpgGFfVSCaJT+PDxokofqcIVi2wJJH09BASXsggfISIJkFWH2TS
Gcb34fT7rUtbVIjjaIVp9A/fN7bG5O1c+i7tbbtXesTLgIvJqDF7BpuX+fJo1PMY
7gbxvV+QKS+1H/73CIozCMb08UIFmj7SgGFxxCgtg9ZFbud4rX6Uw8PfQdG+0Xid
GX2kMyt/z/m6+4+3uqix3c4pjOSa80cBOCGrU/ZEZKSg6XE8w6dB9i9uRvRIdcAz
5v19Ig0Nn/eVwPQCvck3DL+BF3wY4TyAVPxhzg8z0ZzNEGQdUyAotwCoWY/SmqIl
FaPJBQhYCyOa8tZRQq5doJ6n0VnJ+rZw5EA2NsueXEB+ZeS5591fupNJP2oenWPM
mACKAjHAzTm21ezNPoHi5b+Sq3Ogz83JdXW5VZV7kLNtL6QuTXZL1LnVs1UXGbFR
R5pHpvDB+TRzgEzRB88HnLzsIwK8rW/w/HYl6s9YtXsEOL6OoSiQ0ZXmvy56jWkc
GD5Uz8uvqJAn+RoKlgubajePuNtFTtDnr3lOpefoiiv16tNZQu0Ns0TPVFBToXpY
n2lctcH6LpjGudbaY01eCj/DAo/i3fQYyGeFNCgitXbSRZcsNJoVnrDI8irdrghA
S5zEMAJhJG1LP+nL+xfFdJmWZOXJC6Rjp0tPogJETH3QOaU4IOwnglYhH7J3GYv0
8tgGX/DJpRJjRc9H5gcOLw4JPD/R5+3Qp5Z0ltThPs/+AMyHJSip96lwAD7U9b8L
LfwB0PboeGpOdOeCUsNaM0IdmMbPOM3v33c9z/VDej84AA2Jx3jKl3eX0AcMwHtK
OwYMm9dvYBh5BI/kUMha1HbDY/EM7q6+n8fcXcnRQ2qSvw9qC//Cxo+rmPuq0XLK
g6mD2f64qBoTilK1jC03XrKkeMGSdntqEFrRaO5Bo5ZFgC8GcPQ2NSU+Quw27Qb/
W73f25vY/u7qL9Vw2eR/uxIGdBKsDsC8TKfP9zKCt6SB7zmMR+HaIXvM4MwMIWzj
M+ee10CrAhc84/fns7riFWXSI4N8DHzJ1wMu+dlyTa0E4PN9KRShiZjlyJ7Fe+wD
EwaSz4FV1hLi81bZjOOGV8ibH2iN7jXbGf/YqjgbDO8TOzfS+avAYdB5YdxFsOkZ
pMpnpTK+XEblTy+P2w6QL5xNu/Z1cjhqjAt5v14oWGUzOzHQTB/EWZp/zhGQHNOj
r6fTICYx19NutJHjKshiCbOIQZRvD3GrULQrA0K+HugwQenz4Su3Tr3h2RWhgMzT
bIgyJhGJ891bbwKxf4Xbm+od7hEMoxcSy6aJ4k5z/e9aWilTuiepHtIx2L7juP3j
lXRzfkw1FnemILwbrXz3K+gLvuPJXfAlYTWBPgpVBSrzKkE3S7p6BUJJw1DwZfJW
RLh1NXxE7HxNjgg5G4Y9aETkLNz0bmOV3uK5veMS5OBuJ/0qZT6w85PbL18dk0ir
cHTNsh7byLKF9u1hzh4fPXuG5kRNuzL3EaPC5jlQIIux/YDvMtJrvpxepqyTx4kU
z7FKm4hHL2SVpHk5VGEH3prVlatEPnKgYIUduYCJqDOrg78lgcP+isQ1eaz0aeQ1
cUA89VgSUuOHxMfSXSr5sxsHFtDFKyw0nEh3F8DpuwCFrNajskyPg7Qm1xx+lwpf
HPS683PUHCZ9VCAC7sdT3M9ewnZUEa65pm8WI4vCFMDSc1vNbfwZ24oRlA1V1DwZ
kjbpcV/YPJ9oxFS2SjWf9x2UGJlyvK30W/1GpFw+gP19nWjzz18i43tLn/cvVHI2
FyrNhq3QuQAcM8J4j5XwPICQhCRTKvE6Nczqw5Qtq7fVZJlg2SWKlx3G3RotyLu9
CuEPsbq2rMZZBljXbSn7ZmlS0EaoDtuyd22eAvAI1NVANw93NrNFYXKCzPy7BAoh
SJpCC2bSjVEfcz6MC5Sj+ULY+0BlrkxUMvVuTfXo9bc7aWj7qBGxEI+sSy3bPxVE
cwdnFm5FIzY7+5j560s6LOGyXtr8VFtjaDpli+WuegjR14ZL3w495G/VW11ljVso
M64B0cbJ6c3yot7HpNdmhk+oTGBebq5cA09QXmU/ePmsYowyVrixfyD6YD9OaEbv
RmTwGqQFyATDH95THxPHMD9rrMnsE6UGf67VENa48EzWtwYCQai7t76SpfY6ina4
NjRGHBp7gHQuPDczmSnE5HdQpcL5aPEiL1JUkBfrn8Vsg3mLdFXzMi1ioNWDemTU
a2ogSIM1xRya3VX+btCyk2QCAeIAM0bhUSoOVzdJ/0BhrGzIiTWHGJNx42aIWFMr
/JH69Wog7cRDKQhKCF728SNSd4bBJ/I1xSDajlROCXXw4aCNcbOpKJHnzl/MBELc
g0yJPvf2yN0khac2VYnzxDshCqeLarNTCySsyAcqA8Y0KeBpXXxOtWo7DjEvMUOA
GMzLcDIQo1QxKUxeDF6m4jlVy/wq0jbJScTkE2r7YyH3pY8PJDjR6MMn5AWcAdAZ
m8ZNhyKZjezBfcrha5fVO+T1xkXLuP0VxRsU5STSrwO4oTZR/7O8t70IOeZYgHgc
N5C60Unc8vQ2n1FEsnEyFNXD3qxR4mnWl2wW1we0anpY5igb64NYimLqNcDwlFbZ
o+p+m4XP0iGZWO/Y43/bezKV5lp2f9nU4pxL4SgKAsPuos/tl4BAPy9jJmBOhD05
enpeDeLBL1jYFf3kGNEF8g/ZhQs0p8eNFRSxhbWQ8ZCaky/YsuP4OThc4OGcBLZK
mpEUo0U8HuOUjavnKuwW3QbJ43Ge3B2gzMGEs4xxghWcU7L9eHuKRF/36Ec5eSt9
ukWG4WP6dZG/d7bBelMXCaveSGsd6SuA1LaRo4uhTwiFZPb0plsCkyVjlhiQsKqn
W3SlnD1DnjDW+V1cH4T0ia+joMhvRorO3PbQj7QKao9bBBOtA3ee06xugHbZa3XQ
EYfQJTwwcKztN7opvvFBfbjnLYVG2fQPvNsaGW8P9zXpXmoReIPrfVcXVNdCnVPG
lZ3wKp39YExaHl6S4VzIqMzk6UDKrIdNEVLUaWJ5fIIAqo4ACliIUs3RUVbI7cSf
aQpfBhLWawsI1qgNtMq0fRhNVPY5fF/GGUWCmhOeL5iWmfazVKg2SzOvvGgoB5og
AGSIfPf68I1+fa6GrERmKtBUQ7LYe1GNkqs8nfLTbVCtXUhVGvb4qadcq5z0rcAJ
etMg5LvYk/npm6mJ9/93LD7Uk6tFE0WRzza0OSlbaI6o75EP2Nt6QyKlgwLWQA5S
TEUOIztemDk7kSNh1Ha6fN5hVwE8Tn3AkWLztpl95/jA6Gj+Y7mbms85Qi0TDNR7
69s/VxOhV4aEVWNDeCMZRmO4/NX3t57hj3rfc27ZRDgnFtcK6Eb8urJMezvkBL26
lQeF+yst+MLQ7pTweql9crtSQpbX5rKAYmZBfjOycaGSpX/V5LULEpljRxdd3FXx
0ESjMYLxbOQxyHGtN1simWj4yD8VuoRMAxKbkvqN9+lfqofgrORpaOI6KQgl7LAE
tmdIa2xQ0O45SjoSHobtHU28tEmQtodJChgehnqI0UTvwfMXyaWK/kYtK3H6hCO/
WJzGE0u5cy2O8fQ1qgv+gIG9Gc4VLQFoDoCUOHVPvOEOOtwNfLyWyfzgNrJ7rP6k
FdDBjg9uCHpCVUBYcM1ShvuapmXJgg692OHsOyUJ5xEYrQOj7f0THMqjbJkHvOS6
Ex2jBDsFOR08ESVJDy30tdBG7Pl7dsIhScEPvmu4mdePtGn1IPHtktZIZWUzmgvc
k4hbP3zf8sJdJaE9Vq4QghXE73RGtLL08paRx9nLoyKSGNDbPSkFe+wyqcxmPNEg
ACuWKZoq8Ml+0SHBLajzEGbi0AIg17ca55OHCjw2qVHFBAUauRtXaJXmAlw3tN2E
/OlnOvFrXOyJceMIfR4x6xyy8uo2QuiMCuBywi1Hkdkqla5f7wl860do7hWaowGi
NQ6EI/YdqbU65R28xqZP+zRiJIABKVP4mrNVQG8LNjx7i9fT24Jty8ZbiAmXcPwX
MABjMPPf1m53Zj1IRHP5hnrG9t733j7NYKn/XCCnA85zzr8te1QoKF3mFp7xRsGf
j2XL+WfPgajCNv1Jln23bPFpNFwbGvQfcJDE0V0jnSXFfJGdsDu1FLlzt+gUa1L0
ctEb8VsQb4ZGtYoxyoq8PiVze/ydH9ihv3saWfYAoA6nHgSLqX3k4DZdIlKLLlHT
ptfkONmm84b7Ls2xfnAl9QbAGdkz01VCL/rheXjTUw+l0iXplZZGSoEoxu3hkYAj
LewpJTqVWlL0LvytqpH7Y3wYVHPfDLvhrspo+yPSW6WhMswlYfEFUCZ3ZQkhjwjH
uiaM5Y7y8+0Wq7W7siOMFPoCrdaSweFvjwlffG9Khi8iTy3IACrOqumWdmjgH27L
ZaG1k6HqdE4rbC0XIkfDRcX+53SrzCobb6ZCM9OXOXSYg5nEHggdAnRBPuIcnttB
Qp+oMOpF7hw2gH8lGhNRuTymIFBpsVe+zPagTwlJKfXJgdzFxyIa7BW/FnOMqYPu
SgcKBHRsyyLuDRD6hIiVatupVcWz204CpeW++AOx5lcKy6cun+HtT3MLbyHXL0P3
B9jrJkU8f+zXuxD476AvPu4vcY2tvD8mewcLs7zq5+m0A8a/8lnfj6IQK5OvXGjN
2nwNPn8N92WbZ3pPJuBiKFQ7TSQVROvYiswDPNdf/XvQiY4FpkaO00WLI3H9aIyj
YhACMm6FyrX2rfgJZYiPhhfGYkbfZKvO7QAHy0gQ1QqvhTvrDcu42dw56XDskLxp
YiAIeiKqkzZoNdubUHmhy/hpUDZnubqzthixFgYpmYbcyqu4J6fKu2UDKf7aVPzW
c94+bkU9lG+RYNKndOQAFHM0O76yQRVCA//ebygcGPHbMajasZsVT4Z1MRNBgSZW
GaPUegwNIPTJTVtWjuOHreAgij3Bv4t/MbQVmS3kiq2QUUQT5L1hD5lOkNUn3aW0
2UQEQGuygbl8lC8Ss4quTQqJNs9bZ2cmRkmnrAo6EEQBeXKtt6EHvS0bk5mwzdNG
Ij+eot4JSauNFINjlTIu/j5PyHmcEb3SkQinQeg8Dt+XPX4eSSWuRW6n2y5lDKoy
xqzCxEeCj5yKYIvxCi1Oe1Fmll53D4f9lXLRvnGx2MsR9sWz7zDTY1RoZ0+B8mA3
aG0ePUW7HJbNliOF3zsQl+f0XC2wmdNfm/z3ktH7kVU+ZBTupESZryI81wkibYAY
RzrWb+xXa1uM/JDPkt2S0Q+j5MnLcNgJRwqLUGF0RuKyjJF7BtDJqBCAkhobOLGv
1du9I+573qULbyHGB3rNRuTXm0Cr4s7bqqcIYG0tz34jJDxeDB+HFf/WeXYMmYfU
S1WKNBDW3UnyQYimpuqo0z+d8K+LtWvE74yoWuFpB4MbXtZ/9Vs2EykPuELKoGkU
VqbRRwelrH1jZ9DlPO6iJZLOScJW0ehYUAbZPaFRkA+a8kc1IRNz2VJZf3QMLM7h
+3KIrVoh1hngZ7AHwnMzJgueRRFCPJuFq2gibt5mHG6pmno4AtbMe4yyhRmy9fFl
D3JUmdvG+3zN8mVRjEaWJxAaxLD0sXgetQZl24W40sGsWB3D7Km86HXcCGd4cxaq
o6dSlAHjAk4EmtW6hRbO2EvLboY4GGGQ9YxIRyo2jScu89DZg1mwzmyhGxsy2OxM
x+IGMV53oVw6RxNigNDdB2F74mhz7J8GcsURsJRMcmenVvutQQew7IJr/izE5ceL
/Tj9LvjpIROh8eg4NdWOmYOgaoJSB118+2qL2WMEfTXsfQ+Pcdx1+854UK2m8Gs7
DCsbMyAMvc60ONuIsodpAAV1qqq9m4Deit6L59ozfnDmnsWdP/7Q1AeLgn5i9tYR
5Z/Dt8Qz+2trkjSKiUlbymXZzSKRplmyUMTrwWzpJ4ITFuhYrq7RkD9gHeTKgWOt
zYUaC2PU3Qz9xnVVe9/HizHsyy0MBsGdVTMsI8JERZbmRXrN/D2FTw3Nve/O2TCl
rTaepvhq+1fF1CbA56Sz8nPkbONuqdkgw3A1AIc0sq8XWuRocseq92Aw83UXHz3+
OisnHbxM46lw/ErGEkktjNq5lyx7zVQnbcccGzseiT6sL6KC1/WwPkycVV6MOWui
+6YP2slugwJRFzGHXX4NR1kZfDMrEP4k8rqNeoOrCQjnHjD3ZsrBGuNtH4xXXKUp
vkF1pPYWRjos5p+4DfRuT/1hHA2mWRXN3tvzum3lUOoe7eBNgzz/adXuT+yS5Awh
MeSfhtQ7UgggONjXtJsgAXT55Cf6r2kRfhfdTADfG8jRgfbO45b6fWDdaq2vxpqd
/3NHJ6YXu/S+O+nZtJVF5SSzlFl2T7CysEcKu2ngUm6CNYMz6b9RurkYERoAzeEC
ZkdkYYbq3CVNEaHpFcYsQU2eddDGip+ovy+MJSJjRtvklysh6TkbwOm1V9f0P8K7
rFV8sIP8P6v+sh6T9hcRGzRz9Ull1XrTXzt3rNyg7X1nwAw+ZQ8sM4+ev95pzYgT
m1yQ8EiX2V2fsst1h2SPMNDatFdQdhF763VQBjZfvRHAlm2A67YUYLMWQm+dQ/TU
t5Z+Rkgb6dJ/iRVyp+d5YSLbjkVm0kFcCwshPd+HvIU/JWiwOv+iIN6PrgCoUeDL
raExQySrMqP6gvIAbqRgzkpgJSUIRvdW2NtSNXRW2++pMi1v/fqGb/f5il3RtHQ8
mO1RJ75smDqipkOOP2FJl63PrAKnCCCJJ22StDP+6rzyaHMFCHAHrx/ZX6UNEuI4
qMLCSVM/FoYI0L378nO6F0o6KcUAU5iNBwYPxIa6OGS0dlHzpV3JuEAP7eIJSLSS
9d+kj7+iK3Rb9Ur5D3uwRQtmT4f+XgARcWhr/wYkuvsgA+T0pC7+VV6MFW5B/18q
suFZOLscAa0vm8rGhY8lntTIQjz9aZBc7HW22df4m9bmz9pAwXUSmEX0W7ywAho6
EU0BjvW4MmomdzCIqPcm22EZB/9aM91tTuosD31sb+XKDfquEAmC0LzxDclGEN9t
Swaywieagdr4DH2rkqIP/AlRlzMmUABhEllo190icIOL+aQDEmUwJK8DWDLGs/fr
e85XLpw6h7DWO57VTsutNUR+YnlpimEseMPLcYAIz8TFHkfk9Eelnpr+aqm/cbdE
iQZwlLMR8K9YJiUXj0JpLthTjutSiA/MO2rX2Y2WEcSp3mbMtlWEaWGj5N7UPXvg
xpTgvDopPnU0CRTqbEKpxoH3epEFs8OxvlSXatAgGuWfq/a0XCcTQxKpeO7TpomV
CEOfcMbbRM6fF4t/msroG3XMc8gYbe5bUT00//YZnENZ2lox4Fy8X2iPOpAN55rQ
sASmv49Pz/j/syFiSnLtZLGyXVHt4mx5Le+2lBA6+SMMBCerWeM40I2y/yJBKwAV
HbBLPsqdQdR3pTYMpDNUDVVQgwpDVnIjFhpKNM8YM5Yk2RUv8QeNXCOImBqGev5c
/IFNWYhq8HwgWqwejUfDUrmytHIKhx7zjLAsEV7F6rlQ0cix/L1CF63r/+rPxqfv
N+ltqul+Jr0ckMEf5PBBGvvcnxcKWt/CVV7CL/gj5n4BE9uTcT4gyh4iHRo+S93h
8rK57IBLR3yua8fkqhO/qzyYBkmXEQ+z9bs+q3rODXlQG11weHc/7lAzZzrn0SLN
CVeznFW0OPEFWC6PlXqwP+B7ibwxoKRLSqp8yGJiMiCmqxMJoaiHOExZEOWoLuWI
fc0un41pRCvXsxLtvqW418pQMPxJpwKiW8GlXsyY4flfPOhQKizy8Uc84VXhGLaH
SPnU3XW9jf5ES+vPVoXdyM43rZbeNiGDtVVdXJ6IhwNd0vIlhWPJeIJXCytEud7t
p6BveA2CS3cGgqopzpaH0Vzx3g+pDNhd9M1CkTarmKp9/JNfR+eyOe7vmjJj++xo
BO5aQ6JVn89LfzCIebTe0bRBNSIOjDuqialuyF57Wp+PlXJ2zY3XZ5wZOBe/h9Kw
URHEE0zGn3FthEUEgbVStlfrAscuAmU699N1xNbA3mk8IZM0Y19OZEVxf2+9TY0S
Od8FLWEZfrKtHGWqt7SEpfu4AVQuK4i7pQwW5yOjKhX9bD2DweHKkP/hYYJ655rd
YNLFs2N0mlu+2T0Gp7YTn7c/+UBP6e/JqWIIZ6sy8ocsjsM9aA5lTxhZzHnVhYxf
itbhQMHaK8FDp4I1HjiGJ3bxKzNLHFLWKo+MPDfCtW8r1aNoBmuRQWz/kK1dVYVw
DTOI5tMrBm53jTESFHOZSs/Qiq7S9vf4XnG+YC4V1IFEuchJ87orReYOrWMYIRc+
uE35ZSFFxEIB5Afsa3yaCw1ExKVOS6LgD3XXmqHv2Dhug4e/9diH4c+jksg2cKFu
cVFxqDh/L/KJaUXbacmsEaLX0UkvxnlA7/7XHMo6UlwFgIoq3nvddEMSKkKL11Jb
yM+G2rUCQQ2xm9MlTi0nkKBLR8aC6B9Hr+ApKkxc3iJSSFTdUf/B0DlE0PcFgAWO
NCyNDfBuNUmqqxPOFi2Fpn74S4ttPp31FpDjlx4gPjKigzCZcUPazR1AGK2d0+Yx
01ZV1RZegidY6YNbPEVsuyix+IhXtS3SqmLi9dtakD20nBsI2fDdDDA0Z4aRk6+4
8+iGIerB8iiPsESrb2btqIief9AvRWF+Vhr9lyAAgEYcfYeRH1YA/6qnLoylAbKt
3ioEE2BkfZzEK/joYiaw7pCFFdEIQ0Yi1jL6osUWsbvMYwoV7OkSJJ+aU4PYAMP2
d6CRlVBaLNlgYC0q1AAlwTxMcvXsMa9eUtL4tD5+9T59HFpueqUWikFo0PkmUEl/
RspPP6I0xFF41XGd3wofuxV7l4l6tcMbL25rriO1nxzl822OerkeW4kVsxV1/kvW
KJHFunX6ZEM5g9QRmEy0vTfgYzzVPskkAf9HZUvJDTw5ehOV5+0Uaew6MejRBss4
wkQ2Vp6sJUsTRli9LiSPpHavJmj8/vsgoFUrLAIl0evSgWqHIyc336HwjolsbY7V
U0ipF3xOGIX6zrr5O3ofNCjSdgEUDv76B0UC0OJSIO9Qfjw2RxryLV1jd0/JUIG8
ccE+wCEyBR/Iuj2bjcEZbXR8f7/Ocut/5rNQcpJxLkDcReqokJB140iqMq/t+eP7
1JXufpYE+zCigAukOnwM4e+LlICrJx7mOcGlbiUIr3RmWyHzfJCJWh6IjQYkqcFv
0xF+IjBxMqWqWazP5zPYJpHn81hqo1s0avWDDMm8V8d1DJGYQkDd2i5c2NmfZEm9
YEn6btFxoDU3rfiJVnfcTycA0NM4f0Ec5IQkwzz+c7sEYF7+dw5gHx90NpPIH63e
oXPPj3aX48pHkLNtfE8V+trBxEKeLKA7Wt5e61NA8m8mWUDmDsMEBTiDZt9s/fyb
lC75TdSRPLEt/t/oYNuvPu+b43O5kcZI7gbl1ewHlkn65hFONiD8iYbZRRO1J+JH
gHSxLwfrfdjUkisx0uSrNzudNOY8mcnpzIeyOw+1ivUeqcqxOICSD1okopUhZQIf
8y0A3kkD8e6PNs8yfR+Jb5tr/iSiST78H9Q5wb1vU5xZwFvWTdECgas4MB8+joRc
g5dtrsBnPDy0SWaMAIOwvUd7o8T3IR+JNcFG7yrr+95jlVluoJnsA2C2K16z5tv7
cz4iFX4nf/d2/rJ/cfSdIweoV94TRnxWeL5s90kVr9pHRZb4lo8AM9OKUKldGYfJ
fr7DbkN9X+4I2uQwCTqv/0jYAxFLMkIC4Pk/CGY2ag5/jHk1HeyZONHt9Lasyrge
hN0d/225786xqqjF/RJkA4T0fxFo2578Qc8oXrSardYvEMebLwpv7DV2SxmDihBu
//uueq+AwpWJg5quGV2yFomTNe+BX9s0za4UheVQFdZnUpCNU1u/AftugD13yTfA
HsYmAaI0PXNZUeZM6TEGY6uOSHecU0AXCKHSWA++NV4kgRBWF7VZ36rvrSaEiheF
Cl+b1+zycIwiNtBzyWp1overKh8SfSlN+Uz1+svkzFe9+7Ox4DhRiQrRaheBaaMF
u0Mp6V5AZDbk60kshknGVcKjkdEwT6PUcmD5h1RxfuNZVOOMsIlFucwmD1E1L7y0
1sy+VrOaYVntTSto3ML+MhXcP0YHMnpkF8YUb5JddWu8+8yWKxGw69cCDgQ1Nl8b
AhUb2EkLb/io9MIJFKvyb8m2mI9E47MzYolCsKQyBzbXkTzQa6RR52IMJk9VWVDy
yKwM47y4syQ/kx0/b/Gy+8Rf9EIBGeOlj2DuzoXOa0nqR8ip7JNbPu0qq51fDkdA
oXJ4nL5pVY2l0c9ud9LsMaUcZ7qb9jUChjgfAvAb3Xl1ifBiMPM9OYO3AlGMsWyd
k3xp2QSS+rXAtKO5Q2dUu7N8pTDyRqqNXw9fZ/1sv0H9U8QeKPxZlXnnN8uE+9NB
SjjomwRV9x02kxcTbmEI4qSOx6kDpAp/VWW29kH1nsCBD25Fdc/A2CegHg07cgpw
au3v02hRm3RL4QGhC68OS/AhgPZcvrlvvMVLcinxcYpGetS7MyD5xg8OX5/NakBE
9QEu0vSuYTfCjEIALuk8HQtZLwNbqAohGxQKQoRBTUl/Qbp8/EfY9pZHKCfOtonG
2w6fwyU9mxZiogqKmFtxMGVHJ5f+joJ07hwLCytrLamDFOSaj7q4xQ/xY9IBnTOh
Bw13aVW9QxCuhdCK3dVskqrrRCgw68bGBDKq8IFYpT24/6yzii1P9IohIr6rMmCT
BqK+Mp4MZnYUmaHsfubzGEA3dsysBsMivf4e9GyQ+S/nZqNlxBMDEld47l2LO8Ic
V1kp85YozSy+O+JmONha/+blMTyLeQMbgL6wjzjBitoyic5WqcltxB+ZQfZGliIw
le8UYDEj9F3Xv7VLDQkTAsXKyLkBB0XSR1PafsZRtoKNcRITrZJo2uoSJqCgBxeU
AkH+/1XjiOei8AOMBvhvBWtDl/ONq6yn4djsiVgAJQ9d0Ki7B+d1MjROHZoyiXFz
6TkIs+JLgjyDlTQnA82Vxobvql7hkeE06z1UeP5sugQ5++zwfaDJRAk3DBbXNFim
lh0NbyevvJf91XBe5ahgytpiFdAk51ot22ZTAFqO40TKJP6oduM54KDgLmMfGmoh
QDZ6KQHGBgVTKmuWlwItuQljIo+eoIc6Ifk69T9pN0omeXIYsKAfUSwttWXtkSqu
VAH92pU26n6gxXptwdkupwTU7BVp97hTfz7Cq1/rhuyWOrTc6/gdk9RkqAknM3o7
r7SGqbRklmzrxeY4FD9Fe7MeIIkvIZJfMblFkR2/4E+Zed33rNUqLh2k/qqwYFql
8Ci4kj8a46LTpXrLEXBQnytNcoU+5Xe7OiMSZIwUXDYZJxk8o5ONYuCwFr32r6AY
Ae1oba46ylo8w+qIwLOXX2DtkA2v23pphX+8pGd6rCoY2ymViyCYKQDMGBdLUa4v
xclkafZwQ0aURuUgAsdfFSl7qX2hADQSmbvTq3uHj7xTR6isc0KkD0HPhfKgnAWm
/DPCe28xw3Uk+Lfr9rtnKuW6cCiSEePKXTLoqVSHIFKPVSo/l/nb7vFap5yXUaFS
Gk01XAIN0jG0Ac1ZvXKkSyBDS0+PF6kd41qMECFJRB6+9Yq6/EIuZNa7VeDM5z7Q
CUIy/Xuvf/IDF0NLvcy37ElTHP7vVeW5kkup+0Q8sx3ik+C+fJJrR6ryM82Lm3VY
zMEK1FQkRTBVes4IrARXPfnIuhc72vW27eMeljNJL33W7CmfTtA9vSFvZq9SYQHv
SlFeNeHNh14pKXzdIYZlGwp+1E37l+oijgyX35577MGB+KL2wUCh+IrTDT3mhpq2
5r8OuEnj1FAyrX2lNXqh8aRSQFxUZfw1jDUDOKPhNlEyre1C0+5TWUIhAh3wulIq
RAzwTe2SAc8KaA4NA6ellT77ExszUNIjgVhDij/J/b0bs6jENED5nJBPiXwnTSt2
mkPkPLkF0nfPqJ6fa7c970oYmBJQ7H71MypyPm05/TvuxFrWUqTp6zCoQDEhixW8
d6Cx3POrScnrSgE3TyI+Nir8oDNM5Zk+ph2PRe0x7H8lekbVlHvo54AQyPFvd9Gg
0Gi4XhT+9QVKnxzrCl0tWULN3cM6MaEl1N3VdRxz6PoxikzSkQl+vDOvQOZ4nJF4
+gok05HIxs+Vkv7605NKvOog7Y3NvQAZQ0IZludW2UlX1rRzEzkvEPB+y/pRLNZP
K8yZ3A453FUPGzN2lB7gl6H2lzk4UxrcjSOM7C1OQVYuGkbb/ii+2iKboevnhTgd
w0tsKgpa3aM3T1ym8iHDEx3bQf6363oQvhANwUqDweQaiRPw/GtjWDto9bodniyJ
ATXjmWqZ2cXCMEPzLUFq7ICu+RHhQoe8+52orXus1xdFljSNBKXLMlrR3PI6aBqU
v224y1R03xkJeJCyaeMCm7ILPcDyxA1YB8P4y3idYiQXCh5hdP2ZKl5ozwuxNPFs
dkdifCxxXpY2Dj1bbDROTaI9ACt1of+PK2EuokDi/7zJBse2g8418J0y+spRJyBF
+/YK5z9Mo2qYumNCGKoBGGOEoWFc/ya8UxGHLqrcijnqfxFu3SqSgAtgpdgwX2fE
MCeC5W/ZlLQIfHNe3XjtYyUhtMu/qV3NkoxZWG7lSRI+xRgz2GdU6JUp1ebKxzgZ
q+HPL+SkAYN2We39tTWGEDk+Z5Rbh+onJlmwWAZB4RAkzRq3rA4yFcRSgPhhsLZ7
OvuyPyNwG+sE0w5Z9/9ljPYhu9ugHOr7mMKbYKsfv70R5PKQ48hJCi2x2VVzinBE
K7ZOHOwVZhMJHm1+k1ppgAbOdzWv9pLL1hA3rmL1qzDVvTQiwliJQpc2jAvCIHp4
ODETYqVj16pwTj9WfplOAL2BqcNsKuR/5qa71bgDpvBUfDfnhWA5DdB16A8iW0DS
nXlcdjUsrW4PV/8jYOdkQ3lJktoKvw9ik2RbLGtz+p8hHRf3o0myh0+DfuzUS/Fu
31waktx9cWgFUI/OEMTWm8T+nso+FwRgpgnf8MbzJRI7BX+gjWlYLL37pDRUh7es
FAcMEmOE6VVZCFGV1YA0qrGFgAUDVceiw1KKwasw6KkrXsMQt6FjfY8XoobLGpxk
P+DcUnIQwXpAM0R1ov00LZ4tJvBJYywqRHJemfwF5PVv5NT8RkjixOVssyBzwYSx
BJ5crNJzPlwLrqXcmKEwooIXZOuVvwQ3KylLm3MexpiKL5aK6F1jym/vnvgKb27j
g+xdLVQpuaEG90XKyJbXlBISwqcp3/NDAmSvt36CdCm7nx2rVz7oKREsoTUYwGt7
yEhVBAiIgeXHRUGwiv46jgog2B2RyRDiI1g3rX1+/h5PEDZgXRKAKjE1jhhGshYN
S45AxzBUErViBu4o3+pmhONbgvlCJNx6OrAU45W+acAuJISaHyzVuZLxtdVH+Th3
khEI2m7fvz1vhn33bgKn1oJcXZHw7UIkwF4FWWNGCpamOZSdFdDCCMAARgo9GYBD
SJNmrCqLxH+VVODAR/p7gE+4fu5uOAW5OA6VZgtOvsbIgbCeRyTUvr2noZ+YGfRD
UaBCrMjJsINKw9Bw6x5OZ595xis7yzk7jytFHrRqK04oPbLPS6QMkBOyKBU648x+
ES5h7q8w7bu7yOt6AL2wKIP1l1fczhzZOPonm6An2zszbTpWBNRTKeVBzw2/VMsr
V2xKN1SdG6+9HkLHObsa2kmqyh1Hatz33DKHY21ggghmTpyTgcW5ppOnpciBADb9
Pn2Ft+TFYbCfmx3CPAiYRWvIRRXRB9QMSu6eTrsxhxa0JspwKc/bMRUSJ0q38GZI
bOcJuFN+ArByp2gFw95J0L9QhhxqhCle21Fw50CcMNk/o2tW58fGggLOmup4/+JV
D5E7WQXQI9k9B4fXWKU+yuRqQZw+QM+HaSn+Q0253/jP0inN/LX1iI8HszRFK0wa
gyhdqNy3mX/Ot1zuICuw6Ns8MXxYo9wTXZRON9eJrSMeAIW2Djq9hBMUz8XP2uYD
V9ysKecDkkj6zIANU0bzI62RlUHkizHLsHz3ia2mstcRmGcqbHIuhNGIeWPGUwFt
FyhKXflCo7Zy2c/at68XsSgjJXJR7/dHRviWXg6dq1lZpWHyGzzw5wdwjN6RNmuK
eij35nW5PuRawrcFzAyqz1snFRdK0x9NjSzZX7tBlgugaCNz6QF35a04tbLLZVbI
QOobgmQdAlq6oZfDbQB2eplQfnVRoTfwfbP/b3R/TnakbR56uxwPe/3VKxNNVUky
Jf77+4zS1GCSRhxMaRRPPHynIVyxsi4BSmvkjVdFa22yUt+gSpElv1uSyXMS/g6Q
Ol2hX8Ja+IMNM0/2JAk7BT375+YQQjL9BJO/ig4EO8oSzKHuhBBEhLleS1c+ivun
8gF/o9DZ+RSn6dBfXT0ID3pckeuaK9F7fRkvuiga7ft1wKYCv4bbIG6/xA/bdvTn
IshzPuDyUZ12k6fFpBbd1ySoMqpyK9K84sqIrhly6iWqHkwtSICxeH5axaovAgYo
o5glOkpZgDCXGYT1+uuW6dPucbhS0mxBeBlhbj2/SByZSJRpoScP/PaMqkRZFRob
45myRO61hIQnQEgdVzDlcanXI5lCEP8PYR4JNHiyCNHwWPOT3Jl++RsrH5idWASa
q3OrGaVAVzVBgzfCPDvGhb5OEVNAvFNUdx4N/BWB3Z68sXE892986bJfGxl9xpmH
A+lCWC3364IcIpeov1AvmrhlO0k5nfYnaT0cckZK7rTrUsRYaiAu03eD6/KnOUAe
acTawPREkyShGgHZiFv/7aAeGQr+LpJ/siQhsmvuYsmu+/hecNemg14yAeJvC8jV
xbh8Bc25jmmBBYrtBw4lh3nz0LNqJxH8ns+fOfC3nrmWzof8a2MIFQDZwnUBBTVe
xu/TaiZqHg5hbtBubCB8vRA+4XrC+t6DEeDl2onJtkzvpivuqpUVrzmurhEuFJv2
xqJh3aObw+Pp97pyXYSrh0DTIcbhw+Dqy/79D1N6IvbRMSep3IerOKQ+npAiLVKs
bnSuqKBo+3pB3WQjzl6EOZ/WRFm0aQImEY1zfjVLjB/UjFDwjTNMNecR5zPYqcQH
hDB7Z7J46a+XNgUm6P4TwRK19uk0BCPh0jzJU60AYy8BVyzOz6NrmVdE0dLi/zP6
OdQIzjcVKa+VFuSzBr+7+ooA8gqUMB2Iu4/+FkDoICbF2qd5YhBniES2kJ62cr8I
EivQ1gnlTmyofbexF2BF5celL+0F8TXiRgnAgvRhYY7U1ZCZUVc9xeW+rFAjOQSz
OFmQ84JUkZ4azillSfo/90bu7Yud81u71TxiZ+XXwuDc12jUEEK2OCv4FzI2KKFS
5dTTTQAEb5scnXrzYukr0E5ml75yn0Xitn9wSpCrl2pdpqlJzFhZbSXM9Sugsy9v
0MgB0yU298I+qsMugalLDHdffllblUIwT7dvyJpBmQ4WjCmUDV1I2dzxeSexiIUP
YbhpOh4e+mvoAPvjBN3qn/Em+w7nqC1dPXxfQ8KMaT8hhwiBF1SoQqEyIGV+2l84
shLmxVytdbbrjSIRc6gc+oN7aWY3k1qjF/7hgmlzSOBgJ1zyOSmltn57NEDKY0lm
TF33GScAPqxLeF9tLkQfSFw/ZB1+HZRGbDE6FOw/LCEllxzBRj81ZMfUG7U/zTLU
FxbZHNr0dZj2KtSF5EooIPAVyF9r270StXQDxOFyAQqHcuPNbGps2vDu+Sr571hc
G7PaoxqJBGfUvJWleJZza9gxbFurHnqu+dyWIlH8qKpUxy+E10tbew81hCt65ZF2
Fhf2oP2fzNrkUa0sVtzhIhOS/jxuu4LTIQ+CTCTnk6qANQZ7Ma6qe/jbQMT7kS/n
Yk4c9I0PywUWjKs1kRHrL9C0/p4mZKpDY7nyDjKbds3Zeme3ObxTJp1BWrVf7Qvk
NSFhHhX/wQzS1tHf31Vt1g==
`protect END_PROTECTED