��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F��������n�BJ�F���U�FW9d����T�+�wt3��^��r�q;\��af�י,��9NL���ٴ�[�Z��^��Jy���0�T����l|�x�5#B�o* ��J/�CO������|�)6b,P;����t��ew�u��5�v�u�E�8����R�oIk�����Wb�A1���5��r�5Hڜ �r�n+��MS5��n��þ�|R1��������E�%��0E���;%�6�׸ۈ�6��:�!�#��L�jT�a�S�N�LS�[�&Ϫ���]/��nm� 8K� 7�H�be��
@��1>��?���X�U��&��P4
��J��tz�6�^�O�A��S�������EjS�V�6�$�g)�H!�uA�����.����c:k���:J�G�y�*aio������6M�pʫ��QZkw5~��ΰ <�z���i����Y�T�w-�q$��k�d�V�5i��[�r6t�`?�.�^�v�
��l�;�y/��y6�]*T�۔"N��d�V۬����/S[�B�U��7 a��p~q������~�5�LPؐ�V�T��?*�ؓ�C�r�����	�].o������߽o8+\i+�`K��+darwEi�JI��4?�}͍�<<�,�j��'��u��K�C���=a�X̉��37�Z?�(ȣ�$��Yl\e���=~�Xa��s	 -~����w�N���,v-�xa��$a2��hA$]��g���[\�7�x���{�MO|���1Wc���C��e,m�"��$�O��
	��M_O�~���jCL�"����V��P�h�Jm�_E��HaT0CS��&�L1<LJ�ګg 9Tp���N�Hm�}r�NBa<��9����-L��s�/�ap6@^߇T��!�3��`�[�� [ݭ��O�>F��� ���&�	��A�A��.V�Sk^�%�M������P ���v׮���w���>��!S��'ho)�ˆ�v󃜎�u�G�E?! ^�ZY�����m���<˨[S���t�sp#�5	�(1���{���ݶb ���Z���������q������Eő�-U���V�||J���F�7 ���gD���ș��-'�^��Qt�N�?���Zu�ܲ;pULJ.ku;�8h���nô�q	�Zk�[^Q�s ŀo_�-����H|��\C7}:)NLQ�Ծ��w�r(@���-�l�N�5*�q��-��KR+�]wN��
h�rtu�d���g<��YO���.[��6��ތ!���R��yNE��D�I�Γ(��Z �Q�b[��o`r~Q�"Z�j�x��+�L��G���Q ��c�_W,�t�E��`H��W�k
I~g��%ß�!)Y�
"��0���k�[]�3,���Jb����Xsp�2c�(���E�������J�G���n�z-�r-s/_�"��0�l�G��%�y0�=�}TΜ��O_ҹ�ĉ8u�Q��Î��z�ge��9;�)�N|q��"��Fx������'LpP��SS?����tX96/��S�<�����)	�<e(�]7�3�b�ѝ�Ӈk�1��x:H.�{0�/�J��MR+��ֿ�����|������V�c�?{lP�yլ��Q�H�ߍ�;�Q���p)�U���\D�LExO-��c�nh�{�[b8���~��\�!�������mD�s�l����B��4����R��٘ f����`r4����-
P�X�|���8��#в���V�s3�YIk�i������f��������k��3&Qޢ�:^Z�����O|���烛a��6[�I���B���D9`ͻ����!��鎄����f)�-%t�6IPy9C�0������1��*P�Q��b���lI#�oF$�4�և���uk]�u9*���_Y�[����3!�#q�{�����@N�"G��g,}�v
:����c�{���+eTuX�:�%����Ǡд�CY�v��5���0OOi�s��.�I�Pz+.�K��%��\�2m\��+��؊Z ���{Y_���Us��g�4D�#}�XJ^��4��5G�v�h���� 	��]��Nߋ�L��j��.m�|����틮��=@�Ҧk�⤞Q�C����K!v�1�x�gBo��zZ.��ɛfz/c�4��.��Y�^��~zC�׷Z��]�+�s;�!��8
�ݍS��Q~�����]�1�����9m�	Az���|:�/30c.�!j�;�[2趯�ȢAH}4?/b������	�����<)]��Gwݻt~��a��K{|�BH�"�F�T�r��x��:��ݏM@�&<�ݱ�O�,\�������� ��!;N���X+��2�p��@��r�5V�$pb�]�2)�my'���r$y�����u�%[����6If�0+*K��Z�F>��	������Q�/�f��Ꚃ�<}��7��jI5Nw�p�J�#�H��p�"TJbɺ���%I�Bз3�$�>�Z�_�,;uó�Oߩrw%T��O�N��S��/<Q0{f���G�������jL�j��aUL�a���`kk>��.���͈�Zm|'�\���e�6Tt�����1�llG7�j2ݲ)+!�=��?<��8דF�L���\�w�ʫ?i�.
� �cz����Ĉ\���Aj����'���o���K�p�D�(�]���}���*���~�'�`���˟���h`����}�!��{H�؊������ƣ�H���#�H�cN���ٍ&c, �%�\F���7�ֹ�l��&Άz{�v,��-*D�W��I�t#�-����2D%�b`D�<+V�!_�*X�a��Ph����G��[<�۠*S#��⩄�vvF��VQ
[S���ú'O�ԋ��k��VkK9b_��� �\���L5k4 䨴kQB��.�F�?GV�r�1�L~6��� ���`�3}Q2ԖSb��)ZVY�����Qw`�:/�=o�g��l84y}�ݐ���f!�k�����e%%��uAot��5M��Qk��"�RC��9�3�I�i����g!H�������r�P73�	|���%0U�_j������y��$^���֪�jJ��fu�_�w̚(oħ1���>
�)l--�9�\��N(Fi+�� D��QQ�b��U�_^�.G}�����#�s��$OW�T�>��pN����C�7��5z��5&�A]�����Q�):�7"�����}rHuκ(�kǞ�����,�1��h�4m  �I�����^�;XcF뽌\�Į�X9�q*�kTB��$��Z�al�R��:�NA�ñ�)\���Ht�9�`)Y�5x���T����Hտ�s�#j@�Y�C0�����n]W�b����COk譒yTʱ�iH����j�( s�ƴ^���.�|)�4��jI�9�7S�f����U	�
�����$"��L���7��PM�P��R&������^����T�%�9�磤�~����@������J�J��e�gU!�h���GU9�	Y+.m�$�&��y��T(	R�@��I��D;�"G�}C��L���%㚥���z����ax��fzɨ�Y����V+�jş����+����5
�E�ϛfi���{�����t�(�I�oBo�W��"�_I�e���oi��>q5f%����tW�Hc���'Q�@l	Q�!�{!�I���!��dx�Q�
�Vc�ɁO�z(Ł�U���P�-0��!_�/
��ԪQ�ը=��x���Gm���JOu��y�u�Hm��gT@���BV��⹙��N�{)µD�!s��+���e]��il'��(�gy�u *Ml�r�[O��S�O*��hX"Pw�������L7t��^O�V<��IO���S(�qD�CC�2bXEI��`�v�6���!��3�ʃy�L��Q�$(�\8E����R �Pw�/��p���x&>> ��Q�����HWAw�]�kn��Iωy�@&��4k_�rie~�����.�������yQcH�_����	s�f\���$���ֱ�@�Nf��}��Q�P����%�b��:Կ�i-I�Y]Y��F7Iڜ{�؞�i��5 .v��dU+�0����ݾ5��$'A���'�z%�ƀ��f���<�=5]"����V���W�';_"��C�=9�3o����.A�z<��x������ڗDp������M$�Z��Q����X��2��G�rd�`�w��_b�q�^4�O��?�	�9{���o�x��cq�H�g��8;:�4���0��om���
��h��e��uo>j�r�G{����}{4�m�ۛp]nA��\����|��ʙ?4�>�Hvq��]W���=5\vC���Q�)�'S(:�'��>����n��+�|��=@O�i�"^>W]�q�Ռ��������Y�,��qi�tf1F<=�ݽ�%��TP���W$��d8���(Փ�qXa`����q�r:��.j���bi�;kI��+Z֦�K� ����T�q~���R>�?"��]֟�4/�f�0���&##�6<���Gu����`�O��,h�稟�*�Vr�8�M�8:)*1r�[�"�^R���;-�0��7#j���Ǧ~���[��v��
<'���!�K�;h8��	��V�`�6�