-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
LsGRibhJjCkEIs9phXLKEw4anzmYUJTN2KuXSlAvkw5l2DhiwdRAHuF3YZzwcIH8xr2XE0HsMji5
lK3tswid+BUCkv/2UK3s8t8vsv7SWDQKlAJ7p/k+gkNsQs/0EGYtpGXJoo2K/R+BgmI6CFbzvvwO
F4ZvNoHa4WlzfpXrrRHv51nxAzE10ryNbCq/BY08yTia4fpQj4sXrbVloVRtE9OzWiJyBM7+EDbe
4ix4eAL9/TUV5A/17NBeXuJaZBL6nrrNWuiKPGVdJ77zeYxMbyL3+/hhnL1X5QBfaSpmXyJupqZ9
hHoDcja2nrePzjtoXfOp8C61EJgl/3YboaATJQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 24704)
`protect data_block
thDVDV+3BwSLgwEfaIf6Nj3WbPVbrFFBxxey9ENrs6vx4t3BMxCvLdYxQ23Xii5772V8kyBwnRB6
I+ZkAUjEC/F4kOlNKHzRuQ0kmdU3y6tNQoMazIlU23ALN5es/kc4QB6QTMcqgkGiattjYm4QgZC0
IhH3NB/Z3ljBnvBeBRYZISMNhiD1EHuHujlAhBhCfRvZVJct2Ps6oBZ8DvS+qJAB6FQ/c+Y9F0rg
oOp0NAk3Cf0O+UJLqaNUfIH1TKmbCZaf9frgGimZPR4zg5GmGVC/2rhdMsR1oMA6CWP1w6V9PSZN
MwJ8JPnlTZYVplaVKqOfoyGBAzMrDEXMJWeiK5oWTAjs8q8o5HLcULsm0McMTLUNWbIM9wynF+ov
cvgXkYKhtHFU6pCnQKQW5N7AHlXzZWyGSeH+aZBQrXAO7UwsuqHZU0WAtbJnnuDH5FT6zaJsQPEa
OjI2C+Krj6YXXB0Tw0MSJNfiolMPNXVg0WCarclt5EEYgeePivcSDicV/7W0MYi4xDCF3CE3ueIV
QAFwIAKWGW2/3TLQfhbo1K9o3ft0ypxk4dZsJ2Et0NMS1ardRTrNhGKLJwwyT4JXnGmCr7abxNbt
wwaVXUK/q6GWy5/PGm6lfqSCkEBG7KQ37WcQzGye8Zjsc50i4fvD0WVFaFwyBs/bN9N28eiCui4c
rC2WMpGC8WzDLF8VYcYsoqgeIsIjwu7MZycwe1zkwQRajjEs1Ljg0TehDrM9T4Fa9ACsqc1jkgxV
dwZFl5t7kJ2Ua7CTqStoxVk3/MvKr3FvEq8D+zWeinUUW9nH2YZEZNEre4Gem++2Z2ofS4Nol38z
oRW1COeVRf9JUSweyH1DUvraj+krN4ovfs/oftAy7ARjOckIbevvBHDG+Qx/BKwBPjzONsVX8pVZ
cwXgIds7l31XQEuP47yLzW1Fv5RI8r90u27BE5eYHeTA/mxwgIj1mBkPLkO66McLz6/DFR8Oyt+P
byLhhbK1VK7isFHu1wFE6yk1lXxfeUh5uGlLA6Ig+jPLzmsS1rSTz+E2+oYab4R64Rle70o1OocT
apS/k5uMYqPWP9uj6l7cGpINjIRV+3QgB5hE0ADyBhJEPNzjgfkGJA8PgcVpgrCPqalhTTDLtP31
n1U+94XwvhpUYl5B+lRP0x2pDKsVgOnh64V0la8BJl1xOhMTvxLUlCHDCA7F6b2hnAsLxbRuKPAv
iRgjiXewT1gHs9A4i3Tgb7dIs8joq8B/Dl617sVCzl/XLS/m511MzKGXhNEReLGkiqu8RafO4yZC
s//5drZRj//Qb/HMqkflDNy+wU4lu8X8jzWKT84q+NSZgMRUufxRYUr+JB8ar8/XNQlLv10QZ9IE
XV+bWVaYl6QRkWNeZ5UaiDtqGhnLGtJm7K6hlklPqBLW1YWzoc/+bF/0EvUFActgHjZHIDtDi6S5
0WxlDNii4g1VwPFgMHnyVE/l7Q+wuCAmS66qixhijOlTzV9sXHq5guIR4bwWQ1Ml4qpIBJkA9KAT
il4Px6Y+LVEXbM5KqKwKslBMx0K6DU6/xT34JKSwOD2+Iq1awlJi91mStj5n6wr3Ck9EWW7rWK0T
DmiFJpkxLBr63QNA5mL6WGM6KFWZGen9S8GaM8xhQCi+syVmFOlPIi2kmuvEd0SK5khWofAWd0kM
jkg9zcGbu4DKotaykg5w9bMyclW1tSwFIbyUQeXH4mBU4A/8Zodm6zqbAwGiRiaFLLWCwMtMzs86
C4WPOQM29Ixleo4LAhR68xRKf4hL9klKhbBM1XGPpLNbdcITg8UuOcTKPFqxJX62jYO0V2XIqsvX
u+Tl3cNS2I3CoSWeP2UyIfQW9kG9S5JxzOua93gw6LEIksVLx7r59ScDpl8fykKmKgUHTPk8kNqT
otF7fN/dLOd3iGjpsN5XOgcNDzT8dhI2hZN19i0uh7T6LA8NdB1RjT48XyznQwU92tfa4MAzCZmX
D3C2IyYspGbbRk6XkNfvi6JdH5vyRPVDGyjl9pyTxLJTdxmdo4BpSH0r6Ikd+6yyrrzDa5CN7sZ9
iLJBplpm6IsSpgGm33DuhyjrlpxGC6IoBSIMngf/7YEFEc6Q72mwdWveUc0lzPUSLDa0V5L+zw8C
XPait/RW1oDIn3WJp6Vj5gfXicS2+PRWiaKkk7qFDNOOvA45mgO9Nlju2YRH4BKl2O7GriksMdYR
HY7YgStpAzOOhrlrd3RfLnfKKxnqSjvl95lL7qPxoO2pepftV0r+4ZFm4rR2WnrlcQaW0til4+0o
8kYx/qvaZrMmaPUEycIck2d0vjeQvqenQE90zAVqcKiThiqlHnwsKZyzfE4DPBcFIMpJ9Xw8n4gm
sYDdTdeQJiihqeJsqvjcnBJxfYdvvu3sgUu0Z/NnDab+eHwyITOAwJfLE+b6g1dcILHBkgAm68gT
4uzUo4dfONvmuYbQkRfeE7Gu/Z4sMZLx76jTIT7bAhmeY+V7vq/wR20/bXH6xErpenfkHIM3EEnu
Cwgb0YJ4z8DsWB7lWlTRHa9arzvq2mIRn6JsdrkoTrJSvI/FjlVPcfgQHTtq4+Mn5WKNTpKd31PG
ZYuLb7dhJLsFj4xi/JrI/BKN++rz9VDjf4Oyz6cMKTOLgpWQ4VWBr8PigG23VLyVELUO7Ji9XDYv
Zjw7mHmBNfi8CwSfqcm9xC3KqMg1PPdleJ2vS5te0ATFJnfwxnnVTdp7xhCnu9c1U09QwehBLnDG
5ExPqCIkzq2BLGFwvBvwIlTAkysX7nmw/Eem9MFA5KPuHLZJHuWpkOiv/IWfpEPyAATFKkMGmK+Z
Bq6tpKhTUEPUHJSCVN3YfvR+hKXxmlNtuhL4A38FIAHSF4DtBcgW2wVyALpQL445KIqdHtRwYIa2
87NCrzYejbYWyI7b92BAQan5DXiYirI4EG1a+FXPejblPs3dJuRBdKigkmvO/+BO8ktUcNI0Vm/Z
jbbVXClDv676Dup/Xl7pzCbUc2ALIszvUYlr2dZkov+sCaRg36rlJjEhfbjigrmkg7gFAUivlgie
V71qI3BM6IAWlSbE9+rpKIL6oIlFkP2yxJMuCAsrmfHo1NxY1Bc2pT8Zsydc6cYm+A58VbdjZQjy
4CGpoINR3O9xdIKJHa4JK3RuoGYljud0C1cbZ+ENL/eS5O2qPx4WfpXnSBGY2IcgBpGmIPxZrVTW
QNwEiHUuyn0iLkOG2GSeWr/tOtG78OLOB87qJKz9pY0FzF1BA4dkYDBXNxFutR6nMsEpS97kK2Re
Iv9XHgxhNBnVkE0SUvLKzhSSes3xl/480SShRdjnFmjNbO0ORggTvWhnCfjvGKWYBkdBEIPmpRii
FmJfnkHQlptalXTzpc5fNbKlP7VNh6xLBHWwmGCaH47BApOD84yn/GzvyVu9SSHjWeAxoSKpDwbU
vG6MPLs8x9enUulsFaHVbbfImONJGCcMNJ0NR5h66ICT7DH2d0NHhjRp6sBCr29YWiJkmMFJ3UNu
FpLIHQuvNBN0m5k0/nFH0ecHOUZsB4Ot7MQo7PSZe/vnVQEPp2Ftw4HHeab0XH0KpVfWNMhadEIx
qZQLjM2/3qbRQ/fM/lFpZgyJGl4dQv10cYwww/K2quT0CIvjgz5WcJu9tQSovgGFD09aepAv2Mvs
1FcIc0aJBVpvbrFDQfms9SssL8BhaB+Bah6f+3S61G4m3U3cZD06BRLxFLDhPQmVVfJZbu7ExVJz
Pth8W+8zalbmVV6QRSwKsXsZ4oVfNbWQNNNL8CDfftUi1KlZiyttxQsKf6us1B4j3xCLmzYGaVfg
R20kK6sLdvEcJVUJmkjgUNurIuQi1GHCAhs7p+yCgaESVc6CsAxpgfZpSJsgEjhYFPDW99OcKWCZ
ENr97DLgXo/rEYsBynp3fMlxcX3t+1TzpCAVJqeY/MB5Ob8ualvT6Xj1ZW4qLtd70EjCLhvOHGaY
z6mjEGEzDDYjj9u29PXRux6YoSNAzA5eOK3nedkRmJypoWI9TdvsRQ89yiFukPar5wtJ7/UlTeOB
HztxXWHCWbOvi8ztCIqmBfOas3pqSY6EutTpTHZEKKDyKxlSAZN4DT+9kVhsSNRrJi8kwIvIbfiN
uxdUDAHGl1qutjHw438Y5Cdmgo7w1nr948ekVWI7XKtjeqRT9O/T9eM5rdTK2V7a114tfqHsdWG5
8ozyO6Gov8dUzu2CUWw8UIyafxL0Ibbd8fia1IePljwY5f3exx2NzuP/kzxFVlTdf+o8d6xx32nb
WJ764Wj/vaZXo7SGr200Ul1zXnVyIrFwbxyEVkOAy+kK7DdVzroy//HzmVjrRwERu176r6vu/4wq
l2u8TUiJVXAc831JrB1bxbVcrhLRcOunhudHXvgzD1rM7/ItVY6ot/4QptDygsTS6tKt4FqPnBBT
6dzJILWNkvAhFKgy3qBxUkEC/GW3jn7nIbP4r7wwjhLbH3TIwxPKfnzmpEyh/WYzXUcPNyxhwzM0
nnH8BXepHkjgEb29SxTdXHd6gOd0rsgCZA/9ohdADtZMHwbXrTW6cPdGRN4BEZ7Mr1Vg0+G4wA4L
ILYH5wMEZECnSiMgTjK1LRAj20Nea+dj7FazTUfx8Z6BpN7w1epV2DdeQYOR1Hs8VASEtNa2e035
FIHZiQ/QZjo9yfuEAm8LklwDL+v77Ox6KqvrQVGBcbU0ZMCYh2laaTyp3NcZu1ni5GFSll39DTY6
NHAPVlsazb6RJZ6iNSBDoC0qSZwfQx5u4BHkCi8dyp40PMQIguIP+FJEAG0JAf663iFmVCdKuvP3
zm3HbuIuYxfqH6HmfUdL7TVp91R7JejERY/W/+ZoswlTObC6LAabOoaHtuqxjjloiz4O9tqNhhHu
FnfpXaUEBHebQm5jUXai+vW6CB0UveBKqkqPL7ZJ0T5Gxi8ffxXhAybhXTuoNyipvjScKS0AWQLm
Gf/aXJqcY+Ph/Tm7j66OKt4hksGtvwx7i6QDsV6dxvZWWiUpg2wley/MGKL/8NoqJ+SCJA0GZXZ0
ex3pZOzm8lYNuh6XQWxCKXcIkHQ58DKpltPebKs8whLPpAjfXuthQqC60lhkxoUKFl2FYAXLXUkk
ipYRkDkgzgwlgwHC+zu0WTlIQJ3yKz6GVaFHW4rvllvi7JKDx0QrlYTs8ib8WvDK1NK1Ipahc8A2
EVP1YSnXxcdbi+zPgZ5j2nKWt7/hlpzWCErjmcnvnQOAk68hFsUq+KWdFDsX7C95eK6G17ar1VVR
OthPKAN7q7g7F5eVdgo18vq6URotKDF85bbG5Yrt63J3kXNWwxxpmdDzbfTQ9ZzrMfc+CIfkf6Ws
7FtM9R52NIxRNhZaLW7IWYvsajIvoEHH4UDiVOpLnZ/qa2qbJjpBe7S5iXy+UJ2pItQ+BxoXlQ/U
Bt+C2ZgDtN+1fUWAprKjx/ZGZtMmdfmlbpSzBECGfbCTtnLilmAk0Q3/xf4Y8rUZBDy8vN26bKyh
NS1XR0NMvjOjfkYRxYjTisza+rfZaqnmBC5TWk2av4niYnoEGzI0K+Ru0U8j12pd5YGUMg8CDHXz
t8rca38o4uTM9c4+l1uZrXPuHMjxR4sF3ys4kFO/EKQiO6VT8Ptn466fRzp8CB6uZlCn2V16SD43
pXB+xag7Nw9jP6GnRj5eYGUv3MeB6ozVp6l6vB3WSNNwaUziPv/L4a+36qJj+Ub7DhXF2drDRseU
5nKY8MEBW7lOxwmJJzn1DPqbdZ+tto2EHVYyD2KtkPRUh+nEW/fqyLb5VIK7RJCfwQOONd8ru/Qp
6zf/ktlGpFTaoqBfEnu4VH2yifmUjw1zX7eOTKTksLMz88yhEuRRo+HzHIOgnhv24MfjtGLOOM5n
HtVvV9KJovIvjB7JP75qmdtCc4NvKW3GCOn825qj6o+ITo6oDXr/x/RWSJzaxDnRSicsEU0PDbLa
cDP5cEoCp8YBwr+CfSfZuRK8RDdDtLJqHDPFt7DzKhgn5o03oRhZP6RqcGHrvXyz09CY2QCK0exN
VXg6vAx20e9ErslpAHFIhiLxTFSEkeejILPvgmP8zE0h0INZxouVC48Ckr9IRUVazREWv4NTd+OR
8gfoi6EFP5pca7CQfWRopHa4V1vBFkh3D13M6Enj/1CxZoNvW39ddvqQJlYlQtc9/kqWu2PczPce
6gRByBIcU8MfSFy7j7t/sfmDrheI9Q0jg08HL/EE1I+YR04kCbBYFCOyS3gN0Rh8Ba70ul9s67PR
AKS0txogeGQa/9P1kIpS90FyL3YFbmr+f5KWNZReMngJwRIhmmdiQds3DTxm537XYl3cUB1CWwFp
SNaIf+UXdnVtZ/fqpyNbUyIx+xvyvFh0q974ePsEsitnLsBEorAYwW2BZDB7kgIHeu00R6pXoKN+
IBtSguqCwraUmkEXGsDZWP1ZD6NyL0I1HXoWobnCyWuXGJdVZC8xJmZpRdfjw12xr2kA5T3eBt6S
AmK5RhXwiYFR4J79yLUhqtIaS3XtKKn/Qdr9xELIQD2tS+5vPeHnBKPx1BB6UWYQYG1VG20O2SO1
XwXwNB/yq79I9RQudvc4hpG7/d2LpBHykdflB7JHiVeYtpqJ67tIUmSlg7e2ZVboYzZCaIVmpM7x
1DtrBynSi0MVlLUG97nlOl8cX55ffm5C0umFQmgfpDogGYuMfP7qSfP7iR/2CsNqCPYSthFOB/KO
E5N77U6GiFeKhEFvJoX44y7Zwww8MDxJTt+rDYVfIwDTuaDpyBwfLIEeH4WXrtRRV2dXqWsApnXe
K8wrxzydcDSFNvq0UO59V/BLxjCE9wRJgrWRttd0FdNIvdTCzdFyUeXJTaAQMIxfNp8RGrQabH7N
Val4O98gN1/Qv476PS+4d0TwMux+Ap6jFrvs2hMqqUtSbREBh8sPRCtT1bt42IacmHc3rUXXnbN/
pprbfCBiVWrgGQFlvo0GudGXcLv8u5om4bzu0BAda1jQ1gA+Ab81KeXd73Dl6dradjifHP0rXCQg
wr3Kt2qxzM3gESXRSYVZMu90G2Le2wJGFJIjo9uDyuLKFT9cPGEp4t1NbppT8Htw2ED3jEa/cOLf
GKyYZGuwX9Xbk3N6BfMuaA2I2vs+ggYXQN2R//Anf0nABrEd++qmIajkM/2ziEzwgjnXOdEQW30E
GlF22GwPtDzvdKfv38+pQWiyojFh88LBzRFTFsDMnAk6GBDh4a2JBJPa1cEStyd33Wc2aNFBjFti
nXMshhTYjkRDF2t7QhFsnKw0R7RFTxhJl0thDhAs+U1coa8vYdB4erR/4koivAJgfXJwive3Zsi9
RLEqFmtqIMAGS2Ptu1rZBh6odwixw7KYvFQ5iRh0F8zF2dG0JN+TUzamjxpo0fTSBWPqMSHc4JaF
NTnYcnwUXTNDVcTSYG+hL1dapebrEQXcLS1O7c3L2Tq2Cz7qfr7AU379LiqZqWyq9D0xGhd+Iqbf
tQOMfbWfE51xld/aJ/cEaw2ehp/6E2zLv1CUkudguzyafKGloQ6ygEwnK3VZAUIZTzyG1hW1pJ1G
r3oOKYjbVIek4kt2o3URmcrWaBLZkcr12up3/o5vKlc6COUcjyLwfcmDWyZmkvlrgYy1e1rcLiF9
XQ4jqKSphrDQLb0HrxbgpWyV1NsUjMwLFRbQrnocAvDGIdqLWFPUaKTbIiMD5GJa1yoHfqPlo+tj
kl2idxN9KHBVyAwKuxaAChpLCyc22hYkyy4HfznPrq3SQh4V5fHQ3ZF/LkQFwEQeD+X30MLWbb1O
367MwQ7pQ2AsdDMU/3WV2pKKD0j/mH9RmOo1ef+4ZMw/VjPuAb0YynSbeczrlO0SVgefbm+5KRjn
E9Ci+5gKqePNWV1FBGqYqguH641JWJls3LVZ0gYlVAMs6gwnUHbLUIiGqpxTB/SxSBTQZDIpcxT6
VMC9fxpY0raO94/x756fiF1nDFpeCFmRZRPbg4ipQZPI9FfUKPoJ3Penn4Cer0uEe7thVO5K73jz
rBDWu9SAHtnXe69cpbFbiHrk1g/3OZS+DrXH6BBbqgJCuM/3fA/KulG8Et2y/uyRzeW2+wcucI/g
mmVTBVHioQeSxUlxnGz/3gW0TZYtl98JnVyku4fp55RzoiJTF+iupLfPdKiQL00ptRM//3UN7cLG
unN/2E0gbDENrjQuRlYYi49mZWZLPc3LVYUk7mbmgdGQIQkahy6Z3uMIxGTVLICs+ApJR8XtMjeT
O25x9zDfxyNrHcrG0DlZ0hTxiL4Xp/8AKYBphhnugQRTAPFIgKmlny08HLb2YP4YDklNwnDGlGio
n2ccqxL79P3uLILK13TNXd7IVEts3IC1vl+yhya0nY2gHwywz0mOYOZJr8ofipgLvY35ek6eIbEX
m343VyZVFTSq0km5pYm8MS/0yeoP3Ni8VKaY7/JUPDgM4v+2q3S+Kvj+b2t1/rHWt5UfB3H87rEV
tmwPLOuti/wWP7I4IgQfYvsIfN0qnIRG/ChsPrLlCT/Dl+mOKyWOykkXbTMxaBtSUKteNNQMw8Go
k1dEg73sSQJRTdQZRxNCaKKmRtKq2QAz6CizXMeL0E8SiP68W8cvOT1F3mqzTF1Q9Gq8HlnImZn9
mkX9h72nMkIWvOJWh3L3/0pMscy/TmjBzfuYyRt/hOU9KK7zDEULZoKdkzTZ0HmGfnXAYWkmop2q
rs2R5f77f6rAGTxSyvAKihvwYhTfm1uM8gH4eOF1g35aJcd6Y8G3dbLQe8AB7Ujg3S7XHJ7M913V
wwhclWiv+y6Wie5QVmzuBlptzelnUAco57HzSWm9qlI7aElwlXPcxvlxhiQsyktLzLH3EieD9RVw
evCbap/fjmwQz5tKUHHFrg5hCr+6XkWE79MFYeAV6iSVSs9wQf2V2m8+lA9iSRohdgZIUrOmBcGn
RaeJqK03MwwF9Ik58nfaxeS6W1BATms8elP226NHN75ngJSoIdM6+iX6slZCr13p4WTayE/4BmLw
RG2P2XsVv4DQHqb4Sz883EQf5wwQZ6or6WXslnhP5BjbTHeDOTuh8YykYxZkj8JiQ//gVMDSh6If
VufuItCq9qsZ5+eNoxhNqXfifd9ZMwgHkpcnN7vibpdAaOfqMYIb9bI1ITLxKBsDkUt8G/Ul5wpb
23rNY2YI0AksQrABwlKxOKC/Iuq0D3ClEre5uIZsIvsMzzlI+aJEhgzio6aV5/xzV7uv2IcQF12d
s+qVpF34mw21jucAO5rOCavc9NcCCfn0VsuxZg9MS5aUZtiLga0nMjgIwCkjikYhAFCc2Bpmwy94
KDObFnnSGmlOE2pfP65VpM3+vdzV/1uwHUKux5udMKTWDe9E76gJknEmHQBnldeVqZpnp3VzAY75
sXN07v5iULrHdC7txOFhlzEgjb7v76dVn5YK0oK9OyxLVWWBhGf+MfLWQkIHTXcnSveK8j8BQcNn
mh1TgYxhAaXv6lxST2a/uZ/O77m6EVQ1yPChIWR5/EqNdMOkGReOofd7XFC0+4TC4H2miJL0m0FD
hybPsyoQEj7jyQzSWmkCW0NOXACGUQOmR3yVUK++IHTbBjmhsmEwWkzL8ZQz+emDNgVYn8GRuJ59
JOTF6sOfhcLL5seYKZV2xYA5OqZpcR9n3+mdWnCxK5ML2HoCUsEMX3N4SrwbQgfYRRTv6aVMUvC7
OXvb7hNU8bBoH6eH8RXyvJDLY/K4BQry6GGmrWXLV66S7f/bs+7Q6tkxQBlQpk9JXZCnmf+81p4L
iwuoK7mAy07ffayvOmrAcDeBFu0/X8TW72WxOyAi+rzvTWsvKkXXXjoWPFfXaAl+e9eqerNs3Rzy
DAnevMWNt3bgMCfRwT2lpzBB9V+XxSOjFF24FYfXSqFS2IGKKLt7keDC7iLnfzoeLWK2l79r5W9e
MQ5nIBFJjqEh9ilnCmvDSb008YlBANYbAdfvut51MA4zEqTbLn2n9A4JS89w/XAoIryO6W0/Oqc2
YemCTJMmFr5CC2KGYznF6c8qXsos6r85Qvu6AqBeTrbTIZjWjgr9EW7oq1b76wlhzG9SlAvBPStj
hpTDVyOwDBRXEF5L1BaS9Xem1n5+KNvYc3kXjoTkYRjpXj7l7gLh5ZBP7a0QpPTVMmma15/Rxvp9
xl6jMMRFIfenBHCdF9bjQ7T/tU4Addd/yX0QxUZveD+dIsJHqyHzNqmwmUCOuWpCT5kI2q36qbdO
58RK4QR4VPsq+gsL0lIHssgQXLPYcrKJVWQQPn5qM/l91QopiKdF7xyWOVV1Nwp5nYS1HRAdXMgA
7eYj82KvwpW7KorDIpBzSzMV+/9fOXIktbhv/guIfwUlF5GmUgNWtw+bdJCGIeahA9tAKAFKTesj
Nczz1HLWGb1P8d1fC8u6mP8zC5BO5KhgxvHXKahQ73E2BODa8IN51kyg7lbeaKHVNee7phVMGj0Y
shaSqFfLHbN5jieF80Sa60RFbkxJKgEfAcPNYBwdZwjEHlPwx4hGgSEEE8lbKt02FDlUq99+6C5p
sxDnWFf+XvQqAzJ6dTZJo6YQPeIzu1fvMSg3jv1QidNbzixcEZCwF/2pnVd+Y6fsFXmyAFB4Y7nn
1W20nrHZBaYA++Gc2rOw7iBBGtXvBXuvvNd4V9+EnTQDLtIpcO+nSdKNnNJqwDE64UD5TUOKoD3R
LyxNYSZGyHaaOm9pmPAj0x5ctbJtVsMl5TjPhGV44/SDCK/TKRwy3rwOqLiCzdRnBatN5uIYgDG6
vpwSdsuD6aAauhsucIflLCRk0AH40vZIdpXmRpgx6tpmc9gBe9A3zAnYMt7jllC7NXlwg4UpPoRe
3VZ67T8enG0j4w3rC16hi5ud6sXUNVH4mo9NqMI5bXRBc9L6wjriYKnsCmawH560iWEjgDAK0dZR
GHydmTvDok3wIgjqu6K9jnvboUa7L0n3R1aEFFV6JvhvZ3dCSsUzNV4b3OM5dIyFAk+XV9+5WjAI
ino0D7EmiW9mzFrgcTMC6B8AL8/DSxGGChk3Z9K8XPx52ypuoQVIovKTKhkbS9i2onkl35Yosrxd
ntIwxFxk6e443mAxLBzD5YdQVCPyGho5NEi9uVtSlQm4iedIM3dtscmgTW4EOudY9YqTb2dYm4a/
/NVl2Gfpd5lfjzVXHvxb6pAsqARFOcbQFbZybGoHoM7BKjQkJKiZdwM1/A1iBqdTy5JmRQ7b5dKK
kfyu/oLUgUrbIAP/HUCW/OCByRi/mIulqNLQQCkQP1L+5I+WTmFR7r9r8wCjm7QKQUNaPa3IRrd7
ytsKJtA1LvPLO/bnWpNxPEUhOq7+eymHzSUveS8TXnEQfsn6eGIbDX2KTOeXrslHz6x9Og13lYTB
orbog+R3AOnv3V112ngaUiC4yY6JBvZJQGS7rK9ZC++XPE5ioIQOQlNuk7bsoCy1d30Ra0FFlfOQ
rMQIfdJ9VJcXKJT38Ng90lrWpkVuovnzN41gGktB7+Thn14eGCWP5IudQcSN/YBei/Hkwo0r1Iok
f7e8yiAhpqOpjE2VN5ndrEjvkVKpVeQD2Is9bSc8ESBs+ND1ldewa+knJ5xJUHOujm/cRodStmqm
pAKIcIaqMP34+E0qW3WTkOI9Wvby4u/IbDpVN6DKr7KrQRaUebi8TI1D1zuBYSixzxLBUZqXMrQQ
iLXag4EpYlZkrffJ3fnlDvDG+3a0S1kjgl3ZSiJ8U47NJgVTm3ArG+fgSHyplLCEV5qvKZx8YpE0
1e9wbANbdbL//Dsn+Cyp4xi+VJsGH7WNPG/XqMi8s98kunNSIXqUfi6xpGjCwGEnUNa1zb0CJtDq
2sIXU/VuoD/nz+ZhKDPPM50AAYWPcR8ClVtVCiLX6sjG/qfuag0ejMtXbUOL4YqB4/JZ0PDapWKt
FIdRVveHUXSpVdRsoSTDGzUJCBdpDM2/WbhOjBDlWXPVS3QpkJtk9PQttyOY5ZSovRn4HfGj7T2f
vW7ZVKzR8idvt+DjMjX5oLdF0MGsSG4/xHMMcBwpcabebMl3coCw9X8bwCrOS3IrwwfJu99Q63pi
3vFdfUPDJQGW9V1nglFlX1JagOtadid8qmVifOHZD0jnoqC650quuKfGlNP0DXHSlbCF6kwuICCb
MLprxhMt7XE/d+IfkzZA0OgDFUWHzdTgu9tobmxRC3ENYaAsxegoZcs9flqdJWp4MnFMChyMmvbL
ToaIJ0fI0mJLoEBxQc+2xwFoRTSGVJSDEEQzXFXavw926orQT8D2eaPgZWJfA2TDr4GjdWLQIie5
xPMKW3VoY0JbE3pCHhnRvyxwsk95SoKJ0lTLEgULlZA4nomSDRpGsFdchOFqQpn/51NOvrxUtYMz
6Uugu8bSk9+527Hzy4nrt3K7qmRtifeXN4YhU1JXUW+Pq3LZmjoeOig0K39ecHxXYX1bjZzc4VUX
BkgS4+vCu2UDNzOLpLlP6EcmfTVrQjVgeTrwomO1SSUNVMKWjN1BIEuT7PveBhUsTKQ4S2gdKcir
K8N6/3PwotmbzktzQcafV3dBB6IdIK5H0J6KphPB8DVWsLYvDRnx2i+2J7MymfBwIPilDV1KckFh
mMgU9c+S+bYh3ieliu5/DgPf7qxsv878TRbEho519SXQNIZ9bqOw1oRULgE+o7721Wx5GGfwzrcx
2SjR37/bGzbbTirh5TmjZPe4lzq5iFLnbs/VXXq6WDhSN/Y2JL0xZpWusEE+U6WLNSgrHNRr+rEE
QJ5VL+ODm6sjPA/GDMM5uJUq48pnBVqkcIOfsAmGwq0L3Dc8PSJ2HtoUk7Q5WLx2mwBsrXZRu6M2
hKRT+asBpeNr5DQLBgtlXPXqCLfTphsu4KhekG7PvR1T2gQi7mzHIBq73NCxZI7/wRsisKQ87fQA
xDLNy4uPuc2kJlSN/upClXhjOR/02fhux9yKhELVjYHkWVB234qFIq3YdvCNUnf9bA7FUuvNFUd0
9O3pESC3LQUIKqmeD3xje9Qkv1jg/TzDZTMERard7V5ZDZwbYGKQeHxqmrKLtxujQqqj6aqvygG9
my+bqlP9Prn+G9IOiJXsbJknJsFRD1OUHJANGmFBYH9qt/S/38Y+2yj0ypiyCWP1bHClHWSwUsBO
48Zp48jvki4Mjaulf9k2t0cGPmKr91mbB+E/yZd5U+t2kktxFexB75uiYtHzLSAIKq+ThzhPAx6P
HaNrC89fdKTEh0X/45F6uMh+yPKZY2roQkH0rI7ISFw5kD5Q45YGCet6kPuELwjkgCsismmnGDyZ
TpDWGYOVEzGFZOtBlreBuRBVM3NzN/yJg8yCNZtKJmTLnDpO6uSc2vufPMRRRSoYZ94HtoWOWOBV
gsUj+z8qI6dhqXByooPdG8VWvgOeGRnnlJAZMxwvBA0aUddRZNgBYGj9I7QG9aQOZTbLh8f+1LI0
HXj26d2Gr5dm18C4m23utcJtGhN+ig06lx+qLSGmEydMasZo0c1p6j4mnyQSzzCxNo/5R68FBvY3
xtfnm2F70na13Z9lX3zoqk7fF+9S3p4fQ2DCCnvyfc4ZYGc/9lar5qcNZU7tsVoqXxxtPf2j2LDm
Ixly93gGEsRUNiXWdFtexctCR4yPPFDT1FIeqzfCl6PNLMlIscCwSa0w+pfn0qiRBAspq6VU0OqU
cKnHvm2bzEl3FHRqpwUcPJ/CgpwGSeA22PmnZD4Q/7dbRcy7tHzE386008Y/5TwNhwaOF1pap4nG
RQYq2gaSKuIiyHsRgniAv0gTmJZJRmXNMa5fgOqND+CjXdEgl/JIlhXvi1en+8x8Rj92WUcfe0xQ
XyIiRoCxOsKiVmFdWbXZTKcnkIfBch8UU2ndCvJNMLEUcPO5L7xQRDtSRRqgeV1dejB9/9eAzBtE
B98wW/zBRyIbNQeoadUu1raN5zITYZtPzvw39Dw0GaBY6zZ6FKDlwF/9sKVoj/LqgbQrB1Dq/cr4
7ekreVLyrsTtVwcBqZnsR2o8iUSk0AusDo8x5Q96lw+OaPcIrEI9fdD8GTH72ZRjfHN4koW81xxQ
bRvcWYHHdC4+RMI4JXDZRBktShyT5wWPFi04RAFwIaGUEEUMYJxDNITZueYIKhte8y2VDWXF/Zb0
HvaCAHZrXm9v57BB+o3DrP4q6kvuCpbQoQMhSVnU8hxVd7rgroC8IDG1KsHCXvrWdAQeEgJQKuwx
FE7lar5pU/RX7KR6BEbkGqA86OwbSeOZqELEW2hvlMNWcn+Kir5bEdCSC94I9c89P4oj7YJVCq3j
OAu7g+YM8Cd+M4O+1BFRx/Xtp37WKUxsHAn+b9ABQ0rTWv0QL7lHbSUxCewhnZGKpSr+nurCMqZH
lu1ne0G0eCfi7oClrmvALcsSKjZhhKePgdLX2bzmz4ioL18+HNKuoVGOegEwrrjhA1LagKkH5Zdw
M9M11IKGJzTw7tKSRV3SwGj7XBktBIm5hua4VMDFF1bRFWPmMv8Tt5Ip3SSvhU2DVtke4xz/Ddw/
pjzTzxptbzVSxaM/4CqOm4yi9H/TXvp0/i4sH15LBAMK/FpUwZxIcbMdTd+hmqhUZ99xwmTNmaQ9
5zaf2I+tpFf/TfUe2ovC8pzIwMkq2kUqwV/U0n6969KTmKPVtYnFSzFgTBWloZProg9rRr1z1Vww
LVfJ+J53WqMAsfzG5z17XM3CbxPe/DN25aN/vqLgwbtVe8vvxFMSNgr5InvHYK483Afv7dzcjYMP
A30ZzP33/+HtI7PoXFzbsUctJ11pHTBsCNFkZ4kFFLJuNEUJM8kMdJUladBkQLSRgv+hGf8XdV3j
YH2hRKT2ujit4oB20Ym05IldbLsmRLgBJBHn/HMD9xfh4YSke1ud+M577gSLGIfCl3x/VD1HfL/7
wNG9vU74dMDiFDSE4yiCQMVfOQKEIix9lvykomrTydY6E2oQ5v6axnfHXapFAMLTDO1pKsrVAJ8M
FdHScUOpcHwj0zOM83ssDLgZHl1rlto7AmlnfTLfDFhgnhKtJ5B8Eg9v0bR0YE9zQHTJ7uYmMHet
To+5X35VTjYYCQMrUKzO4OM0L0j1EHzVIHNsU3JhiZtupFvi0yWAm9m/xqqXUFKK5y9GOYHDzBmp
ZKDQpJ0wAY4/b42KxSoqT39vMBh0H9mKfn3pbQnlDaanREBgsIudzWt4eWOu8NZe12qB0reFIjTO
dt/dK/4o3PRoQBrub53rwq1F6uwREx5w+tU6mVgRHSZzaykX+J4RSblh4JZxD8IhctnWKQFlw0A5
Ai/L1FAJQTOWDgbKm7WKu9BEtdbH8NTfFjxwr3TiHEDY5URghaB4/DuvH44QJolTayqukwTC8DmK
dXBYe3yJQza2lIOUDvz3ICiAR/sR4iC4dmolO4ttsiq1E75ANzSyU63rA0peib8Jh5U7hWJBSero
1ZfxHNRRIy51ReLCgwiOaaNPztTaNmXF2/2TTgDl6PgdKBKEqAulZaNHxRlYKT7u/vJT2I9cCno9
N/mPfje/x0gNqkWNbNtiNaquKgsHGCNdZozVQSN9ErSJPrbRZ4ANGttX+Zq+leJB6ohe3aDv8S8H
ICupr8VI6rbkK7rTyJYU5gnQ6mELNxUY6DXUbawzQdUKko+Wo7rM8SHMhTDsf0wF0e+yvQx+QZvF
Y2sOzHxLoaIKUDRMGBqsUoRcUlN4SYjHYerk2IO+9IunJvkiK7Ssk1ZPKQgc3VJofEImBhYdfDDA
Hcrc/tes2mn+vq+kcWeCM4lNDK39XzUjXDHPSjxhiAPptJ2U7zb1hzyiR2KdLG9rUltE0zOwqzHa
fg6+HX6/3Rzjf+dpP+yuBVzptpN7nFPiY72/CQrmRony3Iqq6KdF6mbVffUD1+0pVPmYE1NgijJx
PBHSMoVVwJEaUWAhpS/oVSac7jEDDtwJ4AszPl9/TXLN2dPFX6yr0W9lBc0lZ7OvZjaHUFuNzHgJ
VTnMzvpDahyCBu5BkMGpfGLBTHn20N8jZQ98weIBhB2lKgEOESWG1uMk5OnT0iOJfxT16woBWDJf
s1LmCnCT3VvbQ5dmDPNU8Z+w3MUcWoMGUhsBDRYiXEvqt4XDELKG+wOkpt0Ic+UEbIUUqykylZx3
cveqrR/i6+xqc/gSu9eZKEVsOT+z+5Z7/Xsn6AJKAmz/ezIkaOiHI9v7jj3dROX7SgDm6KqFLjiK
JKhw+j4yz9kYJYzkhUaR2YCgc3Mzlh58AxReWp6+KV9vIZ6+5AtKNcqRvQ4YOEUukoYwsWt9IwWP
TpBdNvutJzjyS3qqh21LOY8ZsYfSGeWllaRpWO2UL8OFnQV9aAaZZq73WkbeBmTB6B9pbMIB7JBN
aAicEC+rX/5distR4EC5K1XJ5cuDwmvqtnSh7+CII6Xk6UIyT5i2ia17B4ghnL+Gc1mNDn/sUdme
LtDzBDsOyOyLAGQx1IlPzNAfAvliks+dhsOzlwwwI95uWSGvuPvNPg4KfeT9f/eZvkhbG3Fg5qLr
pahqSE9u9BY2KjKPuOndM3EAkXrGU9eRmHQbh/fu82HdNYsr3yMNkEHRj0Q96cWloPD42cxRGpei
3VWMJstBf50I3nUCFpQxe8jCqY1LB7DifBJpUgavEUnGV4CCOZZOFj/RwNW03RipMheWKq+NZnkE
wg1JYAUi1B22+i/w33XozMH6bVtRpSNkTDRi3WKhIxN99iYqobXTY4aDSqefI/ytv4G9eUDNp7EV
cjrI7zsup1w2ExWUNGSfr0/jiI8df8k3etrjLYY8iE9KxiwLcxOoXUV201cFzF8kUDIxp3VzVtGS
E+gJj3yKognvkNt2FBxx1awp29w7BJOo07OE8+xCm1fwfYhxbJsYh6hsO7yu/z6UvnhVFymfNLfR
qZce3S/13MyYRIrIBxlMJwJPhVZDeXJ9enUH3B8G/DYVOilDGZN8hTXZRa2w3ZkAvtQ7ho3t+BTq
vHG6VrwIwiCTUFPOL91IFWz+q8hu3R/ypGTOo288JFmIR0wDu0vfI2vkvcOkhg5sD4qzdrslwTEP
/N/QDuHUOdRZThpl5s8ReGm5HEYdGESz9wU09NtfbiUFxKZbkzjPbVDnur0ABRF5by178ZeOz8bJ
euv38mazyJxvdjyXlUfXMeQkWZXPz+BHCe8scWkGH8gXzWkBAO0pi5YdEweVQoknznwD9HoloBwu
XAgCmhH2gO3dDVqS33lVcaKwQZQjCDITCwVwxi226rqq9zTKY1WAlqG+l2e/KuydPS2GQtq/8U22
clQDkNPDiQ7zg2aQA1oMO/rFMOlmvj/hLP3TDRi/lujXb4N5gV4W9JeVrhBl9ccgglWDf1CCBWEM
FbRjRQ1l5jp4dokhtsKEN95IYQOqSpWbH3/JsdmzOuHcBUnBCg+anh01j5RGMFj+WBms7b6zYO7U
liJaVbR70LVM56K4bN0Ex4OvEPWMPtSFt8Vvtm2TVfbRM6QZF0MryIYWT2aMDDfUDiT8vKyzCJmV
i1WfCDDQe0hbl0dT8wmI1IrwLGmAD7EXbFe55okKx4WXkRhA+6HFbswIB5UEP7FQIm4d7zCNjPir
8Wu/qnIsThkNlVj2pjk+veQf65MF8xZ87HBVWsrfCy/+w1T4yvsh7yYJR/lkJeYVxD47sE+/EqH0
EOr+kgDc0NoIxI8hGqgYfUL3leZceqrhZgirPMCdl/kdn69J2TcFNggfEOW4SYWLHndVQ/0g4HRE
qDZ+mqYS6AMLHq88QATZNC7ZDZN67/Bhe+VCksoRQgJlo6Cf4Re/Zijo+sOvy9RT3GcP5ge/9i97
ct/EpvPt7/H/V77ZJ3iPa9NA4qXZZ0/HdqLhjcNoZk1y7p1OoKVe/Stc5/owPzxvb6VEjhfZR5gq
r0A7hD6dPdeKgw+iWeF8hNDKpZgSGokhD/OaiKAnoiCzan/gObHGzLXLEB1IIug6ZPOGnVz07cC0
T1JeoCMq1MjTDFJxCtgQdhsBdmr7NO/I099z0lmzEu5oe+fouCVLgb3FfVMItCzAXpmy/vmAAC8s
NEPIPzvvlPEv1ibqUYFZSRv7K4+wy/r9EIJJp2aXKRWGIsI1fuNjpTlGeR25vM57YuOhlhChLALU
8I2VKGOZufiJnbIwCK7ZBFw739ds2SiVLGapHU//EV8MYEvQCitSLMZEDtT1sB8RLCpI1X6BN5Ww
JW0LBrdQRhqt1UPPnAuFXR+sA40AAmGrxWVHd0L2OAHqQlHYNHcCgYKV0nqvbt/YagRK7PpB6F6s
aLYrGtdN5juqQqU9b3a4lpGlBZD8VWUObnG2DSauEFFcLYn/Nz8qJB95J/6GMlIPYxPOncY+adXJ
nywlRtkTZEcgSYPe/13/SeIpGMiIgrSiDttFpcOFRKQEkat+CHjpLS0ewVVuFE3zUZL/NIy5xFjd
frrOBPTlvcXqZD5HY5SybTJZfe3r/86Q5IKhY47GICYW/umaYgAGsNXzYSzBF5lnP3t7pzM4Fz3k
2oi9FE1sera5GTHg+j9LDfWARogbHPOg46s0PwN5K8NkYSFsvHfH+ocuExDky2EP9jA1grjcIzSW
HOakjMFf3xH81zhATetAaEoHIECYOeDe6WOQ1YsoVu/6EcblPuJKhluxDvCfHN5Ee5xHIhvFRSb1
M0/eegR8HRkM6Qs6+Bk8S8jztnHepItYN385p4a5O6VurvPX4y2V/zF17hOv2JMeLaQBG0IzYydL
bHhgO0K8R5f6vfI6lugudkQrsMhkCvg7Ts+BiJV5B9GHkez0VfCCugbpzQEarD8MbjAwmtGH77eY
c5MG/P24JWAwt+CbCsJiEPck4aBmUNyRv0qHq1vTgtrie5iwJAJJOqJrv+Vnp5NFZ6IRc4v1P6Rm
lBlS86Tb18cbclpC7VCXtlsQZOj1TtP1KLuOw6VafqTgiwGjgZ4qkzhzlKFPPf2yCjDbsUHIt3M8
1EU57G6cd3h2I2jDDQqZrXJzWfG4CMKlBc7gSGj9CP6IAVbRPHrpdhCTIiSbXjUgs1Go0YZXU/D6
6p6uVmz26WHrwLY6HYDbqMgijQm1MEFl7aZkex5oUP2ZgXzFb4X9Lq/+qeekbkRwt67CfDsuu+c1
KJGmMbbUeXPVfEdPiwWPrPxGjI9hFnHleRNzX7P43aP3QH7lThjggGdw4kCq7H9L/88+EJFQQ/Xn
B+TJk9Fpb6X+tNNpC3pfBb43YiEkMoba4ZS4myGfYGJqW4NrNiQ8aShle01vLSiOlWGUEaKoCh33
heOcuZ6mXzxTUhzwWOikcIST+BeIzeXm2oyDmZnVI71B1mjCbDcsBdoKsuzA2Po+z7fDzXvrK+KS
z0Ycsm1loWi7o6edJC6s3I5S/Hcyq9dunTcTP1mZasYgBAszZ6qSKTFBrdMQnrfCZdv25H7CZA0m
+zG3mJUIscU4XgM2zZaIcrZYt7/oNRziahXSXdiaPwz1FPsAgTZBuvgOWBrqUJpUTC4m1K67/DG8
96Wkw04jvgwTNfexaJbdxagIBQyLulZsX8DcaXz7IsBduHTV5zGAiXiBNLxQoWpqhFkPRZ2mhRb6
XLxAVp+GzCAizs+6nBGEWGq7VAQrjnK95fNdr/q+wfAMekCaJiOo+uh4Tdl5vd+amVt7JGVEX7c4
KYqGop48r8T8hNWOGSj67rV54CdQKe9UQsb6JyVlRAshmBx32D7cMZ71AcS4gRg9ma3KhQnVrwma
Lttnu3el4i4cIBU0KNOZWdyVlABA46NpC+CK97/AQiQWhE91tzbJCMpndhm+3V/n34lMRb4qV7gi
VXehnOXgfEGbMeTfbWxkKrYXP2Q1A6K1NxGdZAejZp+h8YdSMR26YrqbfbU2t/xRVUsTpuG2JFGf
2p1wM0lh5MG+Q6uuAHgdNaYvTcw4Ig06zJ7e1M9O8gm0O63L7+fr2pDXaj6Oo2NeCyPvfzPXa9mT
Uo6pM86IMn320PEdP/sF7pgtbavgMc6lF/YS7c2nLceA0iESr6LSrS7vcqS3JOSHlhWsvFs3W8db
hXDyB0K5k5GIc34tpXrLZhWBAOaiu2K4NqXZ6I0vjeFv4GDz4AuQQvr7HM51JFQoEYnA91ppjpJr
vJqt5bCPVa1G0TjrLiHxmrumu8agKjfCLI0FRt707RA585jk6TCkwOciUktsOc+X0Fg0vR3icP1+
8OLMWzyqF0zoQBimmSmunMy+bPFa0yLXaSedIudf5vhmfMt9SntgLeHKYpGDaUOd8ByuGicyj9Xz
GX/BKpfY2bJPnd7fB+Ag2XJhUW9br7NVLzBWMOv7SC10Tuag9gOhLf8DC8XjPAuxTxlRBthXCW+9
+DtWIyBuJjT5PpkapLA5ImtbMzk6nftKlbRV7iYysuerUvR0sgCoBglp1ifzSKxxyAJFEnd0g133
2HJmb860G/1w7cx5dVB6kjeMKovXdmQRtW4hrTCM/5NOCNwPlGJgN593lUYBHxTYgLMd89JR+VB/
8LFb5hGeUrZ2t8yGju//DqTmlGOFz5TbWyT8ueQ+h8b+nD9otn2JOSCx/NwA/pIOf5I4IXe1J6Ic
Gi+KmeyjGttAaZX9wg24WkxyW8H8EReNrSPyudj0WT7koCgbompM+TL0I3rbHHGf5mFRv9VQfNCs
NUxdE2NnYqEU7SMhF8QAQv42Xts0YrFB8VRQhdfR5aGPr9URwbVyxdQKuMa2/xN18yb9PkbYv9ny
GVxUtfaCmaDQ4OYfTGA6tJBGhjaRmWjlU9u6s9K9i+Dtp5JjXn13RpCLI1SbEv1JIYoLko9XI2qw
t+nn8aA5hYoYqMm+UzcQjaSYeouuaAkLq5VwKCjPsH/jL3b9b8EX2Uhg8z94c/3z8LL4xbchuZ5c
8GJfMB+35TOelbMQ2EbroO8b3F3AT7EPYbJPn26rHwMnUfs0hqV1loNf5qUnqci6WDpJWqrnxRk5
G+niDXXWD70BvBIr5TqcpWWHNe/vYRQ/fQGZGWmfBnVE2Yl5v6Lgs3lc2aqTRYO6H/nbNGtjsv3H
6vB46+7z8kzpP0Z15Bl56RJCJVRzFR89ZWIGVEbkKOcqAih8DyHJaMbHBa1jcgB1mRh5DArrJfXd
y5Qdb6BPbHj9OfZiXSTbdfMv8H+PUaF8eVhFdHzoOutlitjuAuAoJLTlf1i34d+3UJ5MnZIFlShh
v+zKDeMM3c2h+LCn4DWhQfj+5ghbS44wQSKEdLLJmn9ip18ppd5ZdFHOR2CI7/8riy8W06jOmzgy
VyAkKZJiIFILh/HGfwJmc7axFttufB2p7WM15Cn2BJ+lQCUezrReRdwC/y6n8UlwlJZM48bjE2f7
VhmE05Qts7URfiK9Lxkjq0Lv/0K63ehYjWAGuqEIZVJqJmml4MjKx5Q7zrVEQZ9W9inHg9a3x32v
spLCYKnoJCYfQy7m/13utFiGzBvSGAcjtS8xinaouEAQ/GhSEsF8d5k5tlmoxkYNBX1/5ifpH6KE
8SgJWsRYEX1JubT475tTK4l8OdEtOgdyJmqnqx3/O+p1SGJyAoftapvuCZSKrBOEtCWpsl1Zlddz
n0ff6pQdOPkokZDC7bWd9awbGMgWGSFFqg5bjzpPFbnOE++7rex5yHiVgo/pay2JhgkBlK+Nbib4
dr/6HdeyxgLY/0IS7AOajOjMc2J3IoC/+UlqvURWFgmTQBZycTV1GxBi40OxvXA1oT9VNfiPY/Qp
h0DkuLTTfmgCholNNln3n6A6ULkf4nJlFcIPTEiArlWS2E/eNpeokC4OlPXEZ62ih4xM6/eLi7hZ
aYFwtHK0SH97/a4PQqPP98IY4BA7+No+Z6T001Ze6OazDAP9KpuFGNHNodYwrq38jHZ4nDbqIYpc
QT6XBRdCRnBh4/As4vaqR2dZz0IxLUZWpErkqQ5PcDC8Nyw6EwPO60TZTsbnxGzcAa1Yj7LAPkL5
518oiXaHx2zqO2Sn2Y0EHwnn1SvHXHqRT9dGXWYKzrHAEH29GGWI0ixYGSj/zp0GXm6GWhMLqUgp
mPULKmTG2BFHgiQlZA0YTTYk2WP4gd2T3nU/LHmuZpqjWQSJ5VIKBjEysz7jRMFKZaHTH5HksbYs
gc50ikyn6rkYpe79C6/iab5YUpSOnvB8vvKS2O79TLHAN3fp0xkz9vqUWEgBbGPvfFA4NM2ipGEm
fJT947Ovw+Q/gRZAQ773W/3YLPTrMQyPTGTu6/5spixNV74vAqTKvTP07gnQPKis7FtSmTiRM7jU
Ystb3vrvbaNyWjlfdtcaGk9dHJWpQy2+M2Qkp2+TgxFdccFsudC6e7uLyAiJaK9N2XYqcqzcxvYk
Sd5XKKxkfE6soo6Vmgl1Q4BQVwKnNwDsNuqolaPWWk7UhSsuyyF1+rnRfcQNFFKrg4Rze6F+lqRa
ygHsFZhFYt+lewU9NSybhTxtKi6mdDmDbnIOYExiCOzcxYL7AGmr2VaRuqatJ0WUh5Lm1doWAq7o
lYLJ/QePRdlLPR53i4FuCuv02KJWTndVOwFL9murusu4buDvmLf5ztpFWvbm/AJub96UWFPvhNkr
FmbI6/kRzux+f8BVtfsV9j44P+Hfk6y0GsaBNv8bBCKoYeh/K5BjhpeRjvSlmYGSq5JNNjTffPb5
JFFtcoJf8urdFJtvMEvVU7/kJ2z3OMd9S1yHYh0UHy/eKBJbWxlTO3EKdc4w3WqaiCN12JbeEizW
ZOJ/QpHejMuFsqon58zHnde5mCeH2DmBMsqZWdIWwS8vXwgf9avksSHHWzbOXxZ8F4Nyu5jRBOGu
brAbgYix9EiXwELA2SoLGFE+BEjcmkk3nFSLwlDpcDuvBeyITchl/gP2qsG297BgN6zaMlu3NOvA
inv6croNQlanX9Z93hyKjN1X7UNu8+2jCApeFHxAyEji/pfAmfueZ1cCIRlLk0lXKqhL9OEFr9bH
oUDItZSXC4eDh55li6Tey9KhYzBWig8BNPDUrsl9O026pDqOM/weqEpqjHqy4NBLmTzVNdOthv4D
+5WtPGilwvX3cbbMGtJdHT2XZlk9aJp69wYBBBFLCPDIaCPbVNOOaFcVSSxYFNHc3yEONpqssToS
B4h+lVyMVMzfUn7pY4ao+gpuShM+JcmFgod7zn8FhCdTRM+F4DcQkRjj7DxPYKAzTgOF97eOISgC
Uwwc/XquPg5v8IiUCW6w1eLpZpVaox2c6Iz4MC8B8R2zbvP9VmUpxPZAPLpn0aQVywPUzVaAEbqb
hJQfJSX1KyqIx9CLhaWptk/KQtm9MvZFJWGTK3m28Y9Z7424BxV3knD/5RzzPMS55lnX7wlcPe+k
FFxr8VNL7ku3EbYjCdERi+1EvqTDpPppSv2dw4Hy8nSURdGhrfTQmBIV5pHXAUK/r0aYD6KmBwyY
cNyii+m57hoTTzBLyWYw6uZTKevC/LkBH+lY/X9ovv46qOkL/BFFQSW6XLDHvTLgRSgJUAPPLeyl
j81u5CRELQ5yXRu6wuMDutLg070FxNHzsy9RxyvlmeEHBi+U41bKlJTaKoLzAvlcC3lzhLY2madN
8qJ9nDXKfvlX6ABgGqhaDHG2UmzKg9hwW8L97MwcAScacyiOm/ZmsMpX14nyS/kiYQsBfPh79eIv
+e5+LbYDSJGLpolgURuEl9k5Gwb7misZVk9pvh8iXzc1UaoUFz3mghz3X0vHQ0XvedKKW6bs4JaB
QbFt7SJBzWCW0j6AzteWhNndIu4MYyTPduVvPkrDKCCapxp310KlfRdYgh4K+aanm6TLv/LGLCGC
aXJWIoy+FelnEMyk09xNFvuh8WNSTz5xqoIiD4kjIG+spVzhJ0DxFTsvOzMFkuLvIUH0UnvvFKaG
xy7pOUrkNkWD5vKR0x/jvzbkz2uGek0VcQOV4cXceB4JqT+kED1zSpEu3go0jugMh5amj5AKNI9d
3eqY3YnZrSPEPMlYRQX5KcEq+mpadg4vRCCFBwtWd7CqRrNXm771sc/BmV/kD2nPuCUMV3gqYM51
wJ+XogbFmQppunMqxLcyC2/ZQ8VOe+gxBLEkpZ/nUZZ+6AUKejC08oFnhB59Q9kLi0sKhlr88Msk
fFxwh0MUFo8D4B8nkXDRjRzHAgAHkU+MBEE+2gJejVxOllfIAt0aXLGIo5lH54NAlDhdlEwiNpho
zVPkSk1nQCSnKgd1QAAfcMOTmpIffl14CEnL72FAxSWx1ANcRjkpOhVXbbhrMG2FzYnEBZFAG8kb
Q3ULvrC7EQqJ0TAt1YgG2PsZV9wuw2S9LctTgXyQ2iloRumkP3m8FweHW5zGUuAijuBH+7r542mI
1BokULzpvHaz33U3AwUaFGLYv95aBlX/evLos7VXUZCzFMoc+hUTbwaCZxQdoWiLDKG2+sYMvLJJ
aOdt2MBb9OWg090M/iPF+TlLDAIPF9Hd0C80VObSIbIJpo5BNXZY3BzkAkPm/PjXv4T6/XrtpOHE
CeWyl3PaJ9vI8NnmqwuubLhxbFtz6/lCmsQ7B4yf4oU7OPAIO0OHLsCswMZx7Ebl/JDoxT9XJDK1
BccdTi8mjxciZYnRQBRAaZg+h7RAiUW5d1hxiVMviPW5z2d7Z7cqD/OC/GKiXQw9Iyab6FDuJBAe
OTZZuFW/v5XAriL0Zarlo0eUeOQBImqZ9AlVD21T3IY/KFY4kITpqdk/0TDZ3fTxHyTjpVyDeoPw
3vhwuy4OVByPUMd2nd3w65AwxXXyVkJ8Bm9pRdUokLgSlSRbhZBPiso5pRtUfs9Y2dZLn5KCeCis
kFo7tpU1C2oxwQkEwwSuIz/OH/H5mFn5NBbGUfOGYNOqhBw+stcx8p/7q8uox3nkVoFpY/eyJzNN
NtHx6lkYow6iVUDZNhEMmR9DP7DfZ4ST3ngQpT+DflJbPudxEWAaTto3q1RsRu+IdfRp+opn+FWr
f3xImc3BK7uVsZUZ9nrkYVCIY43x8vTVd5elVvl0WVJ5+xRmGRAYtmxz9ALNUGS40RO/Rk8bu6X4
1FOtXNLwvYXttw1SgitnMK1/sjBQbN4M5eq8hK/GtdX1iCRzND5tN29FR81EY9FAg1Sbz2i6jm1V
192b/nS3dLKZ0/CkVH+9V0gB004O/E1chtp3VzxXvCBSfQqPXDkJjbMUG1jt/cStl6b3nKxSLEHH
tzXWvc/Qi7/dQzpbYKl0bzolekS1PaNK3djlc+dDdZQxWKsxymQmorcVkoa9NbrdRxq6rm+fojpe
TBuU5inIi+2n6ZQx1qulf0ODMizU25+e70L7Yv5phz6zwmD0qnhfDnMgol5dvm/w0ZlOdsGv1PvT
qHE8k1Nx658IrScjB2+nqSxNr53C9icmZ5lFZCjh4bVlFSQhRTXuDg4GlnKX+yWtinjyUR9Ha7h8
p/6DD8i6kbDE3sWmUKcc4VxHT3rslWpj+VhTXKLIsBxeS0SkiTNRthjQ1kCqBMUioKuo8mo8544R
uyzdYr3mFSNn93UgCNG8SUtSYt0fR7BCNj1j/uEdjMjBa01+9gdHqqDTR8CFy/ANxLCaVYkJZkkP
OZXzvFJGPVgIXN5kpf9J6njInpmmTKEBy/60KcHSRKggj+/iLuYOzaU1RRQlZE3m29BMPs8yApdg
1n92Um+5eHQ7vbuBx2hDip2P8v/2C1v3DK/q/MXJGz///RO7+spyDwXz4xekCyJ5MGM12+2voiAj
Nx12fOl1X5J6POSEBu6oEW6kzJ7tTCDa1XzBD0LKO6+a33Q5xxEbU/ftxs6Ov0U5Y+wbBgGNyZXf
tBQg9gPwgFwG4GeKJDEQBa9CjmYWGkalbijwgfbC1ZpYClxBdZgTg6dztANbmqDcKreSStNC0U8z
vY37GEab7WSdTlT4iTrLYVgNk++tgcEn1fplsEV7b+CzGlC9fCoJFwgFVYYT5JlM5GNAnBDuJ/Do
6EOb4MrcxdF09Tw23kC+RzAA9n1Iz38Ebz3pTwgmpSmZQHJcOJ9OIn8ZVh7Tg2Ff+Q+wx7kTlp8q
RMoqMY8PGjvEzwW5yS6JqS2HNrADdn3DO5v+rQANWAJ51QTM2Hs/GywCov+nemHUgooKEjh3ipGu
uWN9cldcdPOBQVz9HzYl9b5/qVpbpziI6KKzfbixyWD/rb+vZCC3+NYy54p3Wz7fOehoL0Csls0k
ANlFowLyonRfqGXe6W9CNaqhnEiuj3nBR957Wn5fQr9UO/e3es+NIendsrAjMiRZDoo7tFme2yCE
rBvJYjMOcnvmxkJsqV6HNZ6Zha4NCkRcNPgLeGMu7w5VZ4OTPCi8frpuJFebPmydH+ztlIjfSUDs
scb4Xtb3yyzrDIgwYgqY9NBvcKFWsKmTgdKrXnOxHmbViybg66hCwN6mbySR4D3BVqLs3UnK+aLB
xHCrk9d86YBnfghIudL7jzd4CydHa+6wkeIQ5e3wSgsaQs7bJLFKSUBCsUCjzx8H74lBsgiQwpQF
8PAbfFSiJkBAlY4AGNMssFoPE9AWPVSq4WvV6YmIV+fLRUG5FcU0OheuYWWjtav2h33zTwAXgFUL
w1tWZm+eVXPpL/mHQIdfHp3cTm62nNWnwKAxqhvh49FbH3zQBMv9BKbCz2mNgxPNe7yxOAkVvnSX
PYvuLB7u+k0NmCZpMUrWUuV0l247tmnHq9KEg8mexkBxopTEBGPJNP91SClQNj58k69J+Mm9YFTx
C8xgqb9U3MWl74ZFhZyQ884Qj/jtUcZqjT9TszNXDzQNG/hFLkb60mN5Kg4AbbcNq8yDzFieKzpX
flgZ62Iu72rRuY1bJZZtdUN6ZN38TilRr9Qb7dGPwAhLHh9uESMwmhSwcD6dhWFMSZjHvnpnR6Zc
zpp1tgR6rXDuZju8i7Md1Hn2D5AkL9RU0VaSzI2lBfeX9NhoznP6UUPUqfMJglJ94zOCQ/bnPuVv
NNUWKT/JeJFv37QIuxxjNHcPqglRuOLYpev6AaOzLYBh0M2H/Bc6M6REuoj+MNK7ikxtDfNwIGeq
DwMVU3Odxmmo4Aps5WxnSMD/toN065QSaviLB5trcrWiwnqQsw6cYDO4i+ig+8uuZK9lI+CZ+iMG
tf4uNjXXbiP4Fb7S1JQBRw48dhMScIBw2zVwe17KRKRBLU/PdZAvnqLhmcEkePvrrv4NcDC7cPd1
qvXCRCltGQjPme6QN+acmSo5CTp+yL/njYqmsalzVHw9lnJJK1qQZG/zx9zPLlFUJTV0yvFGQUgE
35ZPk5a08UlkofNJnDUY7jJ1cFgnDfb8fxbYFx8airbAg1XbCv9Yp6i+542yOK3Yizb288yzxCPy
W2F7kwimVu3wOSGF9c6o3OIn5Hm7hqnMLb5X9PhMqBwDI12IeZmHOUHDQuMcAQ2xMz6kyvmIN9Jf
K/Y/sQ5OhyUHxc5cjt70fyHwt4B6O/WSFqUSUJdBcJ6rQ1umSfd+pOLpfPKb71XuiRXIHY9FYU6n
QfYAMTb9QOF6GEPHU3PlDtA0uOoKJXz3Y/iI13IcGsAAQkgMfNSi5RYGtKFdnWhskhUaIsB8L1ZM
tKpENFTPx3dyHADZzwZemaSV8rLdbzS2LUKFcl9mmtmpwmJqAGCJdtHODO4UzWA7ZLv8aWOm1poi
X3NNDmZiQhOXJ8zAKpAjXEgKh6jcm00bOTIZo5CtKmuE73+m1WkX7zkHeEXME6yKXdReb+Ed3ucd
SzHYtft2zifpQiilVCBevJYG+gonpJ5GewAxSjQUsKO3SYluXL9PifcIluwScOqHnkezfLxtaHij
xh4Enz89hxir6zuDFA+o3cck6Niwv1p0iMtXrIGcwkedBsY/bV/0G0KYmvUKZUbmuAhTejvMIud8
cIsY5+DTackPR+X0akloaLOjGH7KyK5BRJeS2pqFqwk4mLx0X8OSHZTc12O4jofkdQh3dGtm4NzW
ujdG3690HANBowHUgVIptwUdlk+sxONcN/V07Bx/uDLI0z8moEP5U7dtk+KHrd8HbJTT6eLwD0aT
0cypzVq0Q2/1j2esmvGzYdivpl9h6gdyWj53+GsLyCKWevw/PGDHDUu0bVmKJR8S2Eitp/v//btK
KAwAG7Rq0NDmBM9XS+CfeNDjcaRM/bLmY/LFDibKQ/5hmmf5yFNNU7Sz8QGeM80sTIL0K0hIxhn4
It5QmTGFAYU6JkRCDLo1oaS6YU0brCoILNt0m2h6Q3ugQbTuArU0wgtyp2cBfmp0tWDU+YeUMszD
csAQWhtNmb/QaqcGzro+pU+WVUJGs5axIwyqGGzD264kqNXscRwdsQu9yaaF4dzA6PL6bGprfv8D
gX/2aLnzcWvOqLVtGkvY6tgCikIsuq/VDYHKCjTmLh5ijWi6R3BN58o5CsepXBYp7pdlZkLraKBY
eFCNJrpNYWBNESBS9cZtfxijtj9C2UIKu8GhxsUTROCF1wa11g1gmZgFIN9scFVmr5HCrQ16tCa0
/pnrQ0GjJR0yVle9aQEuZs45n/F0eq6HJ/AQ0zYit+VPMRnbcvfcl/OD6Mr23rJVXhqn8IjzD87Q
njAoeTUJe3GModkbHBQZQxDbsl4pmsI13T4ZpYVMzdn6QFLSAIlhqgsWsrXj9czQhjPimMAvDCgg
tXo7fVHRh7N04Xi7z0CTp6GRe8vcduNcpFfnqUPBMMzGvlcTnSPUSqehGktVnG5s99JyooVFf9hT
1mK4/cCSSGkdt/0QJgw+AQ7iFyJVrxqCQNCvwYlhZgSVIha8/rxjwytqtgo0BvSmJvoWJ8YaH9iv
mC66yKmaAVebHv1CJ1JE6NGWTIzew4UW6mopOdNSkqBDLP5uOgWAROdGa00WZNYc9Nu5Zbb/MYrX
G4Bs5cqtEIxXdpWM6U5nCVMk1L+mS8s4U/LkxsSZzS7O7jmHqR4QpvrZj1K/Qga1vofapLD6ojsV
JQ2QIJKQGTV+noaEnc46I40NmwTN3t6twubQp8RRKCSlX4vIQAOwWKmE7obABPhknIsmWz5wsdMQ
Jebyyd48pvulCBGZBByEztpkrulzS86Dl7mE8F2gB615Zxb8zC50EiyY8ztjru96G7R2pf/gtbrm
FBc8F/i83bm7GLeVkhg2ACKDSCn94BSBW835hmy33sWG/Ru+nt+o3e7//DaxREvio2NSDFWkvoM0
HxeW9fsomvEMZ1hZ4Kc77H1Kb+TedMMoljDz9zz1JZCDT62yXqcVxP71Cxqcx7OS3JP+mwab+0GA
nIeY6D5AVgwDuamiXmdgASCKJ9D5y6cMHLF0d9/M2xrLFtt/gfLK8TvNocHNxTW+GcaG0gJwQbDp
8EcsJBcDl5hy+7khxqxhOsd5AeYE8D4NsX09ib4wI4At5CT5+8gixiY3+fWXOcadE1vt5nkgZfRk
bLJ435fGoqbcKacyZj6+MNOOtbKnz5/bb57TrquO5mOUH1AatZKvI3TtRyhU/mpkpSwtJmwxPuH3
caXpL6n+MDXwTZsDvQxr2y7dwqPqMkMpgr+opqZ0gAMtgU5Sqvvsj3Tg9dNGqUGk3oc0rRlB+SH+
cfJMva/jgRApj9+Eun3BKXEXwOVz0gIybsMqOzJcy41zaRSff4c26WNUvN+mStD+oQjGlAk+KmMw
Xmx4f8St/zayiDvOs8jQxQJtR+i1mJmK/9x2IPREYR91womjbmoCVBkZDLK2SU7UiMPp71JO09zd
owUafmhN/p/qV7TC06LcRTXZDax+moPmDKRTUwbeIGU4UMoRbC3jSs4PyJoM3czB1Qh8MePjdpuX
AAo+Uk5S4W1cELFLRFTsezC+MO0iJbS9B1HBQ2AP6fVWbGCOdli8c7SWBrc1uAs3VoyBFIpsUKn6
v9C+c2r7VDkgsgM3iW0B/2anO1JMEuJ4/+fC09EZdKUNTVUFA2Bu8liNklqIhjbwWRVJIf5UVXvR
76DQpDJkIj+Mao6cuAWXRmKgCl0SpcHbuCGMfE146Jk5ky+zudgneqFZ80UgMilvF3w3sico8u10
mD353gOV5em/ckIIv6LedyMSkQUlocBPg6GXPugiARvqOJ+pz/l33b2SIaoWRVHS/FwcFXpj/JC9
lNfikbD3ECjbH5Nrgu91rf7pH8+1PzddT+98Cm0WlBnBAVeTMdTuqUHJ2V2PBqmzVt/kBcGTQAh/
WhiMhKryYmNHk+SIlk4/C3HVFu0FTRce4gghg9CVMfS8ynQ+AWFEofnKQcrPdE84dijiINVCXZlj
ldiBNv/LTZ5dvSiRa7jTJnKpyiFJyAxAEu6gu7F94W/KW4Lbv3/szDHE7nZ/X2jxTfzxfWGwNeEU
0743r5ssNR+1cMhzM15QElHVbviEJ9vWDGDOW56yrK7gm7AMPa3QqgAAu5uzQr9yVI5xYkltPfoK
tB/w272Jv6V0B0TfxpbyM7ljEkmDBPQPK7YD7asqdF+MI/x4PU/g7Q84BgRU6XltRIkye2cARx3e
o1xnKlF5D+KYhhheJzsriuYrYx27hqDCIkTn05+Vkn7+fVV7a5Sx0/RV8EJCADqokl2GXXdFS9uu
gHhADULusEF9TBZDLts0aZIpPfk6S+GCFrZm8a9sSAOxq2Sr2i91XROWq5JPj1ApUzei9Qtz2DjP
70iv7IrlWOrIbJlqx0zAV4/xpy0IT5NAy603l8HapesnBjHdgL11NsjZaGzHbZZGo3RkRcUH+bSH
mOv9tKDbJ4/9TxSQoSViFGltTbl5EOgqnibiMUGsa3jAaF/jRuUoxMa9zdLVmI/bKefnELL7SC7t
fBaUTfpsoUyWKFsTQSRS5mPT0EKAIZkUpTUdlSG4zZwCnGF2YmGk8WP7AFj8qDYradfOVY59PdDl
XSPEw0siCkmLJX03S0KCHk8UUGoipacI4TAmcihT/+5JNCIh5k1jGqFvf/dGJW0JE9MHSbstSofW
TJ4x+er+jQ+lqXsZW9/HVdFmvAEuv6KIXoKiycXxU1sRjneePP/pY98GEi36YKR02hdenHpZKJ+6
HDqMEjtop9O9oMfdnQVqrTPAaV88PT62CDNHHq6KKW3b6Yx8I3oI5tPcZ9XAZ7KcFafvchL5I+gX
T03FjW7GBUM5rqADAnY41R/2h2D0JTdHET/rIAqDIWTz4XDEwNZIcpsikDmYsaP2PV5UZ3e9IFKD
J8pjYbIEphOAjiBQywn+Dn3gBiZzN5OpZ/fmH3+Z9bSMaolopJNwRJx9CEid+NNKDPJ9hOilAjj0
+YTBzzuVgsUZrePSzB9TOo9Js6pafWcuA2dyrAmzpfnbk1Gy7mURqyqfP5J/8R4NFAhXrYmRIP3G
5qhzjf6q3ELRK1PSxZgDNgsr9q7eZ+hXc4AlG8+rmDi4lJARWL0ZKHodtUHE9CvKIao+HYxdGjuR
b9EYtiFUHqKFzj8bDmQnllObUvCbGRjyAcSDWvJzwG2Qsbu5JaGTqDJfqzjWhDClbve/dl8EMFUw
1q8ADDjxS0dvBruQ8x3YxaZO5kAL602y4XIxKx0n3Yod3SQCiPDHDRl43XIQHIwku29uwViL+ogD
Fcz82oFXRTIiWtx8aM8ub2xN3ji9K+IxIqwdAP+qv7YwH2O1MDOccmmQYvqwhZQ9hQwLAdCl+Sds
Zb5YuIcS15X8qewcp9pfpBQz5HkFxxOflseNg7RflVNbLYX1PxMPligtbQTPPJYT4rLWypFejwuv
hJWW0h/oLyHolDPR5j+LBHxHjk6Adw934dYpUh4i3gt/70M1cNyE1N/vNjiIVn8Mk/7VgFsIWYXM
2DEToBdv3MdDjsV06LyTipGewWb9s2y3yWWwYOgFbvyLyPssV94Y6u10ukteEPPvs4FVyg/mtEqn
pBs2fCX1aX2s23WSTpUTf0oB4Q67ycqJB5TIPFjBwkGNZ3gxO5qRMU1CFeDnooks6csJimBSuqet
MqzRRAUUn+y4xY+cpy9OgAk6qbmcbLCnmeSoqabKSqdFy78RDY6nyYv6byJHHlnrZkJ9ooFBQTKQ
a/4dCeyvVZkHUobogXvHQbDSkCFBhY3XEVLEH2Ru9fvxT/I300CCpRb16eS7y21pD6z8mbUvcWHv
jFUNxIhCpHoDMpQ9EssjINLiU1VuLe+wT6ZCcdA6fWX+LYEhK1K12QdZJTtZG/XaZHVCDEMtk/y2
5tWgP3/ejZkzQXFD8YuJwNhyyU9Mc5nj4zw+PBrikQGvBj2ybwXGXQ4JRWXjoMBnNiTGh0QL+tVY
VuMUKGZqQXmZ/nYHPA0nZFRKStcWMrWdlLoH+Y1FAU2Bn2J1ZSy8b8CggTSAn1shk0kKIn6qMeAw
1w4ExIVBAvHMleNNfU2BtLcNr4erkwAjyqMHShGygG6lLjG6BHkHLAttXz5MjTiGc1PO3JaDwTfB
3DIRGXTNqNL9f+iHt6ppdn3kpOXgdANOE7HViFjRjt/9u6C1xNeHcXoi3/qvhVxezaY24vjMDduW
d6aNG+qm9BCsUAbKGMo9189Etcwc2G6Ykb39OrPTbEjOdOEmrMIHBPagj+kTrUmIkGafb+x/l+Lr
yajtiNDbXoVuTuz0oG3unRRSLTV31oT0H0CTpXB4HrCKA9zx5UbNDaMTL2SLf2aPg9MaToZnxm4G
s8ekwrdDXiambOlsXHGMc0lA9YEz5KdIvpttLKFPYapugA2eqGTC9VoSiZKntyc2c+G4+RC6ZWXe
U/zyraqyHCSDCoRUoOHcErIqEzl5096DYxBHwOWdmbaGwRdYZAuJOQruqJmJE4qvqQwSU2HFfXle
JxC4XVEP2yKBbnc1nONPVIPN12CMf17pcvtiuej8B8MzX8kqtq67I1qUHTw8vUhwHSp2M7SD+FHm
ORQ7G01thTfaYN0UG5OrDnrD+kOmqIj/CMSndvWjFBu/TRlbaavy4pLLkmjRWt/PNklcwBBqXGov
QbMXZg8MgjicQejT65UjyOaelOFdtCWRKYon+D3dS9Jo29jF1RkdjpL+ETIoDoj+h1zuE7FaIZx3
g53QxEDnu2nJ9Az3ushwcLKN7PZD3oiXdPfU113driEWbMKqZhWe7JB3QVQ/+wNmcAMA4W61qqEn
4ilThYD5xF80E32TqEm9eohbO2i+ePGzcehyDp86OUxotTKIAWxkHsj+OyWfxIDt5hPCn/cvFGsh
k/5aomR7nrQxZhAN/WWNiZWy/2IZhwg=
`protect end_protected
