��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���=��;u�#��� hH����<�C�l�1��9��� ��;��*~�~� �B𨰹TPvd��w0����Bm�`�~:����&�������d�6�.�����&[�R&MK��MU �
V0mc*�9���v�kո�p���@?�+���O��p���U[��?,^!���0�^�E�CMY��&���7B)�P��f�ꅿ08��h�Zx�~�����O+���B�s��s��p [��#�{�2+d4u8�Hd���F9�C�����t�����pǰz�>; e����w�S�I=�x��eנ�3�x�ۗ�=���)��'�0ge��R���Ph*r��Պ�1�����F��ܯ�Xx�W1���d�u(����m�O�Xb�P�`9K���Z�j��-(2m4u���YP�.N���*^n���ޢ��b��K�TMai&s�f� Nf=��Nȗi6���թ��uG����䊕��f�� (a�X߇��/���Q��Cv{��u� ��F�gH0���F-�{�_Q
��S��oG7p��x2�;�`�/��vZp�sHu5��y�0k<'�Y���J4*��{u�C}5�I�vn���%~�9��8�8;����߻ �����E�&<��.P^���D�9�y�yy��죨�~�΍��'A&AKZ��e��0�u�SE�nM��w1]�bAG��f�7����Wf���I�q؎�h4��>�����PhTa�,���&W�0�����3�b|��i�|ă0�A��F�:������W�Z*��N��MR������0S�*gI� �[��1K��X��o�S{�F��v�K_�TW��Hr��!��@�~�&T��J^�~��wA�R�T�cIj���_�͔�J��5�>z�Æ[[���-�+�=8c�Npk}�c����Q���D{��T�5=ͭ�����}�#Ӓ�w�0�_@?`�n,�e��[�M#��J����ܩΧ��
|PGm�L��0��apJ�����0��b��cs�]_�󴇆���Z)Ȳˮ�A;��*ٴJ�B�7�������n�;Q6�8�4��#ǅ?��!������w�<���&�Tõ�C��I�̀S�D��c�e~�/6��� ���y?},�e�`�;�]�%tYڜ�!�|�����Ri���޴�v�t�b��ב��=��YQV�z�5@o/���2��3r���X<����/Z_��@���>}���3��ᡫ7��͡�|��q�RΙn\�I%�hw��)@�>�D�|τ�����&��`؅�L��~���f&ͅG(�k��i�ClS���H)�ѿk�{�$��-�����_���%�����=c���gy�v��>��g5ݦ���m*L˔q��hj�ٸ�^��vD7���:m\�v��L��u���蛷�1��}���;H�D��%I͹C��d�Z�Q)f����wX��0s��>�:%��ժ3ɾ���3�q󓦶6*�т��_�Tb����b�D�N���n}>1��r���RV��.�XW6�J�,.�����"?��� �7�ί��⪦������{����/_���ŕ��Pq;$fA�O��y�L�2v�gC ��A��u]���Y/M�ױ���m���+�m@,A¤�W�h�$ん�1@�I�Bk�[
�'����'n�W&�%��K��OIV�7(�TY1��}wm�p� rB�@v�,��bz/e�FF�;���+	�Jp��<��e"�=��8H��w�]�2�����.�1E��0ׁ�М���#�`�c7�'�=n�}�0�&��6w���7�WmKCn�ﻌ�_�@��1��6	�H��W�H���3���<�ا�(o�%�֠M6>���'�LLN�T��x�'�E�G�b0w��[	����k���J��2�Z��z�)�h��ω�]�lO�!� ͊)S4��w�i�V���<e�v�ҫVS��b�ٶM}�v���8��d��n������ځ.��!�W�>H�뗍Q��wd���$<?�]}*�������]#��)��FϺYE�����h��%@M1~}�s
��}nȞS��J��؋��a'mfL���h	�F��ep��6��+K����X��+��u���,e4��}��T�S��,��:�X��f��K���-���/ȘA�C� ǳ�@�꓇"c��+X� 4�8�5S}�2�js��x�����'�(�)p zDy07��0�G�1[��_�8;J��K9>l�蛫S��>�[�턣um���Z�)���{BlD������ s���ly\A�����l��#�;��Ȁ�G
�ݜ^�������8Qq�~��O�V[��ͼ6��`K�
!'�J�∨3�E��42�0,8��t�����Ϧ8sL�qiT��x&-�`$J]\
�gqO�9D� ��G��ma��ca����6�,�F>������<?+�:��J�08����+Y��� �Р�ѭ�<��(yk(-�.�r�13D+���ro�AyA��?3<2��W�_�mlM2yQq��%i1B$��]$N����7=����'���S��@�����*$w+?��5��U1��puuqmW�0�@`#f�pw�M��5yI��S)M&�Ġ��^�&�����-��m��<z�I�TD��ݦ6�N�٢��3o+� �)+׽�˃���i��װ!(w4J��NpￜV.Q���?=�?#8�;�#4}�8=�!�B({)7�Sa�)���<	��!�UF��uK5];��
����\ ����wN�h��\�0Zx!�BS!|-@�eL�ŋ
����t��x�&�l���!�]��>�_%��Y�!�ɧ����#ӳ�lZˌf5��h�QU+l�z��q�o��hs��'�y�=hصMV��̏g�X�=�W�i�nV��bI�/����9��`�nګ0a���C����"
M��^��8{=O��y�,A#��~$ڎ���"_x�ܫ(���ã��(�ꉪ6��� 1py��u���&ŷ�k��l^��͟QY���S�;3�G=�,ր7c{���U�=�l���,�ёS�e�E'������̻9�����|Ʈ�T��A�a���w�I!�����#���EDY�<gOztB=l!Oj���1lb��EJL|P��q� K�\	p���2�L`(�2���d��݀t��%�ʹbR%�C�*t v�!%�ZJ#���d�s���>����ZJ��Upܯ>� -�;D2t�>o�x��q�H���(��LH�"2eB��zY�xx�p���@Z}�`�ې�2d���%FV�-�ps"c���&�A¹]I��:���՝�D$q�k�S���Jzx�&�MZ����Eo�������:�Ȋ�f*�J�����'^X3��"�$�$��S6?v�k�x�P�1p"���`Q�R��ߌ�-Y�RP�+9�(�e'�{b��5sDAB����Km���e�R���3'�M&!��=i�.�|Q�������^ڷU/���#��L�G���c�9I�?�OK#0���Lb�4�Z��ΓT�yż&u�p좹�s	^o�<��s��y��==maM��g�W�^VN���dM
P��0��ƪ�k!�&SI[j���1�A�m~�������������tL-Dx��:D��Q�ۊho	yV�I�>�G�P�"<|ۂ�[2/�V!Ϟ��<���n�\��=3�Wr�˹���geDdҎ��L����(4��Y��KȢ5VǗ�h3��B숯�p����Bp���������]Yw�x=��ʿq�O,k��Zk0�ʡt ʵ�$�O�䒿�7"����t9��\�[�a�/p=^'ټd�2i�e�����'��:�r�r>L��Ѿ�Iʜ�8�TL����&jMy���/�ZaB�%��f�Y�=��ӵ����S0�	z�C��8�Y�����u�6+��������.���1ʚدP�b� �gW���l��BI|�ž�S���<��7�d�߄jl��9;�z�u��a5R�(��T��߁�1X:"o�ߋ^\f@�p$�]op+((�%�w<La�D��#�<��Zg�����<�'��ਮ����I��j���vp:���	۟�&�C�Cf���.ߪ�B�ܝ[�U�G�A{b���ۙԚ�M\����x	h�B�e�pBe &D���o\�;��O:�*�GEV���@��\c�	9��4B|KS+�FQ���W5�����T�/�6W��ݒ�ߚ� u���T4�erJ��Gd�|��!3{"��>��\ ��Ϙ�Lt�ϥ�����%�����'0m��m��d%B�A}���R.��Iۡ�9�����Eh���ج
8�B2\ќ*�/�0k��χx9�$�V����mQ����k�Y�"8�H�}XΗ.�$�O�_��<�妼�6 �.��5�>�5��k�&�w�83
��|���)�i�<ԗ%��J�1���B�C��d'6�=J�@��c*WJmg2-y4�ЕT��g2���f:����'����ٮÎ�_���`c[X�1~���ބ,bZ�K6��D�>�X ݒ�L],E~�Q�F��s�%ʤ�e�����LOn%�����x��#ᅗ�q9����h��.��� R-(�� � ����+���Ku�s�V2�B�f7R��n�%�Ȫ}���-�'ef��pi��q���*�����A�C"��5��0�{������XHp�ޝyfH�� ���퍝6�ݠ�%G���nBٿ�X��E�X@N	=��[�61�ٹ�dR��9���,>��qE�TL�= ,��A���5����F����Uk�u�"8R�� ��dM	
�
���αe_�V̞���[3����_�0�:�0�TU��v����۪�b�F;9������+O�7P-♪_�d.�o�V�����ua�����,����n^��9\���,S����,�������jFaZ*qx�c������Eʉ��O�*�S&6���W$St�ȶo�i��=���%ڎ�p �����P@��%��tP<1����xLU��`8�=eX+V�^Kt[$R��F�-�U�7�{>�x3p�G��n� �ٵ���$�N�-V�]����VI$����-:[ݏ�y�͕��b�A�WQ�:�����Mv}a�� ��z��Y����&�aes� u�f~SաI��L0������_�q�/f�����T���͢�1������WŒ~gj�,��V�j;�u��w���m��D����Zce���O=�L��W�H��_I�s�h�A>��ĳ�_� U�{���o�<?�y� /a�������fF�^XC��q�]o�d��7�8B��D�,��,���x2Y�/Z�T�a�d�gi�u�����Vg���W�	��´���Ldŉv(l�
�8	,��Z_�,&Z'8���HWz�lA���J��wHAJ�W�s��zf�Ws�����J�4�-��g��+�9J��h�G�{M�<Z�L%����6���x��-���nQ�Hs6�R ]��i�2+Z�2�����bhb�0�@ֹƒ(:%�~9�Iz�mǓ�O�5�F���R��C�E�}_���-�����{�/2
Y�����Q�d� �ba��k�A  �t�W���8[^��*)�=�F�eAv��D%�e�D&ޠ-$�� 0��4^���L�Q��U�۽���P�t7	n�-�3����D�t�8w-Ñ-��kp���ã���q�;��lQ�ã�Y�<�ol�b�o��1�.fZ��J�P�H�h�6�z�^���U�g�2��Q����H���^���La'_[����;���܏h��<`g޲c�j������8�\cN,��ϵ݇�(�)��亲(��\zI�f[#]���L(�*�[��D��`;�����f����=����;\�N6�����3����]�]i�����K�NqD�t .���U!c:'�O����@��_��ڣ��U,*�U�a�5 _fm��y��G��\�:G������TQ-$d��#�@����s�=v��HM8��Q�q�Op(}a��M'��M��]����ѥ!a2҇�!�ݼ��ٗ����3������T�����͈X�^K~=J!�ꏀ�pk�cN��z֯{�Dl�b�����he=� �!ɏH����=����
{�Y��6�Wl��ݺ"��}i,��0��Nro,C��=�9���}YJ���lc�P���߆-1�V���D{�'��u��̠a>P�ÓPT���؞��^�B�'���^�F�c����Ǔd������5>*G�fnf���H9,[���*��F����o)u@B��ɷ�Ĩ��{ϰ�B�)̱YC	Bl��6_�>�67#w���HHo��\�;����I�TO��7����
����pU��>�k^l�5 ������E]̥��>�a�ƻY�	V�G�6���Ѷ�U��ވ�,Yc�0X���F�ui�"DZ�9a��\�09�gYO�9Á+��6�����ϭ�r��#���b��%���,w��*�5!�qq#��?N�]3r[F8�`'w5�x��*͠
��;��0T}�~�k׉Bb<�fq���4p�a�$5a�� ��*��&r�����|6�`���� �]�g���.x����O4����F��H�tܓr��|��u(�-y|Ä(�[p�.RaG\��l |���|�B�����6��U�y�I,��HvO���0��o��?D70g�A'_����S6������|�������ݧ�r�޳�(��:�S|�0��Ē�esN���Wn��tvЩ�7�*�������,r
��yy���C8���.}�7�*=;�'Ƀ�o���8��eO�|8̾B�M�
".{U��n��u�����B�����R#%w�m#G��U�����=2�/��%2�V�pШn���v�M7YTZF�b�un�٣�(>3F�u���¨4J��`��2�@�\@~wzr��(*��%�b�A��UW�T�p��]x�K���Ҿ`E4�C������F(yË]�1���߻���["*%��gg�u�쪌L�����Ӷ����  �Ӊ��a��'S�%
��t���b1>_v�_��}n�T0�u�Ƶk��,�8�Oc����(Njqn��hɄz8�b��R�D�K�A�.��B�b}U�q�����O��YM}Mcq17Ep�(d�U�+C��C��K��X`�^*���O��u�rjZ��Q�]�4K�O\��!�=�š_]���.��*���3e_��S?�
'Y5��6�i{�Y�:��<������"p�H��{�	Ҩv�z{��ĳ���:����;�M���3�E�}X�����I)�;�x|:�n^c�d����|��px}�I��Zrdo\:��3��B�J�;�����#��+��5��^U/ǉϚ�V�{���l� �1Q/�\��T�u�v�BJQK9g(�re&��]7��Жo��S\�j/"�Hf�VP?�; d����@D$g(+	�Q ��^�|W(��Z��+Kde𫉑�L��/[:^�)��N�H|q$\�M�!�Go��3���o�c=�VG3p&�C�*�xRP�`�9�l0Cy	\UiQ
Y�xi^Dr����}�G/���^���������?��}@�&�%����io}T�)D8��u�G�֬� ��s����I��=�֎" PK�7^}CD�9s�������S�#erՇ�����J"�0�h
�9�c�81ưzv�D5�~�RV3	�N0�`���A+��m��x`1��|4abg�*��F���wp�_Q��ylIF���5�r�sE�9�b��Ŏ���#!���Q�#��A�2��g��D���1/'$YH��_��Λ ]Wut�S�COv�qF��?*r��k��	�2��i$Q�n4�FUC�ʉ�
M^r3�t���0 ��RR2������.����B��w�	�ǖ�L��:���~�]89э�18w"2������/�ɱF�V����,n��V��7�؋��>���}l���B����$�$�
x;.jXC=w3�V֐#Wsqg�����m0a�N���턎(l�U#�;&f�c��g�oN8�y/(�}H�LQ�(ْ<q* ���gy�j�[���&Oql�~k�`�[���H�����%�ˆp�x~�Q1ZG&l~��A��^�z�kgb,��
<qm�8UލY�Ve-i�]1�8j�CQ.����\�l㆑LFs��s0�Rޘ,���DË{�S"]��R/t(t�9հ_�U�����%�$݂]�f���yy�[>�$����c������)�%d�<���a��1�����O����i�)	�f�UY�&�9�i���,�ϲ%�3n �FK?�Ɖ��d��w�X��7�N��P��"[�-P� �ª���K$�#�E��QޙL��h�z����r�Q��1�U�6�2z��q��Hl���A�}��QYɟeZ��2�)�zȆüΛ� �lL���A4r�]s�J&�%���x]�Bv�c�WC�;�+�G)+t���/7=�-�c �Z�F����]-P�E��[�(�m�1cxU��*�Oe_6��:Bl{[�RIit<ʛ/*o\s=��D��'�R������1��WUy�c��ɍ�E�qr�WY��<���I>��T	�˩!3�sW�R%-21Ô�"�,E��.߂ �ҼdN���qMK��'j��z�e	��_/�%)�U�����V�K���i�<��%ғN��ն�2���F;p��z����
7x��Y�
�{����T�Vf� Z�܁�&9yAR�.@Z,0�g-����wЫ \����<vf��*�|�(_uN;zLZfH�Y�9.*<��:�/%�@������x�p<��8_����������6�kI)K��c�L �F�AX��2���ˆ�$D�`��
��|��__����2U���84@QN�s���]��2���,�c5�l�bl��G�6��&�"B�w����\����2���������`{�����)QK%n����� Qnul���k���ⲛ�Ĕ>YT�� �8b�l��H�%��g#�Ȩq�M``���EL��[,�� �f;��M(��S�7�C��=9�TS%���Jg�0-�"�D�z�	�������דX���`���À���Dx�D�9��%S�;�{ܼε�y1�%�ew9�?��+�M�چ����J�~ܙvv��%x�J��	��٧��%��B2I�z�s+��S��ˈu�7���G&j{�]/d���Z�����q�M�+�z�9�4������.3V	Hъ,*WV}A0����z�K:�з��6Q�_��y�%�s�4D)�]J3l�6[��<�N�L[��W�A��_������s��RouX��q��d[9a*�*Z��:�kfvV��(���[9�j*����8+y",<k��N��ւ�L�[P-d�����HR��(���l'�C!w2�E��G�V�/m��,�%��ʤ·��?��� �(s���u�#		?M���-��huʠ],�%�"�3h���\�w�GBB||��	Z�v�~H����vdQ�Xlm�_�l�
�=���]&Ď=<x��A��P�`(���^��9��'	v�:c�TIM)��@,N�҈��翇A��q��o�}����KRrT0z��I���R���e�㱭�9` ��hn9��d�]C\�\�P��{�c��`�Np���s��ա����m��9�������ʪ��>��RL�h��&:p�#�Ɍf*��Ѕ�7��G�V~�F3��o�a9�P�;p����=���X��40 ���\����sn�;��A�0�L�i8'�U�!���������H��a^t4	2��1��W���\���jC=}��s����C����vnE�CˁÀ��j�PK��g+���h����I�
�U���F��jA�u�WR��cy{:�X��q|4�Y��1���|�PѮZw��[3�!t����(^.�<�t#<6i����x��+a_�9-��;�೭Hb�f"x=�6��%$����QR��%��~��?� ��������M;v�v���H~@��Ģ\|�cyn��n��)�ul���')��	?��.�B9c[�����2J�"�q�`���%<�T�#���F�_+	T]s4�GB�k7�^Sd�	_�7tw�LH�~���V�GZ� ^��_%=f@"��Pb�)�`�]5;��h	�����l;��+�p(�<��N�����p8b�ic8(��d��2��\�p���h��㻐�P���zkb; ���:f�ˁ���W��>[W����8�JӍW�8����W��c]�h���,�A��٧*�D�fss��X`r%t�́R���M
n���)�r-���Wu^bq���L��i�x����y�������ga�q��^G��q�����s��q}g�$6�P?�\���"����������Mi�\�M��k_��H�#�(ԫ�J��?,.Y	�էJ���8g�HM��q7�3����QZ��8��/|�R���vR���'2�>|EŞ�h�>��z��6"-���%�q��f��ݝ��4�0:�_�}�*�%�뷹��a�E)�[�Lk��� ��#���[.8�U��ՙ�B���ص��������>���_�`#�������ǼDPwE��ӟ�ʼ*�fn+���3wX��*��]'Qa
�l��ώ`�&�<��gQG�i-��#K��eߺ��j�ζ�DI&�	?�a���13Oj����m��2(rY?�^qȅT��qAWn���
J�ȵ��iA)�CW��u[�6E�1���(MzX� �X�ǂ5u��?��A����]��ATB$$�)��?����i�4� ��Y�t���w��db �Y��=�^Q����Ii�Bjznb�h�c��T�b�jڙ\����Ե�=�v�e��b[��Z�_Хz�#9
X�&�mV�U�Q��UU�ѝj0�ι�G�	]��f(� i{.��;����/����l��;m��+�6��ީ�\c�8��`���@�'\V�F�r�cי3�O�|��P��Ձ��]�]�' @E�RF�{�s�Rb}�T=�b�o��6P���Ĺ�_F��ɮ��������"�_H�+�����L��db<-0,��,��p�lmi��?8q���HQ��m-u�G���.�D���ѷ�kA��zo~�6��Z�'S,X��f�/|�8P�������xF���	d�qUǛ)�X6�������bǳ�� ���y�j��}i��o�0��B�����s/l��U�$U�-��Zg��+Z�CV;�M���R���/[���
 2���/�ߡ	e��)���uZ�����@�M=�������r��^0����]�2�<1�w]�B��búH�I.̬�MY/���ϬMc�D�8��Щd��pR�`�/�еd*�4=���hP��P��h:��f����]*{ʶZ����iZ��:O/� �h��ߑd8D�P��p��C%2v�)`����7�7�Q��w����)���߂�M��SXb�yq[Zi(��((&��Gٗ�ډ"Ӻ��1D��l��f9�b��%�ћ���x�
T.DL��jW�3W֕�]He.b��&.;��g��JOx�*%�#��C�_�,��:5
F��N�k^c̃�|
�5{�bKn5�(v�u�w��Ů�����Ў��Z$ݴ�=��Ս��^L��;���a�],����"m��J�4�?�3O�n2���Ŕ�3�Й�y/�����L���w�]�3�>�y�I�A�
����x�v��S�d�OOS�4�!������:�K�#����˲����[sIW����{'�H�$.�o�UwWݪnڨ�^��4�7:�y�x3��44ǫ�=<�P-Fl2�VY��a�gI�p6��_�ד�^����U��jn�\t�ю%;������[�No~+��l��� =�`1s��g��y�{�E���#/�n�]P�&�@OL����/���%�r��"�X^���ޔ���u[h�k�o�І �-�te�V��K�IC�\���%w�p�8�ɽUb�W$E��h�!ϫ�����+��?�u�x:0��RӠg#Z1�V��0<nc���O��f�2Z���6l<1�����<��"�,���_�mh)�Xk�_�5���g��tT��}�X)��.��r<�����f��$���>���1�^������VL�����D����d M�|��%42��c���(<�� �=<.�I��h��'������G9���3^����f!�l���*��"E9�p��J*/�Y�
=b�v�Ah� E�¾@������-^�R��ac�=―9�΢-7��V!�cnԍ��]�I������M"��6�n@_8r�&:ab��J6�����ǆ�(��t5%�[��.׼:a�����#rsWSM���K[l�^i�6O�F���?�V��1��<8���#i���񫞠�+��|P8�{Xâ���Dc�H�>������J� �Fa��j��^�}ĵש�߰@��%Iu��?A˧#)����rC�4����a.Ƃ�2�	�{�?O�.��YG��2㎵;�iY���A�uZ�&�MP�������J��ͫ�9��2��;k�C�+��sc�Ŵ��Σ#L��	�a�1މ���h]�=������M�P�w���x��τ�'���xW�=�3�N�vK��"�K^��%�~&��wI�!�^��wj���Q�ݱ�.�l� �}��������?��=J��H='Gv�]��2+��v��(~;���0��k��R�2���x��:�[$H���΀���+3��%���Y";i�d8�kK�)�'Z�ɍf�u�B �S�^	�������K��$a.���:>���}���3䰸��������/���ۇtb�<}@��A�h�:���e|I������fmX�Ԧ����66Y�Y�����BhF���{��Z�y�TP\	��yV��3ֶ(���M\�!��?&�� WxJk�k^ޓ%lA� b/
��l49�K��w����_E�G�*�y5E��'���y��J���V �_�`}yg��B�X��X�"M>!s.�
wȫ�y�������@�]�mlbj � D��a�7��8����'���A���3��[T�=+�J=H?I�n��~>BF��`Y�S%4�`�C�r��9`�rQ�����E;�)%�ܲEC�`oM��~���e��͇���s$78j����P��S�U�����yQ��6�FF4���@ChS�f1vӋ����S�w^p	���jI��ͺ]j��b����a��}p��̇Th;�O�/��}U�H_W=�"�[4R�S��'0�@ͳ2� nA�N��3SN�l����a��%VP)B��-��Kץ3�ʴ����<�ma�Ď*	Б�cEb�ޘ6F�Զq!�s�i�j�l�۵=��/�>��� �	UǠ�^'`V�V5/1��/#����6��y�,����pB6�y�BD���rYx��JK�e��8��>�qÂ�Kd��Z_04��CY@�K�\��p��f�+{�?�jĒ\	��X���Z�Z��d�Md9w��I�m���礇�us-vJ���|Ka)����\���u�/�o�����]��G��z5@�PZU��@s��1�z4��v����Й8�-�w�b.�(?m�7"�����
�ˑ��Oއ��ӑəd�
����VR�=�4t��td��e�-rlӍ���{��/ؠ��K:޴J�\�X`��ޖ���+[�6���K�,j�:d0���}Cy�	�6���c*M�a#����|��+���ŋ\�}M��%ȚV��A� `�kt������]���R�N��rh`T%��T�/�0�a�s�o�E7�jt�}�k�!-�����@T�ІN��L�88"߸\50aZ�H�X˶��cbUӠ��fM:���8���)	A�7�3���n9��"O�,
 Q��A�h���(3�;,��5pۯ����W����wؒ�@Tx��^<]��u�l��;WR�����O�J#C��up�,�W£9�b#X{��O�!�4�����WmHe~�)g0�c"곕��^`L]\�@�jNm8j 0�m*QB��
C4��l��?�M�]�V7�+!H������Ӱ�(A�o��gh�Q$w��E�+�z��m`�!�v��B�_�(|s���ˣ���	N  ��	"C,���C:��ӥ����c>4�cD��"]��W)�x�D)OgVCU��uJ��B�WD�^u�!f[���]G�~����U߃���Q���d��4xe�w���(?�v�j[��)��1R�YT��J%����H�@H� iDDKhv*��h�����֚���C����u�}z�2�vl�␋�!
!L	�T�9�W�rЌ~�i	Bh���~RkV���y����Ѝ�9e���(�3+?�k�A�K`?-O�����v���N�p�L�#��lE^PЗ���ߍ��Dh�4@X�^�٨~A�y#��o{����d��iB�;&'������o�_��Of��� ��:��cc���	���d��=����ɮX>�ܩP��E�h&�n�2�ۥPҭ˳8�v��ŅB�c��<SF)e�'3��Ss����n����܃��JK<�n=SY+�w~[T �^��ߕm@�	��B�o����͑5����?_8Ŝl��#u�w�_H_?�d/��|���1�fy@��6β�:�6;����n�:"�H��F \'�q��/]H�B�X�v_a'���!0�!�t���Ƽ	�>I�'<�K&�ء�o��?�5��OƇalA3?ǍBe� �X����$srү4JRWbA7�]��j
AW')?��0��'*��x�U��sԱ9�vE()����`\׎�e��`��Țb����Wx���t�M����:'A�̾b~j&%]@���>���Y���'.��:�Z�d
�	R��fލ��m�:���^��fb��� ���ʥ&�0�6��n��%d��s�d��a��I^�s�j8�b�u��&���/����=�P���ɦI �h�B=��JK�1�,���<$̊�	c���MR3���Q�L#�,$I�ò��z,�Np=h��2� �r�%x"�g�����n��͈�hL�)[xX��*��${���9��A�p^Vˠ�����(��Hh]�1V��<|{u
��<�u�G6�G����A�Lj�����;:�,���,N��pp�r2� }6
*���Z�-W>��;�Mo!�*6xo�}=Nݲ���6E'��67J4#ȟX����v��7��ia�_o��,C�*�C`ɿ�tG_o�Z�a��֭�8�N�e�Җb��)w��.��(P�V��}�#�B��d !v�%�TƴX �x�(X\��~=F�Y��i.��+0�u�;A�_b-��vݰE5'h�M~B�m�������L��Qt .O�$��/c{�vM	��z`3�	:&��8\4��f��C�&���諪��ڮ՘r�&���r1��'r�|հ,A���'M��D�	͟� t��Mq�vp+>i��и;�u�a��dZ9�(d��#���e��5s�Rq�Hnj��P���F���:	�#�I��ɶ,�W�^^�H��\`dڟ���V1b6D��L<u�0��^&+��v��tI�q�����t�3�BQ9�� ��=U��%�����4���)��C�(��l�N������"�Wg{��=�5���j�|�2��f	�|�Ҙ]�J�eV��s&%�S������Ipc1x���z��'��jo��V�7�K3�a�N5H�h��Y�=�[}��Ť&=�K�+���z^�_{[���z�>TcXA؄�p�3����ߍC�{C��4:b�3�I,����j�ۙ���.Ƭ�c�][��g��3��4�g*V2OD������.5���,��YZU3�֦��gE�{Ϗ��TAGB�j��ʩ՜%(��Vdz�T�DH����7�o{���5?$X�]~���3�v:i��\�>��>�i��u���& jB<�ir����G�<�S�IOk՟���֡j���%��n(o�x�N[� �D�!����x��� J���j�
���&d����u+l�c�d�ĺ�A_����)�ȋ��ڪ,*�̍?�nX���o?�:'F������3CS7;`Rl�	y݌��N�N ���wն�'�)>#lG��,�4rL����|/ʑ[���'�g��s�T�X8��+d�rS���K�.�v?T9U�+Es�(C�Giv�6&W����	1����������F�;���^��a�*u��y�b�W?C��T?�F1�}�%~`r]`�`�Me��ŗ����t��l�Z�����ET�?�s��(ַ�fݫh\yX�< �~++FYc�&��̕Cq,��x���Z���x�q>���,X���B���:��2O�kUk�����O| ��+�I�5|	tK�����������m�6�WG��n�/'Y��@hQ1�X�6�-�W*�Z&Z�[�{�����"��*��0�!��д�����I4b���(=�0�R���G9����y�z��&���%��D'�Ma�D��_)h��A0�7ʜ UE�����K�"*���ҙ��Ь�w&k�0UÙ��\TV�}$�cםq)S<� &���.AW���b4D"WXh��bx��ϩ�2Y�rq�5;�h@_��ѕ�NFr�CimV�!?Z�}���D4����Ǆ�S*�	��Al�|d����h��0�)�.�a/&������)�.K�E�K�]�	�♿S|���<[!	w��G!J���[~Rڗ*�+h���2��{d_�+XA�P��F�z�;IQ�>Z-�=�P�Hqr�t�U4��T�k�k����E�Z�[�g�𽝢C�i��z��!��m���u������η�4�h�<�{Ś�{��� ��1���䌬�G�k�;+�I��&`o4�ʲ��<�����T�`ʲ���n|<`Ŗd�cA�`<�R뢡X
P��\��W��<�{tݢJ��p��@�o�'c��H��I܅��l��լ�s��Y��H�w��"v)�G��5j��vB4("�u
S��t�Y
�G77LVX���_�(b�+��Z�0�H6T9r�2p����K���ڠ�뾷*��p�T���~�����ܑ1ֶ�o���L뼠%˯3��~8e�3N�*��8��v�)m=³�=�Z��qי}�2�1��5BE�%B�Y�����?��؀��%3CĨJ�~�y��ܭ�������N��𙓇p�<	����S����p�N>��l��w�̤�}�^�U*d��F�«�/\A�J��j,j�36�~^��[��K�"v�gνNV��؈Hx*ѽp�s��:@�{q6T�X�m�t>9�}>�iʧ����c6�lC�$y����s�����%����٢�{y��U�sD�1]�?;@���8D�ˎ�*�|�"����'(LFp?���%��Ѐ�F*����G���-�=@%��<����B�ځ���=����$��`�~[5�\.�E��_��j�T�4Ghaö�v'�������?%�2�0�2|�������X����𬝰~'�̳!�E�h��س�
� �R{Cc�V'��J��>����vIn��������K���<�)���w��>1�M��M-����%>��@��A*_x���F�
�%-�{fp�.��lݿ9̆���=�������j	�����wk�s�S�n5�Tt<�Yg�d.�V�?�Dd�����vPl�a�@Ø̧Z1�N�+sj�����O�w�"�0�����Xkk>�%!�HS"��}j�h��ĥ�i���^ׇ�6%,���^"iP��_��	��X£�WD����^���9�����|�ұ)v+�=�.#�Uv�(�M�{f�|�݇�h�M]��>S���;���Ơ�9.Z��zG2�F�c�6"�c�0�'+����̸g� 3���l���� �:�1�����Zl4.�ӪJ��x��K���V��aò���y�֪c���)� \�.�G��6�i����v���8s3�r�~Z���Q�J�O��ɟ���ڰ\'���G�,�I,wBY�������9� 4+��-"�;CM�R����!���r � 3E�;yo�>� �RS��0_	B�\�W�!�;�IC��g���y�����%���05��!�ݷ$s�^��<�r�d��r�Wb.�@�s��u��w��8��XgA��%JĮ�i皲*ڒ��"``GO��\�Н�abֱ��,("�ܩK�i��~�缺�#�T�0S <^�XMdeۤh�!Љ.Y�e'��BS�u����U�<7���e�;t�7wT�p�3dk�P��,�3��ꮚ^�v+�p|��]d���BL� :JY�Őh	4�#�Y�(�S}�^W*�}4��ԑ�����9@*'��n���6ྪ	��gH��'�,x{��L�ߨ�Q2�W�x�9�8���?4{��z��@�0%ి�^����T��:����=�R��CavN`kˎ�K�>�b��j�47AMohu&u~A9n�P��>:m�U1_��Q	�b�냁���#�!�Sk�������|7\mt�����Y���(^b�
�d	���w�V(��SZ�`��m=�D�>j�i���ǳG�f\x��[��_՚A��SIr���c[0G,�}�% ��c��fo��1�y}��Vw@�d�m,Ü��Q�@S�=�4�(-B	�S��<���kwcpS�unT�?�	��	ҏ#�mw���Y���e�:��>���'�{�S%��B�#b]Z'��C�G�mi�:��@_s.T�fK
տT��o�v�]�P�qH>#!�i�}3�lT�R9e����х��B��~��e�@���.fQ�paG�Hci�7�S[3��E��)��X�FCvew�7�j�F�/-� g���p�w�����Uj��*G#�Ad��١`�������ŊՐ��G�H���j���ۀ7��L�:l�նSC'� �"�N�����	ڋ�@,�M,����3hn}_k���'�ݴ�p`����N(��V`<���%��h��U[�����Ȅ�!���kU#��G>�FM٧5��6�]�*�]�X6������L��v:��d�8�W����8��-�LP+��D�{���=U����@V�T���y�|�P�q���~)��l�4AY�>��8��5!	q���fw�~��Z�ڮ���,ت�ѐ`m���$�U� yWT1{;�؎�C��W=l��/�h�����V@�{��/�5<C&d9̃dJ߀1�G|�A��&7RK���F����}�|��{�J�BRY`b�L�Z@�yl�f��ٿ�8��;�����OD�qw{�M� F���~SO�j���?s�D�ň�+�)I=u9����c�[���g����I�P�cp0c��bT�ENd���(f����ȶ?$H D�w����+����v-�!ȩO
���1t*^��fg�-p�F;�j�?�t�b���2�=�<[�nh�`��X���W)�o>�,}��-Q�%1]xęj�U?X��*ok~2:}����L �4;�:2+0nR��ĉ	��r��jcm��w�Y�R�t#.Qj39W�h�iZ�k���)��u�Re_Q�T���@y��=YF������8�٘��M~�^�<C2�V[�5lľi�4�����C�����d2RZFd?T���wڟ�o���^Mw_��VQ~���;rKv���Z�0�6y�����3/���_��r04��ԅ���h��z�����5I ��żo�9P������r0�>jYU��:���Hæ'6���ۧ&�C�1�D��M�ŋ�߫w���v�}s�1ns?ؑ���i�ͧ�!�-���<
�zqy�s2-��s�A � {�U��Zi�2�VV�r֏|?���Ĺ�&y��$�2�?	IP?�Oz߻���3�X��x;h'� �Z=��&�ݺ���F>��a[TO�/pu��X��+R�)�e^N�L�P��b���x��ۅc��2�e�������@����m���&g5��ȇ�����^���t�mj�UT���?7�:��d(	Y���i<����+}=i>Ϲ=�q��q�q��n���1$s�J����b��)�x�Q/�ʓ��?�ѽ���E}�0���aQ7Knt�*�
V�U�Sr��y'��TT���o�!S˵<�'�Y7��	��"E�'z��m�ѮQ����G�˷�,���4n�J\��Go�]��V@�:sZl���Z��5��Ć��R��P���>�g�$�ԉ��FM�Bj�B��T�0� Vu᫼r�� ���k		X����S����v�̫�gе�'2ɉTY]��ĝalx+�7��Z�cq�LP� �?����P�Q��5C�(��:^xoI�����A�k�:W�� `�X!���~���ќ2�i�g��큙���m�
����'���C�T���}�����\�u*�FۄMܗ�� ���(��u#�͛�bӱ���/���Q�pho.���\��+B���)���e�!(I��5'�����>L�1�L|�sq���~�a[���Eޙ�#6�TQ��Aq�AB�"7%��QM�7�5�����V!N�
f��r%]�D��Ƕ�guN+ ��ՊÒ.�|W�	 �w�w^ b�tHT� 4�� �S~� y�!��VB�:ɾ�y�#��{���|-wF���u�O���	������:�V-O	��kma�W��롿����ۢ�����u!!��rz��q�#e%l�\b�p��D�r�d��|z�(<��4s�]mZ���M���V�4듨�+6rLh�5�Y,ݲ^<A�p�c]zz/�h3X��N�^\g��o=�}�l�so�+��y�?m"69�6�v�/���\�8"�L�����2E�U>cZ�ܹ,qz�!�bN3���cb��8Y�}�i�ԁ�>�
�ev|Ɩ_M�r�J;�"@"��z�k;sb�H+�yD����R��[��@�ʷQ� +�ag=e��iNz<tP?�U�ɣ�M)wtxn=O��O&JR7j���P�:�F�'�ڑ�>�j���ӳgV�+�Bfcbz� '�-���k���i��(v�'�_��o!�z7���Fk��k�iN�\ړ?�#ۖ�[Ϸ�xU&Cn��=�uJ(`�=�&���2W��lr.P-����<+�D�XY��i�Z��t���3�M�ʴH��Y%]ᴡ��uX�*2�h�U?���OA�u�Z��VӁx�CyYJ��-�4��d��G%:C8^!s���e̤-��L�Wă��y����M�oy}McYi�6���
諨���yc-��f�6S;���>�m*��!�Nl�KF��>W�W��椽#�;�L*����*m��:=��p�I��4�+�)M��*�)�&�hN&�:�.�rn�apL����_���0]�����b��W��<,_�&� 嶱I�W��%��� K�zL�b�J��y䙕R8�Gs�mg��o+|���i����"ħ��]oAm:�Z�U��I�rEf������T�Vt��n	�'<&��5"rp������ʔ��EW�d���o}����@��0��uH�@u�+��^�M��*�.�uK���g]��'��~��԰���q|3wJ��rZ`$G}_L��bӼ~��	����m~���i�n��6�v��P8�2��������b��W��4�E��Pq@���G>P:LI��"[�vBF��GV�-
@�����:>'��Pp!y�ܺ+UG�jbo�O����� X�+�	��rw�Ƙ$T�٫_b��a<��ש���A��6\\� "eYb��íX�l��b|v\G	���$�vy�-_Ie>
H����J����Θ8*n�SF�:�����t�k���&gŠ}A����r��L(���TlʶrS:Y�#b��,�2sd�=ܧ���o���I�2`Ո8�l9�T�,��5��ѹʬhuίG)e�'�%ul�^���l%|MK��()�[>Pm.>��ڃq�y2eL�t��e��ZI��W��g<��9�e�Q� �"��r=�3���§K�)q(��p�.=�S2m7w�@->8����T�W�19�5�s�繓�]0uAL�h�dZ��]���gc8����LZ���`[@�wK#<�*��xE�L}0���E���� {�Ō^F?#���eFK���nz�؈�����r������];ac�J�c1�cq(��z� ��v��χ��%���%��'	;<b^��<S�&�5�����1�3��P��9���[֋|-d�"�>�=ƛ"�^V.'Ͷ��C�+P���l	KR~Fu�Я;HE�n�ܘ�:������uL>,�.(E��/P� �r�8�H����o$���R�F�O�/�e����So����#\I�D����
b�Z����z��y�5AA�	p�v���>%�PDۘQ�֖�!�,E�-��nO��*P�4���b�����y-qG��uAF��dk�3|a1x��m���c����,1�.���.�u��5Zߞ����˦�I�Y���x�>�L6��R��r_�>T�*�ML~�4��y�t=�	%�
!��~J;�:O��Ҋ$��H�϶��\�I�G�T�uz�b������sG�k��s� �!r�1��%2��pi�ϳw�j4�Lr�[�=g��5�}Ү��*�ن���.�0�bM/Z�86Eq~>�M����˛ء�)cߵ}���u���>�ֱf�� D�e�L"�}t�p *����u���ũG�3�fګ�w��NM~F���)�P���"����o�����fG(����P=���cH(�+]n�k����~�u���>�$�`��B˄�}�Ɯc(��ęy!bfo\�2��I8�m&�+ra4��ft��,��F��F͟���JEГ/%�ƅ�؃��N�f�|��Ɯ�U�Őʥrf�̟4/�,&	���<�,>����C��߅(��7$��^.�R=/P㾰�섡�	kӐ��29�?�c{We�4bƉ�αݕ�'��
W��1���Rd�
���'��/�h �r��a^vVKG�?*B�tQ�4K7�&�~Fٝ�2�@ű�6�\C�����6���.�~��y:����1��p�������ӭ+*���2]���,d&�pMl��'�G����1u��v�,��2%�0D.��� �/�����7�<W0��լ�s�/&�� b����<�rg���`�3�4�_��s��M��K��������~+����0��Í�i�O0���G|��m���@�6KuN�z����IyT�9�G�sG�MR=Ҕ���h�P 	A�`��M�K��nuI��L�O�yӝ[vG�[cHՉ:�E�K�e��N�0�6��|��Ȍ}���o�+� L�Xf�o	7�L��Y�i�+�~�j�A�H$t@��΋��F6g����_��5?l����4\��zOb�>fcN�`���*�[{o!�%�f-T���P��R�W�B�o"�_�R�x(!��?����jSX�F(ۖ��5�Q��#�e	F�ϑ/k�*ƈ��mkJL�w���]�����ݮ��o"�����C�H���Y;�(�������k�pqgW��*�GAJ[.���tRpF��5�'<_F'����
��$P=�P�C(w{�̇�
�#zf�Nj㳦��c�!Y�Vn|��l�P��]�#PN�Ũ��6���5t�k�)f�Y��+��Ǝ��������is�/� S8R�=o?4�N�� _�Ԛ%�Ǥ�����z��c]���%�q�DGC�Vi�XuXv�R�8O>e��f !}"gT��wN�k���ng�N쟕�a,���.�h��ך��Zf$� �6�;���Y4y��X��I�8�n��v�͉�P�8�߾i��_��H��Xv�G�K{���U$�C��(ݖq��E�}{|��8�H��3��8�.,���[
�A��Յ����3�EYNF�	�
$�ƽ��
���F����Է8[�ⶠ{�DIhmd�hL�,7�ޑ�~L�jW�#���]X�V�a�����3鑗��S��Ջ��H>�zY�e�҂r��������t���f`�7e� |�.����W�҃c�&���|�r⿁u��eޫ�t?��q t�6j���������ҋ7��I��WD&T���i6*��?0��AȔ������o�������7�[��0Q2%燘S�y�!���Y�a���^��,��b�����Ǵܨi�Xm���6��/sC�|���rI��,���kXWQ���^�X|BY������˿��[��@���y�K�����2WQHKX�*Rm�aEiN�L2�XO�@��m-����	Cκ?v�9�1�����en�|c鎌��%�fP��+��?�?��w�%��=R�Vy10��-jN?��պ2&���k\z��Sv��&-�ɴT�N���S��ƦR��E�q�&�RE][�1���z1�s��2fxt|��2�ߐ9��x�E�U6ނ�E{���@ǀK&�Zxp��2Vym��z0�2�S�F_߾w��������
_[����n0 �%͝Lp��Ǝq���Żsm���$Tz�	|��%⯃�C�N@�|�)m 5�C�[�<M�������]��}O���K2oZ]�[��oُL� ��~�,ۮm��1@ca�����2u��/Y�X�Y[��Ttz|S�H�A�t�k;}�P�;�o2�N�)����xS�>qC��xDA�0[�k�챉P�������v�������l�xț�;Pd�G�1��N�ԕ�Xܰ� H�2�����u�iR3�L�{�|� ���<V}�\�����!�
��F�8��T�BU���8�����
�?�9�IX,p��,�"{v���о��,�_�=W�x�Dbn����a {�$;���m,-�=R#�Cr5��)���]\s|z�w����Bp>E�R�	AF�:��+��KAo�gQ�=G�jyC�q@G����ϡ�P�� |��.�̟�K���dDZ���V%&�ژk;7��N�K�|���S���#"h�}�F7+���+'8l��x'_�nM����)�0ߎ>���e���L�6�lݒWO�L���~��"D�_O�E&R��
`4�>+es�Ƽ�קJYM�erXw�ݠ_h��G-�*"ڤ@ot\c=��᧮`g��_A��G�!�J�Zkϵ���5�u)�l:�Ը��6��AƟ\a�v_����I��M����i_Y,�-=pm�h)-����g��Ǜ��NO#���4�1
p͍���'7.�	S�P���䣗���c��h�S_W����rZ�淅���]z|0���9MJ�BWB5*�"3x+�n7���`1�a�=�g��h�J���Q��qV���axߊ��x��뀗��g@������2>�Ir:�%���
Ì�	}���܌���F��C�H̓��7e|Km �l�A�W�{Bٖ��R�\�Y��TЪީ�+h��Ì�YT�\�q�6�1
$�d)t��L��݂f������3~Q�_�%�%j����C�+ W3"�T덭!�����(�#R�+$��z�����˵��0���-R��3�g�v	�q������uR�J�ͮ�4D�@���q�)��y5��
������-�4Ζj	>�fJIo�I�����C��s�b�
з$
9a��|�;��EuG$Cl s�g���tO���tJ�ks��$i�]�a.���3��4����_��b��._�h�n�Q�-�����e9bK�9
�jm�m�Τ�Po�[�Dۍe���죤L���`M4%��{��^���	�E�ө'G�|�v,QP��5o���ԼĦS�}n���z��Uo_��tZ-�"�ݑ�D����Ti�\ҁ�37b�ф�*�'����Eq�ő/�	�K�,q�jq�o���j�)��3v E/s�`T�_�
GK�X#N�y���n�3}�Z։�k$���V��ؤ�"��yy���ݺ�^�Ѐ(����D=`Ɖ��E�E	i)z�D������@�2N�:����,�ޑB��BHSi/���Pv��:��ؔJ1C+�������m<��ߤ�|> ��S��PT�FOA��K���|,���P+�w��{��S��W $�]hs�'�c�l"Jk���ɡ���L�������K�g�=�4��,��&�ԭ����[Ne�0�o��Y�M����e6�~�}�RS�?|+�X�m@�HNCό��#��Ơ�\��̜�]h��q���!3��8�Jl������:/��c��H��Wʝr�&`^���OW�8��;K�W{] �Q-��<.�H(�ʴ���-/H��$17�)7(0�Iҡg�!$��3�p[�v��Z�*6;K���>%�+�҆��6M@&l%;��h��,����wT�l�̴0��;��v}��ز�F��)|u�)7rA����>gM}n��!�xtt}g��ɸ� d�B������1�I�
ѺF�%Vi��2a�Q�G�!P`?:��2�g!��k'�);(�bŮ�!���j-�왥��&*+#W�lMi'�ႭF����Lq�6�?��^,�4����4�~��OEpP@"�9�:�w�?7ط���orQ0�w�ft�K�`��Im�}()�`sHfr���Icv^��ڙP�Ф5�ׇWqQ���&H��r��b�"���8�M�'�#��c��d(<h�=�o~j2پU�6��	Y�T}���0�������� ��ګW�ؙE��^�Ȉ�{i���@��Uy�a 2 ��})��1u�2�w\�e1v=E0�t�а����FMz����1	~H
����A~��F&V���r$�?D�(�+��������1f$�E�頝����c�>��EQ��]y�[٪aP�J���:xݧ��f�7dXl�G�+���iE�����Y� �]���W�[̸��D/�*����FR���x���j��U��+�v� �֕6�ܔ��l���v�4Dһ�{P[Ë���$�XaD��5	�[�	�gÒb��	-Ma'�R�8|UY�}HXK0�EJ D~�����g��>�I^��&��A��.�d�Y�>�$;��g�\۹&~c9o�O�)���kW�[ �s�>�:�!�������o�Z͈Q#��w��)���z�����D����C�"�r��,v��	dG������0I�gz07�@�Z؏#]�3Wf���b(kÎ�Z��a=l���|��Q�ҰS�(x��µh���E�����!���f��t��t�Y���|�-'��
Uaȗd嘨�d���n,��@�-s:Xv����

����o�դ�c&��T��/�;J�.>d�f. dq�73���y�����D����Z0p�ٝ΁ez�X�T�1C06���9��/��D}Mwr���%�-C��0L���3U�y��~��1�����-�qk�1}�sLg�AR�FK�=X+����Os�a�m�ĕ�H��s )�������a�\Ts�����e,6Y٦,�T��j�	��//_zΥE�4x�_�S�IC��SJ
�	|�߼b��������'H���2��W��%�"m��֮1ϛ�)��P�j�&�``f�-3��:��@���C��b�*�Bq	�g ����	tw�ӥ?��
�'D�{ֶT�H�)�����|<n��l���C�k�'���'j�2�`PO�JO�ݜ/��CT����,���"c\A��<`�=j&��5�2Ko*�)�C���l�k�@�.up?��eA�$��Z��*����'���;Y�]3��c��{��T�$"�"~�K�����TX�Ƶ�]H��1�	�Y��H/=���� Z��6�8�7���~~����_Gq����;�2��즜6�(�����®���(����[�Z)�W]){��Oq�,^�4��E�=N+ϴ��&�ȶ�'�6#\|W�MM���g�H���N�6c� ��~m����Q�z�='�o�ylӥ�@�G�[@5x�"R��J�����݇(2�"ڌ�- �ku�����W!9{(!K�V�`�ޮ�u��T8��s���F�@��D��!M�&a~}l MT�/1��6{F2쳆<�d�Mܦ4١z͢.t�������Ͳ9�5=N�����yT�	N�[�9�0�ed�Ǡc�`~�wD�:(����X����1$�pt4�"���jm<��m����k���b^���͈��X'8��> �!2nWl-$]v�	l��?v?�E}��\��RO��l�G@���4�M*ӊ8�XQ���������啙���&P'��79�AJ�{�����y�J$5P�$^��H��_ﴸ]D�`���fisM���<��3����krd�2��u��0��H�[k��8T\�ljR�����>i��d/�\ӯ���tu��f�E��2?I{k�Ƹ�#�G�èaI�>�ݏ�["�����"��ޮ�8S&܎��!G�����3HM�?Е�I��sd"B!�ӖЛ8u�8 ^��`��c�ja#��ݩn���{�̖��S��3��<	�I��+�і�6|��W<���$M<T�CB�3��	�b��Y�ZŕN��(��zʳ�z�b<��w�݄3���1��`��̷[�M�|p��p�korY��w��i@�-�xL{�O���V�����ӽE0��5wYI�V�=�Rⵤw��5�閃aj�ʕ%�A�j$a�@&;Ƃ�����3���qèP��>k�� <�M޴�y��S'��<D�U����s��,�w/�}�|������Uű����Ky��i�j@8��;�M������N��8�FJ�d���c�P����:�&�JW�����6'ﯟ�!v��D���3���b䣆Jc������ac����
���M=J�P]��&�����p33:4
|��Hִ��Qx��O���
�k��J�U��R76���[cX��af�����q�y�W}�2�0o	K�4��4P�����G%FkJ��kMf��-���Ζ�F��4�E���	Z���e�.�~�2t�ًD��qxs?�?��4��[�c�u�����Q�D��Rt�ַ_�<7�$B��Em`��ME�s�y��g�4��d�x{�v�)jgQ�Y�
Ϡ�#�!�l�`x��Z`V4�-��YQd�:1���qꥠw�]����,`=��IL%�(tx�LH��>8�slڮ���mb�c�gL+V�*�ٹ�g���ō��fxC�dZ�׳�a%,)xtCT�L:e���TR��c(�rf�{q�X�I.��wٱ���>����%�y���tq�6+���gl�ѹcG�@���o�M#�]ɿC[y-�#fj���
��]@#���U7�����i��&�)���5�i ���6�hW��l���F��ö�aY����}%O߄:�%����,M��c�v�R�ItB&�WL�Hpf��ˌ�R�����W�$�&@'�؈ ���qZ�����������VF�M���)ք��j�}s��C�Cؐe"�H��<yx	P׆RS����2� ��x\�{,���%����������~t��=��n.����$�ڛ�r���*�{H��ӑ� OؑD���T�bo��9e!M�2�VA��Q�� R�v�\x�,����U�U�3?���@��K�,�F����7o�_�&ۿ��	-�Pzh���ƺ�Q��2Y��`_���;���'��p�tލ��n-6X���]�� ���^`X t�@WΤ�)�*5F�6�����5#Z���,o��7�~f�@���H5Sr� G�{�j�C�cw��|�8r@MoꢫK\u��I�G�V�N���KF�󲭀]@��)҅�%9�z ��L�%�
,wh�8*��;�����u��(��p����[�<�kKmL7.��R؛I��q�8N�S<1�	�K�vi���NѠ^�5[!-͖��|�D���U�ۺm��:w4�����:�z��"�. tJ�_���m����ߩ���*�ï�6V�?ȏ~.̮G�#(�i��V`]�z%�|����<'R�����iʗ3U�����v��>�6��9���xĕ�p��4S���U�Ch�`�4�o�B�'v�;�%��� ̺�F��|��H���ߎ�]#�o��]X\b���=މ�T����ʠ�3#���F�G'�'�HO�)��rA�l=�M���t�;!�����A)�<9�����{9A]~�I�z�pr�����Λӽ�|�aﶚv��1���<�X�Tլe��X�Ύ�q���C�B&�n�%Kŀ+�.'M���2��o(��.ƭ� ��M4��H�!��^k�ޫB�S�E��<O	�ͯ+�gk]��(��w�J�rh�&�g�:i��ܡzt/T�Lb�h!,�OC��z8� ��#�?�W5�m*�[\
��w8�"��0}��P%(��sRwx��iN4�Xv�P�
O�<?E6޿�'O�n�����6��Ytʺ?�o���k���T��\~�&�쟹��(�_E�N�NIX/��#59+��q�����t$��˺N_Ӟ�=�,�������J0�*����q �
#�b�]e�%w�&|��#�K���^%�E�����������!`%ǟ�Y'07�P���W��G�3g���❟;+�n.��}YT��ώ-��2������Ƌ	b�+������b��?ЍO�J�N�YCUC�fD@�bg��H��>��G�K��Z^>�V5�gx5'"Sy�~�i�����,[H�dA@�-v��:��Q�6x]zb��i�U>	�q��3'ς/f�,�����kFD�!��lS�0��j�V+y"{�Q� ���R�N��:��ၺs�
��Jr>�.����T����u���j��rR�0�����@Z�IpH���Q�Wǆ�6O������[�m��V;� D` ����?����d���+�h���e�=��4:��uG��~�~}���
I�|��n�D��+�?�H<���&�臛��Ψ��oW�bv���V���aJH�������?�(�E���&�Y�U5Ԟ4*��P�Jigx ��(�}�E�'�$�|�T0��/{mCH�r�Gǲ�r`�V��v��iPO����*��d�zg�)&�,�@��c�3ˁX~`I�A��&]1��7X���#�1��p|T3H��;���������\����z)]�.��L�Ǝ��x�7�Yvۙ��E�7x�/P���td{ӂ9!�6���<x�/:'��릺`��U*�R��^����#��r lC.�|<�K���g��v9�X.�V.�����f���Z��a,[��䊦�1S�Ί3���D^(���;Ҍ�qs������T�ymḛ�x\32:��~�P��ۇFB��H����v�\й�~����$����= �=�.�����J[�9����Q��=�[ˊz\�J9�i[��j��P��Z9|��#γ@@IހzX���?:,�~���1,H^ﵸ�B�ݼ:�JB�eڭ|'�(_��f�1OJL���B�����9��Mٿ2P��SXѭ���\�f2��'�]��U"���W\�V�e�ݭ]X�%�>�)�﷊��5�k|%�2��i����VɬS+����V3p�	���`m�1d�y�I����O%Q�/@�\C@�5����F ��n\��=g������[���*g����Ł���lܢS�3 q!�γK[�|A�����H�GW<�����g�����H��JW��
�7p:�(�K�ǩ�,D���6��y�D�G�T���bj�`�C�ޥ���e��^�µ��G�2&E�?y��	�i�EC<E�#���x��s񬢪�ot�����R��������[��y�r�AF�<��[�/H_��Q�����4�7�]��Ԟ.�pͱ��t���j�݉�6��t�����/Q��zgg`�L�GܺcPDA5n�'�F�6《	z5)�Y[*݅׸4��܉���_�8�R�d�4�TJ�N2h����\gg(U$�Xo��N����+���� ��2���<�/�9���'�	�r��ҩCӔN�/�ɀ��ǳ���j����F��ű~4:$v�U���	Kҩ��>�m�Ǎ��)��Ȉ���ل��L��\۶y�^)h2_�ŵ�jJ�>�i5}Z��Bs��}�u6v���9�, ��>��5F� ���}���
�yC�,�c2d%��EKNYiw��m��Y;�� �{u�;�6�PJ����D-\����7�&_Ka�������f���a����o�a��<��RG�9O�1����l�I%��(a�ҁ��W�i����+)-�$d�	h`���9�:W|�<�2^v5�ɳ���p5��Y��$���F��4h��Ă��`�?�\�:�{s���u������O]+�z���B;���u��`��N�A��
�b�;T�+�:2Ѣۧ��`j*�l^$5�u��K�[�<�J�zH�{�Z�G���=(
3R��~�y���ѽ�P"4�v`�Z��(���K}��ԛ��J��8_���otEG*��tP,��׸��N�A���3v�Q�R���%�����,�b,�n:�'�e��|�!`y��U�%�f��;��T|��@�
�^��r�c;�ҳ�hee>��
��U_H8/�xN.�\�:6�j���� ��ڻ.��8r�wηcH|�!�L�v:��J�`����ٵ�`$`K.�C��^���:�g�ܠl��\&�2Uꦛ;�m 
7ߛ�!Ӷ[�ߩ��r��K1y���� NϢ=&7�i,�6ǚ��
���H����N4����6R!V���6ʶ�m������P��Q��g�j���'ɘ��̐?���jZ�o�|��q�}}az�a��)�PX�YB�����8ζ�z�Cq-��ʡ+�fTצ�=��O>Ȋ�)��сGXO��
G���P'��W&#���Gێ^���TMn���Y��x���a���������~�bl�4�{�"?_�,�d@��d#n�ȶݵ	�S��*PY?�߿~5����Feh*�X4.�|��CY͂�'	�m������2~FY9�6�1!�q����]��׹U��g~_/¨�]|}sw��\l�����UUI%�,�{�Nkf9'tX�t7�U}x�pUi��RJMY���d��G�A`��e=)^$'PG�w#�.�`�$A=��/4]ń1��%�	�t*쳍,@�*�1m��h� ��$Du�MZ�z�K@�9��HFpPR��ل-��ڴ\��]�(��Z��t�'E��m�R)1�Ү�]MK��> j��sڠO��فv����V���9$HyX��t�>>5�)�Z�y�OՍ���w{[�����@"�
V�O�������Y�+�E����y���C�|������!C[�}�Eψxl����e�8���o���[�x��S]֬�{�KRJ��q!���r�yE���%�7���\����Rl�C �=�Մ���< ��i9+�����>lG�4?7ڍ�s�٤�ƞ����RJxq�(��]9���nh(ȃ�Wk(��&���$X��J��/�&�b�ƍ�{�i7`��>h��'+Ʀ �[	~8�=ŗo��S�Ⱥ�t��^����;^t��K=W�W�cMӾX��R��F=�:7y�ਲ਼�~��G�������+�zɓY;z�$�HR���T����*�,���"�!�n4�2�0Zƥ���;����@�����Pɯ)��W�l����ψ�"E���H"���*�Q-��V�����p�oR���r�EbK�A����Qgg�@��(�ϡ�tP�÷Nk/I�����J�SӘe�~g���q�F�6�3l���c��Й|�?Զ]��D9�[]n^����p#�oPl}��ET`�N� ���@$&Mq|�P)7��"�d�5�����8�0^.����؃��xo�3�C���p��xГ�	��r�!h�{�Y�FqR\�Ux��(�]k�NK8���(t�ܫ�������T��Q�e��������$t.6dm�F��9�?�q0��|��Q�Ra�0��:���ֲ'�ʈ���>�Ҋ5��_�DoP�_�q�J!_B��7"@@b+�Q��5Y�7w���&�� *�<K�:Z�=䇃�$p�\�J����l* ����~��4#�".���¦Y�:xB�a)i0����H�.�Z�񷊘��y� ����R�OK�%f��$Q�����h��O+�/ya��F_7J�,�̻1��P�����8:lh��F<�����h@hN|5~rEp͠F�~���ƨ��]�}S�j���_�L��DQ�p�}`Eq��b��܋iQ��P*�5[ ����s%B@�Ӣog���=��e��I
�aZ�"��a`$C�R|��={iW�.>����"�����'�ޝ�W{�f��>����U�{��}�҄q�k�D�$\�0�斲X;�6���}*e�����k4�/��9�5A�������G|��l�U�� �p�F�+(�]ȁ�����~��|�m`�lY�s�?��m�P�a��TF��m-u~޳���]J����$���bm���Ly�ViN����DZ��w��w4����������&�!��1׸Ja	����iY�m�v����Gy����{x]��$ǉVZl�B�
r\*"y�7���#^ҿH$d&h|�i��.R�i$��5�z�D�Ķ2ڹGv ~��I�9��7��g����(k�E/#�Q���͞��UQ��N�J�?��T�Q��H�'�ELZ�M$�If��lD��K�5y)�kH�y��4,�w�ݰ7�������yuo��-Gl`��a��yy�G���G�_ ��|G~�k��s&�'L�Y[� ��9�8MۃxP�Ar�D�+�I���xt�$\#&��-j}���`�!R��y��z����`L��t�1����KGjO�s���}���k������w��T����ڽ+fr�2��4NO/���GSP���uÝ|_0���SN�!(�a9o��m,�����y�c{�I=]�Cuub${����T�VN׌����Ȉ=j�l��Y��_�4c(}RG0d��3�t�|��]�"�.G�����1��î���_�.ǅv]l1))A���7�Luh����v�ƣ�<[k�,��5���*���]�w�F[�M���3�� Jt��&�����7��[��������H�Gq�4j�%ə*��Jhkj�\У��D<�����h![.e֮9�C$�x�[������o���%:����.6�41���"i�=�y�.����-��0x�i�hu���X��
18/�MZ�����P�E&�`_��f�]��|jj�q�y	�F���]1�*x:C��զǦχ X����}�Mk��E�O���T%<�uN��-��Қ�:>�E�l�M$���Ne��2�%Kԍ-�q�mi�b��Q��GKwNEb�6Xa.ڼu�u`f�-i��GA�=V3c��?9��ǩ�oy��K!FFC�[ܝ[���_�n�Z:Q#G�T����������.�~i_ �8�⃙GƋ��x������Of��E�K�&�տ!6ӝ��YYloTn>�6���R�������5�1��>��; -V��0�(���q�PjJ����\ľ�:���Z--�c�4��! _\y�|�C�!S����az�I�r/j��v��ĨMh"�/���˳�F��0��a-���߶��xv���p,�$�r\+L�ٺ�
\��px*���n ��٨ս0u�1����d�l���Hn<W>�K��>���.=�h;���\����!�c��g�	���X�w�V��A�Ccc1��1'��J($��5su.n��c9�/Ζ\�I��;����t�����6�-|��b�`N�Jg��&��+94��zY�tQ
6��]d�NH�m�eH�ѹ>��$V��!�e�4
����M��
8r��C�D��Q���'��g�b�h�mD��Y�Л ۲ݱn����8@2Q�_򡷽���wԮh0┩�H8%����n$��F��*)f������б���J�Q�ۑg��hx��q�Aj&�E#s�v���6��G���uPB���Nzs[ߍ�9��y��uv��1��@Ɔ�QD�XH[W�^�o,�ߒn9λ�V�ǧ[����Z��Di[����a�������Y^�۟ᶆdy�Zgq���u㯎�:M���Gc8v�D�!c�4Q-ԗ�L�#;���Ozd�&��6�ȧ4)�s�Xl�pt�hnO Sp���+��#�ϊ��E���_�ϫ�߱r�'o)�T����]���q�bh��#ޚM�<Lo���Ԭe���ޖ����Mw� 24.�<�9�G;/�b����B���	x��{���C�|��f�s��/��gڄʰ]�Y�&���P�S� #`Zu;N�3?c)�a�F�x��Rn��z�Ô�;���v'�ص*y_E�I���>��qF~7�xa��$P]��%�6�<���((�*3�Gu�A�ƚZ�����c?�MV�Hc~�5����H�>?��X4+x�pwc�+�
��#ʹ�U�h9�.��������u%�mM����g��2~��s���yr}�R����*�p;4�oR��|�6��F� �������$��)28�;-2[�AHK-�7��$�!P �%I6�_��7�o��z3���LS���%�w6����A�4��|�{�x]�ۡ��'>cR	�tH�n�C���ϫR�iL���c�3�pY']Y�����x#��9NK�H�6>l���~�j��U�r�c���E�z���|�U��[��=!����W)�9$m��s�T4�`	�g�{�/����Z�'��m+�~�vl�����f:w �}�͚z��}�I]�Ť���o����7F�	�^��;W�i���fM�q^�e�`�8l �y�����/��X~��AS�y��V���@�ҹ�	���iF;(��]ͪ�(ʂ8�)w�P�n�K{���\�9�mB�H��$��HC%�ԁ����d��Ka�������y�����z,m�BuVSO��'�ԑ*���_+�f��4"M����q�i�L��F�^Y��s¥���R2,Gm��O�&� ��@��_��@Z�pZ!^V�����nW)�[��T���a�Q'�>�
��<�6����uE���]T��b�[��~�8��}D!�#0s��ң`�rl�H1�U���|�g�����]��H ��V�!�6Q����(��w�ke{
!sAkzr�:�J�,�[�î�R����5ٶ�G_A�u�߁�5I��m��m=����1p�*X��M�3�lp/��eRV��诜�`�C}��X�պc����@��x�7{T��Tg��n�@����{d��>+'V�|y�֊g_��(�q��`����V��U�m6�y����_j�Q��T��,#�5�y#�A�d����$�`D8gׇ)4)-�F�(��������,�E_ȠG�QT	�^"�Y׆���7^�A.W������ݏ&:��&�{~�k�#p����I�/;K����G&�rX� �����jd��z�豴R��d��[�d��z�-���Y�"~�rL���0f�9�|���r�*9���&�8�����Q�����V�Q3��u+3<��M66Ù_.L*�M��=�x��줬M0����͞�}��������k5?*�a7����}o�BY��km��B�����줊�@uWU�uW��\���p������_��jZ4N2�"r�y̟���"�R���Ŀ�EMoȲ6-���~E��I���4C:�|sn��h4*Jy�O	�>k�IӰ6h���y�gvz���0�!ɨ;��k�p�	y�-4[�":4U��=V.��=#'9K�*'*�:��:5,��5m`�Y�#gm�+���t�QR\���\�I�!5�]cx��nɴcʺ):�2ݘ4��楱���S/����}�Z�*�v�@_�C��S�[Z���h��&QL�<���Q�)��#�X���A��ß� 7�%(�r�%�)o�j�r4�j�>�΅|Q4���ɭ�7��G�Pf��v.�m:ş�Ԯ6Bm��%��C��ú��
��s�f��*؊�����<E���SkY�d�/��<tB$�$�s)
C��넜 ]��� �1���uqNGZ/�Uv>���������� ���MF�5/�):I�\�x�MKE|���Iw-ݗC���o� U��_ aT8��3�(��?I8���f������~����m��6��ʛ��ϴ?g��@�FE]z�,to�'}ͨ*���)���o�"��,Ц~��7�$y�:�j� E�q�����i	R��0�h����h��.��?�h.���F�\9V�l��y{EE^<�Jk���6�����˭�%�zkP�Ԋdm�J0Yh�U�U?w�kY��D�R�au�L�޽t�j^|�D�{P�{!��O �N������4x�J�A��X��č�s��.���؇��� ����0~w���VC$5�%�%��C���מU�Y��DX76��0��Ssy�P�~��Mʰ\l��"�)��27������(��8����cQ��J� �>Y�%u������|5����2�C�c7��� 1���%����	SΪ����Mi��w�)p������b'�Y["ǎ�������`��,��wOP2�H���S�y�ܰh�9#�˕ڦ�z��-�n�����0ɦ��y����+�R����sZ��	t�� ��h��1��h�a�.C/6�e'���A��;c�Z�W%̚L��W(k8�Y�l�������^�!\�m�lsD����?R�ݱ�V���J�O�f�����:��Уm�ٚ��.�/�h|���x�oNL�v7�9�[�;��d_��U��ٹ�!އDBv'��nsR��J�AcfV,���Kb)4Ȳ=�G�cN:�S|�1	F����r��%a"�,s���
	��:?&�БT�ȵ$J�=s�)0�ZS^B�zD1��	��8��ֽ6�U}��&z��$�	��g!W(���Im���={?M%���=| ����Q"W�7�|N��	�3y�l�1�GKRWH��L'$�$�#[O��ZjwȾ�z�t�%�����=ғ<���yƑP��npȰ*�S��ɱ������?.fK8j^��D�V^�2Y�)@(:�r|����[N�-��&���0������}֭_��j��|��iYN�����=6�z��)9L��q�Gs�%$�T ���ק��Dۺ�H�;$����e	�����[ڢ�(TNO��U*�,�?=��+�g���w���`�ⴓFH�>�4Yl��"$|�0�a�ڄdl�Dr��^���ݚ���Y&��$��e�"����R���G��+�9ò�?x�o�1׽RTBm�w�:�F��{d����Qcu)�Kn�������G_R�i��5��I�6�a*��$�s�t'�x�i:��ࢗ�k�����3��&Y�&����:��������᫕�'s�� <��ӧi��l�|�l��>2��M�)���dt�l+}�F�+���]\@�_��A
��{U��ӓЃ(��hrxƎ�m�������`@Y�1�H��5��B����d�n]��QU��}���2�%��J�X���ۤq[w��tu6������B�Y�[nRl��S1u�T��~���щM9e�g6,R�JZ���@ ��Q�,��x��*��	��#G��� �V���QԖ�W	V�'��W���'�����8��#f�L|z���Df�fH�qeKN��1����_��̻������'5�����ƭf��2��G:���2QS\��	+�	i�+��BZ��u�w*cd��|-&|s��5�'�,�(�)�X^l"jB�z�)�V���P���x����x'�.�O�m��{J�Z��}v���\��Gh�X�ۼ����$�$~G��O��Y��2�ډ�6��A��˂]�>�vƑ�\�ˤ��vj�a�xGQcB��w{���1+�J�o�:S��L�|˴(q�ZSI�P8�X��iB\��T"L�_������$��T�3�z�u4x^2*Ȩ���22���C�����y;�QkFs�IHm����F3�W�:vK�3؝D�f��O�6W�r�+�7¨`%$i�������
��������-4��	Xq+�Ŕ��A��g$(�����%9����A-�y5F�1������ELMT�(ZF�EܯNʖ��cRP`ڶ��n���G$�v����%~y$&�1�M�?О�5�9�~(��O���6�$u�x\��	���l�$��p����(�������S�t�G=����y���t~�2�pF��a㡫Q����|>�ǁ���ȍF�>2�Kwd�@m�b�H��20��;��T�L�=��x�j�v"} ��f�W_(K���Z��^>��3%�Wي�&Բ� n��d�7_��n�-cp�F=��k~(7)wP�tZ��l��T�\U7���"iƛ��錟���pW�
V��ClF��e*u����9��L�J�K�)L��l�>���}�i������u��4aK�m)݃����<�ZQ��A�54�暣���Jc�կ�,u-A�����T���6�n9�(��.}^�cB�I�6��>W7~J��|�m0d�S�e�K���G�	��~&��TB�	�_;�h0���H��U8�MMZ��Z�2-V���.�x֞������4�Wh`��<��=���f��l��n�zĽL��l|�)�����$�|Ӧ:�Q�w|S�~�V������X�%^�D�@�����k#�u�!_	��T�1�NT�k�e���q�L?CTi�bԊ��G�]I���qv
���-D�ܫ���/_%�\��H�o�̠	EU��QU��+/�Т������	�����#n�$y�y=��d���8��`
�k)�D�Y��J��
��Y�,��p�����?�uC v��6#M�c^0T�g�"FF�ɑ�:�����y�-`m,j�Y�>��Jכ������5���\5ے�>��
�1gqA
�#�SѰ���Q��/�NՀS�&�U����L���@H#:����mÙo�9��.z=��b(��a���ވ�}�:�*M$���WFX 't&Ns��h�1kqhg״L�d3�\S�j|���3�X��M!�Itz��Ť_evD�]��X4�* �l�=���k%��E�X�_`�b��/�P����9I6��f�#�ı�y��Q���y58j�W�##����Q��G�$�x҃���&���S���I��E�7sS߻�ȥ�)�& ���6@�ÏFys�({Z�<f�<�o��H�hN�VoiUUY���Ĭ��_,��[2O��5/p� l�?ji�R�/֩h��V���l�0P:�\�k6�-j�̸��1�L�a�Y*�z�Rn��/�@ �t6�\g֌�8^	��χ$Ͱ��o��H��o;K���55�`�h�1��k���%H#�i�R��F�ht�* �*�FW��{1��J�\"�4lUGu�Iu>v�l��}�u+��s<v���X������x�_j\#��㹁
.�i`1r�_#��mda>'V~�����P@��/�)�'�9 �Z`H�&A�1�Ln�sZ�in��1�R���t�Qw��#�Ie�n$U�]Z��4� g�M��*��<�m�,��X�D��3�<(�ہeJc#�x��ߵYd�Pl+����v��*O|���{�N��$�v�)Ҟ�Z�E2���C��1�o�[Yթ�ٞ��h���S�_�t���פN�)�U{��z�ϗ�DYZ���.T�C,��Z����ŧ���7@Ɗ,�ː١#B�Ɇ̀��*S�4�k�U��Y��dC�+7|D��i��OK���<[w�rw�:f�Q6* 숞BZ�޼���`;�pRO�P-�4��L��{������}���Yv0���#���^�|*�U����^z�P��M
��vAֿg�!�J
��&k6��oQ�ŋ�����