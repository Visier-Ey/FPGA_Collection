��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���d�v����0�i�=\��A��?��� (��1_B�f�	�Ѻ+|n��y��Q4�]�aY�����*2�y%����>��������K������ �
�D��z�z��C�y�B����
_�U��hkF<�~x�ܕ�c�	?G�I ���&r���r�,	7=���b�ĝ�#�*�aØ��ο�H�x/�-�R�o5���u�6%�~����kq��yW�9i�ф���rH� �����|"�9	U#�'�iͿ`,�,]7�����3n���1:�c�s�ju�B��Zx㭹��,V���^����kpӏ���(1T��"~k�i�B�̫��� �%+F��F-��;�S҅�/�d%�շ&�I�����U��4w�Lxv�y�����`_�_'K6*M���>܃�(��������Y�H����w��4@/A�M����K���b3�Y@�%��JU'�8�}�����c}Q��dL���4NC��V~j�\����fa��Cg�2L%��f�w��d�{=/��s�O6�!
!>^Q�������Bi5��ěk�e��i�6�]�-U�'�;-�{�b��*�;8�16n�VkЍe'@�c3�������V�S��u��/�[)��Αݎ�Yt�3�W�'jC��y� ��k)�Ӷ��g��7d%�_	�.��x�A�ȇ�h=g�Z��g�}���2���S��>�
y���E<�Ҙ��d>����=�aCT��[������ �c\�#�u�W̶~�I���IpC��:Y~����m�������	���Sd,n�-|'d,hO&�W��}m-��-\���ఞ�N,kC��f +�q��!��j����kAa�p7ޚ�=�<>���5K�~��F$��$��b�N��9
�:H��%��1PG���A4RgLu���ӅVnD1L��16X��e�ː^�~��{I�x#mY����DtE9Pә�ZgZ�`��q\��]7�D{n�G��¼m���ZbG����w8�ݔ@��m">D���v$B�F	�3�LI�n�Q
����c��h��ߋ����u�ϫ6��V��y�(�Q+�i�U�"�.�)�2ckbH����X� �(璱̟�=�����DV0����a�R(�#v3��!i�1�`8foR.��nЅ���2��O��Vh�b�����?
�jZ�-BR��%����6i�yA��<�Ky\�2�֩r�k���9�%���!u5vx���x��ҭ@#l5OKykHL^��E���P
/N����B�w�Yg!�YQT>z]�V�Q��r#dC>��gu&����P�ΐɌ�if,�qs���,��|�	u�8�A��Az=����(^*�ws�0�L�V��@��ULGR����5�^�����C�[�����`&�;e�F��C\�"��	Gp�*��z}�w��9�3?�S�V���m�t�:5�N6�����iW���'��)��?���P������%M�5?�D�D�N���P�s9c*��IQ�E�T=�ytgwٶ�Տ�d�dN���ъ�:{�`Y��7�weR���׹��l
Q�c�s���c�r�#���WE�'9����iE�!y28�7�A�:�6#)~��@xg��D/醠Y9�����ž��X˲V��p{3��T�< �e���·�oZ�J!�!��=�z�L�A��HLw�O��F:�O� �*�!���9�DS�Fֻ$�?R�bQ��L��/c�Л�~(:Є!�֝��rtK���޾��YKx���>LsI��m���q�|���������pk4$���l���C����-�\_m��Ȋ�XM���x��X�]�v�P��?=6��wn�70�	�H^7	[�������kr2?��=�O�\]C��QZ�f*�!_P�}$x�{+����ŭg[�boO��?}�7g��G"�G(2��k�Ѡ�Z�OS�ɫ"��O���{G���i[���6��@m�]�*�#�MД�|W�H����z�-��P�Z<t���$���;zI��6�!�J�=���i�W�uq�L5�Y[;��}2*�R������A>r��t��7D���i\�|Ci3��.n��� �h��q���r<|`'PI�C��5�w�{D�7[�<5p�]烏:�Ֆڟ�Ԏڑy����+b!�&�V:v/X#�A���Z�[�xCÚ��E8ْE����X*�6�˹y���Q�SjH���k��뢱�Lq�k�p)��F�\��Ơ�ELb ����tes���"�W�uߔ@�j",�U�?)�Q��7ML/i�I�Ѯ�պ﵂ن �ů�ൌx`�� 8ɲ|�ZLcR MR_uO���r��r��P����B�+��z [:M"��w��5���$�#n��ϗ�+�O+2cDQ[+\���U#oo8�eb�]�@�,�<`���V�6S�����U���a-�|wQ^�\F�:�`5k���ӽ"d:N(����]�j�9��#�-Q�:�v� $9Cʿ����1�aF;������[t��8��,�9W���0���}������Z� ��G�%�9�M���h�Z�-���MG�ODiDn���A��Xf���X�Y3/�O��D:���οe
1��t&�i5��������}�l�hy�4�k74����	.,U2��pi�)a��Eo�41�6\.���l�O�6%�h�������B��in�x�Rk�6�a}��M�Y���?&7��rQ����X)�@�F��:G��%��ߺ�E��6�Y8�w �N�Q����U���N��>?MbJ�CoV��C��Ѯz��)��>n}FM�1�+:c���a�jOy��EX�Iz�Q�eY���d�"�(s���<��t��TW���f�I�~��*H�.������&;�9�����4%X�a(*���oʟ�h]A�:��ꀘv}(���ZU�@à6���{l�kja�<O�IoF�(l8|���T��*���&�-��`PH�T���x��;K��[���`�n=�>�U?��'fޝ�O�L����q����"���	D�J�|C�ׄ%��H���b�/��^	p��\u�c��˨6���+.N���*���n=�<�B����f0����ڎ��!}��_��&J�5��g�x{�\C�s�]� ������q=�q�J���9&2)��*���`콗Y��()9�[�T�& �a6Iڒ0s_��5����gJ�ü#Z���s�8/��%S�L#��@k����r\ߗ�`����:)�M�\�,�f��dG�3��n��6�>
KM�ɧ�:�]dLbSÉ�3VA���Q��iltEN�p�c����!3�W]�D�+\bP�
:eF�Н�⠟�"��rrNZ��5�.�P�����W-��5��X�N0;���bawNNW:%8�����[>=�Xj�i:�PK40+T��u��P4
���=�k���M1.W�,���<�.�T��^�.}T�H�Hu�)���F`��7о�@���*`��3�q���s�-��9S�j��q���:cv��4U$>A���κA�&�}��������Yҋ�w���nesr����0m�H�-�mV���L$�2��n�0�E	����υ/FDeK�bm$(x]E*t̄��R�Ӟ��u;�f�l�]e�� ��+ܸ�m��8�����@�+�劔�M����(ȣ��
�ZW�����d~>�M�G�v�;!��\�5�֖5^��Q��aN�'*���|�t,�n-�d���I�S����Ί0;&��!&��aK�L̹$)�8_Y�2V_��_�I�=��,�����F��(.N�����j�4$�_�YGr�<��׸�m�s!��Z�{��Cjm+��\���_���b���=I���w��T	.��(��g�W���Ī��̈���T(�bcO��GP���t�Ŝ��Pp}�*���o��U���.n�!�11[�
}xG3�%�І�+�
��u�D
��x�,
N{�Xm>��bz241�=��x��ͯIXq��.���� �^ M@C��?*�~u�O �}����t+#�~���ʜn�ٷ�� ���^����Hh`Z-���_S<0�e�0?�C����#���S?���DC��d���G�eb�q��!�R;Tr��ZJ�$:���o�&�8��]��S��VY���~�E+CT0�ڗ�8P�VSNV��@�؉���4L9�e|<]�����m����a���X��v�(�V�Y���ll_o���ljl=)tM���|'B)�l�Qa�W�Uq���$H��qM����	�h���%=��4��Ԡ�[�i���&����X����ؕ$c/�����v��Ѳ̂��(��ϡ����r�a^��y^����U7br�l\��n�1g-�w'�M����%z���, L)��*s��z�C��ϋ�ckS��c����=ܦI�Qz]������i�" 
�/���^�c��z��`t6���Ÿr)>mN�@�c�8[)I�G��R�M�0��f����ݲ!�8��d�a� �!��ȍ�@ ��6�_�5���#�B��П�����cc��y5I�D�c�GX��F9J�#B-WY�0�i��E�� _��_���a9�D���Hġ���H�C非h^s�l@ѥ(���~CJ� G������F��`g�E�罁��b)?��m-�dE�U���j8qO�2���V�"�����⁮����p:X1�I���{�8��"�0DO��2`�}�#挤<W�PЪ:
R���ۻ!�w�9��e+�eV�G83�r;p˧�,f��D9�&V�������.ʢ�^P/D�G��Bаۨ!��܎��1��>J&uj��-���Y{%���e�<{��Ȟm-B��*�΄�vA�׋�?�[�+���"&Q�����<!a���J<Y�۲���\��Jp�UMWP�K���JgUd����&�)��f��h��D
�hD����ٰ��t�oR�����1��N#V�@�M��E:�K<�'mk�n~�!kLH����x��po}�{�7#RDnj�l�!��5��L��N�>ط�#� �����K�b�P"�����_F��JJ�>��B�����G�8%�i� 1�����~��>I�h 
ۮ@h��X�A˥;��IK�/�V&�bкZ�ץ��D6UV�T��o�1����a�8�zRց/���4��c
ІY�q�D_�IV|u��f��`���65I�O��)G��:�)�ٖsj��W�V��ǋ|X7e�ݾ��U��(.��8��u8os����@��nl�9f��]������)�Ϻ��4I�-��9�ڶ!��5 *Uj|a����耙+���D��أ�����F�WL]�]F]:
IɽI�#��r�4��m&V���3<��ZU�^s�������W&��I�����~��%	2�I	���_$�c��捡��Mp`�\����v��9T�΍x�^���ר1��r�U����p��K`��lRN�0��l���c���J��~�'�gHd��|�6�).�$�`:�٢�ý#�Ʒ����y?&o� N�t��ua`��`��zg9"����14�X�oܘ�ꚓG�9�C���u�,}.'h#HD;g}3��{K�jC����5�@�p>K�/��N�a�J����/xZr�.A��3B�Nw�\}�AH����%����n���ͼ��,jV]/��iv��)1y�T}&I-I�r�_�t�,װD?@��"s��xr �(d8`Kq$Xp�d�V��]��mp���l=G�}(�������*�VZNE��q����Z�.p���)�%7a�p8�?��t97.Z�0Ix���BT�M]����H󀩎���V2F����/d]�dY}���e-n6��U�}��=�vC��&���s�_�(a�x>/���	CL�/"'����/���̤��v�!82�j y׵S��ou�2��v��	��nrj�dݪ�n����o�|�DUJ����X���\�YK��Q�H~uV��������&ݞ��m��Ǥh6�Jƶ%~u �j`)Gq����r���[4i�"�v��^	ǃ�_�J��$V\am��Ă�Ӝ��3,��p��[c�������A�Ӿ�ݐ��B�Hf�"�c� 9m�|jx�$��qGE!��)%1�bqoQ�'�������ўm=Nuߋ���xP��%?TJ<?"�_sFl���t���/��6mZb�a��\��z��Ӕ�Z�2ޝڦ�G:PY˰�I�g���G��:��!�%�\��� wx�Tk>�I��:k�ʘ�p.+��r��N�k<(K5v�22[>��(�$I�uc2�Q.�2���<PU ӥ�>��!���;�k��(���ژ�+�QI��N�F-���2��r�x5��'ί�טx"��\sz*�Џ b�y��ub�#���0��h[�7����1�9����"�Z=�e@�4�"� @j������tɽ't�h��m�V]���|�Jׇ��i[qY�%`�Zph�'j?Ko"x:Ķ�_t��)f�|�p�%�ZS�"ݩR�R���1��r3Q�"G���NR#�JB��B��^0gaPX�v�L穠��U������v�X�m���ؿZ�v��UC�uE�/���f��HM	�ZK���gU�Zb�����ǂ[�kZT.�t��Qn��Zn�;�J�lc���M?:���)�["����D�������P-'���>�j�6�Z�ީ:�3JW7h5!2��������=����&�N_R�s�[#��'~tk�>}Ɔ�wN�Ǔ!���J�r�L�<
7��`�F�%ծ�9�Љbܡ��Z��3���gS^l�I���Ag�Z#iĠj�V��\���&�B�L���b#�� ��B�C1.�k��!���0sc�:�)B.J�`8��҄'�3����	d%þ@�&-T\�-�0�⏘��-T�\Y��j� �͍��I>Y�̙��"U�V�R��� oþ!r��Kcv�&K���+@���90D�0"��|�Y�Ao����cb�_�dJ7��r�]����^Ol�:���8��:?��[C�Í��I���"��oJʢ���G��Mm0�d�?���`����
9���
R8g��d"���`��ꔲ	���p۩$[#���G%�GT�e��L�Q��ۨO���Xe��^�=�F!E�k5'�'���[�J�,�Y�a�˝�~��^�O�L�'u�r����t����gv��%}<Wg�ܳ�gRs��xF8s��$=����j�T�[k���8��'���gl��9�f�<�]ı�Iy�b��i�pc:*��u�Y�5��Wv��^t.}���(>���B.u6dn`�g�(�o��p�չJW��.�%�����\�R�n�ɫ�ԛ$ӄ�H�]���3"�o֊!�/�B���x�Y'E��8�׿9+wAt@j�@�T�1�}Z*7'�`�
�]?��#0L��U�&�諫��~�r��f5����"#\"��D�¯�����QG%��e%q�K�M�r5���vo3@��	,G|��u�����Umhe���z7�9g%ϋ�8�etx�+�!�Hh��5��e�$�5���2���C���YK�G��^���4�����i����T�}�m�믒����As��='ƫުy>����x!\��i��;X,���J�Ɂ��	��I?�1b9��T'P�߆݉{b?�E-�	_���ˋ�L��
)���9$r�u`�����f۳>[��@W�/�S]��`=�&�E����\��B�S-Ry�7І^�:k�g���AqϹ�j��PzBp��C���`�h�9BAvNٛϷM�F&V׌d9crFc��Zqww�p�6�� �����r�THL~����AK��#���A^�D����_��B:)�=m}ɢ�5�P�m���']��X���m+�5r��Hغ�H Eue�Q��n[)Y�V����7��BӦY^�9��f/��h��<����z���E�A�v��金�� �pCP)��sQ$�2��2�[�+��#���v9m�F��>�3>�z�B���]�;O�����7�}4������ܗ�I�.��`'�9��_)vC�}��g����fC+� ����|��2���cEc�͡������=׍5�ؑ�C����kGPn�������E��0�k��)nF� �,��N �wm��
�R���!$�gtն���q�a֫��ٴ)���[r�+���)��Kn
�fv�,��^ֽ��$P��-Z�./kn�$���y5�ȡ}�ĥ���xQN�F�E#��0x�@1�9�������u��T�:W��L���K�t@���ƄVJ4��Orc���S�8
Y�_*�7��*9�3��c�-�d���ȫ�S6p�h�[�?���<V�g{��r�Õp٩�l5�g�L	 �]���P�.���U[dj�q<�7얳�ROv�Lb?��J�����2��U'fv{��PO��K[#�QL�GQ�f)��Hb�P�e����"�����g�I̝��ȸu�6���/���E!@��0�����4Rw�I�FA�fc�D%5 7@�)�$Ui�}{p,�i��P��oP?<�Λ,�1��@��"��(k���R)JI������Mqt��$�����9H��Xߊ]��7�@ߞ�A֣�Xd���܂Z����\v���?�ٰ:�x���I�a�;��\n\!L�y:U�P�� �Yawh|8MP # 2^C	�D�ڒS�"�&��3Z��S�Cu������p�I�����읦�g��Z�<�,үk�+�	�C��Ɨ�8�zM�պ�7I<Bʞ�V� ?����hܪI���=��d5�y�\���[�Cܭ��1�����넄�v;s���/��~�DPN��$C�(Q8U�ڌl�P��y)��}��qƵ����Ӹ9�崢���N� ե9!�NQ�iƤ��G�:m��!�9��0zh1<��T���`)��*�F�i�N�����J�A���^��8�	V!h|Ҋk����=�#�f-ÕZ/D�0W��������LH��=y�CLC3t�PE:��;_����� i?�o��L��6���vʓ��%���ٌxp%3�ܦ�k��=xml)���*�9�V!p�˼e�̾A=	���l~2�Qw=�ql�*����053�q��_�T ���T��<��C)���U�H�����-�a�<�e�U����j��j���<�&⩭U,�X>��4���Ӌd+vm&�S5 �)�^���.1̌7��]�!y�p�k�hDb�-���z�k�+�NΆ/B]�\�h0v�d�þz8
5DI[�h� S8���d�8,�,�Qn�Dh�ҷ�:�%F��M_������Fu�77?���#?�-�,V�C�G�U?C�V]	�[�p��&�N
y��h'�2��J��g�Q(����>�Sp:v@i@~��PTU���2�L�ہ�d��<��\���B����cKX t������&D��O	ίiDj`_;d����籛3��&�&r����H��� ��}�z�~��f�}��Q��������5��,{�F�i����h�x���o���V���3��ߊe'����7&�2�].�ww��9���Ц~]�0�_II�:%��W�?�30e(��B�d࢟LNd���Qƥ��3Q�! \m�W:��s�#z�+�<|_f��j�HY��E1�8_�d|=�0j��]?5�s��Sa�֒Co�DBRe�rED�w������O�S�I�Ń$�����b��?k��A=��"�A�A_��9��ǯ�cpD}��m�&ڪ=\�>ׄ����|���YtY�	��3�Dˊ�/W�x�m�+-=�(
t����8z1���/�k1i��AGo;1ps�1�	"������)���Q�]3���[���"B�H.X��}s\bl�`���.C5�?��m���yAi��y2�£�}��[��A�*<#��x���%������2J�b7�x?�,�q۪C�I�B�7��������p��4�h}|I�"���7�X�H�R@��se�Q�%$!a�|&�_ϭ�ph8qj�+ 
aҚQ���]$7o-%����i\���'� d4�»쬁t����ҍhT�*��ß�����:I���<�Z� ��o	9���V������Jxi�6��\�E��G��Yk�V(�⑼aw�#�c��`,D�������a�^9����z�wY�)�e��@����)��\x�{MWf�NlQK�$d9�$s�3!�5��T�n�1���l`���z|�΃�����Icw�#�.^Ҡ�)n � џ�Mk����w,4o�x���{�L���u�����N�0���I�H��F�ؙ,��O������%���3"��A��h��7��%��.1��?�%��Å���,�b��z��'���r?]�bJ��+y�����C[��
�+e���n�_�l�Ӣ��(>z5�H�`n���ْ�F�̿m�W҃mMz*�r��T���(ӑ�C:�[<Z�}-�̋\�����o�}��c����;D�]��Ƞ�9�4Uj:P����7���ׇ>p��� t'7�U*���_у�i�t�F��o��k�L^�cO��)rƳW��q�]���L�=j�pv��5�W���́6�i�|�IgӬm���"8z�L����)��3gq����y|!���ݜC�1#
$%�����s��{C��PnPwf�y����E1S�n�ڧ~�1��K!u��|�8�U��V��Ӷk�)������=9x�XW04:+�X}LE��!oS�K���f�V���`Ҕ����Q��L!r2������I;�P����k��A��5�))��1�4eO���~?�r��ZOS?\9�����N�g����w!��t�D�:�%��Ot_z$�8ZB��tm���U�{����O�eYlb}_��I[b��.*nF��D��
}x�;*����\KL�?�"i`IC0Y���&c�Z�{<Չ��e�T��OF��ʇV�$��+ݪ��l��O#�?�ٔA�'iBD�M��"�
���W�0�#bt���RW�ԎГ|�0~���ʉ�h]��R��x����X_�M��32eZ�������a�:����_/��U�%?�ȱ���k�V� �0���1�sE:���E��v�;=^k���XQ�I4�ۄ^u#a?����H*�f (h�y����2��{
u�9��w��M>�Z@~�	=�&�X �,x�8e�ȏ������٤��J{��{��N\�	�iU��3��e���a�Qr�����`��~I���ƀ�yJ˃�c�v��'���O��_�B'�8���W�5z��CZ����g�5̽_>�pvK�����uNy��z++HB`k����U*l��/�߈����W� �-+�.��s՛m�H�#�h�D��jTV�������%��h@�}�\��ʐ�;o ���*�'�� U�(�&�uZj��1���|�(��5^(3�9e
�r�G�����^�����ڬ�{�+���Z�ڬ�N�{�����N�O)���i��?h�L}'B�P~32�j�N^Z��ڤd��^�8�װY���B����TZ!�#�ۚ�Q� ��~r��lu|"�N�%�޶$a�+������e�A�SUp�:�ڗ�z�{)����B�N	��ɩ�m��l���OP�:�����,����bP�Ծ�h�\-��������can����u_Q��9Ϟ�� :{�%��6�]���Xҝ� 8M�+2���YZT�疻��r|T��dd�%�9~�p�d� @��2�у��`x��S�z2ڕ_C�� l��O�?���G̿�K�]|n�"��܃���D�ߪC%>��t�܏1L��t�'\����&7gXA���(���1ИR�DͰ1�+�䪩�C{�~�\}�s.D�����@`5XpI&�W��P�5�ݓ��hG�A���[������Uw:[�3����q�8UJ8�5.�֜Hz2#,�{��p�Y9Rr�T������R�����5wd��%�pa����Ve@��`у�]�E4)a���[lސ<��IIz}���\
]O����5k �|*��
\i�M�Δ�7уh�l���6Πc��r!ݏ~��H�{���d-/�[$�b,b���`�Zⵙ�d���~��*�$�H��X��_*F	��z�.�t��b���nT��x_X�^D���L�xAcx��)ڧ�K����I eW����-���?�;�Pɠ;����������~�����P'���N�7��"9pyjރ&�����N�p8ti�������؝��D����1�qEI�r��:4�&p��J�ݩ�=�N����Ol��d�%ϖr
��"���:�&nXea5��D�ϴ�w1���]ٿ�pϋ;/"`��w�����bC�k˸��~L��d�BYK�W��]0�e?S�\���hЩjx0r����۟0����:��'{�V���jڂt5��b�>�z�v�c��w�����01�v�M�@�Ҽen0�V�y�0��.+{$��5��#_��S1�Y�G�9&�92�=H�[��b��ކ�N�Q�o������.}�& �jO�wF2���/5��*Ȍ�(�|�˟�;�J)��JOd%��v��:Q ��Bp�Xz�6����?�~������'�*���t��(�؁T��[�Jϑ��>-VOk��LWO��-�-�I��S���9�>���b?�&��vq58k��M20u=�t�z$� �ٷs���/�J� A���aC�F&�^ w�9�$�}���;�����,�a,R)b�b��]��t�C�&��d4�M�@o�]72Z�N~�ϭ�.%C*��E�/d��WT���u�6-E�u���@��l�E���g4�}sf���<;�D}��2$b���ꊑ%e1�sD�68��U;u�2���� �`96b����n�w��T6p�Tnm�K�l��U����g���j��%uya�t�uk-����������Fv����}�J�
]]Ms�T50gޑ:�H,)m�E�q��pr���-:c�m?^�ѩFA����;��M0�&/i�d���Ǩ풺�N�ۼC쒥��΂�ǿ�Y^@�N�ݿ+04{^���#�?{b.�D�t��Y��v���U�����k�B E��T����$V/�{�_L�91%�wYs�U�����^�J�(݈��:i�����D�BQgs	��%52��\��}�!�7i��@�����}�U��å����$a�|n�x;>�
p��H��+5s6�w���,�z4f�!_׸�̀�7(�YԘ����o����7��1��F��6}nrZ�p|��4[��?���)�*|АIiML��K^�L��e��?
`�2�ѥ[8�纗 t㧴I��6��{K���7��?X��O6!�BK�S���7T	���?����y�܇�.hE����S$�-��+D<�u���zk�0��js
��� Dph�KY�t�nG.M����6  H$˫k�@������G�v�8����N9P��7��bP-���\2�4Otț�2�-M������~$pO�8H��<;4�SX�,T#ڶ��MJ���xB��U��&
��1wa&)��(�r)�n2w."�4d���V�k�k«��J:wW�R�8�+�̥�h�]\q�;������#��W�^��m��9N��H`��1bR�e�����>���a���Q!�Xp�`A�M4V�_1�|W"�=�Z�w��sҳ"N��o]@>r�������h���3ʟ�APcs��U����-Y/�S�'�\�˔@F�20�E:�},�B�'mY0��<3�hz`[y���V9��T_]�Y��U`
��V����-Ҽ+w��������wLkrn��}��p��۾ϚqI�o����3k�d��h�,X2�g�����\�?m��eΤ<?pL|�PJ�Ș��po!�Їgì���T㫀ϲ��(򔱦*ܤ�Y�rXn�27�P������$���7q/��)ݸ�AK]A�ߛ�j[\ Ǳ�S��4��ƞ�q#����C(��:�FP�z���}�ʷ��5\܃Eyi��� J4����ԢN�����\�0M� ]2��Z���#
�[��H��}hJ�y��|�_2�G��C�� 0ge���Gq����i�|ey�;j4r����5�b����<���+���2%��j�`����r�G��U�v�'�KZ	�
������3N�Y��sQ̲����dse	Co�����V+c�9܏�y���yU�z����SS<U���-sQ|���\���H����7T�US�q�\���	hU����348f���b֤���^~y�A�j��C4e����X��m�;ti��Ĩ�8����|\��"�� /I�Ŕ7�<�ޚg
U��9Z��B���n_A-��C���Y�0'�ũ�y+��wO�;�h�V�˺�Լț�A����:t����.�÷s'�6��U�7�g��t>S�MYt:؉�l�>��LK�b�
�6$�J�b�x ���,��	i�h
i���EB]�7Xi�!&�O��W���0�T?�:�
p��dԎ����X���6���T�(��Ҫ�7܎��$?�iNa��	ր)ȫ<�7u�p'D��Ȇ8X��{�����oM9���&#0��z{|a�J��v?7�(�5d�*Yx(a�fta�0Y�ob��Vx��$5`���J7�!%����[�WL�i8����luH�"+;:e=|�>��ٗ������mW,�r+�^�Z�l���; �3�WkC'?�/lڱJt��w_�"Ǡ�u� �[��.�j�Z��F��+1.�Zg����1guD�T������,�d��d��	�Y#�Wv��~�bw�b�V@�����]i�&@�Sךީ��u�7j/��_2mω��V�u����J���#��6ɸ���w���D��4%Vݜ(�;��kn��:Y���_ʵ�RCh��H��t��^JH���QR�"=�qɧ9����G������-�n`�|k�'�d�Mq2n2���½�"��f�G9Wsc�����E�a�)ZM+Ҽ �e��B���"�9�}b-�8����F�oTY����6���s]�s�bML��=o,`��\T�!!�G�TY��X}�i&�p�ks�{b5��~�n%�H��u� ��ȉ�۪ �~
��0�0Hl��ȫ��]Ȃ�Cn�S�X��tJ����S;�E��K�j���	��!��!K�=:!g�(��/�W�m�q��5�OP�69)�X��m�e�n�F�:}��r��/�����rd3��i]��Xs�`�[n��D�@��g�$n�K�\�j��L���1.�Vͻ*�" ~��=��фP;S@
>kCI֋_�C�wΣ	X_A��\Λ�ǔ�>�J��%��U>W��u�ԡ[���G$��I6�'
�wjo#���en^�5i�ܾ�Q9"W L��� e٘��U�۳*̪�֦&�#��<Uv��֒p�T�2�tL�pk�� �أ-����{��O����t�d��\��Ph屰&��ə�	�ct���(u�����H����ba��6Z*T>��V�x��7�SJs
��蕗�_��)+jY?�:�D3j��q*{=}�5���PN,F�8���#j�A_��N��pJ@i��<8,H���뮇��LKï�Q�zf�S:as�(��cP�:@f�� ��2�E� `��{|�@�+��%�G.�%g��E�.����x�e�:����w";��B��<�y�hn�q��u�T��z:�u���"2Z[����.�Ix�����X d�ܝV-� �칑���?I��Qǧ �z ��bذF�WgZlf�bz�ZY�uo���y�ձ76��ʙ�\�4�G��\�݊���`�x�H,���U$�[ Z}�(����G��� J��J���s�;�$��h.L]H����Yqx�YkؠYa���GmN���4@elu����^�� ��]^���Lc��ha�A�<��)m~>/P��^�iOn^�H��Q�����ku�#�6I��Q���4���l�J�?n���B��b)��ge*�L�u���~)�Z	 &��E��揸n��m���o���D�o&��G�ե�����{�r6{% F���?��<�# r5X�]ZJؙ��HD�5#2成�T��-/�00A�ժǗ���=B}۶�7�̿�E���s��=6or|�.� �F�yF�a�%���� ��+Ah�Q�~F��q��*"-�
����8~X��$�`*��M��0=���Jx!�C�;��,֮۠�h7��aGF�I����$5���=�<��AL �aR+;ҧ�+r�R���@	�]��[�;!.L�j�*�P�9�i�q�(��X�^��ڄ@��	�-]�hH�}U=�;��P�v�
6����m2�D��-��+��Е^q��h����X�w�ÉA���lLT�K�2
��-*G�7���_B��#Բ���u鵽ovC]B�V�!`�`��[Rn>����x�&��GU��v]N�5iĒx���6lʵ�� uf貆���l=��D ȼ {yU$B|��``|���YنwP�i���i�2Fd�9}1D����L�84L�>��юç�#�i�eŴ���.a_BPVΨk��s}�,��;��)ր:{����Qm�0l�	Ƞ֞Z���p�9�_S�v�:$�e�	QۆKc�Ш�O���~�M�	u����2�����)�����u��^e���9'�Z²c,P&�Apc)3�X�x8�s���u`5u�����PAsT�^^@y�e%ۨ0��,<��$�RX���[b��'�-=���ꇦu�]HC���x�:y����/x��$>[T�Qr���/K�<����j�K����h\��H�*HA�h�mj�^e�[����-j/�
��$^6Sa�+孑CW���]�U�
^#���n)$��Q,�ݠW�z��F���E�ՅG��G�D�=t/r܍	'��)|[6^�?F|��݆�:7稶���z����zȹq��Е�e1�xSkG��ai��<��ጜMX)�g�9*(6���G>,����	os��ts8{�B�$#���]�:�)��S��ߜ��4�$=*������$��-F�^��[Bb�Z��̀�5���/����� 
�D��~�L�`P�C�=�b0|��g��� 齃�d "J`�����jET>"�;G���[�C�ـD�)��tز,~v �	�Q�)~yD�1��L�ژ�b_u�ˠ5�OU��e潌��fh��7����GN��D7b$��>c��DH��U��{�g�d�t��i��y}�,/!��ku�������7��#s�6>yP��Y�-��s���LnO�r�ԛc��E�X��v�:���%��X��Z��ݧ��;q9K��t%��|�a�NCM�d䶉l�R�r��r25���I*�U�ȃ�
���L�8�nZ�lPSP |�(��V�eY�Z��$�"�պ$�yn�Bh��؃-d��I�(�_�만�tU����s�,W�=��/�T��=��0ئ# ���@�6��Y���LEפN[�ŻB����j<�<)��wz�2�J�	+SP3��� ���|/�Bk�Y�?�Zѽ�Ĕx���y}i�Y��'��Idx)�� �ԋ�M�cW��z���yas�bx�Iv����m�s�j'W���l)R�.���:����݉���k�'/p�hr�3O_� ��Wl�H��p��.b}췫���O@\涚lD��������_/�1*�#J?� ,^Rd���Bva�ㅑ�~`�mwfzV�^-ŕ��{�w�e�v����;�Y/�,[�� i����!��Q4N}��yʳ"�e�����m������Z�x�{K+�C�Wqz�R�ڢ�>\Y	���[F����B��!�M��:1��5)yQYY���yw*x��V�߹����Pzk��lY/�Bƌ']�6��?rM����q�"�N ���&VnRt�ʋ��u�{$7
��W��!7�g��P�M笍�{nƃv#XN��oT@��k|x��YW0��h-ͨ�G�'or��t�sD4V���_'߻�#���M�Y~ޖ�$���U�E���/���2�ޜ���Q�����LN�T}����A���ܿ��I�!�(�L<���0}�R��C���P���5c�ԍ�9���b.ROǰR�-Rc����:[�w��7oM��zn?��Au�o��bC�o�
"�����ϮW^���֍e}u�I�c���"�����y�8�ڶ�:�AI�S�����/C6�|������$<���D��*_ݸF��>0o�Q�bK�BǮ0E�E��#�V'+��������[c ��	+�sx�y�'��ƎhJ�$�t�V�U}�A�4�cXH'�iF�	\��,|�f�	x.���C�o��k�#Ea�/#��d�W�2�[<�5+�\����sT�3[J�?1�;��eO�U�'�WҴ�f��R�پ|("u��I��~�����������s�~3��d�*��U^.V�y2YXE��ҡ�:�!��9��gٱ��U�u��6��h����@�����<�5!i��'"͘��^e�D�ʙҩ��Y�L5l�[j�fO�v�ۏ��U8vD��@e���I��M)I(�Y�tG���R9��{Ń���(�7����A��p�Q'=�ȳ��'��Z�"x=,�mANd6�9٥F��½e�${��hg���ԡ)7��a�r�H�!ge��Y�n����v�,�����P���gk9�2Ĉ���Ann}ZU�_V���f���]��V�C�����t���KT0��ˆ�b����	M�mK4q���l�;v�yq=:��<��ؘ��X�I�M���2���H����H8��I��&�B����j4N�,���Z!c�
e��W��P�x��к�=�ƃ��s�$�1I/*��>��`�q}_�8'�������֨���΋��F ��7��UE?�2��1��e�I'��B�[A{&���Ȉ�� g�g L�+��S��AK�� r�����\X=�3�ڹ�F��~�7�O����#]��^R���?*�n�?JO�s�KH[��c��w
�	"��d��B�J7"o?!�#iKA`NM&�;�@��Ac���-�&Q��]��rm��p!}�&7@�N��tF%ؘ�a1�8o�Ds9\� ���8��8�dQ��vX�F� _뫟�����u��W�q����\�����Lfy����S��>E`r]͛L���z"�<%�MD�$q>O�̛<�4~� ��,og�-"�N��Jٖ\��n2�d=�ֵ����3?�����/���_[�̓�KcƧ_�]���QS�� =�!��o�6�\�P�u!������ӓ>�+@�0ޮ�ᝮ�D�����*����XAN��Rv=�A*�/��8P,F�CgGQ��-c����O_���Bh�Y���l�E���VB�]bK��!�L'_�',����j�;t���,�c95W��P{�Tuzɳ�����t��Z�LDPγ���݀�=�O�hs�G�Q[)Ew����V�\�Fy�:��f��jl>���u\`��O�5ĮDy����dTFүȅ��4��&`�9����ӼC8�HQK��AW�qs��݄;�8{���;,$�a�0��~�%�yr~�yMZ5,}�VI��A�r��Zn5�hY���D��Ibc��U'�R�Vd�I���V��6��������*�J�b�7z~U�?>����0���
MG����p�2�d���6��͐��A���g'�\H�����n����D��i�dr�Wm!^a>Gf�J���QI�51�Tp�����:���E�4ձ�_�8�ɭ��;&$ %��^9���{���im���H��1��{{=s���Ni��?j�g���'�MU����HfΑI��۫/y�i�Ԉ��f~ya�d��hþ$�뫫��51ƽdb��ܦ��)�qԒlt�1��u6GfZ ����M6ٕm]ܬ�����������%&�f�� R�X�N���qx����A�Ez*�
��iLi��.�ۧ��߈�,w%�����j��o;o�\�������P�B	"�L{�m��N�=jM�g�2��Ō�Nl�!����/�k��C�ۺ�f&/�F�n���|õ�*7�B_.�����6珨�#�D.^\jD`���(Eܗ!�v~�-�:\˖�*�U�s�ϡ��bl�O��د��g�vbXOv��QL����x򉺈[d>��-�S���L�P%Q���c6~#�T/7���4����XJ3�I�������}���`T w}��\E*���vI�((�Mi6th�����#���_t@Oz�S���k8���e1�ɤV�f��>����f�U=rt����x�(���N�5�0�*f<��o�?�޽3`���|$#nw�O��f��^izgA���o$+�2p�fV"� �?����{�Q�K�~q]?7�I 1Ңr�>��O�{�%����?؋�~^�1��膧~����.
���=�P��v��xg]���e|Ӗ��(#Ga�b	�K�����ö�p��<� ������9&�ҳ"b��ɐ�|u����HD���86����w�z;�'(#aZ?�9o����Nd���.W����Xnݣ�2Y,9���^�KZ��Aͭ�j����C��: ��i�­�z�߸n2tA7�A���>��^\�g�����Z�+�����v��'r�<��+X/�]�^��]JVyW٦�$�tr��H#c�!H�U+�}x?qaŤmq�Y��)bqB`l`��ӧ|�Rz�����&�߳A��L-����Ɠ�~�����{n��9�M]`1�w��Dܝ��-*28��?#>�;�M� �\.���#���h�[��'��x�Y���>���Ud�/	{�{��
y�i��x1��zZz�_��S�1����'�E�( ^����IRP�Ht9�-s�7\����v�����],��xg�y K���8�R�A�a~��� ׯlq����he���6s��*WI�h4�4� ���v�cH���U�Q�=&rL������m@ޣ�t-!X���A��c��̿¶&��jK����Ogs����.�uS�����W*c���y'�� _[WmeA�w��Pb#~���a�g���I	�C��.�"N�7�A�T����bX��z�%������P&����.�R�\瓇�\~����|۔v]j��<Q#�Ud���^�{�������Q9���z��{VJ���χ[�g|��}����N��r�"�C&��r��git&�_�	��:��W�EN���l9�l��|U�]A.b��<��t�����o�9W��@�*O&V(�$�AS�2�� �	~S��Z~�љu�9��sY*
q�"�N*��k�yˣ�?��<�嵊�E���N��������vK��r
`I��2aZ�zD�ƛ�t�P��S|_tC5"η�i(�sx}C�[< =9ҡ!
�����׾�f�χ�N�a=#{l7P�̲�:�(���lk�lDK%ʈ�Dgi�K !S��Z�J9}𹩲7��>m[&�5A7�(o��q�"��B�!�no�����8ܥd�W�����沶H;>(��o��(3��#6h$n��7�,���˪���#�u�':0��˼�~��l��E��a��ۭ�f녏G���gp͘�[��iē�^����o�����l�a0̊l��'��^S�ߚ��wHJ^�a�R�QJz�7�1�iJw�����%s&�h2"�**T],YSJ��A�����s�;7�����1A�Rɜ<�y�E�����KF�{1\�(|[w��g�
 ��l'�;���1m������d��J����צ��3��YFIq��cr_�X��:c�	�q-3YWb	j�[���*0�W���U�Ea#�jx���JUM�j���^���0�lp��+H>j�V��T)�z��2J�1�/��g�a��?�����$�Y�p�^�6@m�f�=T����vb��N���z0����ra�= mn����͠�Y2d*6W����V�D��.W��kf�t��	��cBҩ�&� |e��+3��⻂��]݆�} +�BTxY�dsw��6Zbk�x��:_O&���A��fnI%�,�f��G�*���<6���e�ES�����<\�*�W��n0l�(��jz�ʸ���ƌa&ouk�<B�!��@�I�_S�Xn�)/��x�J�4�3��!���2�YhMH�e��/;�}J��i��x�qVv�B>�ju��v��հ�H���9��4���n�����KO�`��<��Y"z�Dq�����:^�G�HHz˻I��Е8�D�`$QԖxn�O/~Ԃ'�9�I�$��el�t�'��@T���HGڳbL�W�4,��C���#������_f'��ֲ�M�ʔ3�x% �OZ�P![��L.����8̯d�ԵXU |�g�T#�) z�$�auKzX�����l�WCN�?�p�3�b�d.r� /
(�
�݉�����L�y���Y^]������G\0�>Z���q~=��������SH˃�%����c��[?\�@:	蠲&(w��ǫ�ߧ�@E9�Δ`v��h�O�_@�!�aU��'�6f�����r��