��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F��������n�oJ7���ˇfΡ�%��貑��n��FF��^�T���HFd,���0bzڏvA7��Z�u�f���T�Pk��%����ý�/^^�� �����_U4ʴ�n���z�_���q�����Mp'���l(q��e5�>��]����>$96ƿ�	g��'q���#�z��o���FB+�o�ۚ�w�fJ;b�AS�|�j�O�
�8��Xc%J@�ٮtxp8��Ʉʈ��"�"�a�4���V`%�"Qe��0����o�=p������:����ٹ҆��~��}^l���v��U�"_[����x�L�M}
��>v�/N�����#�k#�ɑ#Q��/��V��m|H��	�m�������n�[Q���@�蓸�*�☛�r@�=�A\б��t�_Z���gU�ִj�Nw��GE4��� ]z��|l���yKs�¬̱�o��!� ��q�'z�bi����!��
x��y�"�C5Ǡ�������M�����o�G,�*�_�;�=I�p�xw{��հ�j46o�a�,S]���F���ב�pZ���R�����S8�����ǐY����n�[ C$2v��Q�Բ�@B�Ͱ����
Kzb�����5��ʈ�{����ه7�^m��V�Zl���$J{$�^�f~}g���O2�UE�1�Nb������@��3�
CT�ub���|+������@xJP1�L�Kv�)�y�u:�_�ч �-�>�8������Z��˾�;"E�f�q�1�7Y��^�j/�N �%
�׀��nʽT������y�T#����wխFP
������;��[�#��=�.m0N�p�M� x��V�󢠯n�wtsm�;���?�=C�XV\�L�+�Ι!IdX/�ou��3�)��#P1�-f�W1<>�P��;����v�k�.�
=�=�_�3���3h?��vY���HbaS\�C3N��!�,�����iKm]�\S�����k�c]|�G�7ubv;N�~�x��ק� D&m˜��j��q��mm0�� =���b!�f� ��?ՏR�ĝdd[=�IeAAY�衉1�T��������(���R�>�������v��#�[��� P,���2А�	���̗_��H$���K�m��W�zt�����L��w�N��*IOY�9ɪ�S���{&\n��~�]nk���
cΗ\��y1q8v�f��ȯ"Ej��&u�E�U�t�lOܓ� $V����
G�9�C�"5K�Ͻ65V�o�ݽ��a]�a�P|��%��p�B��>rWk����������\�+�=/��� >$���od�I�$F�-���H?��8��=|���\P���S7w�wib��GD�I��&�h���gB��mwv�p�	�Y�9ݫV��~-����N�qE��m�uE] I��l���erfi�6ý�onFa�ځM��eң�B-/-�
r-/kt6OC8��Z#@-��Tr����5�J'�T���_Ƀ ����� �#4;PP�n�K�`�y���'��h�bR_o�,��D��[5P�1��A�x���x���'�		e9�=ʙ�2���/��/L�ah;\�[6��I*���q�Dr�ǖ�+$Y��7,�<]�eB����77�g/c�b�R?]k=���^�	!�~A��(\��_Jw�~�����٢鲽ٌ�Y�����3<b����)����xщ��D�ŧ���ڬO?4k�*��r�z��;��R��Y	�O�Bcp����2Me��d�ϸ_5��!�p�{P�l�@�LS���X�B:�Y	�ˮ��d"�"_�^����)�U�E�!���6(�\��26,���<]�\�7`;+��ex^7��E�~g�-��u�-�����r3;i��?�<�BF6@�==���>�4�gD���Jo�90kO�y~y��!,�7�A�&�bU�Ev3������yY��@/�յ��E9C\�6�ԯ�S��.|xH�x`~w$�Ǒ^Z�F3�J�An����I�'��K�)�)gfb��c�eDގ6v�	7�3�E#!��U�tǣs�,�N��'/�
��+��Nm���9 ��Y:��5�5;Y�z�����GX�^ �}�7�k��wň͙�hs"��Eo�ާ�x����I��cw�	K�d�$Eh�	#�o��"���!��E���MM��$	�~G�aZ5��P�����nu�?�v�(qو=Ѿ���E��-�+:G�@@�#W�~�䵓e�UHS��@7�m}��4�>6Ͽ�S�YANb�:>�^�[ �M^_!0[����}m���:(����Z���J_".����5z"�%A�΄v�1��R���i�ǭyy[WҐb��ܱ��P�W$տ���g�߹8�`�BuR�9/���7�9�څ�'S����ڼQ���v�������%�	�8^NE��pS_r�.�����O@�HK��(�^̝kQk�ܼh��-/K�xo��IX��'-(��]��w���tw;az�w�E��� �'k���y���u�'~�t��*�3[�֯���l>�?da�|���0����N��[�H�����-��`�2m���� Zy[�M^�,>�m��̶g6�fr?#+2������0؏K�8܃�&^"[��!�f� �3^�
`�����v�?��u��?��M�K8Y<�gs�� �"��~������?�/��A��3�/%����؛#����A '<��{��Õ�^5q������p1��:����C���!j,2�kݱ#`QjpwO-i~������F�:�쉌K� ���i���j/�>GXWY�#�?B!�d�������K�C|ߪ8G���f3Z����!/���c~��]&��"�ߊ��&׸�n�z�(_��}ᇦF����>�A���F�C9��\7�꫏��X`w��&û���W�̄#���  a{=�!f_��U��P��r` -��.���.�J?�N:FE�DI�s��d�'Y�֒ e{U��x�� +���~:��}����$_�x�����'I�VNf�M���o�*E~�c6,ѳYkZ����}HlC#31v�4���"�4!{ize�x}1,�g<ph���t��ҍ9��J?9���L'��6�n)�B[4H׭�Rs�����q}sSBN'��4=�Y�;��d�2_�_Ka
S���y
��]M*o ��qp�:9S�O��p�BS|
�b`�r������4 �<	�@G}L�j���\�}����^�:&棰��a����q�Ϗ��e)s�S�FR*,�J$tT�2���uE#Uj���ߐ��Z�3��&[;�����o�y4�p�r���{._�р��2 #�>Y
�۲����ƀ����vK�0]|�	���w���t���7���t\��'��8m�W4U+�W�4�G��f��2�|��}� [��:��ъv��P����{��(�Q����4�ԍQO��������Xw��k�!����������,��l�j	����]xѠ���^`�)*��9�#֠�.��eڙ��]��;t�'=�V	L
�#P�Q�����;b�G�Eɠ|
�~[��"}_ip&h�-2�7�օ�|�7\�y����_�o6V}(*�]����Vp�bP�[��[b��{�K��{�.�s_�.�26�!Ġ�6uE��u[��yl���\��-�y�p�3�G��Oᬝ '��_$��Ɏ`�V���)�[Еb%����.d��)30W�VЕl��tB$�L]����p������`���@�|	�F�n0�/��o��x���醂5W�^�F4P��8P
Ի�3���he�?��vS��G�U�Q���S��o�Z�y�:��f�f��o�E�%~+]�" �Ý��l���T�
���E�}ڜ�L�V�\��p3H[OҸ�>���xb_%����I�T-�s	I����"�#�k?�J8�7*��`�EY
�����y[hS5�Niվ��6�;		Ȱ��$ْ-ك��:>��8GD�E�I�ڸ�lￊ7��h	���Bǿ�#�t*���Aa`;�/sɄ�z!{����'!��5�� Z_Z��]��@��Fp[Tƒ�ʨ�7���3eu	{6�o7�(���#Q|�^0a�\?� )Bs��
qC���p�~���jjf����"�;�����󦇚c̝�����kJ�,l���xx.����V[[�/��/�����L1^C�x���� ����{*JƟ�[9TV���շA���s[�۽�N�T�x:~}�O��{ ���ɍ��M��N���s�PV�O���0�9y�a�<���-���\S �jd&^\ƨP��Ea��%)jmQ,��	N���c�� q�\NϊF�-�V��S���D��(EY���j�v �Ӗ�Y8g�
=X��.*̊-�"�pހy�μ��1/����<�c�Pj�#�S��idCh�w߈Yl�R��+3`�pm�6��L�6�ք[��[���=%�Y�+b�[���ۜ�9m�`�_m���)M+�_hF��+�s�FW����@OMm��Y��1~	��0���b�fI���)ڠ�1�Vd���4�t!���Z;=�ד��K+OT��a�r��Ƣ�=��5Rz�<�DHn��0,��l��-:�(j.�Ђ���b�i	 �&�6�ٮ����g�a�O'��I-4t�����cC}%2f��61r-?������+�<xD�.���p��s���/�)݊A	cl��V�]Xċce��K���zh?�w̤(�/�?7��//��;�,��4�n����k	"L'�ds���	55�`;���> �q�e���y0}�gOxg" �<M%�6��g����-��B|��������;���/����/;���x���O��ɐT)�Tp��1ا�n�6���a>n7�_<�''�G|Uƌ�UbyJ���@A(��bfJ�ٔ�\��n����Ԯ�L#̆����hR0�]��Q���+�$gt����|GyݟI*�f��rE�h9�r̺��!���^`FC���a���F��f�ӛ��}��oY�X�Q�?aEt"»�$�=�c|D6Τ�]*k�����0���f��?A�H8���nn�h;R��Q!�%-z*:ȋ�O
�ZE�R�\F��A2q�%>1ߨ�����!���-��ٻ�Ȗ�q�u�����:�C�\��Af$a|r��Ԛ�$C��ᕄD0;kb���p�T��i��
z�	�L��=�sO�y��I�vE��D��[�.����.jA����
H�eIp:�)���q��i�|�`�[�Mq������$�K���"�-Xi��-UO����4���@��o�B�r�;�������D���U���k`�����]7�:ps��z�$�<��lu�%W=U��CA������'8r�(o�x���Rx_ڲ�Gnl%�9���b)'�R�g�d�9)�8���3�q��p�*��U���:�L�u'�w4ՖUM�h�@��vl�'��D��)����+̑�byBt��7�������y�̏���vEI�C��~���^�I���++	����@l��Y��2��9�I	�%�&k]�Fd+�� �Q���h�}ey��e
lJ��fP�u�����7L>@n���ug+#BZ7�f�2@ ��4�_�ѽG������5?�WjG�Z���������篟����5H�J<��L�aZbw45�֌�_knVY��*����?@a7@��*f2w��δ�əq���:��F�H�	xq��At=K���
сf#��[��y��kf;�iU2�iLI�/ ���'n��x�q$Ԗ'c_VS�,^$������z�B���7��sBf�Rf��A�
�[t`LO�u�K�bғ�=(���A6�[�j��R�1V}����P�6��A+�V)�1��tE���7��ZxW�%�&~;�dt	���'��z����2(�^�9���[.�[�<��yN�qt5���qs�ƹ�Nf�U�>O�|����a�',����|5�e��LQxj��0�C�4C%�!�}�oB��wT� 耡�_T�Rg^˚�k�GQ2�_��ane���&����z7�K�Bt��A�s�ӌ�sߣ��r����[)
`���\B�q�@�L�=�_����'y:��wX�|B�'��X���$�~�ץ�jj�������ˬ�)_��hwD���#y]Y���v���`%�yH�b�iV����z0��Ŏ��؟ҍ��%���_�}�ZYz�Û���$�/pD#ԏ
���h~0�͞��'��d�? 9�K���p墏O�׽��$:$��S�Wj&���h��#媍�o}JHG�-pe,�"�W�5����[�n�kµ�J�� ����fL�­�F!���=�^��U��i���x��q�N��
��݃��YX]��\0ڲ�x�1���r^�3̧�����7��� -�`��)�7��Ϣ�����L��W��^el��]�2"��\�>��l?���b����m�vz��A;�2ˇ{�[��T��)���I�	>��p�3���������R:BV�WJ.ǭ|L�+='��TF�iW���U��G�Ԉ��[�t�e�.��Ǝ���"X�6�Z�RX�K��l�o�tޚ%���:h�H�Bu��ݍv�3��%�~�&�I(����ݔy�,O��%��2dE�M����'pD8\{�������>��S]鼾����SN���tz5�F�Y�4$���Ӫ���ЋXq!�e�z3��e��3	�H�HB���u��"7M�R���S��8I~����>���B$d��ƞBҼ��?�p_E7��:O�r���"\�
��;��P"K���h�[��A�כ|:{��¿rUA2�X��e��_�?D���A�S�)�4�~o�S�+lw��ЪS���Th�z�Ȉ2��n��rlo������il[����@�	e%[zY+ô,�e�<���+�1�Z���Ջ��q�*k8�9`�af�e5isK� O�3ߒ�{�+*7��P���"녕�o٠�����u�N�?<� �&�	S�D7q剦�!�;�u�u��*��.����l��u��K��p�����C`F0]:l