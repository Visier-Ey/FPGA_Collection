-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
--pragma protect begin_protected
--pragma protect encrypt_agent="NCPROTECT"
--pragma protect encrypt_agent_info="Encrypted using API"
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
--pragma protect key_method=RSA
--pragma protect key_block
kp3XwK+4EIhmN3wSsYbIWaRMrOGH8QElTAKL3/8pzfxBi9bjFH/24UbmUY963GTK
Vt7Yn1YyQy7+3eITfmUuTifCdrepjJLiJ2H0f8Z5RO6MP8X5w/L/4D3x3jvlFd7q
2Cm2kgzaUexYd9KBdOLIrngxYo2VgEVexPQwYFsdlEbgkmu6AMKf9p65ddBBFIJe
jqWYVw4gYW+zD6ZB66xNrv7FWrGeK/7gSImxLMhqZsPxFsfhFQw5yppGi1xV4A4o
xTfg6vwU44GZ7YIWEO+m4Q+kj+w7FeFbJFMUnkA3J/IVcS9S/uXhI/CvhYtcq+w0
ZpXEceYSqScEJ1zqHj7Hkw==
--pragma protect end_key_block
--pragma protect digest_block
KEWxhRCmXJx6ugMQEmBH9CXTZbw=
--pragma protect end_digest_block
--pragma protect data_block
3fYsPEKw9CzpUJaPblXrkReLnF0GF4XN7YA55qusRZcJuM4S0w4R7VkqK56O1lQL
kZ2vbPc2V5wK5uqvxiBB9RGbl2LRObOX637jd/WZ+WtLlqSUwdEYw5CP9CdTmd00
UDRLNT3+SpC1h7Im6wW47LcwBvtjpM3yeEeTLCzSBwoczaHdnwIXSre8+kZtMQ1g
pQ5cV2DewNGkwbkoaEkju5oLTsA+f0TUQX3Xwjiwba+R7bygUNItNlEryzrutf+C
arwXGBRcQZo498RxvWn/8GDx9v2Wn6NKL30TXrMfFqcF9qjGJSHUIkExfHpl0iD4
x7HgH0H3zOSCZ1yW8qFObGWQUlIX6pSSoeIlANwiCg7vfRZUAPlyZ4W6pp/nR+jE
tpw6b9EVA7dhGFJKzn28DOxaWLdW3yr1ksCZUgyVeuuCJKsvIDrUQmbXt7+nv51A
4Vn2yh2jgqStrNMg/qqW5kwhO+nf8MhCwHM6F7DzB0v8q4A1caSPlIVW9/pDj/SD
L9cN4ZAob71+LUupBsA9jAIZlh7VsbyxTpBxHDgjgX7jzSsn3N2BVY7c+32m2Tx2
f/RuZhR56d/1DjoycpmTZLGdR7V3Uit7hyjtG1ApkfPWksgVMjHIPNWrvb1+ohFf
DWQHuJ++DRuxqyjZ3c8cFR5wcPXxTId/AO85UBc+XPPLHzLVsC228NmY22DceJm3
Q1a11NR4Bcu0sLtLMXlB1D2CF/Op9zWFBod/TWNpip+ShUK3swTxVUGujHFrONNv
OlEkIWGojtP7sY2U0/mGChSujZjQFLMBTfUBONYsyglFzeAJVBpF7pFyAIviht3L
msqFIYp4w9uG6OYZvD5HpzK9d9lsBkvVS2K+/zBauddeb2IRKJiGgorO1x8XuxiI
n7R1djtXitJ0fC7+2DDH1E+0i9mpf3+P0z2BGKi9zVRliElHG4YyhzRzjKZI4VWX
h2jzwEVTSQtWIUidVPuOZm5yqQa8WB2okWZdP1yIO3FzB/tN+kI3tRA4nCeFj2g2
hE6TDehNnvy1Nt+sa+2u7c6JUKYcmNhDlM3zQdhgT9j5K0yjYxGN3xA5vbSa/DVC
Hwbj/Qpuhdbm201cEAYuXRq/RIccI0a+7cM4ZukwDSaJ9UQa9otAY5cZwE4TW5P4
fc+i7aM6Vg9BY9WVLIKqJxmWQ/NmoWG3Zb/od9uV+VMNFRQ6hTrAdMd0d/aRNsez
BCYNKTe0gpwqyWbsH81+OGwWcV9IV0BnCuOuWki4I5RmNcdMM4he/bAkTQWDNLTx
hthT3Cevq+Z/YPnVAvVwW/YctZGKuEFInTrHhf+KzZFDOdQWUMji8XFchqf6zcVv
wmUZZ/u8DwoUSJAyXKUDMeD0UgFFb/t3CG6ZCrZv5PP/bt8mX3ZSCmWv1nnamVMW
6pK6wZ+rruGBAh7PqDNfdTbmrNkw6g3eD3RzSz30vpYuZy+zeakxDemNQ+kbsVs+
pN5Ck1lsaEDWNVLDOHBUxgAyVKmnc/wmnw1wERbht9yc9t33lJA0TfM7LPPiaPBS
3xBPHJ0Fynpujlxrdz8bbrGKTumfH6ko8xJOR5/IcSCuyzQl/sEqGp13XqoipPoQ
mSPzSsca5LUZ/Hl2ZaAWe0Ygjnn+F58WO7zaMf07uUP8zUqlTig5IVj0wvVSHnC/
Gc4t8yJa5hILdoWoUOuD9wWI3Hg2F8dVj7pe7OhIhdwDOoeHeVn8MIo9aRrvSsr6
tf5B1vCyvJy/5M+q4vq350p48kpAhqHuKoVxK1qzgPcSA8TMd9gi9id4W77qCgJR
o4hKZwhytJ1XXroGV2yJ3n+cWeB+pFZOZ63iLHSR80XzmBIB43XyQHA0DyEyF+Bb
Ojyta1s2UUawgcZ/99gq9FxeTodTwBLHCLnxOAhweNHiQbvLJNA9hJzeP3qmVmlk
S49VZbmoyAXbbApUMmbr6F+zLURdRmyIQvY5lgRlKGM+xN9GUhFjo1Qv6v3SQbLt
Umpq5olgCGrhsLOgcfjcSlaQJoX9k8cgy0IOcb97k+JPW4jP7MinS2SA47lQuE6X
PuV3eRwTWd4GULR8pwDcrasHFsH16IjAVnqYgMcdqevYwcEtR9X/QvfV+HpMZZpz
WjBxvfJaMNPz+ndxRZwCM+Vm+AUr0NTaz28663d6ondpLR+mU5SjLSa/NaviVoKM
YdXo7Za+rOYEQjLYkkJ2vQ6C/WUe1Y9rHWhM5HolakpFSAmAJA4oMjxT8Jn5lpei
4JbA1eV3Sb94ERsVfBZtf2AZUy3HJzzM/3mDvaciyITT9yvKvcM9JBrUuhYr/Syr
0pigzQIM3J7jTqBlFFzWx15F2sKweuV4h3MPKlsOy8EImbm/D2CT6BdleaGwH3ze
qRdJWJX3b4SU2vR0nCeTMwxOrQXBx0mRfyQdDgciPkV5Q5fclL6GhkP0DvAQKOzt
KsJTskjYjY7lSe9+jYijyUQWVvy/48h6rfZQaqqo/JAzeKAXGNft84FTMaxd0fIe
WCO6nFevMusJHYA304gopteUqEkP9D9bfNVaTUN9X8YHJtC8KJ3T7uQ0yFsMmF06
ml9FmXbI+iOxheuYC/zJ568ZsXv3SdPyTCwrVUDb4nQuEJXj6n+4gUKlWaN6CGbH
NMsx6qSZvpDZKnhWKHozBStE6MKC7F7gY6XDnR7ZUGtsfWeSCuxugzh6VKqggLrF
hKsoYKxuIHl/VzaKSEUkOrgdlB5VTW0bmzBSyQY1VoQBOt2ClRCAW3a+t1XIw1MS
rsW/vpCiA6GT/Z920t/04CT0khUKsq2G0wFfqhbpMxS3GaOdgjONPiAzGLLfx8um
MLBTnBJjAo9sexpV5YhERXB1+Ejox7cHsAzBwJ6nuTgVO+aYdk421Zc5qCZgKNf9
ZVspIo/s7Sh8D4p39ABX1UJJP2zPs4wBLa8iBOjG01ONaK30UYVfmEf0heyeL1tR
S091/vBizIpHAYQ9EQ0IXt4aXLndOAaCh14EpI/O+/A1hD+2DEib+pCN0BI7gvuO
J0uaMumujsQpOxQki3VX3ZVj66Z0zfAdTUdBV7TZ/j/otOXhfjes46LRfk4dLc/f
9WdQJQvNHrmNLUkyVCu2aTQRm0R2Xb1JqfmyeoTKiZKKiHitEy2XMtwmKGbQ0wh9
ny+41rk3+VI4jwtcBtz2TxrAgz4AUdsRqVHBsGYxi341PyBiVYIOxaIzecKOFSbZ
H1SuU6sdyDuhgSdB+EmZrUdjIvdQinMK9gbw7SOnlC9Yxcbz+pUm4fGlvOVKntyT
ahyWdGjKMnCr/WOVuCTXJPREVisicWddkz/YXncKhrOzd/FhxsBSo75lBhmCznNF
fJTOqLr18LZ4RQbrlkq3mnAzNe3ofGxb/W8Q9lCkOjBXrNaEVBOdLI+uT8rn96SQ
yy1xMjv6toSx06Nx/Xh9i9HcFzadI+095bIpn4M0xU7SiUzY+wqpK7zsJ+UjF5tb
mB3ckUk3UlMKz30BrL58Vl31TJuIZ/pfVban2Cd+prW0HU8AfJYpu1xHlh6fz/AQ
5DxMNs7tPCG456Pl4h2dG41GoMhg0vi5NNMXkx+h2d7y96hopZgqwSllYXwx/5AL
6V4xGBM4GPTB6Hevc29OIOdVC+YNH7auO+fsZ/b31D4kth5rAzj3dfhkHG3Ch5fs
0OB+SvH76qhNQb0o1WVQJwaIt9ElFT9W1WkpvVRXvgxQsihcdocOa7NvuZZ7aC2R
qPkmERIiB41Zdm1YSeorNWCo0qnXk5oMCJgykXYwJaSw0Qm2yrhT/IcdcZie8qH9
ZocXJb1O3FubwwKa9SIRu3iSj6ZX54zzGAfSw2uMKfIsdkdBTA1HSastam317tpc
mRIP6JqJFLvH8fgwnM8dYXw7UKJomGmegSb/n8ktAAzdswkuc5yr87XhZYmxP1C0
relHnWHO82bTPxw4CU1Bzay13uoRGXhcDf2ONOZyj7QvaBV612/5u6p2aUohPEdb
FbRpoinP6cWNjWFSlSdyQ0OUueZJ9GdxeA/iGWH2+uALC7qi+fPhbUlB8SQk1e8+
auUngsL8AlXLEGdT/ylVKA1RqOt7VaZD82Pe7b6J9aMfPxxVwAxPUd7ZdaC4xrI/
2D0L8Ytxu9LWS6MU/SMyO5AACAvjAQn5d+hxlEoGUfpeN10k9x9BHXE17zC2l5+o
OP86wdcA6FmQAwF5HIQSKdd36nVOMl/8+puK3gybYD3EBsQk9AYUQkJikpldeD0T
/dE6zRp7+N7dWl9g+GqALJ6joDtztHgWB8najTslSNKefkO+wcLoKLRbTnqBvzs7
ZSRbC2/6m/K9TJd32y3rEDl78yntP2lzZ8wWjmqZ/o9Is9axpH0R9lux51aeCF7Z
RkqVL4Uh+9LNFwc63gWIiHrojlgWWhl4GjTIC2n7WUIuhlXNvtUC2G8n0nIQ2VTT
LXJ7Ue4TyjScgG8hia6+lAQXFLKU2Er2X9YQGERstEME1OjyfadEAuS77upIwYGu
odQiFNcbUughnZbK06KRYmUxU4WFpU9CPjlC7DcGPGNjH4uRfNWNPhwsAslO3FAU
gjQcM9BS74rDp0MWhylPIJblvduFZR0/jBB/xgFwA0XuBa4D+0XZ+yeuXQUmJyOh
U9RSGgT05xOpXgTDPZBiWt5dwIN5RLua0DNJv4HawRtE15pn3EElGoVvflAsC7C4
L2IycBiE0oVfAYL7fHCdPyWn7IBZjwLDJZjjgNbICL3iy4QS2PUtmt2zX3z7KcY1
OWu2fHohXf9bzcinixaPFYBSNnz2/NYK4LAVjWO5qdsqvxaV5eqBIjeiZI1SdL4U
TiYNF4l6zVcpLKCupvEO2iebwfSwu4bx5VEaw4TpwpRJfOrWOCqtYRLdqQyPqLaB
KCMKf9NofC1QRjv/w5rQ6mEZuVSTgrgk4XoMWyfQLoNzua+qDmE2s1nhCu3oms+f
1xYjqLOd0HS/rGoaxwJWRGi+kIPf7D4wl5tiXrycTjoMNgwlnMgA6EEcjZTYZLhz
2J+knXcERd5GMVuoEowK6Qfv9O0q9lMzBhgtIA82Ch0rzmouplDjTa4vkBxTkL9E
OuiO4tena2q1ksi2tZGAVRgqrCohWmRrA5Zazpfegh6dp8ikFw2VFCM6MxJmgPK4
7sPjri3DLB9poZGxFs35FuJW1ryNXh4o/sF85oqC72nix3XscgK2nHQsjZM0Td/t
wyFZC/M+w7KragF5Zw3UAfL4StNXn+fZaSsLjaJrtYFzsJMMW1/hLZr30IhVsdmM
xNfpUOmGMS5B68htubr9nc0mbp8V60m+holpVIAEeLl1Wl0gZ3PLPsOrTLif8a66
15izZoXzzIZlV1CSm67EJd9o++aM0YlSMakAuYMYqejwme2t/VM/E+3lY6pOIqZs
sDOZWnALhdTkxTvNZn/5haMrUIG5wCMMoQTNmQB6LO7rceAUCOaEq8Jknxw0GEwe
5ehBtqZU7Rw3R8kG8L5Fzptu74ePTwYFY1Q6GdEvzb2leDaAW0GgKWYg593ntL6G
LeGVMY2ySogHmNHAzjggMCkz62Ne8Cblqc7OcghyjVnUG3yJnsx9j4AUKJ7fZkVz
lc1n19Jp74iPfIZArN/9v6+xuvcP8YIcpvefdsO7VyUqiDSGx9HGFXQgTjBCt2iS
+4LnmPYavINkwdvTDmsl47xtkLqdNw5iNWOf8gZwyfv3GVZIZpn1gKksdovdh7NC
JBuOL/UIcakjF6Zs8w5zID+7sCdu6KKGZAJDk2wtRTV2BsN3Iuu4RjBRNxO/ClsL
OwEwnXnppSVoGWX68tZWxOJ7CyYzWmB1HbTDTkcv9GjTlGm6+fg0TjHD+sxQsdJv
PxSnf50U2mjg+5pdNTDrm8f50Mdx3bnxNxJU7ctLjU4qUZAwYwnHrBI6vhNaDX91
r1JmuJ+3+7BwXHPPLjaLVrTyDdlCotYuwYNv2a7k1658YmOv3MJdA/OF2aBdnpKK
5lM69f2LgsdA+cyP8rg8cge8AZXDkgQVf6pb+FkSD+g1WJaQfYRnih8OOSYZDF/I
bkWkuaCTVNAQJD98LLIpu8uBlAeXQ2XCaHO5d1NnwZW/9rzBQ7UpkVE2jpIerZaY
TDjMc29pkseT/ztcA9qXOvZEGZV7m8Z3yDDpXEG9Gj4qBavnuA3V1YkaHCkgWIQq
t5XgUuTDSNGkkTj+9AhRPhXhSLF8Ak1RwReWWH+rJianw8KMXCX4DB+H0uJn8wbM
O1QuZo1IbbK3PTDVXJ8T+8wnFAZ+/gBwS0XTLUFnQ1a5GqDQ1UpjUxXE7SaxTnR3
zsUPT1EDDF6kaLiXc8XENES3WyDpUAjSFw6v4rXWTJKfW1xBD6XyFOdgPKcbTCrk
tlZ6jqJc1JjfwXQRRG0GnsE1rMhGdL8Ljzh3OE7f/XDc3oy+5o0LPze6ts1qzSrS
J3FRdlZ9iRhJ8qlY7UYgT44+DP9YozekpNYwKk/buT36WHZPLNLO1lmaA/+kYbXh
0MgpVZNuY0riMzZqU1kDI03W34E9KJ49GOVY+V6MdnOnpzOdrYoZ9Ot8wQedAqrQ
grYIVvjdQD5ZuLx0LBkC/8kRJCq9D0p9apyZxtruT0SRAYY3jPm9Dv8r9NpzMpt4
O2GsfMGlTSweF4uB1QOG/SpMqdMuz1smALUYhCga9nzqKSuX/dfP0Aqf4L3Q/eC1
6nu9MZCWno3yDji4caiySrVnJo6neienmJikwmDnmQXaeHZT5WWtNlvSGpumCAQP
Ala4jD1dV3lT2rtn1Bv03tl/VceJTV5W5MbKN+tjyt5o1hpkGqvKUfEUI2y/E6Yh
Ghu9GqXKV2yxoUipvLwfpReOpqC7PvTlQQdLWc0FzqhsGVlyLyW45CJMw4JUXbBv
Zq4MITqu0rOZUOcQM5iaCLjRPjO1SPmQqdaFZ35K60dhOysVjt4NVEiX3XRNdAh1
ac+taKw1iG+s4WFtXtewipeKMY9XI5rIpjrOT1H4Gd6ap3nSXuJ/Lcm8ySLRTAF9
7jdIa3KQP6qKibdXPoq/PkGPCxxtMhb8IjU5Q8CT/hiR/yW6VarT1JwUSibjcmbu
ZrAQ1GhdxDpuaTudm23vxJBhArvYEJTOJnqyBcb8VIDO7OtCxkgYhqxpQDBRmzYy
I0oKgJMq/nLdZVWbbVFsTSCErSOogzYeNc+1HP6zlzYH2qxU7VXOZZj3h1ZE1/Ka
reZR02Dg8EayQ9XGPOzLrg0tlc4OFR956iwx64nJH/DrJg6TD2UySQivCB5VriEC
3eiyn7cICcLwqBADcsV3mHUVSLOAchMU4pBTc/MWAXAGWRc4gjyrSE8BO12Cy7es
1FRUxHkd0q7uQleuRmzmGHQ0IsiV9bwuLlnX392dW9YTXJb20p9grtRNPt8CY93T
GqJCZNdGng4B/VA3ZwsLNQlLkHUy18WoZHStQCNe4GrV5OQJm54qnw6F8aHd04DE
rMbeDw/nj9NO2XudaM+XAyO9lDjIdEF+hdv4ELYwx50/egMzKWP8xdR0c4BxCXOt
xz8af9J+ohlJQjvW/O8L76z57ws8fSpArgrcezlEFcsedmUpe+x3tlOFIeSnk+a1
Mb19VucySzaN6LF+0zjlYrjqU5I329TAZ+4jlkFtbUkHqLzQh3PQxqlXO9CaUa9q
yq+SmLJGelWQpY+CvmTf5L3bmjC23M+GillSA0mYWc5Vdg37gH680jaiERH9d9D8
dcj5KQdHJUunBWAVi0C4YYUI+70kHL+olMTAK9adk2Z/zz13fMHI+kMK6Z3+I4T2
DP16628yzxNw5FERuQdNF3s+ItubJJjxnMHkYxBx/FOD2dizpxOruNG+V/ZellAE
z32y/fPN/wvH3J6Mykh5+c73YblPlqNV23UUB2wD0/X4CfRAfoRKLGFGjfMQG24r
zjTvd0lpcALRZq88BqI3lsn47lEUwqmSUQ6OoD8Uy5aim4CxUMMcSWXuiWXkRHxO
IqATIISxW62CKQiKe+W9kBmPBthzXhoi8qBCQFzSeqwPbk7y5J/ebEFKsgXEP7zj
9hn7bTtLkPMKkPpBoHc04++FCOJZpboC6LKWIw6XrafbhGd3OpQS7/aaOnKjcWrQ
gZK0kpF1pFq276nlE3EZFUZb6wY1IYsSW9buK2MWHsZ22Qg3x7s0BTYG3GxozRn/
s6SyzHPoDTpHOEgwDFCR+UL7E2B+2IX5ZOqTsNE9V+dzpFI2GXzoI3ExMl5blFnS
dnQFEgdqnLSEdoYO4gA11D1vmZpuwT1O+uZ+VyRSKIVrHy5NEIA5z8hr2Ij8Le1v
6ZSVrAfFTzAvoiCy+bbxMdusKBeqH3NuzSYUnmisFs52Et2oY1NylrTvUoi1qnix
fZBJvUO0k2qznA06LMM+4p/7AMYo8NPlbtP/b9/R66aobAxRMpN44OZHpBBFwUYr
3C7K8aMr5+Fvc0jtjgnSaaeQdK93pg4S2xi1+GkAZFcPoh8qRTKv+1WORp7l2lMC
jYf7PhTdq5Se80CjOHGP8n8ba3rM/qGHRnheCYfvXjHqgxw2JJHKIfmWs1dLbFtj
Cqg3RUG0OImqmXYyt093pMX4HnD+UpxqdApNq7dN5BGjydxZFn8nLMUA1QwuQ0bt
KJ1HvX+VjaownVOas5ySZkNQa0E887cBhAIAbVhY3QbcLHE162+1PZx3EtK/fkCp
f/QblHVwXFRAnuHfyprbG1+ARxi6mYYUtqtqQwti5m+JvqcUOFLUDphj6oTSVpx0
csq1IxIMpb9Lo1wnjiKziJQPxWftY9h7CaEXlJy7LI/EU+FB9ylO4ZPnfXicLZRv
iI8cqC4cBZHXcH4CO44m0DAgwcMxrIeVJ8r7FvqqIVVzY7d5RUFA9tXTqe0N8Z9d
q0eitprS8nPD3HjISKOQ8036il7xr+kRA0iya0qGO5nAba8biqe+fpBUM69Vd6pq
sK+65cAe73xyNGHEAuhic1iZeUazQm9HikabXMEPW+IQ34mqDBWCOJ1y656yOlS2
XdVp49FA1uNW78U4pWR4nuXdjguz8+n34H/Js0CiI2xJ1l0pXOjjZbZUdumWxMuK
Y5TUi+VCTYDQMM1YhveUCMAMs5xY8YrwrO1idCDwushFF6fXUDv7wEQJblUoiz1M
EYquLA6G86vsIEpYiXUfRroFTOr/+G7rvEF/8DPaLRzLpbmC6uHJ5/nHoKCvVlk/
YkN2x2CLetMWDT1LmqyaZq3Lao3VGVW+emQ/vNF6EfZ1pnTbirzk8j3wAcr8ufPq
6KJxK9EwUVPtKb0D0Tw4286JE6ugS8E9O/Pkm47rRXu77oJ8LoIhk2J7cHGFDg2N
FV83mOgJuMTgclHG/Ah+8sah0dAafMKLLdBk6Z6kQI/MKVJqYC5bSSJF9mUcN1+J
VYgR2bil3AMVzuCfPhwLWfAJv2YKh+At1sa9xt0FB7/tCcpGpB5Ph+nl5xsfNvPG
C5KkvavzZcNyP9o8wfOxtoOljr3OoqjVahjJ8S8CRFF30BMOpMt8cv3MtlxIoVcV
fuxxcgcf/I4HqvD3DwnQaWvoLBJ0ponVVhjalVClLD1jyCOQO9pVF9rBkDOrDGvy
1TZT1Q+codHdD89GzEi8q2wBiSUSXfQOBCXpUJgMZZQCh+UK+KcW3FCdfqX+vbQh
x+a6dHv6dIOQdUglgQL2POd6ZaZ9IzSlQeuBfOMZzUS7XS6kFmfWzLOzgHRlZ0jJ
TTla2UMPFWf7Y1WBMF64QXyvkQ68GA6C6VOptsX9AWEkEX5MCXBZBfovgNHbAgCV
PdgEmEdnbbh4KhDQOmEu0wDb7vhTHp+fwYdUny/Z5UZ/las1QVXfOC9rL4J1SfO2
B99wcbv+q5uKi2TC2ocUqiNHpO+vPu16iUGJ59Z0JMxy7w/Loo1fQgXG58uIzcqK
1y/ymRY17dqrzZsVRt5R8HxkiSD+1UAYq1fUeptMw0Vp19HeTIACytAhoPe8g6I5
a6xBCzxpX8lRS4TkCHIxb0AqFQD3skjla8AMR88XFhvbFrJcUpEw3lMFIpbUPHQz
ixd5z2u0+tWvYBjsxDUakrtaaTvMT8K+u2tsyzWeyyb1te3JX40iYc4PKpngiHXZ
zAzP98Aa25QTbvzrikw36VuFMoRcUzAmlhQVNXDWzHnWnMELUwIzv+V0D6jDx9KC
DbkPXtHP2BlfFgLSJpNYw5jVXzvMuq8nIktqlwHW3RdMOTIGZ1cYTcd/HdCm5vvy
LR30kVZVBKIcFYgkhtsHIy6vaE4ve6mw/E/dM3DDJJOFtuYu0GUQEdpQG5ajmsOJ
m2FDu/IHLHjgJV6d4Fogou01rOwsizSFxcwDStKNxZls1Q8Qb83qjxY4dQJJq9KQ
nwOeSLPM54c0Ryb2dfk10YnZ+Vj9WeIbWlHFb+5hAezr1Uaagi3Y53iM6yOCrOfN
Y+eEvrugkDvPyaeBajc0xpyhPlb5VG+PAU9c54Y7vmjIMZwz+MLU/yjHx+x13ukn
qDJwVtkpgPEuHZxgXA/NVrgK9vxIYjUJiwjeZOH030uIerR7Cwdo3xwxQKl++S0x
DhLQfYSqzGpqh7+jyauy9V0BVjmZmm9IeP/mc3kMLWT6KBFu+cr+cCFJFMop8H6r
lc5jyNdpffIcoq5umiGrqXFb97TQAZLXxMeX/rFL1/k8k+3Yq3/QKbrIVo9J3kTd
oTmUsefr3VytIHweZGzo1y9RkeYpIgKWe5IM6Nl16mPKsIWLLUAZU2wnKnDzVgLG
CTMzvcICrVGBw4hK7ZcqZmObXjDYF2XzRViLKm+3hH33E4XQLMpkgPHEu4sfKiSw
jUhbyIpcBMrvYq3M7YE7DPSN+7sHOPyC/SAXwTkqLfFgZHYBflFIzn/7opjfzuyb
LSIMk5iwxvSBaEDCEdMdc+0WRHdMv9V3qJ/1O70NCJroBQ4PlNiW7/CFR3Mqky2g
IfPtzZXCr05ds3kecr56SaauQ18LCJG153Dh3uKvbSq3UKj/1VQktn2fwmzBPQfO
cyXoQiL7dJPXUnDMUz94q2BoCylMiIHTNAHqiaS/l9cj7KdhxKcFOv940bvyh2bg
5dgSHj6OOQAZH05cd5wuAmvYZezk4h6dmEgjl6lAvfv1AuywXKx0v0HLt6qqroPj
+GHga18+LkYsw1ESv3YNzpqkPCP5SIlBv/tGNUpgJvXWNx0i2hYf+NX1irCmpZt5
ZXui3CIZ8iSs4Hr0XWFr/XoreJkSv9fHfPazfiiwRII0o9r0Nr1mqj4Wvzl8qlVr
eKp+7oZ3OkQcwevKjXcElEQ9075azPC48WmaovwXe8ONIxGldXJqmsIUi8oXYjzq
Q+kOrtByRoxphQfdJEUWD3SDTn1r5FRop53jeQW9aEiTl40Vl2wtHRiuzq3zQ1FL
DigN1wWEgXKSKvPvLqZYrlBSvQminndB1CmffXGgw3vnHqrnEqDrMgkaUPFxU/A0
fY429DpNaHs9cWq6im30ldQ7dekwff8Pr2dbs5cUOYYjXtHkX7StCnnO3+w5TlZ8
sTdY0l+t4PQkc3zg3dDrTDa/Kpem1rOJQbHloQuluNzHqq7ZlZzhzOVTzzSztAwc
rTxfY7C2HZhnhKpYl5r2Ue3KfJ3CBT2CC163MblO6V/A0/3w4OWcO311Xdi2M6Cr
ts2sbPjq8gFAxodFNMTBL307+isOM7gE+b1fyhfMrJOb0Fd0rIbaPdxeHBnoInum
s68KgSE0SUomp0zseeCokwkmYrZwSUh2gGARNA8cT1K8ae65yxfumNDyvkubDdsx
yuEzfhR2uxTGOPtDUxQnyZZSq0YhUbDLz0AN5IzjjOueOulrw+MVoVH2lyMdpX5p
QG3DL43QWio7pL8MylqYFwEk3VCUTudJZfUrlxO3Wukl09p39wH/V+3GwmfRomCi
lmTWEc2RkGjMRqHiUZNtmDwN6QVih2nbaQdAnisdYXQhBfGTP4NUCS2PmoEqvLag
3XAPxmT6EGjTMrmLVu4tvLmMJ/DwR4zhFO4v+Y3PCQPxh+9Hp2Uq13q/DRDpFBEp
57JwfURVlYJ5d5Wvb5duccUVmpy4JsfotkUjFd2WV8TIwppJdNWD0UqiMpSgIvIH
SQvDUc8QjXqMa/JQqMDuT5iFXB5IH0iCISDR47RO3t9W1Av/cjSEVblEP1jAKeO0
WTscXAqjWW8NV33AHf7R+FGldP/a3YsBgfct3HwJzfVavtDmgZJVytvnpTNVeG6Y
cPuv+ubQ5Tnbg26hTgeBSwHr3Nn0MZ+c8uizQIOjrRRG1jviHcLIUUQY8E/fbEkU
wQCJ4I+gTos4FOD4UvxJUH1yrl6zrLUVKJtKz9iM0fWMKhwkz7Jz8Iqz2DJONMey
JIweRQkxqbId1qeYWoYLkUeDroiVSC/ZUdFvgkgYhlDdkSyfmsrrjxG9u0D3Vwcl
4Q4nM2pYlqhaEsvsr3iyldgr7nxqODpY4OrW8qa5zt87oqP9KXtOAJ8mwkujlHT/
35PzoKzMRDH7Zuxz/vGiXnHDlxIt2qDS81FHc144GM5xcRtOuUmfgQPJnnlmJo2N
toBqllOT/MvA0ZKfwyPzuxNcjaeGeU18k/EMtf3wHT2yJR3EvG+iDU8iXl+gHYoD
zbg4/KlLuvOnbgy/dQWluaQJh+qeDgSJ5eLdI22XgbzIRwKmRrTrV7FyFSAbg7D9
QW+NE/IV/cukMpSKNwP9LvofqzJ91oTbmmruYwJrkBezD/Cy0lseMvb5RLWL/x35
Zb/ys5r/nC/tq0HvKAoU1nOS7hOT7/pCn4u+j34C1nK7SI1FXsXa0Jsg2FULpfYp
BTrtD74yKOqth69ndt1LPqV/UkmE8piYqlDAmO30k8+bcEWrzpGNBuP7WiZtNtqU
nm+dT///kiDvRuvkyFU/fC3Y5PH4BmgZzzNVgqUmx77OSN69CYaKCK4g6MqGoZRp
kEvN40+bqo9iCY5md4vS/A+Z+/X4xN0/XmYUEItMcpvSsYoIJZr+4Vjhjg6MVRrR
vS4pwpk3dZ0+J7hGRkD9t28eppazueC8raR4dfuDMcbVbw5PXAGOBxmZFt8ZRDdb
lriXR4u0yHnMBDCZ2qeOkTKVDMusA1LpdDko7eWlPEMthedw2M/YY39Oiheid7cX
AiSw5WG8t1A4wYsmQ0HimeyIKlFVg0dDgTFPjZt11MliSlP1/lkCWzT4ETbOJIr6
HSQALS0Vlpi+C4Mccdl5vbGNaxSzhxvGYIjK8efIh3Vcyt4rkmryXjFj9soT632y
Z2BwHRzwVt7PVvDO8bTSiBjlbOJ7JiYBwkaxRQLASdCN6eoWabFOQlTufH5RTPkw
55tqaUCu1Mds3Drrm+82w6AV0kXukjzl0C+mvuPI0jHB9aatPHo0qdxzCh7IoLjg
3rQnn8njWCc/zmSpxx6YhOi4FKdr0j5PPXNOdEWVzAKps6VQLAYfgT10Q45VHbHv
xQlxbC22h0b07YUADv50AKRpxtnErpSvrIMebEeTcxHfcj2pDiOBbYHI2v8cU9OL
QFz9ycRLj1k8zDQCQ+0vBhrRtgmVb3pNvqzHqiTIuWeWxoBJITNxMI5gooigurVF
Hd5efrejpQV+knAo5aN648AAmwCJA57AYZesQLkX17IYncvnqYBmrlwi2LVVA4oO
bN/5cMms8pS7U/iA0PMMnI71LTa/Y1jGnew6obtXHlbAemcjJ71ILs026NqGDB1b
IruUTie5tTQYW4RFXR/cEkeIcDf+XJaXjGsgR/o7rshv4FDCNtDk8LP98oBPsUPy
4xnM7qCvCWhconIJSUH8CXfZmrdTXElbnC00gTREAxI0UfgQaNW7l7JfCTjHhh5w
+HCrG9IuIgGA65j7l7awbBlO8zsjvPGPDuU6VbTLF9J/Q0YEo6cVj4mcTJIdp0SN
ueDx0WAaKcdIOGuSpR9Cynlut9YLvWgIHvkqOGVhPoksAATxpRz4ux/Mv5hVlPds
Qo+Fq9ZI+FIZMR4dYjtFAmfEPerEASAtEIzu5e1sgdbqgoZfNAgsKrrnT+75X8wF
SaNh5dmQzQBniTjg5wHUR3Y0O+nexXyuMdJzeslR9bCJQL9nqM93/dCKbUruFkxw
B+vBSCsTex6GIaEMCy4j1ft5+vVh2Afu02RwXPTUoykcvP2CXngsHfysJC99Z5rV
QesoiLYMV6P8jUWU67kJw0msyP9QHFuifFzryRO+UgcopdC4LgsgU/gECDwo7IRW
U8u+aBxASDPIwMzNqbo2//x+IZDOSivn0YgwrfN/z3XoX2C9Bt4v6mUUKYTTNehR
uwzJr4Q89ywYjxRViAKXNnZkqCMq7ULzr2Wxar2I6Z+zNmi8a3+arAfgeUvkMlyo
L4Rz7nkb9ovfSzHdh3kpXu0zwuW5MjTl+ZfQedNXVjB/v1LtlUj5Lg7wtgz/grcM
05I02MWlpfvwcIHCi3ECuDCmsr+qAc663AYYsGJbyxjZTGjz2HMnfMFzGhH1Dw4g
EEid+x9idRUODetM+xzkUOryu8qJsUC/qQGCNy7qFH/vSTkqcJjfW8A9aU7O07a7
hBGKYf9pRdFwsiy8jVgD0ygr/4xZNfrXkah9u0y1yOXe8hPJUtxCxiS/ZkRIlYfO
pie9luxttN1NDd9Pj1A1nqr8N8phcehy/saguxfEHeWr6v6djWaeaU5yNZADrhun
KVp4o4WYoNi+RfkEu3VhqLPnoSS5xSu7XZiy74LQJg9A7xNT7oO4WdoLZNbPpuBd
ZhUIMX7Fe/guKmZrR1iQ3tYyS7VePoRz2KZM6O09UbM3eHGxpMSmJcThY5KLLhoG
49FPSWUQN5429WXeTp6IrSIln/pfrtmBRVW+bfOfoDVnoHT4zdmsuQKZan2wSi7C
kl+6190z5UIDbHUQx9jJUvFWgrAvjhKFoiFAJiQ7yVD5DhLErfFk8G+Vzl6zevC/
3n8JU8OkOQ0JSDtjhlF0UB6kjImylor4IE5uXiywijtSD0uwPQS0e5OaLt5xJdHp
J30pVFoQbd/wctWCU7AfRt2M7WDNIB+/gWvPgj7gtgnAE6rqJtlw2qi9Cn7ES7R1
0+mM+5jH/GMpxYNOJ9ez429l0CoPKtGHjuYT4hYtzweb804PmZxUq4Ci/4371Gz9
2aVAZOpTCJ2iRDP3Cps/DJjMNkZm1KLVfLGYIU54m/uAo7hXU3AtBkcTftGQ1PTl
VMmZAFDgqog0LO/zhhB7u+uO5U/Pk0AeIfeZKr5STY9INg+5CmWWz56zv7NRQSpA
KZhCVghyeIr5zxWgRC0pdVbG4YklQuTTEu2ongtjDbQueU9xSmrVJfDuAz4fIwHi
Miv3hgQPqlhjeI1/2UXbU6fEi3DQ7xeiUClUqvCzWdUY/jJ3rfSpKTaAUP55QH4M
ZJnefgK0klVQKPV15JfH41DnmPqx1xoTs+lNvc3CgiLaBKgZ2mTlbhkPxYfkdUgj
EOBpjxkqxovJX/lNbtuSk7O02q1YusGMhN8fsWgtVwpbSYyUGw1idTIXBHTCYVxo
UyNeBatAqbOcVH7DmdxiUckOtrLG69J/y8u/NU+eSiuqSe+FdLvF5vV4W4hAjfzk
N4hsYK9ST8JyWLUNTcpvOFBcVsJZCHLPNtigpKTmmirgu0ijhP4KeRQYonMaDTv/
umhNJXW61luBoSk8s+SxN+NU2u5GER8tiAJKpd5orn9E4oM7u70Nqi/V527ueblx
VLimT8m/by/lAcsV9b5U8MabKgZ+swR+tIwVAeGrdG7aGbGG86tQMCZO2S8I214u
rY02zaGouJqrZNpG/9O6oc/ea+9xkx0QgDgnK5zdF9HWMhiTkLYb13MUNyXqLE11
U6z1p2hOcAMtPvC9KA8LKW/TS3AToUHZVnWOiYQI5L0+qBoMe0Qn7LQzsFlJyOPT
9Fl907+jCEty1hoYgHxaud7pExOw502msJK8ZP0+UR1p9hCVmsszKfQucdvutAIu
b0sOID8TOPHZMMV1Pu7Za6EY7ncJDhGOZXYdfYZKribYfwfggNME4WAwfjxJ6tYs
NlVlOMRU8h1GG0f4DNXXPlrjhlggnGucKB8iwQp4o8ZQ83Im3RerYlr2UPy413+r
RABoDFdzFzH24Y2DVLgyxZoV4BfpJ5hAxSdHom3MrLQRYQ2AElZcuBubw7K13NYk
bUNjPbckwO+OTMuZbV78HSYvbtcTkrCbGCDMgffNbm2Qgwojqtbs8DAORln8weje
hSo5uNnTCHRgDy+3/pR6BhFvgAOb/ejF4HGVrIk0UXG/ftA4IcF8QcuDM9ClQ9lr
95OKxbAUvhN8iBl5SexrjQV/ulrl43+7CslR9e2CJAJYMTL0vYt34TN4dxgSYXur
Ymv8eNuyHDcS3Iiqru6QCzqJGE9XG4/FCDr4exLs+hk9wiBLwyHCvpnvrZ8c1Ipz
49SeoatfBp299d4rLhU1BvcmKsopLiIaT5+9kvjKR4a6J4g6fCqTitZV7SmQgNkQ
widrTZn+xAs7hV9zGZQLxanL7lBN1z5ps1C28GFWN+WnMzCbs83HcJ4mPDAThAc9
W30cOBZngrwYTkIDB/uDHr9Fkb+0IXUnbSUrLf0mgi47DpIIWYPWNSP+Q5jbBrcH
Vxre+bw+jjv3x4A8khRFcLjaaTUlVJURqYepsOVrg6LXFeCMoCitmeqOpgVwDOEX
Xqp4PbGRE4Ajp1pKRGMYprPD1mVY4aEQ5GHf6bZ3qSU+09+zGFXYbdW1Fp2qgid/
gvmMo0I4l9dzbieFKx9MTej57M+jTTpuf61Uij+rRHnWcJUtGvZy8TOyDVpZzz4+
PF2/b9hShJ8pJh8MD9DS0Pxa1eYdYfgLLKYrYMCldIwOc0cl7uruGuOivj8DS1oQ
XJ8OObNMroQLeG1n82HCkrwoxak9LyK61J8cBS2UF7yoDz26+NYOhmvF+nI6IuZd
Ygq60R0UM+e/DAeNKBfu8SefRrB72ZuAAPot1QLBE4N7tktcFBXY3IHMSl+GlF6d
T5OESv2pzOV2qV+zD/2qOJlDypRDEhup8Pn7Rcrojl2bOflaMRMbY0wiogHT1via
/LulOaCsc5q2CfUGD7K34v0z5c1Q9d/xrBoV+G9Ts17HrvF7Dbtl3PhJFQttASDJ
gSSbnjPZzppkguUgJ6Vp4Xhlv+hdECKdvsL2RiRPybe1CNq66pTiKXagJOcDPtQa
zfgco2aLc2QCZasAKgx9k54hD6GECiIvZpt4CiOEhL01uUjlUzMr4uyk7h/5uceg
LUeNmRIYUXxE9A5aeHhZtJV1MVVjBT9a1LMqh/TCrYfWWizmBFVmzKY/1tyOLuzd
uWCZtAHfvgL5JZ4oEZgSpSIB50w0cTmNdIQx2n85YQA0d66uuQWVuENwAlxCZdUh
BHZsAMt60sVXLmnqYxAbIEG/tHc35kdcgIubJjrpAKzu3aQRIvhjkLuZh95y5zjb
0b7MEMZ04B8c20XZvDES/zMFYF2JMj01r8TNlHsSdgLvGJwHRXuGJJuPYeA7Vb64
hWy7fz1GUfWvy00O36jQKIeh288eiOUnu5omH6mgiCVIe2uQ3h9gjB/5mFcR/jfY
Dyp7Amfu9W5Ud75/J310VP378hwUe9tOcbEWF2667TPRhkLWjnX6pcLzgbHBxzeW
m2uzPzCMk+3z/tF+ksVwTgOd7zJOhptS73m0BlVaHjlj2tV2FAHAqAgjODgMzZH2
7gMyKEgEZGlLWmPqCYRVOThNYQ2Wt0NGTqucSxL95cf9bJrJvmrUhQm0S2rKD0rJ
vZdgV/atO+ou/hCwyE63pqwEXcPmbHpSwrwS3USzPLo0wZTSb7pWTLSBoHrEbRvZ
/qEYoglZhUEY7mWP8znTAsiU0ts5+lfM75lX0AbF/jJKTTeUOPA4JlQTnfQPgWAx
mIHtWmrtcyhQK8+CYOs/oL3w0cuzipylKAlsFqjca+bIBPIb5lu2a1y+KUFruOjN
8zyJTYWsCTGhOsJBAiO5aRWbgosZnciIbPBrRBqVotRH4lavIGgoYYQ51q/aL5M4
F3mUDWi4bS7xJYylH/8p0hr2+hACrA3nzlHktxhO6jLqh8nU7agxS42XmxNBqo/p
t8xVUpInDZvGTHFlfn7IBJWTtK9wEPo4XgCWXdiyBTlsrbPtEMD8MpHt1kxNN/5z
0kZ3K+XLIyQ3tp2i1wSW+rKZsXE3MkoLK3S0nWyVwNO3JrFykMu9WhszhvR19uIy
0CzcoDWKF1l/kqWeelDKxeT14y1dLODfQQjSL5uRvgaWPZesb45jAaW8+Bni/NaQ
DRLAnnF2C14zvWSOtOZtyKNLwIXCanRRVmkjMacqYHanDMtyqWPmooHNH1Ulxgsj
kOPMsGwh38SdnJ6WJLTuFwffuXMoscvOYT6xLkkKRFRwrHn9Ut2+Wu46oXU/TGov
YDz9tiav7QkNQUIWg5q881g1fdHT/2LkT0csJjN/5X9b/vPoSewJuVu5lH43HKND
BMKaDcFVTBCGShRyFXd6maqc6j6aUH6GnvzFHhouhCXqnyg7Zl6YSenH0Tkj/DaB
BPh5PRvbpKB+6+jn0+Evk6o5Rb/jVPMkS2A7CIYBnzOGkImoAXBw4o/1uLnD1JS5
GYLhg6GA83YlnQwgeAi0sZHXlkwdcnuNyo1S4l1LyU9pwCM342r/A/CqByCVBA56
wmPZVtD3WhvrySa/Fhj7Cub8MIFubtcwAHTy+Pjh2XuaIrUElBiQ8cui2xdaMTbn
aDq3GHhO7bRXVbFbdXQyJ3lsHpu+zBmOkUfmb5uFbFP885/Hk35viRk/0WrATYdM
Q5V76p67LFtxo0YOGPROpTupQds3cjKtPGYfJiqfYvZfQHftld/vT3XQR7o3wCqU
FP4vimDzRpL+ueYRhHmjD8/uGt8LSJLl58h6HIsZauzSCk5nVWvdKpoL1tH/gM1H
Uofpdgj6vaFXc8dIOHDaWPxHC+IpC9qXe4gHV1E4xwhh1ORSfJFH4HiazRpP98oP
QtE+RgW8d03eEbuaIw8XdznQIzi6jlaSJlyq1XiEPOsVsBccylYGiPSBNpNeJere
Rrf9smfdHsLE20+KbKihKVVdiB3CoJLuVEqVbmkYDyUdCcN7/7w6n0N4dscuAtAX
S7hvOImC1rRVJrlWVBBbxfh9RvGqhoPbQV8RjSfoKv7DfUNNpv9/pwodeicufdUK
mx4+DwSJqNJk9QdJ0hDmtHNj/SUdD3I3+D+i2q86QjApHi/6DadBlktZ8g9Ke7XI
XiOK2uuaIGkeSo9aYjZVJ4WWPm5eaIbg2IKUoHoaGQxWG/uM2V20FZQDMv+XMfX7
7Q6rMhUn5NK6JIAo3ARQ8oLbDUoEvcPBWGvyqCzjdmGDUMmvhNs8o/4f7bZyJEN5
6B47ZW0n7/U9TvYpN1GXVXvN6rnpGK8scIJKtq/eZNlD9ASJ+hhYNj6EWfBDpa4u
XXGdNj7y03RPGfg9KmvIc6yrzGxtH6d81VLgb9W61J+2t5eHwHKT4Q0M35bM/9yx
mZnwoskehbip9BLeZ0GAkLfX0tL8wWXLXx/b2Wq7oNcGYsVn9/swLXKTfhmm9PI3
3CXh8ohjTjxevHXuxLqQVXzGJEA+IBobtJ/rFAsKnJUwJkWdamV5LQfXs309M3fd
jrlKO5RGHBD8rrYGeXWSSE9kSJcrwzGK4fWWbJmvi4zvsyRBMluEXb+ZYpw4XhiS
boIk3+DFkZkB+4zdcS6aH7dPTFuR6/xFZ9SLtGImL6yUre0f5y3CKm6GNJJiZkI5
uAnRF+7LRZ6zWhaSz6+td3Y6cDBYwbqULHy8l65cTg07uEP9/R8hOWTZkzssGrU4
7UXej5vcO0EPGwxEulIDo2DlU6y5SC19D7hV3p1O5z1cBzFgeQNc5Qi/5TNHxu4k
3su7PH+MHOZ8rc9KejQMWTO+XFbjEFXjruA6738GqcLLZOkXkcmPS9mFbjXKiyoW
m7+Yss+IEw1IhNpKqkCcKtavkh7tJwaiMMsGd/lb7zKb3SdP4eNgHtRCmuSVFeJX
2le8NMsLWk2qWXqfnDdybuBUyubJd2GqDhYELh11lFEjW4qclntELAbuVKTyGldi
DoqEcoGcVGe3F2fEOJjK4bHm0TxBMJXl8q8JpeBvBnNDjrMfdXz8GlmYzc2P2SVL
YVVA4wQODLkPFKnqVF26Ey65al1N2Sn12rL0396dC12YI1nplf3Unf7M79JEWD5H
DXD3a8k+aZuGO/+z7E++bbq9ZxTpgnGrE6VK6Wy/6Srn9C1/siu4VtGMxUfvl4gg
MVHdFibbPxWOc25aOJX0XTBLUE0985fUMV77PYy3jpoBfFGT9Il5cNfIDoSxP7pf
FEcWP9R3qtW7N0hQad8iYRJGCv7ureQaDkB6s7yyygxiS2G56FXaPFi+8izxelLX
Y7dYMdj6bNNRdKSTTsQPtqf1f5On/b+tJNkb6t65Gd+h/2Vz7Kza6IQHO4sZhJNS
O5rdkzNf/7530b70gtf0R1SSXqvPSxXEacTaLYKXcQk5r6Y05ufKTbTvo1/ui0Im
bHGm/zOhVoN77SpEHcHaZk3EHf1EP2EkaD4dLg1GfaVwOqwqKmnYULFDNhLHGPWm
LzcshHXK0cCdsD7DidWC2vpVviNwDTofvCYjeafAEg0Q/eYufz3m5GoQd1lrFvUk
7S4dFISwUX5h7t+xf+jbfWr95cMrJbV9y/NR2/Z0M72nYEDGu0BLvo1nII3Kmt1i
aLoeiqQ7Q/j6Dz6XueuGN7prMXiiqEs/P5plWAegLWMlKt4QLbEvAJhW3+EcGHWK
Qnl8w9uTBiMG73+ARum04KVMt9pkMU8roKI6UisbhCm9XLtgZV7MhDm7I4FdTdOr
rYXfstLSTZSCqEudHKletMmcJxkABeVw+DQeO4WbHN3B5jat3oUi2AmBPiviOm9j
GhxeyPQ7pq94hfhUjR/W9QdvLUx2Hx3zC38zL1yLOYqWq2S7cOdqDOLzYgtTYM4d
YgFgOoiE8rz57e3p/vDn3obfi6/mHBm8ADGDjmCsvHdE9brPJKY83Mq3Nbg5Zms+
309sWImkapUvAFavf88CTOhJnQCyouSbvoNxAHiG5nLB4JdnWMeJw3dlsM152GNR
4eQQwZM/nPLd1adluLLRgNhXZZdnLnmCXaBSwvy67tQHhVjGFukTi4+vcp59yXDt
8iBNl44Ito6KLfjf1MEPAYkeVCxjDe5x4g6msOouW8UsjbN5UVA2DazgQlKJRztM
g8sjEsuH0ChLbatNuqw680+qbCfNnvvwWyj8HYlGY4hlCofLBHb8wAZRitkfIQcD
gOYJhAKcB5M2FUci+0Fm82JPlmEYGy8y4XPiahRHtSwnhqoP+OjMZkNKy1Z6pqKQ
PngWfD7RHRM8kxbl1ehhEoDbO/PAUdr9zkHqoS1OPuLj/UVFGSCbsHxtDTAexerU
YC2ONKC9xOhNc5KOWYzsksquBHvFF/ywv6D6AOUH04C5mtXK1hQB3I0mD1a5OvIm
jj0XkJ7dPnuyJT5XwGuboJSnB9lG/Wbwm/dUt96YLxCSInuiwoDlzdQV3HMNK51K
AEljJpg5XFPuApZfoH2rem706WEnGamtFI1JfEro5sYnHbltblDpE95eM90+oENu
CiBpTVu019OT8L6oz4lCgDTRbyqqB99/Jea+CNW5N2ySvP/P8FCQ9L+OKyxUVFdU
6lfzjVk1seWROokgsXwRdsKtBcFuhluYEoZuFyfWoNcsGjEL5vb/D+cAX2+1sLKm
yssjD8UG/3DedWWZiszj2BlnjmNccsuRmY7QL+BQw/8ihQ/o7sYpJ8ykl8JXQsd4
txhAQegAxaCNE1XdVkUHjyA43TBe/kRodq+FFbh3u5HJAhn/wXh5IuCzTyE1+luk
4GPznNkX7biqDFexPWBdrdqIFmiIA3eSy2TGbZ9mFvfhVy7+1qbLetJgxxkbgfBB
vy1Ixf5ZNIJifz/nbzDv4hNWnp16ZR0RHgB5n1v60yqyYVZS5uSGqCk6aeK6lnHQ
fyzeNrKL7R/z2UGQjNHdXGRrTREGuOgJb4GIOr9imhzz6v1NYHXrBcJ7FraZJL6K
znm2Mp1y/eNq4VOgu/YaxL10q46ePVY46buZ/wu7vIITcreD4ECXs2dpWALvmsIB
cAtnFeZIRIxz8EZ1YvNlRgClABSTDzHVJbGOvkjhlqhI9MwE7+tyf29ziqd+wuv7
TL2oLSVykbphoMkqcfjxsVS6yztbiyJ5tF8piR2UshUrYZ+FV0v80SI3BpzGXqL0
zBNWYte+cpZWFwkCAspjvCfzBV9WF1eLHbgGxDOs/V3S7i+aplkO88+B0VgONKhk
uwaAiovYRf8Aoq6fC5sSa3G0TBJeTF+qrQAOvWcSARKkX9DHg5WlUXwdMiqyr61t
HgmEQNr6+gOtw/M4+KBrX6Bix6u/dOX9e9RBCyObic79L5nsIVsfjP1+w4cjrZAZ
kN1q+icaH9zYr113ExuDmQignaM0sx4KaSCQdLM3IFX/Wz229JkGzTwaTb8pXFLm
fIq9Dk/oeci/b9DhR7TV84xeYH6ZuYOs0uSykpAi0qr42qxJPrM1tGm0UbJBtsRT
mqQEHrfYOwaK2biL7bIsseOebt1HdxFL1KNWCseeok4rFu3dtrjlCWAyp/lUhnQs
3vu2Ypn5ocDkL1KcnqO1dAsTjSt3OIIHss0vy0Eb06sQpUn238yBHcSuh6lp3DN8
cRBxLKOq5nZKktSU7ZFLmItES02jF2jUm2l2TOaqyVAzF5o0t0A4nFtRvOXQbqYL
riJC2t5Lw/FdoHD/fR3BE3nSGEAuKrrKMbQUK3PYOdUh7lwlRalK2GhggGl19mEq
yvHgSf+3FrQLMY4yAu8SK6TQ75oJdbLDIySnug2CRMFL0x/RHqhIDeQUAA9NPkn3
aWWbASJa8IWdQKNjoBbvQZ8Q5gpNjLO7EcOOpVYm/X4MuDaiWMQHNgbmvm8XU6sG
qyTi3lHCxR0N0PWf1X9WFQcpwqnh1G++ne08otiqW2O9VyyPqAKKpTkiIa9J8JJ1
cQuPKUZI7q8DR4vpEOQTXhW6rqsIz+7JQlIKbDlbgbhTitd9/mf8cpC4l15VJRMx
vPRJJJa1tX84dGPx4C5L2wW4X9wmXp+fO7MlIoyrcMBenVqN8aLvRMUXJsaVa9O4
YiiipG8lN8kh/+SfoPKBJsQ6Ju5q8X9nJwyCDZAcBxFWmMVB3O54PuRbfhAYtc8Z
xksQiOothIwm8R5z6LmdyXqUYtGhGrfPKh1VB+B9B/cnaT9e0qxoJyyo4ItZ9NOx
nPF64ses8XW9H/9j2KL+exvahg1PcuuwExg6L3fD+CWjTW8YTaRruZfA3qaaAYIq
yov5MEKPFAdzf0lRu6KIi9x1j52x+Ccp6sKvsCVSL9CJaeS8EAsdIR/8s8ji3TtS
ERWxZ6T+pDqUTwCjTLjeKk2jKMeQOr9HPDPU8IpeV+iWYynRnHqpgxOiBhs9Tfxz
73DyxQeD8nW+0DI7uo+ZgbLS82pYJHeCZZPShY6PkXnpWwuF+wyYOFPlLV3a9Fdw
ljKHxBl1nzAb+nyjM609bvAEucWkQlI1t5q7Ry4S3Nn9q3Sqd3sRFUBYViO97gLo
s4CKgeldjhbpoVb1t6rxexflvxQAG7dkiBoEH6CdYx3mqa1WPG4Ze6AfwP7QYdbR
jxJHwOKkyWBvAfXIAgJx1G4fiVddY7F/I5lxHz9jO6T8mnJVzf/9vLCNzNvUs/bR
IQ9oc4OP8FKMMwTL9frSpC+HD32tXqTHjGoa6CQILfO8teAtKsFh0Zn0a1WWgK1e
w/V/KKikTwMhg0Jc11k3y+ddtGqcHJM7L5zZPPpwLDKyEa6xF9vHxSxFrQsZhDbJ
FO8CPEf/86vQv5cf0zDATZMi8tGiLnRKdXu1Vrsa4YDIOdwAESvHc9ExMJJyouLg
q87I+GWlK4doUyPzwphrLtKEAm6PlSc4Btod0cj9hsjwC7Kb/HVTapPLJeU7dJDI
UEcL1KWHAqjcxA0Mv7mdcbGd0XuC0v1V8k8e0OjBUKA98hLuPYoNRM3lIKB3/biY
OoXAOzOFgV/xPaqWYsdwam19niheC43XJSril8+St+VqIiD5KYwvuKHOjnablc/O
S7TEhU9BWOSH9CXAVP6KA+jeiB+Tqmb4JNqj0vNPaFWEhiqmn2Y8ZgJUkGaZpXSo
dX5cnpZUSEro+TVWm8l082NFiszsx/IVdD0Crb3kXwQeEYlfYVDE8ybcumXcQU9x
4Ug1p9RImwRz3e7g+6wVkuSfyL4goyzsxKp44phJb3njVZrbOYydtalmp1p3asoF
1CqSdR1Z7uqUrsFvmkoym8nUBmEIVB5G2DbsOgIguStEcUa5lXonvJApXHg4Rp6N
szL2FlD2cRofUI1U/K999iAxsgVhbIiSewz4mczuBfUqpWRL5jFLs9Q+2cLN40SQ
oIZ7TEp1wp/PyGW53rNQ/LBld5xYTB/Ii6E4OK9GvI3afygPiDyCT15WP/ihTwYu
EY3OI6APuwXws33Nq8WQ4pzPLIJyx3c1S1iqxk+Mw/yf6XWhtJ2uJCfPnlDiFLcx
DtqbyUgBQOuL9yDKcJEoPUHdCPj1sUpWxRXqLpZwObyPAji8840dYhI35gx6884S
L2eiHh42hHj8fGUQG78YlooorbbJY/ecMJproOM+xMPrmdJhbvL/uZenUMDVyLV/
RZuxRtymMd4kOB9wdhKBb+qxu89zRvuonAGTJ6rQYHjUcfbDxLqiFGW5uczu1u2Q
o7+YkWxSgTJkhn8MyDkBqwCs1U18qA0v7BlbRLObrb6UlgWg4duoD8hhBFWL6i+K
SRzphxuQGlcP0DtG5Z6Y3jwd9fCLW3xS8VB8cwQctUaEyAuYADuaA1Ckoyi0gPjY
YF8H+qFsuiS9rA3yV2d0/A1PK3l4YhcBemdFA97hD3FWw92JpiBLMdKt673tVU1U
eiGWnukpFsIbkS7nUa8lyGSbCgnfltNvOgkB4MLRML7UZgulQjaXGUpvn+UpdnEK
GoJxWFBcOHVafU9CBk3nD4jagR7N2fO+8DFDpU26e8B45s80hBTM+0Jgd6nUlfml
5Iv2L77xiHSE809hwjEgCRFHv9yGgcpLPC5pH4S6PeonzbeWWFx/VvC/ImpOdwKn
MzCr013jMe3UWLxk3IbP0yUYBL34qyJLvqve0ZjCPv6Bsoi6jPLaz/+Nk3Gx56nP
YehxfLh+XwP++rzn8On050C+yWQ2GYbXvh92H50zDjqPNrQdYcnmjlbCit7HE5dH
cBoCShlt5F1Z9ZA1OFBzhaRbqOnaFh7CxavhG7Snm+IEtD8xQsF0UhVnM2CYHFdQ
eYyRLCMiAAH3LzONM3utRXNft7D9g3i+AAdtQS/DECYE2wcFbdtzdNYTWuBPdMxy
wuYu6emM62TDVq88hGQNsUsS4C6gB8LR8b/5wNKpwKvZmZs039u8OLOAoqe1t3xE
30RvqvSeIMG/CMy/7d4krrWSDTgKd4Kbgbvcm0bSEXdWTbi3OT+UZv14Dugbxc1g
CN0E1DpikMYYXjIJGfxmoM8kv6L8vQR0duX7c1kkH+G5dtNLnhE8lWdxetjxJp3o
RAgtydECAMMgGyZjnBdv02FPJ+62XRF9LSvCeBQ+F1akBdlFk7j2YUn8mjMO9PZJ
gD0K7Zycywxat1iEwGRYZaMdHKGfrYE2Dpai+blT4feZnQrwM7gvuXAGF80C3hOj
P8CxurMqPH+x8easGwzFb0LtpVeR/hZBTDPm69c5Bd08uK0bBy3etKWEGNFNK9CH
kjWer7duJFg08OBQEZgXmKlgCs6Oi6e1iZzITIjk5P4fzCQRTlZrCxbshyYyjlK9
qDy3nIKM09KJEBUWIstq4G1uTK5GiuszFCSf1qo/FleOQ0YNzQ9O97LBhAZuitBE
9r/MWXjMISlSFlNK3xGfC9wylORFyAr9E5/7i1qZcut0lrVcBjeZDjYHfwXCaZyj
4dlkmXp/hvqbDSdszNzOvDJWEMvr7ryROXJDCvAoEgTLwzEmpbKiThlIlAUmHCFN
lNb5N3GF4A6lZ7o20jhhPwTcm1p6VVkkGeeFm6Kr4xSkHXNdznLTiIZWC3NFUzpb
cRzXO8g2sJwlb3e9UDu0OdtUbs9zwWF4n9YXNhojvwmMJ887+aFu1D5G+SB8o5Ds
C0GfQwRH9mv/6JX688TK6eAjy4PrEQzUDAh5igLEVkxIkWzbp2ekNZkQRIfMSGWR
SXICXNJ23bJ7EDP+reIva6y8o5NItRIzQQVUjOHOf7XNmlvfmi50/ZI/qEvEJKhM
grIPb26WZzjv9HtJuRXOUA9/SAbb5e30igf1OSg6G5c+JSkP5PnILOJXJaa09WAR
KIbNq+Qoh56IdKza7R/O/SMCJ91liF/aGlhdrrw4gGGcPjlvCdAas+wbj9MW5qZU
lpbDHo3UOqd3tUeO5Hxcw836PJD9UPQaIu/le+3zGOZL53GdW7EZKO0XWTvJrU0N
929QxaSjPK+VlRQQw2h45iEmUplruC+l7qWL8FwwkIV0Du1TiAhPIk4azC7PuvXy
N8OfNw1mDtLNBSXdnf7fxuc2pAv8lEY/YLmeRA3NlqURbR/n5RlJTy+oKInOVKxh
U485UnOeo0UW8LUt7vMOcXozPFwqW7Q2cCFPvvO2aa/Ovx1pI+BBYfY7gsVjXrRX
ijTTsH/L4SBmHT80XUf0kLfORBoT86is68qCdovHCpLIY0qd/R6LSfpxy4/4orP7
ba6zSeGtgtTjVu+JyQ5DMFn5zTBjeOGOQp/Om0/U+hmIjwqZ1VSSnqbVlwg44hqa
FsYlDYo1wwSsSKfH2VVJNm9/LvERBZZZiB1S3wPJQHxtwS1Z0Gcwyn+LIqVUjMdi
rg7dxvdgabZozXVFAlR4mPHzAwjsNyJNs1+QzHaR0u565mjZgkKF9LnEBow01tgz
aKVSmI7i7IzrmAwacGTdQAYVSeW0xmLoqgwgH1p21fY3hKAVOhmmcax0RvHFicU9
X381QssKjd9FWyLGcknfrEtwlFkyciIZ9Hi5LNlilWnZoagJUW/RHXEv8G60h2b9
0XjLtnJ7hUuk4eEdhNAbgLdQjt9UH1/HqNcmBrIpqm67Wzhq5WXSnIcNwJgs25Ev
AkxI9Yhzs37oVZ5mpC5t2dCh8Xc09BMfbmzPljyUQV9SBrwwQbeCbSDw3qYW1Vy9
VuiqKxYAKAt6uOh41Ox0SXurmjDiJddtu8/QnT8bwgmQfUlfYayGlWs2ARqZ3tee
nUNsXhoaNScqLQJB99BxwDG14K+vuAT/LzfNO2a4BgnT1YnxS0PkXnh3FGULAKWk
2ejtM7tcds6mQLHTh7XUxurQ9qaXneVgchKqCUzc45Vr7tSnIqUxbFP5gDa+BNLM
x2YYCBfTqu8DUIvGonGjm3KOLgFeZ1cn0fjIY8AEUudeTTqpqLDoZ6NMvWHM9VEY
guust0J4lFs/qfxIqA9UiE3CCh+CxPsT/nZo7ZQXKtnXybYPZZqJpN6Oe5dJo6i8
uzfNxE27Uj+exCeGAfJTBtCvVw+nsjClCOhnWo8YmTAz5e86RSbjHdYTemGWiC4F
QKEVpYoiRFlq79CT2davOIpHm6j6UMOvQdPh85uOKCnznYoP4VLPOXM7BU5UtYNI
1L1y+YvDAog80XPEk8T5xqA+HoWU28zBKLZtwTm+INYBT6r6qEvYELEo8mPb9+9K
Zx0GwExK2pXQ6jJYGfrov+c7q2K8TLHKItapIT7Ppq2ROvDsB6jEpc7RIy3adGjZ
pTWvYGPjTu0Xz06v5ml02Mo/dCF0PrnowbuXC7TPnRTpnOJTnyOwnBVMIv/Msy1s
27XFfWqXHmECkqRdKKLUCnU1XL5NP/vrEwBZbEwdXmgUd6dGaCPS1vI6PF+tSajm
Lnpi1chWZmsVVCMv1mVlCByhdYF396QyER/9Ww/z4NQ6pi8nsmy2eNq4fvw+Bouz
RrHPI4o1UnElyYgSCym92Pso0GHJabMXRIX2AxU8FjPvSz8V3/xsso8N/RqYVlsM
/P0CZdPDRKHSDlOsoi/DIYRhKWWc2EIEis31E14U3Y4+R1jV/gf8QqtlpOFSGpUl
lk69eCi8HvDyLjZPQARyK4+IRKNdfpnmTuCku08rWUeioIbq7Xy1ntR/3eD9NBJD
araH//IXjYNs2LnE5z6M72wjyDqy1dvxXai9rkkHToIcZhgHPwf8l7AZfOs99/Tp
7CHO4gv1LMaU4BC2DUAOBUEEza4eyJX9N4IW7BMSdB5AUZcbNeFChczGynZEf7Ae
+fUBnLLOvI3zJlluoLjE8DQ4sCcAjheyDZQjCBnqUUgkdMWCd7q7ywHRREF+fXTN
azQRGWlpNiKGZgp268LC57a/AVOq/0Wzi+1IOmUkq03IyztrVBVmJMX7WE8wTZ9W
Ipz5PC2imy7ib0HrnBqdtJA2QuihOsnyIMrmpdTDMhUkEHlSVa/pIPKemJJPVG8u
fbnPRLRidCQCHF7ODYT0P7TTTN8FrvkQuFoCr1jEdXov3stw1fdKsIX0MdZ32Kx6
WaAf5Gwkng7//A7tMwAxYKRRIjFPmmMiznUhJJ3qQ8Ri88ziEVmC/gLXcKjA6My8
6oBPtfdBgupnmLK1J/kWbeCvev2NqPO7Be6uPSoRuNJHR380et5d4EeU5nyTIXBY
Oky6RthcdwgssOQjBh1VtU0d8RKDu26DpmNb/SrPy9cf27bcRaprobKnl8fGraiY
riD5/Je4KzGjE3oepQQwmXMYbdv9E5V/b+vUBApTDOZ0/IKv9gHI9m+vq7FIirl9
paccyUceil5f5rd6VSZDctajMtwDgNsMrmTrnUoV5i6Oq10iw52f5JADIRrbCARn
eXzWQhWrPXdOXQLNsOv2AGcUpuoyQlI8K7+dLpFCDlJcvJsIITdXtdmX6wLcnl0H
EzT1+QbG5AuFu3X3qqPybm5MLdRY9PIpIZfSRaoyHmt1YzvOJ162fMWtk8q5vBLy
amXPCRnZQPv38F3ZbDebRMw8ekuratbYB8rSUh8YlZOMxw9cEABuVXnUR2Am37lB
0sXWBzndJ3X0eER3NiDTrAR1bUcAu62hXLijbjCQVqQat7m6KqPdb0pzhIeB8nKH
9JWKeafQ/WpjSNt60YobxRUZDsuT7/R/UGVZAWEFizyswfjoww0QzIhdxbFVqZ2W
EwdfuP8p/zMjbOqXVMGdMCJz0nt128k+/Z9vQQnerNuJQ8jNI+tMirWmY2xEcIqr
uh6arGxA8XzeMd72JVRivDb5uV7NvH7kQGW1E3LMKIDZjTdyvZrgFtWOKIuhxIU1
1WXBYHSjLgQ/+6oUSt592/H3EI5ARSGOmueURP/2ZuCSHDTO0xmgJcicQjIdL2Fm
h7LIeW11MGApnoP2QoPXfzQmQHqk9fLlTZbbOj4Wcaa8rzQGaQCEdB9di3BKuhKF
5ME++160uQXz12c7so2/J953+pDSPpef+wUypKXqAES47occIJTX8kSzoslOddFc
obPK+zLtU2Iwip2r+rCXsZ3nC4qgf7ZiTbAy9YWc3GZecaWlobtM8p/TAqF6yl69
JpEbjPlxcLiO4YbV1hjKsMh/QAonz5cFGBxWuAu5RCxBVgmas/PyRYbt6RkqpTGf
OSN0zvJ9KpAjzjC3GdrbF0DJHPOOIkQcjwkswx1HX/noLlEFTC7q4ram9CgSqd1o
Mg1umqYVJ+9ULht6qkRRG20geI8/zu+uDz+r1r6efqqe/riL4o30ZK19Nk9u9Gum
dim5SEkQ1/5FrJifDo/tPNj00M/JXXTqu2FKRwVzPFDOdOnGP1Xxib0ZH6qe73Ch
E9w8wDxSjROlKrYpym50t3Vogd9XG9n2sBboMTgcOx5BTNB49zi96I94uulDOM8r
Z5Au7vcJMBOdnYTMZbtMgXfhWMeZKza5gOtHZKwzh+UgRW9lE0//L4POtdyK0ua8
VC34VwLa8CbqiqSsGaqyiZ8utWV9DIS+ydtI0FFISW/rrDwb9+SkgnlACCd53Gmh
rr4/hTB5xgPJahph0VEGA+3q19Z64C/fs99eR6K/AuI8aNFJMt9xVH5K0FFkHHyl
08Bmge9VPJVyrXhLAddP6P7bFgg8rm50+vkTs00nnmoQRltYfEtHXJ21C41+2Cx3
+72vanC633RSgCBa+im5nbbphzFQXN1QlYGEGTap51QOa4F1v/SY6r0UtHZgJqpV
tthz5Lmcp2f7r/LWuCantqZqUDvGPw65WuiGdLxruPsw2oC0rbahd8Dwh0mNnG2q
1QyCH0nad4+MHPf+4LYyoHcoSH1pEfpaI/GPNOpPrt31zvogGBCWqdYB6epVzREq
SemKrd201CmF6ebpMmErIaTZcMtP/4XdHtFKXmAA0NxZxtJ20Gis+pRBsvIFyN2X
ICeYD2aVlDevY4VYd+eQotW3j2uB80qCDsl6VSm8cxBcaMwj9mvi0hV+8JFYyGRZ
3hF5Gzrt627rx/zAufAkGaOuK3wZBbucUp6Idg3RsO/bgbPfxcyCm3BviPTtEL5v
WXG2p6mm+7GroaVoY6R3UZxjswMrIkUKwXMiWWpFraiIPAvMOOWsblRYR3+imPNx
/WpHhL3ffaWCLWOUuAp8FwQSMWobR/+joBFxZqAbUsNk9XOEopMFqf/bx45sSPD2
7/BAMaPfcLiexgIwK4uMr2Hzw3l1cTaoNiYFP1Os7FrqklEHDldmfdkdSAcGS+I6
NKTVpVzmfY/OY79scLhOuEZtSygc8CSXE40Wcnn2MtK723HbahbC4+cBSa9ByH1g
ArzBFX/7sDTjLa9YgpBYjK9N/ijeXGIoxpS7aI/gp/tG8VwRIJOqttxUsFSOKd8E
aXQzYQO8ZW4JCU4CR0ELujWQ3GXjZQKhf8o9YSTBrRp5P0ljNWnL6146a5vxn5Ho
gOavNwWHvmATO32wYE9x0aq34/1dOsGzdjtgTLMy/1KNQvklXrq79aRWmvheu6pw
7utcjY7Qqzw23kk+OKZZaql0aGf7LXY4IcoGUH49xhZs8BaQ8jWP6bX9cLJa/a4j
LigFS8CVJfhwDg1ud1y36oBIu5U31bxp474FrwItTh64lYieH0Wswusz5JR7c+6W
P7C1cOVFLbmue5yKSYqKP/gHO6zovhzrs3yfvJwpFikcJ36BLzTvnakM1Fcp89aT
PpFEljwYfh3X9+NEdvu/ukQ4kEvTGWC5NWqBDGDZE1ZjbojpG/5MFOOrZ9z0RXEs
k536LQs6q64Usuod+lcrt9rrBcEQpmP3p73+WgYmhpyWSxUyvIxL82qr/JViEUoS
rvRYG4dTilbwvfJWHgAs35qdzB5v8d9Ggr29gL6rRN4KL51W0kG8kpN/OeR++QaF
Fnoo9+o1Lh3Z1XNQCKPjGGU/D2YBuhS0Yf8uu6fZ1jwOpqySnwMy6LEy37LUZC1R
Nd4J6qI6u0CO5tkXRLOxOEu+/DFL9yWfeU951SmWcqCgFyykSQkKoAVYkzcCs4rx
X+0MXoYpRTg1uyjvIoGUhToaU35885YUNfX1L44LEUnS6DThb20R+oNa7zb2cKoV
gDoV+akPVgQ/fSnmm/Ac2k7JrZz8J1n/gtEXK1oa6QJumM9fuijFz2U1uTVhG6zb
2E27IK75cHzzMJCJcHFyC+i92TGYcX7ACvCHJipdkQGuHlA7+pvrqRb06857MVOq
bFfP1zxIJKZUH4ewt/x6UYlzoIOay+T9AXopYJoHohCTNftb6Xlp7MrtXKMA/7WD
yY6gRgKKKdwQZ3jnGNFjyWWk3fq1E4ZCfp66XHm4b++aFqSTS/b89WGp6Hxw1ZNH
k1G7aAWEaz5xMV5yrQ7hN6Q1Zt+pZq5PNoKxKIFnO/rIs/LrMwYC48Uegkq3Yb8M
V+SAWAAHJH5NcRd8FkYpK82iirWc00JoalvCthvdfIGgJEtOAJk+4/mnT2Annqjv
oKv6+u//sQWgV9xWSwMYY7xOX9F7TqPR95hy9lhf0ceSED42FshYdKOtYVPa1gMf
lZjoi6rMeY4Qi+LUrdaQOWWjA2LzKolyZymIa7iQfArrSmMTdjb0YWYvnYhtYJtA
53zSfY9Mie2Lknt2S/f0EbILH+P0Au5dByGu7oiiRoky4zjoDN1y/Etvk7VYdZjT
++sACjqUSZbXt0MLb/VFYzsNhLN5J2sX3XpFt08Ezd62D4QPA+HVCvZhwZPzxhct
5+NfVhhK3QG9rgAxD272e2aqwhrJH+a5ft3EbNe+lmLX1d/GG35U1yKTqOpHmitg
9P1Xu4xddTQIjQZy1dEWlNd3Ysvn582tpQrQ9KmZSjDJFuhML568J/8AU9nGMpeb
7ifk0nxoTd4LVo0Pz8WxmsGCbiZMNKEuOa+jFkSwSveNLyYFPqXrYOUpZOOv1RBO
zv3YYqSrEkMTUO3sDBQq4+ALPPTe1iOv5EHgzjG6nmOsMVdy9m6zYDCSPl3VKyCH
gePerRe4fwsg2/FBk6Q8xEB+yxS28IiCqEJK71jN7P+EoMF0KpXmku4Cs6NtByDn
iwZlD86soRciOyHHJ7sr0jKuiAeOkoZVf+jFhoPVihOfhgUDH/0q1/DQ6e/3H9J+
0TlFN+qPlV2nDg0DOunCctgERYICz7UU/LippSHZ1Z4jFL5/HhM7FNtgWP8AJMq0
U8sj25TrMJtpnTzVCpsmpfntpT6wyeVKENoAusvctTBXVb9PkTcORfOxCFqGSspK
FET0sIAizffOyUMIwoy3Hgim2R6RXIVd1QgL4+eeX3545+s+NE3htWNMm/pN7GVR
cGCiwOROof0ICDZ885oTS6pxt1nI89oL2ZwofJ1BPJeg/m8utHS7AesbO3fhjeEJ
WUr8lgO2v5srHLnLmOuq8L4JMcgJrV8HzB7k2E4jWGVxip0/jN7f2SPE95zJqfdB
/nV4tti5s8Vahl/5QqJUy7viO08BmFV5FnyDPmIUv/s0QGIw6vScRLucKsaOClSL
XjAvAfflVBw8QbcFA2Dphzd9yG6gvBPj4tQ1hI0yRih2fyw6/QHwZinOgfJCTKoW
TXnLxcSeIGOIxKJlQqO8cixpMqhD8uWtqaqknAff0/UqbYnyz0+kWWqFN3oQvQU3
DDQWk70iNKHJjPM388cJInDiy0aYHsvFbONyzANH0ClYqKD3RU/LsphdNnpGcw3P
MdG1+7VR3hT6i7hCdS7/5oyEOuxmm1W2slUeOGy7wY+UNzVgKjy+zkMBVHAykbHe
pxHdpyugpJGNhF6ZjOjWTB+EkSB6CS4FWARNQ+54FShOZqXA/1MFaxKeOR9/uiRl
1P6dLgq7GYD6lp7QmzjuBO9RqPT1OICfhAFi+kaX1mIiODNdvhGcMWUV99ISA+In
Ee7PXRQQ5UOEcwnRn9KmoZ47UPVu7Mo/PZPljynQR8f3I226Yec5z1KCeEBIieKw
7h04QUyxMDWg8X9WyTgoRFcBg2payMFBTO5qcINEKHggncOl9gDd21ELGQUZeojw
1HRT13PIIkSmHGsDJt2i+Cx8e2ULHH795KR4GsjptfcBPfgrOzkeBJrJ70Cfipyg
dLhZEBi2xesjb8B/E9ph0fkbTv5PAXyYuuMGvEPtmoLcjX6FegwKNP+TaqldKNSP
4pdIF5OUYMjF3E8AlSbIResdnP1HrPcH4S64j5yU609Ja3PqTF6COhUhuJJEGzAd
hp7letFvvu3LnAdQfhfuTNdf4pRbbKSmMoe+jzfq80wJsRd2ObskAFjywyYta1cB
UAJWaO1tuXY08fDD1O3qA9iWNis354jF2NrJ8HsCXNDdPAsp1/CiwPqXDRDwkMJ4
tSrRCearksmNhH+vwWjhMRUjI+35eMhehIr9D4HlUSLfrC9wTCrJO8Se654djyQ9
0EnjE/OwN9FYh9tsOsacQrOlm5gNHveY/Z4K5D/WAP4bTCSFjMy/ncFbLPddFU6F
Pu/6ZNaImdnMah9yoycDIvQ6NbI4hKAvKpH5wVm3nEMDgNTMYEz7Ad0O25LhO4jZ
v/R2sMOvzUznc/pYkRDLxGZ6OoZ3JrDnklsKoDslvD1iHs5cgTPDsW7j0q/bzxom
wjm7yyph9qeG4fU4AE8AIwpHPowtl+SrgGMZRlQTLFn4hkfZi2VBjKF8Llh/dNl/
rb5Gj9JQgwNznTDK+PgGMfzmyMjKLMVJCLDJjA3X8BtON3bzufHdEa+xlXnsdI8M
KiYhXHx9IJZVtBn/sGfgDeH9Y9MFbUgpMzuyI6C7YqvZVznNvt3j/U2L61FiBFkV
26jjtibQDypqZg6XAWhLN1h1U4fKhsRapHORoPeSgmrKmE3ZiIAnC4dPe1YruxiS
14tcTrGlmZJSA3l/LuSX5q+r0I7vmfbMG7ajfqy36ffnii+lYDCd3PybbsfkUS3z
JdUpS4R4XbEBTHjolClCaW2SSSaGg0pgcI7Dof93yK/sHquMW78deC9sjG4Wy1Fm
u69umEJHhq5/+8MwMaW8U/Hs8+bqTRrIZi0kW3cCBGnenmQ8yLBjMYWJFkwZFqi+
momgkKO9GLbxERRmOBkk3OkxpCecLpgN/drQarFRxs19CC4gnWnfHl3KzZEwV7Nb
6uzOVe93XFU5E5UjSFpJV3gNfwOQlF9UNWyCBI+N942Q+FmK2W7FyVqqRWqrKIqa
lLujbGbnE8oe0rE0/chwWqjsbNe41ZWd9x50dG+GLgopo5CLtFpUP5UQt+DwUDxX
SgDDG8nn+F+VPXhCZwc8lggEHyM9b6K15jpNhuOh8/v5wt5ySOPumTtAzT6vblRe
j/jlgqiU64SGym5xlfZDdi+gs79CFvOuf3TaQfmtk1eIwHzJybRjmsPdk5uHm1Ab
vnNIlzGHZ4Ucz3FzcJVuzRC0FtDg5H6n8lSTHkH9WVg9bd8bLBsx8SLEPuFkH4WH
Cy0mu+YohRiuoWXXVwHlt9pkPmj2sCiBebuZul0zBs2qB5Guk23AO7bMe4mdOUO1
777oG7PanLJz0vTUfDmDYmlWb2izFvGg+yc8uDryKJP6SNtAY+48URx4UZBUWZ6W
X3Uco/ip+izqz/G9j+5wFvHVD1Qp1yUFnvDSDmsaPR7q1pInRFZOWRzZWiDPzdBV
ZpVVRODv6tWFcuOkCqCGldjhxgJgea77XD442vsmROjgv9MK/u6TZK937HCkQhMJ
QbM4vnzTx7C+USRuz1KDFOPc8K0SArMAhSbjNurftz0H8drhpT1uVp43gKt8E0+d
zQlfQggcGyjBnTW38+YbcngTaPtxlioh4dw/DPF0okH0WmIyuigrj6iue0BAo+cw
/kNoRamMy6oOpLm/pzU0bi3S/M8uCdfSXTnDbcD0SqWltMZvmf66Uh2k9xnhGwpg
/0spAiOUqUGeEC7Nk55kdj1xVDNKzgTNDacxqCBmSTot87ACia6Bun9QfIXD+YDA
Tgadx1Fsf3tHF8/4GftJZVykRk8PIQ2GQ5cJhslrZdDYxV+26El4ZSa2aoqbRsre
B3CNFP9e0NpI6j8bJHhEYEpg8y0hTZC/6pDZtgWAhM6T2jY/E+BS870eNhhRNs7g
NcIOAY6Y1ikMoKIR4yMrPLg8avfm9DxPSTnDyJGVpV/0CSBzKH3bgmTOg2v8qR39
yZUwbxS4TxGv/O89MCUQsOudu6V5mganv0JEyL43oEPB5BNecj9n1MCJb61YNFvS
eto2VdJ7awpvFFcsSSN6oMrQnewKfTFxjp5q209BBb6KtZaCBZn5OT8YyN20h0To
BB5/2FwsnKQ9jdUh40TAhDWjQk/J9vyDOO3EDDPP6f48vjxLVzTPxPZBfUsvYjDT
DfdGIv3isno0mgZtfJ9MZS1k7+UwIHSmPiVR/konog3Ba+crMy0xLDKKiZtlkR8R
930U5U0D3W4+GeaEbLsQi01KNkj4HZvFkqHPTtZxMisSifyQ2Rb43QE9xS0zq1db
ou3j5vCT3wq27K60cFxBoXzQO3P6CT5v/jbiE9s5ToGn9sWz5VYuLxBDiyyOLwUG
rFO9pMLoYt988D+QeTEnq7d5jcLJ2/CSRq8aUKOu0xTR9cLqXdkDZBU80hs+1Qfx
DapCTKeCKlz9bcoO921MYEae3An1Ei1q7WmBQ0DybNMaaAXFYi0fMk1KOENmCoPg
9onUfuE5Wzz3QUowZC2KAHzKQ18WfFI024RxgYIHxF59xWqDXSIgg+YwSAzH2Puf
9SC6Ws7e6tVkDG/2wLS0Cre2XTwoqUE1aqn+uyek85h4f2ZtvMrQSLQQKLw5iJsY
kr+Z9ZMz6mLkv6/V/e4xOmbqr7foPxmpQloQ7gJIW677i5i0gT/2DQykiLto3Uet
bzMktEoKjHzpOfcyiLbZq/EqjDIjwZZN6IcMBLkn+/S2nINl1eDnd4ncdM7FZLXJ
50QWsZOS5oklz3tVMjGFDCAd5YY9+yMRFyDES7+UAHFwvHns8u0Onw2avN6q35lP
LInR5OGMHVSMGiPellScexEkcmAy46fjkVy6+sG78IpukPZv+Z8O1pTYkUT75g1s
eeG/Uy+iNsYtZQf6tQyVc9yBfrTNciwvn4Mwt1vUuvMz8TF5jmNFpF8KHv6pAerK
F1tFq92zKHPjN6Dso7ABL35khw/JUdq+WiUuTlytPrZ1vF2UoAnNvwuaT6ykjYz8
Ene971illxOAPpaGquajizFqrrS6WAm1kKO847O19wtY62oTzlwu22/QJnkItTgH
OB7a1vI4yx6AYAEy6CfWPE+elJQrXhrQbKJ3CnysyLXg+uN9ryDfrb2EVfCaFotr
uKBpfmiQ+NKx/m9ycmZ5I+Yr/XodAqYzbAEVNkp9J2Mx3qGjdIZY8rgeKHlMHbJa
JLKt16OnR30MmqWU2gVUandBfhQFVY9bFjuYM5qmYl04TDH9hEP+yEg8bYmgPCfN
MZ1MX2m6bDSXaUHJ5KncYRaxtUE5L/s9LJWxEs+JtjRiYh+VSrqByVxXeFp+wqWo
ifhG8ZQuKQTMhlN1qgx/Y2uVyhlI1SfvIeDS5oirwukw6JwnSUZctBzuS7Z1pSSK
+LhAz+1QzYoSr/NgvOHGWEz2JwFoaHjGjALArq9/VPC9Yd6l/oF6FjpZzp9AiWAh
rYX64yMMwHWSBYx3BNUGPjkaChcvTJSWSg5wKtN+mTp0Vah3+nX1woeDa9ABhbqF
RTbq6svtQeDUzoXIW8Ga+TXVUAVfokVVpjlss3xvmCBQX8utESEwRMFllLo6mR2f
Elf/JOHyU359boEeH5X8hoo08NdE+DFmCjqTN2tjdPjC2kNkymN7p+XCX84QRu/F
ZTSC1zSLoAZu0cUbb6PK+2s9ZLvxjyTQJM1Gi1QxS8Mubu3/dUSqbTXRoBm8Bw9w
t6hpgnZD11bnKZqX8OgT2kLKN1U5aMDVY83EEYm+Aj7I4Bq3MBoesCvBwDYrZ0BP
nJ68rmPiZuEgCRnVZSjQXxoZD5svS4yXrCew2DwFUxLCXxx4oVDszjgQ9BfacJCa
nn5w1R1/3wROtH9kA148+ER5xPP43sVdHKrvjb3saGtTSbMD61HBqRgAmyc7g+lS
F2vLGXB6HSf/PAYWUpbwmT1EeH4bBozKkznTAfS9RL+H4LyvAZmHi+hbUTeILHuQ
fJmxT9xA/FTfiT4FLRVj2CiIERi3cDnbHWDCgC/97eeSbmSbBxxc2LSpjdkifYuy
dCtjoXFIR9YJzUlMAJ1LZzgQO74hsQhH44FI7mRqP0YYi8QYNyez5Qg25fpwqoe/
/FZ8teP/GW6uZ2i9pAq1j/IRwhxfKc7LMSxg3qCFGm5c8StHZSeRS/3jm8/uKHuy
EWM8SmLSaMUrEcv1uE6urTFvdgLb7tgVcutKUTESl/gLw7hcM6HpIPIYAfBdYEo7
HNjw2W6Lcn2zw8kKuueiJ3yovjyNcYC9QaPnAVjOnIubcik9cTj2Yl/yv1R9iNKR
VqvfeXZpjU8u7PaMIU4AEEvvvutwVGAqSRcdKx6lAiQknLzrXmSm1pDB7OAHaxkS
ZB8n7smrVxmIh7VTLScRuWRKzso5HOzgDMFPTWX3f9TX5CGjB90QrwcEP2OzdIAz
HChRByJrw7utfQrjjXjZ0gKwu9ENhIt4KEBOY3dig+eP8wSbW1/Z4dWNmmDxlCow
kh6zuqwIcn6qs/dL67b9RLu+rOBgQVXGQAezlcfZ3+oU7B/bxTdHY8ZIB2H0uwWn
qI/NSzBIUAxy8qE+I5opWMWqFZbq0U8zxOEFh+wC52zgCVY8pghtmhAj6hmykBI+
87Q3BVPB5IZRNHUe1Jop9bIsq3PaQ24xd6IRqTuVyMLYVsDmEWPua0PAm4obGAGr
P/3QYWADcXmAuZ4gh2Smm7dW1zB/ghgq/iQPcKBn5fFry+kzXzdv7qlULwmPcOrj
6nG12kEStB6qDDTRhDgVS/CAwTJmzrZ6VVYgU2zwAT64R0GZa4R4O9LZKIpH1SW1
xz+k6JOo8pYaX5zltQX1dAjLyJ3mYV3SO6Wnwu9mc66UZX795kFQ7Ejt7Plf8zWo
2Z0/IYFcQFUh+72LsZJ22lnFe98p1fy3TdQrUd5Dk6e7Uya0GVaYYBME/P2mwsPB
dr7DdSSPsvNvZng8xoYpCnN3q4BlwkHGX5BD5wGba93jYmJ+ocq9yaLIOk+izVRO
EU71rTPzBY4UMmK/AuQiVCo1hrMMNApsrHjnDKax4RgKJnmZMf6AI2wmnFrpY3Bg
1NsciFENjEl1yf72d6Z6IWP0SxMvCWSd7m8Fc3geiC/Gr8k9xV8aiDvfiAzXPoPm
r5+pkVd4Kf1wt3DydfL+qDCV0T+xEuBb7+R/giGL14m1cgdkLebFsWJNzMrwJGPM
2NY/lERvyG0XSCryVf6A0EkgaLBX63AHcEFfyGlvJcuV+6FxYLdHmyiLUffGray/
Ws43ypGZ7AXA0818wBMFIohBcSXLfu2I17LRpIKV553y0zEPWTtP+1IoWzitJ0uJ
owNIYT/18sk1n8TLGhWKffGvPo5A3Tq56CoOt10/ED/W8w+tM/YmK30tRX2ejAAM
AV5J7De3vyQ8KnXjUZN2alEtSyI5Ef3Q0lsjTRttx63N646glnzA4z47xxi/jNoE
6M050SmqlvjmA6f+UaAa5ebaSgBglQ1DqvxYurmDtNFzufNbOjmfwKLVBEaA3RS3
XHtjl9/9D22jJl2E4DhXQ0oj1jBcjH5uOzLHLg2G4ZqB6zPuboRUX1I+lKMLITd6
iygzgfbvOJ4inXoFahQSb5lz0/YMIqDsilHMhiZNTJRBSWYMjnnDSgvkeypS2Hee
uEouvcQGa4JfMazd0PhKCgqyt4mk346BZ40JANtm7mPPITlo25Z8HKqpl+dOBOe5
WuD4r5gIZwPTFqiP5b3k5UG7GIGQhPF944MLiK94Z3VCDl+eyGwopWMH8PIrfl24
njlrAcLWsuQgIgXkvzFadRO4m+P19DKrC3DczUrcwdi01BUmEYVEbp94VDd9M3Fl
7FWA7U9/az3+jXVnEH5cFVpaV+Z2G8YiO8iKMNjwlWmtceJ/kd99/DL8FuMgauMn
wkkNK5/xhPWMCYxmjgQisGeck5X5jtnQ/JvboGS0IrJEOmSbrYlsVkkgLSLS5BJW
1Mo3GiSjWaLPTXK0k6Xjifi2yjqAFdDbc+IzR3lp41zAKhTfQGXk70OUR1nu1FWy
3u+74amt62LgemT/zpetloU1YDxJhhjsiq+W54QoxQe4wRHqcDWy3OLQ+YsvIfr5
SvE1ndrTA6O5KKb2y7sKlLMwdquVYAmCFmFI4Ve85lOoSbHtH0q5l2DkUDEVW0gy
5HZ/UOI1rakNRu6eUmbWFfnPa6TcnBCA0VDBIxHWdiaP0hBVAxy1MXlgNUTKW856
sQ34U9SqES5Zati91g4uJZHczpR7fqVTLIAVDoaxjlQSO6ga6YGREs7ekSxh26sy
XZLi8vPE8LBe7Kv6FP7EAmivK7YS1mBQT5RpiFz2l4/kousqGVDCRxq+pBAymH8+
bb4sJh+BDBO/h0miwg7ibLolJWJfzOgCFGBoy1FHyzL8qGOeurlC75jo8tZDBsKB
1ru9mS3bn6Fn3YaLTjKg+oWwysxUwSHPMm/kz/wfr8vkQcooUEIRzLdU3bMuLtU0
CJCQdZpm8qF4I7xS72aHhxzFNlXmarYdqoV3JyIM7vsObnQsCBCDvTpkrH0spPmV
Nu5NP4vUVC4VaYxLfP/XywIphbfAes5E1D34gggOoZe65JwWNF66K/02NznvL5wE
17rAUWFCifdnAFjCDcHgp3ZEueJynyFwXofZz31TBmjBbbmLv02P5tlKHpHYbu93
1+NBdT/akR7NE8bHml4HkXZU1M9Ie3kgALDBgx0oLzyXSCCZhcFFdYJSX9Pqy/l3
qGXvNk8Fy72xC4xDCQ9ai9BRLxNtxSCJFyr/sGoVMyoqKv556vR9dtTBh6K/U/HT
wXRV1blWvabtARd3jLE55QVo2CFFBYbgsgBpdVm0EIu82gSIG8J7ajiqGgJTzYgL
NbJu2W96OvKcsCS59avv0FwuyyqXu6Itw2gr/X0Y1vBigUq2VYCn1Yb9sroS/vDk
EZCYBBmCz1B4UE9zo6cLJjAvXiTmiz4oMnI0qAlRhYJIejWFQNcZ8+RzXHJ9giNv
5VIuu2OnBgwrBx4UVcvTb6tbTWMC4kJoEWn7xB8w78F4n59DXvOtLkRNfVAKr2RT
NLRlp2OvSTe50DVu3TrX8UrdFGRadBKcYsjxZNkHQzX8ZxuWkNWuH9rNWzMoPUoN
TrgnZCso88umiNhQP+2pkuYX/5CvQQgia9CvRXj5l3VUpCKDFyBSrZFVyYFVRPI+
TkULDYvnEADLEeISoo2JknLayvthjtooAuZJIzpT3/JMj7e9Qr1oUZ5nZSHcQ3XU
tSQZPN4L8NCr1ioUj4eudt5VNbCZps1XSE4wq66YrH5knK+OoENq+PsLIdx6EY7a
yO/vAcQra+xlHxLNHkJD7imIL0+DanLuvTqJG3qNVSTha4uV53P0nGFIPI6xKN6n
l6l3BbMPD8BoE+WVeAuojNRpdLJR4uYmYxMugS6/WUiYsx61I6kUCLstkrEru9BM
n1UJjshZYUIPP8MjqpY/mgyld9zmJoh0BK9Zs1IhFAgD9uE62U773mCkOck5t2hc
S1vTelKSfCKLm/Jqxdamym4LNqRYWceyZ5JaTdrMmlrrSAMpC4oTdWcMrwyf70NH
pPxlwJj2zgn9VF+BTa7rYscGbEXtzoHYwMkJkXSZdc6qn/rSdggBSwEopgT24cDF
AhCp3ezHPGa0Cv9ldj8j6opNacfX9wN8Hwc3lCSb/w+/MfK1Zx3VfPJyKUPHMuQw
Cq/BC34/7H4cR2noyS+bc1tvuzS75y8MvzHQ3O0BKv//X0LyUB8D5isAWeNvrO5y
nknjjMzttCRhHuphYayud2mVAPyL505RjHS34k1MHso0EJ8BLAEXGHCOgjy2s92+
qGb1Xg9wOzzOaIRaV12NX07ETFqTKXCDtsZeJU04T9LPBwshVqQkCx4BZ4BokHA2
a1yZj0090aghb9OMWjXkBOkcE7v8ad2FyO3yqLqXWZBAD7BBNsDK00lahJkAcnD7
Yw/61zYVZgXEbqQoH+t2iEDB984y70gcW3QUE6IjgPWYymLWAXv8ASAzSFxARfG2
FHoJ6MJbpEdyFDfljYcvumBWcdUuLrlXAjF8/Jj/1Stwwqr+BclNTRIpP2ktdym6
QaV4KrZuh2LsBRztBoHU74C+m2snBLgcNkkW8glLRJWNP6RSJqagESZdFQcv+DX8
BpYpo6T2EWqjdmexf2PJ/OKPjSTpurIUg/D04ADsnnla3FCwarqADShudzMaMjFI
2wCQLSCup4WmhyhB6MsVMU0sLDvI8iRqX+OFKOx/3kt+dv72TTxj7LCNSQ3vKciv
aBA4B+kwCelEJti73nUlMQy0VD/nZofx5DluvAAoNuHYJAos0FFIWo/i+XygjonG
RRmtSvxIyH6PaH1FUp2/F7vAfAU7t90hMX39dDYSHsI1KIpFLRsaLDZ+UOgA/yrT
TpeW/ax4laKjBkq66rhE7zIjMrp+kPRyGIziGnKxYJLsHIxcjDBnp7TVjm3ZCL58
dkp+rBrVz1W8kStiCjd5lON6pNuNtH+sM1FLZgHdZIGRExyy2TOvjlJli/mEpERZ
peOj4D6TaIevydGmm6JlNY3q6l7Uji4jFoyY5UWAwSsLQKdzNBPmiZhTxu9A9XeV
xkPtjZ/Ig/LdIBJQtSL0VXRZI/q9usYAf1pJSUFtx4q78YxJqi+1tiNHyp6PT3H5
2tpnkgt+gdB9ifFLZjoa3mSuzjiXatZsQSIva/0bSgwIU/TlJzX6RhYMD7PKy9CC
kGNoTpRiHmffKAAyxCDGKEqMdFnD9w1ZLGujXBC3XsRH71Er0Aht3xiSYbuzuRgp
aRkDOXEjuqgZyGg3i+K2Ax2RagJhSsI2uWETBjaL+G2uQAGU6Kmu0RyZbxDesRh6
k0A7apBCVkme9O7m02pikQjbcNR9c6W4jf3Ttko6bBZE+3nPhebqm9KF18axi77+
ss6PWXA/JXwRO6+DC/dMfErk4XfyHsfCiN3d8NquboWdL1sUSMDOJ0Qk5EKoVr6q
RYfX/abJc3xw003xD3Q693V/vn0u5HuuU8LsvkSXYoQNnbAI67f+jaqG9VWpXfo3
Cet30hv2a90DcC0X8zYRu5GXtaruphJvQm31ONYb1jB6AbB+Hwr0sY1tYuZuj/K7
vyGIPD+yPaPD/JphgIUF/ey6rTlzy03llm4iaoIg9gfPvLA+JRh7iFiWXw95f88z
f1513BNjcVlQsGaCl/79pIiqMGODjuWDCJ68brSJbAhS40OPVNgX4yxiq+ZGvPzR
kVfpnoJ3NR7pk9RNMWV88dke0uVjw5fBAHj11PYP/0pZzNlt5o2Mhex5dMLYwJ3A
ahA3qbrnQrqjL2RBXj3gG13U/LCf9oWPY9HBuYhiM9fHkPNTQoSclmx/vjRMs+4h
ZuH2UjIVEo1YyzYTLbEljPzzcTH/Mc7sl0gIeJ8QoRNE8xXl1PNn+TSmqglMYJVs
ZcynrK8yAbGsH9ROxunpRRJTkewdth+6V0Jk/UcsLx0IdRpyMzZbgtQ0kE6XaD2e
RPX64pBDhM+9HbyvFqIpfDbCx000vx4GzDGHEVFxbB1+Gof0PFYOF1to8+/SV/qB
Yksbfzp+J2Wh2rMvxHFpaHqDWSBqDj4jAj3y/NmdIeqajbL+NcewaamvDGFNfXt/
A2q1lE0JeXssOHCdOVzz1DYgeUYDJXUMU/MNQQIkTBC2rALhVb+kpNVLhleBx+pa
xeHTIVSvFYd+ObLeOEjiydJNmH0FEeZ9XpCsfcQQJG8jY7t29F6loDciIrUukj/Y
aYiV3682SUlIeyd86vAq8aQ+0vJBjtz8MQ+J3S+UWZ38w9A3DTHKnOOEUQHC83Sm
T3PxPdzbDaiNAF9IqrlXO24jTYMj4DH5StoKO5PYcjFKQ90wvQ/KkygIl8RXNNPU
eiMzZGZCD66pfbNtlg49I9O2RlSRUCKPmudnqj6FBWEdXzzxKhD/QVJw6iuLyCnv
Zg7QJgPU8RGqqKyGXY84SoNmylPgltsyNd5vSyBuECkJPCND3mzgBi+QPnfm2awW
xYSxZKtgpsqOu7DojFdAU4miacht0lTOjMEZTkJHPsFEFnYp2ZvOg3WiRAjgsig2
qkR194he9J1zLyvo1vvyulAV416wGCUvzmvO59u3reC8YbUjF0GOrMIfmo/Xt98F
jF8o6qFtbTbx+mMEOpBq7AhClNxkXPKbWC5sma9/qwah3UV3f6+nwRa1sGLNVHyq
q8aRF0+J0ta+6xirwkvIbMRbG5ulOxEd+UtNsholvfKxwtY4Domxzn1eEqgvl91T
UD+CnWtiAlpXLvHFRQcDciAFL3rGzYbn4qrO4vySwGddAe9TOo0BezxRx4j5zAQm
mii+8Y/TqwfjJTX32jVDLfAZEclihI+kU4Jka96kLMVfugWH5uDo+l0JVpvvWZ7R
deXugiIohqNH6uH/x88qUzyTUwF5sY9bX9tWCK+Eohq9BVyK7pz6zHZ2G8duVRX8
+DoVSZcJoqUPq61i20c6xStJYywMI4RgX4efX3MasAm91vaGm0yHmSXB+l+Vq3ei
JPYzTwrx+8CYM2SLXVHtnFXCYMS4O9AzVaSYvSyvj6YmpuW8/BcHU0iE9iIUhynW
OZY8+y+OsJIJylGghig0Upd0T+2lRqb1VgSS5mqSb+iKS6cayAZpgdW8Yoa0JH9o
iPKgt2iEpKqjn+fUt5fYCLvzA/IM23LPEOCRLrxWhHv+pTu6deyuJBsISaAzJO6F
AYDKWMA7h2hluFnrNYz0MAGZhFL5Jix+fStCjBdjothsZQXtq6q+JQaQ1+ijNISp
qsPyg6Sy6WSZQ1aUzebe1++OJs3oW52W21BUB82KFAL6vo/8wFZngqkpP/zTgQh6
lF3VCKdHoDYp9pI4cXvq4fMguifwD2Rz9W0ojvC+V5qp4+NHWEVQLbfs6G7OK/bE
p8PxLJojZXb48zl5Yg3cooqsJoWf/avuXAzBi4eq/xsOl/NRFJXrZsWeX6gO65KZ
tG+rZ2bzx6NlSHW2Z4kGPxSmX7NPg5aEkx1wJ8kPMgHKoiwpwVmGNKRGruGGHl6J
ubZmZPWuDtIQgv2i74T+EtnzrSswbySnNg6ic6OTC/OlvR/8j8IxUjvOWv3rWVLC
OpUAUM8Eauy7JchJSMwsVs52U95yBdbhTHfahAdu7WvjvahEjDSc5hoFskSYQD1h
fDMjh1FTbibsTZk9HDVHDXvIEIEMpxxO4SIRBGwOkMo92nzODTG5IDtKvHSc/uOC
Zt9ZUhGUUx54Re49s4Ely5tSUepVKK/oGh7/D3U++bfsTadcyoXzENaoBaY1zS4q
tCeM9ETk+RndRGxwQPaZK+bp/a4mL7UdBCEXfZCLGu6vm7jjtzBACbUNP7tXRxS1
1hmZOF/yNRj84D67nH+TyBy5YDSVOj+C3M/GjMy2IV0zdt4FXzZcwLmZ3yMH5pav
oSkPO72CYYTGknJoupliR++5+mhTLPw5TIEu47AMpi1yATJ8VcAsg/uq+/k+aYza
Il8YBbeP7TpA/Tb5WDC5oB0zKRkWZsLh3NIK0UzkOXO64UIJsPIkKnpiFj6BwU/M
qcCMfrojAC43zMBtgphcCQPvqB/z20Dz2CbI+L3d8SxDyu13lIEoBToaj1UR1Iwh
YbAxKiDfVSlxRiMWDLNFelhGbagc4tamJwcrkQ0zmlvZJXEnN6mriVQjYnZn1o20
57YNhnCl+SjNO0TEDAfkjZU6c1Lm47OYYgVmmP/nUqJRv/J5K80w2jIg2csfmbcP
IZqcSUfs0t5zQbiY8MAL+4DOJ71glwT3PNXd8QOlmQ77HVh89RclzSwe699vsT10
WnWYjBdDC55qVKoFYZDCsohIifZT7tjnghiukdBcoqpeSDNDvioHLm169jaHIS2x
mC3dS5SNEL8td7lLO9uKTrPkIyE/bvwUZSzbyA64hssCfhQ8MJNXuh3rDognzrv2
k10sH3J4imATdiy+BqmzCKl6gDa9EoeQHd3oDglZJKGniBnu71sQhGtnr6Z1y17i
BHIeMyNGTLnSLHFpoRCL3P6ur/jKp6eRuEVzw4yowR2QH+IdyO9ysu/ntwjxISB7
NkkH3Z5OPHbfwgU8m0jNJrG8WW/GcaF/vUoVyZKd0p2eoz+g8t45mbVgt+Tx8Wqj
J9/Eg3D+oEE7gahiINhJqIQEmB9mllv8jNv9fsk10yqyyRUDpO3QLuTAqLytvWdf
PNn7Y4IP92H8QSZ8NwuNTa9L5pJ5Eudm9zuGN0G+CcC/P5U9CoSK0DePgvJkxnhb
2HsHRjEJ1je9PkZ9SnQZbSP3R3ZybtLR5wmnhcqY2U7WgJORt10cTEw/ZJrc4Ges
4D57jW4ISyx7DaYCCFa1/52PP8aOV7Kf+1pKoVaGCVnTxDK0V9SuZnd73m7ExfYe
y0fsZ3+mPJQTr2HIMUU1HerkpQdq/deJ7lsBtTMqbMmmvR7MLOZx5FYspjsqr+jo
n8GQvMYdJG0kAHa5RK0ddYkDh1wAaTtOfmfQSaipilbvYoY/3oCGIpnjukMff6c7
ebAjzQHAZ79xdxaa2gNLOS40GzIvkZ8St+OCzOGeAWGJccs0MCm49UPFBl82MZ+y
37a9s1cGzAnHPS3K2F0f5al1TOXhw4oDZEITJ0sMUyE0lFWNWC985TM65cufYzuq
W4yL0VN7Auy2Wu6Ye10OBW1Pb1mxd5pGAZy/FHXlbwgCD2YMZ0MeNPAY+EiDc8fe
OL4XT7wDwhpmGBYfIMysy6vY9YyTalWhgDuFkoGUTGd9F08gazzomYXL9DwFeNSi
PaLIm2nWGFXTb9gsx362pCFEaleYt/FZnl2OL84o6RaARIIb1cjiqIPfq5RP0KOI
4LDOAV0SwMmxs1ii8o6riIVtvyw7iARnPk7O3bzzPTZP4nF1vDNtk2rYLXUWNecx
rB8s1OQ5qC31+vfupsmNm+j46k2dQSdOn1w4ajoTFp7AHBHLYlSoh2vd/J5XtpSx
J/Er/Suy3Bdvm6U7trvawoo8yjqMDwnUwsCgbw0eLr58jZ1Pzwn0w0GzDiOUzhD1
70ghMFW0YE0hi0cuTIeHUke1NCbnUR3c4nOEW6avqLPJWAxb7MBOIk63ebRQpVIS
L79QCvFB0XbsfzWQcAR5pzkLw+cJZBpN+TvBDaFiq0mUx1BV6OLK7ie4CrO58e4f
HHoJ9vaixsPfi9fnMLJCKT71P8GkpwS8i9nk6ZwBdFxsl6yTmbazsJMRypEMa6tN
t5/nc4nPCsBHvz7Kx+Bfbie6f1sCrg9dqNxvRrZeYIJ5WU7T5SjmgpMpCde+s/WA
wJHjuJr/e4d92lBRw8aujQXeNThtt0freNEUf/LaUCRgq9pvyAGDMLSsIb948+fU
WG8DXg3ug4g25GVFHk68ymWVk64HA5VBE+yRVtZcpFqk+Zs/QufDBiSEwsYleBxK
FEBEWg5A7xkQU+29aGbTqiG5bM2xXdaJbVhvxuBbNQoUEJhIv6ZkvLfs+gwdVpIi
I4J8+faP7KO9pRvuyS4M4AqPLX0qw818xA/LxO7ahhoMOdqxjT0Tidwn/O0ycdzY
WnqOPaytyhoCnZYwbGTM62V3YouBsVyBd1n4tYqyD1aot85jvcxMcHcYnoR0s7wT
hr/XC5iVpBhG4EcYKnuZTW0+iIwBPKXykLQ1bkYps18PsAyprrveryXK+E6mWzM4
0GomHz45ebc1qk5WJVQK08plcPIgxWR3DXINLkJ11olLAYgJ5mK/K/yuvTXr2l+W
jXzPA5ZD/ICYZqqeZmSNw9c9r7/KtgCf8Teu87lgLciECiaK3Kp+Nw7wD2m31Rll
nWm+JApQxsmAah2yWNno0DrssnlwpSltpIP2s7sKXC63AkU/D2+oqM/issCrrGmU
8HSrMegHzVjdcUZYvIUKdRaAetD/pDe3q7N1gull7YmufBOEAatERNueKSDv3hy1
dcFsNDAE05oXcZg+PEG/niksYPCDT5BS99sXcXZfsFYPrQXYBTxlXdu6+kWORoN0
O8Uui0fM8yk2XgeFEDenisZpHBP2bCr6XWJeyO6fj3l5RFzNI9bn5iQxfaY8DEBY
l2b0hvlI3UkY187L4/qppb0okW+GLPmAiCI5O2UIdyAS1RPrx+7TvJbUDYVa61fY
0mIbTh14dILKp4nRUvEgrQD2o/h6r+xUn3mhmO2C1PSiDSxrbvfbm42SRGyUoCOF
FXisUV6VBS3Jmexvze3BUNkwqUhoZ0kacy9giN2TRFkN0siY1kjHjvkUbkYjrn2n
aVy2KdbREBBRWEf1J8hLp1hxiyndqBA+szuxw2o9xhlWJffoqkkiml0xc+XFPMc2
7uksaZ2S85z9plI3mA40wxr2EzP3Ccmr+4MGSdZn5DzN+gB1hsTe2i0AYCaB0DJy
KuzQeX/QmX9QGgpcTmam5gr9opX0CE53/KAP5btlFoEHM7qhYFAg4IxSZOSL5l/e
k5JCns6enoYv/benZ+ZWh8Lm6xT0cHFbBY76d7FGboab+4RNCZPdRBcVvVWKGm22
rQHtj//IzZ7YtTiBJDOTcF0fvOXTfMc3BXw0qcgNsCIfscYw5DUKkkOkrPEb5kIa
NQH5wDDblWD7hLj6E+NHorPi/fP/X7jN+NbAFD7xbVl/PJhIiFT3ahFOQiGoNCvp
cDoNjyWuwjeL8oPCZ5sDjKKHbUEGe+yEkEPQw/Crhc0rZDpaBccm4ErdrDD9+qul
j0qYPNu2ch4qdVjYRHueiQqBh2dlMzo6kMTypjyCH6gXqbWihJBX1OWHh4FCkg0I
761dXp06g5H4cYJijbqbtbh0ncTaFlirfkYaOkR425BFW/Wv2IcsP1WOp1HZ9mUd
nbz2dlRTBi38gwoJszDWGqRdyuG6vR1H6v0277mWgV0nAUwrYDi6/UIo/xWcOIVc
qgNOZoZznQ45SoIlVV+Wl/3ib4dbU8Yip6Wk+hc7KBhZGe5HKJGOHhFM9LrlnDd9
0Nuo8vzasMnc+5ij/thQCMqlTF9A2zm0hcWnPqikjzC7uVcqaatuXcilecb2298X
nbKR2AVM4uugj+2S/PSFvkUTTsXqlOJ1p2AQzxQctNQbf4KL9sq9hbFWzC8XHDJP
kkT4LlQmJFCps20PeZp5fH3lPghKshPBOO8/Gf7xX1bxN3wqfyqEEGf2vXr3qzR8
4mtdQDRpWF17PBJoWsqZ6O7krOBMWSW2nA9zjjoXA9/XFnkFdpGkL4sEM1gNM6Nt
Bqmq0kfe6SN/W+v1YeMfchBIRc/Cr5zHsR5I6CEelDRf8NS505joEjHenC5WSBok
3TmfL5YP7Cmhnteuk6n+Zrn1osN6AkTdgFbN8bphD1OX7fDPR4gu4mktgdiN08Um
2CGU5+FtB0Y+/3f55fk2NQnRPzWFD+49hLm68L2bXtQU+I8wIc6CdnI4NcJTcyRB
uyiDGf8bsXOGfEPqktDJoEyww+O9gWitQyHS15eypv7ndB08fzyYyYux8TTFVvAU
COSsQ+z+vfEebHpMx4is0/Y9bGl5FIp54m8l98aeYwxmfidO9e5Un4+O3SeMW23v
57imvpaYYdqzTmitlt9QBlMcnB6sn9vpfk5WOhjmT62mMaXC4VfqHhT2M0DZsjyL
0be8TLo0mcd4CKTR6M4Eq86VAsY+n5Sgf8CxwL0NXwA808Bx6Wt9IXZ40sNqrOOE
Yfzh1IFcM8MFGudgRKbNmsPZ8rQ5aIam8GGZm3tWC2FKUblsFrBi35tDamritwoX
t/dW8Udq8rardcsWYcjXZS1zRU5OHONJkqzxP3I46Amt/w90TIK86o6wDJcMuX6E
0kS6letRHr0p7Snx4lEJCmt1fDYX2naiVZAbPX/iFtP2C5GkG4m8sIdrND2KYZD6
OjkZfNrlKg8SDncDM3qF7zjCL5adr4FQ8Z8Eq/9YBQtk2IS9ewBopvc561pp1ioO
u3+rHbAEct3uza8zhhGlMpVK80ed8yQcMigMo8CCPjFbD733fD0VHXPOKJypasoG
pMxOQ2EXczqu0VjwfYXS3aEYrOl/HbM9oeehZ5/ve5PSLU924RpFTjc6n1oY6kbg
tn2BDmcQF/aDbslzrSFs6TNNLTYv7KdgRD9kzPP33PyCKNu0ZkUwpzZLFjMymYkW
2lnAsKs1yeB6gNnkJfxn+hTsGrhDdNnQL4afYiTFxCGzr561K20EFcSifrwAmFUj
JhZhfkrKUclj3KW3KeH7KdhWdjYsLSuNn4rI/b8WHsyDnUsmEsZyC5YkRL/l1XOA
nQpTqxO0D8YWPdfEz/50wVukbaGTZNWasrE8uiffwZxRp0kkwhIV7pkw5AL1WgTw
FIBOC4/3BsC1kbXWE4oXHJjz1jS3oM7TSlYRpOq7nhDmevl6ASzPyNoozWmGtyqm
z1J18NYv9U3wl3it30klmlCrhrpVOJVnAobqxP/wpvqbTrEd11bqFzKTF9N//DwO
+TqPrE9I+t4Kpl06oJZed+dtZSaGJCDsekIf5r7uD4Z8An3mfXP/xHOZv4FrTSlP
TMo77Bh8ZSleG99YvCo4wMkzLPbKQtjr4GJAWjHVWG5ofybZC3bFUAE4jLCSW8tH
ebCrbZfAu8uFx3EWE2Ty5gYLL5BkpLhKCd+1eDxOGD2+ET6PtsshiKmlU8jKTbcd
iW4Hxut+zvn7KcO7PI5Paqh+05A3UWxB0ndi64Wh5CogOFunKNpHA+tUaQAmEGv6
Ao5mQjUUgjE2wBRaytgUBXRsLyQ2N5wisVmJJLoGpk02kyxLDouS1i+KPv2ldAd4
9O/iKxA19l/+LFEtbC16HOIHu2i6qgO7KTv5U09bwx2ijSazPHtHhjBaf/+fJ/M0
drzhlt/9JDK2BfO0VpgCftudSR7QQcEoLWZCpsv1Z1YrXqIVttIl2eS7gdRv25vF
0ySKyuobq1yR3J1/zSTZbdewMWE3dLV3XE+DpIRYFJ62SItx8oreYlnhWSsnsywY
nxz6b2yugu3wnZrGhALo8J/SwgiA00XvSwpeJjKR5l6zvCXQoYdZ87pdpLvSSazP
iRNcKTR/n1Q0zwv4xJF7DOFOCh4OOCb9me5yOyg4rp0GtgugV2TjWRot6uEgiTI2
Gabr8ywvl3Ax5JlVN807TWBV40P/GQixMqMFkVK7CKi6XmRmfycItJzB29HZor5Y
xXyP2apUWAi3h00Vvc37ZR/jdK3qO+u5G0kDDo0+776G1zhZ6+7AnsXkAMPX3Cvf
gLSji4omMBuxjGfQZK99tgNOvfH0TQmaeX/HmnLoeXtNdF1V4W8MI6OtvlLYa2w8
tTBdyYLSbIXPT7M698HG4c9uZcarGajLzXAtevIAVNz7ka+GBvpVtK//IvWGbmzZ
7fVLtZcrBeTdJgsbIEQu6IcIxGDdIz/iXeUAfE3vWxj57+whxVc9nQBp+Mk9oSWk
f5nEuIybvCX9eCpTAO5Ym7GS/gLzU6c5qXOX3d9PBN5APlPGAytpRcn+Hak+MnyG
hOOdp+R6gHx/HUuQQyD4iUZez4AC4xUIbhcmWKQ61YGklK4KppVO98x8wErdlK5c
jViKsW6T+F6Jdu4Vc49noe34DAJznKxBP+KtbQAAkTf5k7dm0t/qMCPnyRFKAZTB
FE3+8fkb7GvyRKnjElwOK56rQVSnUn0J/AQULYzvpwoLhHGCQG56Xs8NAJy09e09
9w3k6WXOBfiTH8eGsE50fTni6GdcdyaPOEKYU8j+ACA5iUIEwcoHdK1QM/Vk7PN9
3jGYmOZdvYPH/mCrvIVPqT9/+L3m1BFP6Z0cvwByuvhsQpsj86AaPK+7xLZmCNkW
LIMWR347V0SIkR2pwV3QU/RKqqn8XUGVS9SWHVPNKNiFg4IXNg2a0bo2QtKbwthn
jm1lp0pnw+SUeq4C+uHxsH6TQqnVgP3Pr6sbAX2kB313FtBkS2hpA49T7oO3mp+H
UAzjAytC3q/DSl7urB+L68t9CYdV9II1blGgQ1dMuWna3kO437+88OLkz3fXtYxv
ER4KQ3RwYNf4eJrOWxrmnNXpTGUXbLcqVURH3jy6C7atv7xQoeh95OyrkpR230XZ
aD/GeCcAxeqhUXYaJQWsMP8LUK52XjarDjyNV3+VwvW8YNJuQyAMq2lWqTZCVYdX
Idwrve8eRXZePRmY3DHGJfUDAPkYPSzR7k3TAG5J479rGaFcMIUwBzhNAqILvruh
5OeHJ4TcT0JMs162sOwHKvqrqSnboC/S06HUg5tP6/x8ZsG/V3BzUQp9EoU0ori9
PUFr6MglWPBvnV1b1+Bwbi6yngn81QaLdkfWB63h+/ZXQBppJg1cDWBb4GSBFuTR
uTCc+2mrQkE8S5GnfVV2diSAVweIyzlRH80amjb1vH+h12QpbAPq5EW5jdFWF/8R
LWA7LDW0kZaIMbytQytgk1DXDZuBYYg6d2hcdZpNwwo+NPPC7wAu+LO+dFiowXlq
xRLeM+oeAGywEHTapobM9lyimCUYkf0mIWr+MlKwCZarfzpCmQWgW+frXQWzz1Fo
ygEiaZPFacbDI3eJDYhQmRQCtmcfR94L/gIeqXu+tI5LbhUcaLBN/mODaLnPsE4A
YVde8pdytFAoNvIXXwyae+r0DqKRvRP1rKN6K8D2vZqYiIxwTIHQEH0r/VPNYwvM
mQ4vjc7Okl9gVqXM+IewP7mQTMm8JFkfQLTfzZEnQrUcpY4f4agPbrZgHi0ELR2x
oTJW4wdVVVLaoE9AX5mw7yszzSZDhARw6BWDGsxhKgyGzofcZPsEzmfZa+yDZkh2
mVYHQueS2V5VDs5YfBUIoQ7Jhqsfk2ZRuVnHC50FSgkX94fpeSO1k/wuDhe3vK3s
O5hfSCi71puLVIgZ8ZYQoKH70DH1wGNfxWb8AiZ0c0FepPF9dRb/uaH2xu8tdydH
NUsw3ds3tJ+rJjyuK/FRYjfZ9NlLtqHfymPONrZiVqS5ghh6mwEzpRKQysAf6Jl5
+E1hTlfKNBNnjmoBqnNLaYZ9r6voXRkIZ75q/aBEZk7Bo94mFIQ4v2398j0j4yLX
Y09gjFAt/l2gE7U11SgZxsrzFbOJXloeoh76/rmmI2wMGLH9DTpyadL4k9NWZ15s
4xwlwkcXAAMoTfw9SxSe5G8wWfpRmXmt5FMdFLl2sacRmABhXRgjdfALjpRutt4G
UHs6kyhqAQ+glY5/m8gfUE4IpUDliRgPbIYDp3029I+ymbXY7f6SrIOqtzNaJL8o
SJS4aVONYFIwwAz1UEloLNe5wGk66IK2etJEKOkUpKLzNvY5byloz43SA3ygg1+i
YcwJPrGwqxqpZZZahLa6yu/zkqZ27/TnaeQv/D4wF1tvx9FZFbUVT4EIIpm+U5Bh
riwdZTepSdY2G0KFGqkGEDgQHd9U5eMRg2BxOQ3oV4jnZ2Kb8DJlzSK443og9Oy8
lDsaVuPNhKMDMo4G2tmW08wqWddYdUDWb2hIg6/ZCng44VmX18CL4hGOaPvgFutf
TntaJM2CUJAdgY3/WjBsY7aM5nbd5kiuD9VD9CFfRsUCWERmQsqMS21mLv6qTkAr
5cAJz+rqsYP7usN3Khlto3e3mt/Zk8j/SgQN/DbgtAycBUVITT799u1SwuDR1wzR
bAaBBf9R3BCNyWdPHTLhzfZ5AgO+l5Zf1LDqW9jVBF2wR1AHzoXFyhh++z6a+cbP
mhAgMnQIS5iqF8lHoVwEfAl8qSQqfqIv/+Z4DG+/TkF4rWvTesfVDMyupfMvBiVI
p0Tf+phund7CNwUMmQSA1WLnF/iEY3pfrcF5gJlaSxin2lO/SgSUpzTimEwTEkxE
b17XfMLGlKKsV+iWd6Da9neFK7z14nhE+exBL1uISdcU1pCVuC6SwnAcQzCB+B/c
5b9f1EjNP9tnZFJOgSDglx/gq6OOhaayV2H7orjPuew3fCPbxZ1Ozdyczi2L10b/
2wGBWavjJX+wDpJaHBXabQcjKQCq6fUaQdIMG6UIQhCxZ0hv2o/l12EjYuhzpHPk
anYjhKdk59yDJETrc8eGEOgruyvJJQhxyi34OeWLixcqhZa/XGHg2GcHJKD8IeDT
QWht/oaq53AEhsMH1rYdiZm0VmC0p5POKG2QsEdB1qt4yAOAf/RKdpCLU/tZJpE4
75mFSj27UeNf98S9+rm3xhXr51c25HR6mCpCKnb5M5uhGkIBmzrRIBq6DzUepvvS
rDNcn3qI01hAUNNl8u9pSeRvF2l5oIJSsazJf1WcrbnK54YN4C83ZWhmBHyhWeNY
TTrfNYkcSXNmpq34RDM4PfpZ9cGnaiT2Rft7SOsPc1LPFLTtmlJMDrw1R7gJyZpn
8FOoB71+zHS+l+75lU3bR4ThVz/4QPmXy+Z91iHDYu9gThCxMW4pOQAsJ5UHv9d3
DmZDF25im6KtJUui6k9gwwnGBxNb8roXNGbSgO6/bLTNJS4YngW8f4YcpQTYBpEh
OnwxlGVCrOpHeEUbchGMpxVRrOMSql1js8wqiCcxVxIGHsvyo0rVqonhUFuIRAqu
+9oAw/e5rwpdaHJ61MUKq9sI/5/pEpibnJ2EqZnt+TqqMBxC+cGDqFHhzOnjZFbz
ZajAdErwvioXI6P4UuJlxbDB4yIPOT+WAn2e4IpXZ2L6JuLyW+AFG1Y98VoD2hYR
eea1Ajcq4M+dZyV9hV7UFrSu9sb6SE2ipf3ctrabtsuDXwQVX6q1JtNnBKvVJx69
ORXDypuORTiW6aV9Iw1QWaHBM306bXZud9bERnP4QPhN/M5SSTnooBHLH/tr9JzN
e794xVbditdDjt4rBmkyqutC0YRkMkLQs+gPAjDSucrTPaehP+v53s8gjJ3d+G70
+5KFAr4xZM8wh3RBPMPIMtEMqDQSjijno/PDTeAi6Ya5mtNRZ/FfiTN4TSxnm98I
tYXRF0999AqaEb2/lhQYetPCKaoIwCLt8h/765PBgQ/Wuobm9wTrENkvpGc+9M/c
+RR0kYeS6iPa+1mMu6OoBzXnnZvMjle4ZTCEwZTBxQWBHYpLXaF3inAn0gtdxepG
0J2wy9FR3mAHYOgfRwYFNWg5ks/RXCDPkWPXCl1O+xKoArafEbuaru3ygeDqu6Vt
O9wc72L/hx2CUkntDAXflKO5zgD+fuHV8fDUc4jUUPEEHNDDjJFi8CHOIwHUWVct
h5d2kgrzbpnlALfI++2Uu+s2n4Hu8I+PLXa7m1I4ei/Qh8y8BAQdxtallXlRXp8T
T7fn+cOf7pADyJJUBQz6nZ4feQW70aSXMxALxxnWmvAvnMz81YsbmaDa4YMwpHdg
Y9tJSsHziAPi5EJ+1IqxhkBGfdjI6GJ6FhpI0dye720LHe3icHvgFfv8y1VIGtwI
f5zzZU1Sv2gi2Fjz9BaQ68LHifRMEE9bgg78Ssy7HGhlDrDPxkKzFp4QeKqsvKo9
wGhp2C0yIoLfR3AGPcVdzKegGR9jV1PpAj4CKPZIMFZoVQ3wq56/+6FMby8+qqve
arGLr3ySknoCRQcfNOdAeRzU8+M4W43f5TRoCbBYlQUcWxe87cZlNadEFouBYlhl
qlTe4NzqSybtqo59CHU5SryE/P5RsjtolaQcFJ8UjlOZtpU2pz9kwu9DZ6iIeNZh
EtlsmAaAXcrGZmiVSxqpS4ycoxTvPD+iIzDjqc8zgRIS1FX4OIkN85aQuAR1wdhC
QmgWKYeu7Nm/R6NOhhCLupSDTdijBWy+vlCDtDlqKREBx+Xa0k7pdUySNkgAq5aM
A7BFSb3yr0TfFFP9Av6XOK3IvKbqxw1yo/y3KHfrywW/M3czy/AtlHk50Xkpt3MS
cLAi01ATgxFFt36UC1xoenTF38N87UHvIl9dQMZWTMdqQ10W0nWY+f0GYYNUiAwW
CnReojDpPGVShpjb4b3H4X3A/PV7ChXdVNZL5olfwzPEe53/YlQGULb2nt9wKZLU
ptnPDNMa2GmLhi6jqrtrjz1MmM9ftO4TQwRo/shn5BbnLZ8iWFTjH2E/kq9JsB7T
7l6VUM7zA2MPmpob2kBq+yXwkbXxgOAkmSjwkIc8/oTDJKZ3kHVlIfKQ32oipsJ6
MdNDAjaDBPtrg5MijExNHfJt69cozcqkOe3zHxVLukw+HmWkKe09Y3Ks6kOIl1xq
Za62LkiTt5R17jY4limL91HBTNRYIIVRsQpRa6ULkscsJ3dDmdcHsrtfqXD43DcM
wSxdrWf6Up4dbxx3UqnzO0udWeipfPXUEd4fFxyvrMFRIUc0lEjYODqx21zhl6Ed
VEKHP47ZAB9mz/kAWfueRzPcysG1F2f2GxmOZurKIyR6GGSktjc118kBNDbBx/p9
tnufT1xjX4zc9lVHtHOPDyHzHvvFQk9ortSfo9uttcrrxX07NJf22Us7viDzrtlm
Ak5/f83Vy+f0dHwkUQxqL+X2VTZbcMRPlk88IuV+/lHzatOFrWZSrhvqoZKpTu3X
RwJxRVCgeReHC41tp3MzY+Qo87T8pRQbvgOSbBcmWFxl24/tJGh2d8P5WwqpgFS1
qwEkh1qUeZsu+nFaJuNWjWGsBAm497CPKiCNj6xom4BnViENd46Z9rsZvGTdzmuo
qR/OEiMfFGGjxrSoihuaxiuG2KDyO6JVCu3dxsHafiJBgRh/YQpxnM+/JQePb4zA
ESQaj4PK2gQ1h/Kiyjwcb8A0Pp/Y7EQVCtev17SQ/dgE84ww541O/8ePsP6Isxtv
I851Q1L5olnADOjo3hLawyPc9O/GPgYaWaFCTcR/MrXN/fRBf3sSMVvlGYD4FFuq
GsHARaGbQ9U5RHzIKutUfioERJgJlN9buSHtvkzx6zng8mmMYmHbqzPJhitj3W4y
JgJr1v2vYvhfOgCplhy7oKPVOm3fJofdbXePDyVJ7bFBs6g/ZfZxT0Zk6mGm5kwj
A8r1hvz00qiLLQ9mGr4np9QhqhwFJSICCj4LUJ5Yffqb3/1yRkdhsCnmnQy5/XfM
Ot8fsZgGEpkwtJO2xENwQna+U1T5Gbk4Kb7E+hiiGmgJUDSgK4usRTtk6sH1CT3O
XxyR6k5fT67wzYMCh6QpxDi5VuFv9LMmS8VBbvPsSmceb5EFFlnBL4QPwiEjZc3J
Wiu9dctcBOte5ML2ZGO8AzJt4uXVdMf9+tNygTfX7zTF7V2OWYUT0Nux1BR1yHt2
95m3Vsp97f88U2vC5XBHX54TVgJxe2PATU+QWRyaFngbP1W7nJdZQGDrQKBGAy2u
irzFde9sj9c+g6pdzjyNmwEGx/iZ3mzam1NFLMrfAcdcsyk8SpOYjKReet0ZUCLV
ULS+IDaJ+/BayQFT5TyLnrZAyCgg93rRxA4GyMHs+MUFmkhgD2fbrZtVHMYRk3Az
hOwR+rOX7UnAEoiIVdoAgfJyeqHd7Z7m+Y0AsiTG8FSjI2IAAWBA2Xm2eDDfojJ/
NP8V/hNUCRMI1ofqMduIOL5Uhv8Oan2UP4I5xPFUFTTvghIC9J9XLkK9JsL7c9Lv
s4ye6HA2RQ0FmyN5wvYyL9bb9myCs92/1U6nm0HgmHxO/VSBuPfQ6177EFNZGlgq
QtjK3nvg6r9+Bp1S5XiwTwrQqiUr3BdUNWeIsLzVbA7DpTG83mD72wbwmpbv5A5R
YE3oCIXvYJlQ9MxGpJfM2pBXUpe7Sy9VXuVrbhB66VWEKtTtZIPe7ZmGerk81+G5
qP9xA0O5oNH5Smuwo02F30PnOxhA8cZJwUGaPK5scfA5tV7E1vZLJV7o8qY+nLdQ
NPqIs1PDweXagf8KWVIX2bvLUCctDRpxYLv+6gXQy1nTinqXl/bHNRbvn/ECDJov
8P2AgUfc1M3O0sSh3fqIzItzCk17CRzhou4HEP2FVh27HASb4BtzAgh5USGFYF5D
2Kf+Dgt+22SbQFYoK3j4LHFNpXIK4pqpWopTLV7iKTCVbKuUoSFmSxYscMhPAWT5
vLAKCnSo+gw5jEtq6EHmwmjLTFKRipBnqgwlVuWqts58tTXm9GlUSxp8OyMbEaQr
9RBBPz2TZYY88o86AKbyprODHbqBxP7a86NfbiOyzHt5YWIWpqiGq7biXZr0C4Rt
EH5kwJKKMfQlbV9j6NLFfBcV+og4tDPOg+li1AgBRuYZhU0WotSm0rgV7RIqxYxb
U0hJdsWv3mDI1y3+B5/CWoZNoz/zXRMTelkAns7Q9+9LrLctpfBEg0k36qH6bCn6
AjPf05elB3HGvxB9hx7MsW9kGE8w9Knfgl96zs3r/GTYtqPshwxwipBS6aeiriE5
9WdR76qy9aNcRm+XHqOpfYGxUm9uD4Zs//OVgMtbTTx0peZuWobHTUEBBAgn+U0i
ibSTisOMoGzyxYSlam9/0r6KxUvUi2/8eTS07bX5ztmTp9kSlmZOowGEm6qOdYQw
xS/hhng9u6I24GUWS4D38zJJt0JIJ2ZEg6eeOCNE1HK39PNbHw+3MKBOy2RtQJFk
hI5k1Ri1xH9B3jiHQZpHbT6g2bvFh5Z2K0ZCRSG7dRwQDjJdOFFRkcekxm+y/IyD
QiC7uU3sEBYf8+B3q0BpavfnVjlMOzS71VjfS73llZJAT+GghQcBFAU/Pr7Zx84f
cRrs1xCjhrn3RtT+5EPfYsRVU68TI8KxL5n7DTrMJkSBJzAUKSyqB5lLIAMIsTII
AtU5KCwNJEmrU2MHYTq3KySW29L4CblGFNX15N4lQn139oKBzksXVRI1DOhM8a73
62Wtwh0kmrM/tziPt3zfJNgx6BccOR5NCKLrJDemvpCzh7kAUFavOr3/4cBHVhdl
h0EUPevCHDp5DvEo7mFmjW63jVFf+Ok/WI1g5P+0ZNAcaRgvTLNI9r6Fi3s7C3GD
fVSzvJ71Icfwjck64oKem3eA9R5+1JAzVSHNR8Pqweo+iddVTc6f/agcVfd7jnbL
jHiWurpgKp4iYfMspOj50bfNdjbaLDOBONvZDOFLD9XkX1GKl2GgUIgpq9XuEoCR
0mJF5duM+G3NmJ19AYF2j6HDFNYjXOknZANTatQAL4jIEyFPQblbdpH9rw3SiOnQ
/ZgIJzU1zWuoWc0YFsNqskyOZJc5P9lBCN1dlF8c0QCkcm03ssAXaItzSDpL5IAP
QJ7k2j7ey6eO6WZuhAt3A65KNrMafDbwLyApioca6Zk/l4utqu83dSCGUe4nOLcA
FhNqlOEt5IbQzvA+oTTmdJOJRk9nvF+q3+nG2mLtYPoX5YnFasyw5D7aOCSe+m0B
PZMO6UasOToAwWmNJYb1QNEeRNvAKn70x5WJZN1XqXh4eT19N4EMWuveYrtUOT/W
1bfePuJmSjRZTBefb9NMoIaQD/IBj2Nl34RItkzvIONgo7WZDVpPOGkUZ24Qc+Z0
lVhfwa2vpa2wTf2SOylccbcCD8wTfWL36uUK6BvbZ//6nPTCTPHR9sV1jT26lZr9
sNk5Y6D/LD280Kc/1dntz1rd45fcWeG7b3R33CsSrisUh5gHZidHrptTRZmPapXN
7CRj7jJESOY7GT8JAyBgHRfat9G5JV/iY5RlLeGD7E6W5T2N48mekWUOsifiFySE
VGhCKsuNVljG5EzJoBjIgGNz5Tra+BKXCpJ2JtVfv2xyeNHXdG7oezxbfc6Z16Io
GyO7ecOC8SYr8LUcyof/RA==
--pragma protect end_data_block
--pragma protect digest_block
auUsyFvZclSGXYbGFVi7QWwX1Tc=
--pragma protect end_digest_block
--pragma protect end_protected
