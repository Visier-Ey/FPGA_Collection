-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
--pragma protect begin_protected
--pragma protect encrypt_agent="NCPROTECT"
--pragma protect encrypt_agent_info="Encrypted using API"
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
--pragma protect key_method=RSA
--pragma protect key_block
J9Rr/ksP1hzZ4yWnkgmFZu86K3kuLVAaZmjJ7KkSgj1ADamSg7epJW8ZDaQ4TkWv
hDgec/67Ygeda7oU4iNYwWIN4agRTogS6va0T9KoZZIKly39YpGp6lztcj6SA77o
dhe4coV41oUCyGAqs5aRYwPFrV/xoVNhNnmBLDdtCEz9gyAR0SNQEJT+sBBElpBB
bwUSNV9TEWzmeDawSr8C2xiFw59bgi7BFVJNshlu9hZ57uGzyW36ofw4qQWzuerm
1kk5XtFG9uRzOG5dplNzpmgggufgTPMx6iQ1DoSNH38/9OPvs9JH0ZmZ9semBeY6
nXxuXjs1LqYwplTPsDwiEw==
--pragma protect end_key_block
--pragma protect digest_block
o5igGm8SBFSz/EhEHE2lGzY5zS0=
--pragma protect end_digest_block
--pragma protect data_block
6vPQ2q7ZPDs7fQfEkA47SyvcQChGdxhqvp4BmfR0Bn17V2+5eMNXxUqMeyLCgZTg
CA4n1QBbGjjfwJEU/nhsr8bz7yVeMgEBUlCRvH0RKCsPmlFOevTU0/qBAT5rkEYE
RXBZ41t/dS5ppV7MTnFApwVB8/eF5fr1ZXFNS3i8StDWSjzH2h4gEj5dO9wxpa8o
ZQgQvWx8JUwjCRv/o3HITcC7rq+WNNxvQf9BpA2f3YP3T44echvOA8ahO8rC8fdv
WEIl6oRXOcjaRZZZORPKz4RhKRiz+mNzxg7Hd3Et8bhU2wBRD0934DWlb5kS6j0F
wz+PNSlnVt96J7AzkYF/Uc8TykF9fLf7wqAi2XZwLex7hDhig/hsv97ZARlcqWJ9
H/S5ksVDIHbqSRlUSDao4GCMN2kxPMdZEyF50IxR27PHGq9ZgHcrqBGolg0UsiJ/
xEdZ/xD1uuak23JnrDsm5ZrU/WT0SQKay1uheSt8ZRJ9D5D0ImMutj/EIP0MU+rb
0S+V4k1sWN51ZipG4k94bkoykZra/E+U1iDrI23qemlJRwg8SVdmXZAvn5PW1vML
yt3xby4Czv/rWg137A17pkXHY/HUJarX3oM8Q3IgveBkjqmai2R19LaUYJ2MYVDj
5pOaz1y4veyfo5jh156UqMLT7v5Ub/G/67pZgdOsItzy3heuwjdzRjkWvPVrQqXS
3jHlawxGnEsmKhvYA+GgQ1LcXuR7YRYSwUGEfZrJTLv0EHyI+sfEp2i6DcRQg41L
UUtkQa3tIjLY3EBGahwsiHOq2UFvBuv0IYS1r4BfMk9u6FLTuQ+5Qv8Ij1hITkA6
8kXSSlW8n/Zuik/ajnd86AJxEt2znQXdj6e9X3f2XWwwHYYf4j4JGDcsgRHcM4L9
Jx0oveQR1zfv0cA/dkVBzcZ9m5iNykPf1GBSShpAgwhzDDIsy/dfZGZK81xIRaW+
hx9QgBTWZw+LHXdRs3FYRShbFZQm0AXevhOAX8f5EZs6V1NoyogPBHVS1a0UM1OW
uMnOFZxW+Hnbc1kZwoE5ZmpzxpauYHnaSQFMnUVDk0qPN1GfqrIbhI/URjbpLf9i
Yv0tlQDcTFT17c+gedqApFJXx3tKpPJjpxAqYPfQzVohcWGz3q7D8zFL0AAynIoK
c2y3oaD8C4MKUz3sQuy1sJZUTC6yacb68JXAaMQE/fsKkixNOHkah0eh+9+/hWu7
uLrlZXNQL5+UN/Vz++9ingfMXFzcQmr+rQIBPhVUX+IQ5fXvnEd7hgurhenjx6A6
FWG7vT+1R9Cmgm+1iRiHl+HY6W31oQ8bORalzjSTPaDjaKqjiGnUpufhjKufObHP
rtrFPkXaIfABGSMK3nn60bhv68JtzTle/aISIeSHToJY7VOASYJ0RmKX2ymNqNb0
91MYfCBXu5UrRKkyUcAiolxL887QD8te2DZ4w2qVoSn2DpckTHDHPSlpbBE58D8V
mv/RvL1O7CUvr9vtU/z46dz2PgQHhKMssZjpEVQ8MCAZMnw42WKHOAgI1ZtuPdy4
54185+toLgX+GpUd0ATM32+BvehIcpJy8Axtevx3Zkf8KJcVF72acC/LYbYxJIXi
EjFCHJverzfnfmf1JpIXJQByPBjShOR3w7iva+fZExD/DMuU47FJp/pO1FlBdTjt
FG8kH7Qq6m3kEEG72AMYbqNmgmmYmrr5yDfrmo+oLM1h2TUB6foY0a7Vpp1zAnxT
d8GqXG63jrCAVWzamC7oPw1wjQ7sCcbOQisWIwDQZPeMPsU2WHiSlihXyDcFq7Gl
6pl4Jyhr/XZLyFzM0VO15qxkgz6RLNeA0TfddeqtkNkT5dMWUqvSlQwvoGkrfhQo
KtxCbhplYNdsHGMI2pBH/VCQ7LKCFFbf8NojSV6lagPNJOgj6u9hIQUzRC1rVIqZ
7+gK8T6VQndD3i/LpmDX+xKnT9exlQLXcEe8KTo4gYXlpzWLIDiV2X7NGS81ox9a
WZrR5QhxTuCpPnnr1cgW5x+YeurNv1yKWrTEqAiaDiORXT1JZagWtRN6EmvVMovl
gR9xG9k8jr7+TIBaC1xOZ8OhmN8iWRXsx008vSfEfpfbfHUIN/MlXz9zbok6qXUO
MMISaFZ1No9OJR2yVmY87RRBlh3ZKySo5joPNaeghEdeW9DWs65yZibsnl+vSVDr
bJ1iCcksx0lUIrYC4dHTbupLfEYci537zC4E/Oukoqm8RtsgdzjLKIPXGwTgMxzT
lmd900Xmq4dsdlxHcKt1r71D3KplHmm64k/V3uyaYTdVw5lYqQhpooeGR5/MHInM
YQBuugXJ1SPJNnhNpRlUMeEd0899KU4cBb3JReqrqV2Eq96SfYC5wc0LF9V+DWaG
cAEnsHxBEt+7fiG2gg7yYev72EiRWtVk5PsEv5oQbycQtCCh2xevMcb/8Qhuf9Bd
yWaia9GhoUbe7ZJFREBtAplSnetQKuvWhIPo7WFv0UlZPH37LVsrMIJTx77gyh8M
RTocSFNs0nbF5Xk8i4pA8U5T4Kolvqv9afzOFhkzWwaM/W31xlxZ3jeCuP7Md7UQ
KZtIJvs0o4vugSC9V3xm1gGfLyUjqvuGVt3dbudx3/EGUATBJw6v5iWLu9DDZ0Bu
ELV+MLdYxCxcRSWM5Dqxyg4NKOZasBXhnMA3k68WHAaMRHOevpbCdugubUuTa8/X
c4Z92H0sgqFGzcwSaJ9uo6lhkKTVZpD0R2qPtfVMOZLuE5jf57UAs8rKcC14gF7m
c0QC2WB/ieXn7bPRwSxGDxc4UX0mPE0VLU76NtNBz/3Syk5+qJz6+xsjJ7EihMnM
nCNqeeUTdtnetwuRqSjw75XHkJx1cxjSZtVE2K3Zr1+I/YZkHBGojqHoEe5S3wbD
q3O1hBJVajPoIWCHQY65raH+TbeV0b8gCQWkEeOyqTmKCfjWZFfQdcPoEzn/PGFG
fEuPTN43u027YxstUt1EkWaWnokkQ6zvoLifPvkaWkV7Tj659B1h43P3Qb5qZuxj
aChWx+4TE/VG4Poo8OWfEFpugtUbc8slMkA9ScQBl4wGlsNqvKThnPzGIyhg4Hxz
on2tT0NSTb7J2yNOKivk1n+As86W3qbVMU3a/GHblCOuVpuT3E9ApfnJZ2k1xBq3
UtGhEQyKPHJNZftOu/xNzqYeliSoPHq6MgCjRPsAhOJ1Y7R1IvrX328Mg1l64Qlw
Bs5Qdvcu8ATXhSlRn00qZyvD7zQkrZkeKi6VO1SfPhE2pT3Kadz2sDO/JDv/0Xdd
gJxYVo1NGlc3dsrPZRW6d2wiVo4pVfuogAo/E+5TbGzimQvfJIfezBy/JuddV9TX
rWMopo1FjlGgfC5ca2Yz1VLs/02j6kaKQ9ttxBSWWQISZ/eCDlvGaorT5aP0QFvW
GQBGxv0Kujr7kugIsd6YPFCn7FYIyTq3uYJGQXGbAFLAo2xsB295TBYbRXk5haJM
gSc4pbYm549e0Ur3+kXGRhix3oZebtFzNQ2/efXzykkMyaSkQTFr2oLdijC8Lef7
WPao/AmguqPQDocYJ5Adhd/4zinzQe4ymIkGfrlOJhCaD1SPgHev7cX/+2yvdny6
XbSKra2zDGUGQg2k3XIyhyvGARtkMbymKp075wWuJQk0dwb+GBUDpjiZlQbWvtM/
WudVi2Bpg+D98w1hwUhAlcyLGx1nnKJPdW/r4iqe4KmSFMNlj8yHaWJw6onG+oWc
o7pXMo4OxAwScpq4L2r0J6jxfDwVITbVuFI+HHzaEMDj5CzfG04HSsumPSeC5XfB
+ih5yzrsCHZrB+kN/y0LaXZiAC8thHF4hWZVELUUPUPKFPw9ohGYx0Y7/AkSZxa+
GWNPtcTLt2244NbGIu5hCR6AMjT/73EawqHixaIqRN0okDmMLe4gU9WOaP84uXyA
TBxUel4rOHoDu1SNa6Y64zYYewQeQLLnmaVDyltSc38CVyMAPQ9wzz05AmMh7Rva
e+oUnnHQnqwCASWPd/lLXH5Ifza+JCZjn4aNvbLlUoPeZbiTJlBj/zNlLoZbwYG3
H+Vwf2gW0YGgdxozq/36kBlZvd7T+EmAyXHE/88TZkiOPxcOhNW2roOffbcrraAj
dEeIfmUDI9l8X2C6kzAErgvn1JS5FxiTO35VhMjDpXA2uBMsHGXOW780QxkGNoBX
2bhxk1FJiCfUhevAyzInd1GYgNS72SGkV77a9FDAkSAb2VJ2Mcp2WPXbyyWTHbFM
HB9Wtxvum3cIbwWeu+vJyoS29l8E4OP95oG3CNproo+OkIX37OljuAoPzDn2QddP
ZjYtOQU8MeMCeTOtMvhaz9Bb4Xq4HmsLmOim8murg00cIHH00Zdim8pa3Eee3hMb
WtfJEnljy/oiIJM2sXldGpPGDblyFAV9Lhk1d/U6j1uM8ATYbciTFGi3twZ40cDr
5EDfKuAGsr2vHVYKOyiV3Hrtr3RXUnl4bs4Efk0p+tFaj6XDvVJDP6rzoJrj1zU2
idVq38iC82sO+rPJgTX7AeyUqs5l9QT64131MNdIRSAmAzqEnH/LbjCoTh20GHBZ
FlS85Sg2lTZVwapdISeCZVI7Z6RSbmUY3P4enD8LsDnYVQu1MmZZ3EHHNC0RTX4C
OU2NUAUlhBaLReZLoOR7Y4cfWvKLH1mNlJP0SLiJ78nhevPkwEN7IQhQrdwkdf5W
V/ECd+DqH1fNF5pRG8f36A3PPrB/gMLsfflLZgKqpKYb8a70On3QGyGk47rBwVWN
kgxI0r+jtGkYSYl/nBjP46A4guAdoi5G3aIDfXEko0aLw80zYixwIfWgYU7n0GCV
liBMlg/1FkuL4QyRhyNHz1hCexfL12m+aLQ+/NPLVU6GuGSV3rBxFCkFPDqqBQE6
VjM6fohtcZ4yRc96A9n8XCUN4KFVPc32pQx7qZGLN6GvJC5zyQhxY2dDJsBm4jI1
wjdqU7uGzb34j/6EOdXy/9SuKLnC72z0/Out4tOK24CfTesUaGzeT6oGH9whRYPi
2Ur4uTp5eJiDPvX3PLnBu+Y+4FJBdK0iKAf102qakKBKHLiIVUgeKNyajm4r4SUC
lBP49TyfMdirLv9BWRHmt1PTJyUzeoDXtorVaue5iYWk2hR/mK0K9w1PPWt4NaQ+
1K52Q6PPuYTsavWnguM4jOdXJsxwCHg0EfLAeZ5oMqHdVdSI8up6LnKklNj5ye3v
dpVUkGHndON2k5KOTHKH8w/TdUg8smj85YfuqnSZwLWmIqqhgS3AtYnH4hSSH7kg
qA5pjH0hcFX2ihsEfIkHRYjjjpeFyCNYxxghX/Q4vw6vWSmyPtRvMm9L1ktMabJA
Mmt0J6jEN6FswLBBP5nMitvzly90xPmm50x/EAOL5b8bpjv577tX0nNST8Og51el
u2brYFjJDK3TfRT5tic81v4It7Ch9LqRe81urqZGTiKEbfgybMqjxVsCGgEbJ9VV
tw4521xsZ53UdgEBo9YDrkudEkMGjElgPJOkAcC7PFjLBCmBth23QMnX7d6iLmAj
gLoy62SiclvjrYQa7WnTfLf9qT/03nb6fA/97+SKsS3wecwZuXShEpKZAimZPPwH
h/V/7+EXwPOuVfSZo2khy7T+8fTDxfQyIg6/yAGiW1R0lUj/zLFXb0oESmGsxIcE
E4dBAUPt0GQfy4HqgF86OH3PE5ctxwaax4r3qGuX86zHBEAFPLt7kgSXsUTgmg3z
iTpgtSdJOBkeRdRWPRsFTLfLjn8Xo2QPoXHZbnWbXAGUueacGyh7KOzlblvLpv1r
xDIvvdFktqM09M+EoPFoRawuDkbjgOC74c3Rqu487wiWM6e4J0bCFBnZxiB5xZWw
j2SCQLwV/h6CVS0vtS/hmz6SGctWanhHlwWwE/BmIbR5FWQtqnDFjbg1Gi99r4Zp
yKu/mCvN+ztoUdZZkXKumFXpk2vlQuB96+cyXcjxKoXuVVoj788pQExFdeUykkJj
GSjpq4Z0IB5BK91+1256k9/22SSel2aa7+sU3Q3GAOmWP+R+nN4DNR2DqcAHn/5q
kCykK4TEgEfCmTRV7y9TpJK+YZMqN0woVbbbVx2ivZauYx4p8mFk6bq+GLwIA12u
Jwb0JytlEZhhplBFH+KMlMcpNqnnOYS4qiKksFUNyLzziR8/7GYBgykpz05w71jr
sqwzc5anIbbph0Bacds5c33XJgMfFpI1teOR0RjAwKEBayWGQfusBnFjb2hngL2X
CdWXTBkkFoJvP51OE0ERuF2T+TQaDJfy1qDavlILHO9hcrtl8tI9Onic1FcKPFgk
WlYBfMpd48FZRHxHdzU8d/d1nqDxWzfp55JzxqkPVnkH0abVVF5/p4dwecn6cr4u
JLSxJwQ8McZYb9354rVVIj5/Gy3uETDrtgyfOcFdYU6UWk9dHa0jcO2+eYBW56hF
uxl9BwsCMwfqV6ba5WP99Kkd0/QGqMqvmCBT5QEea97kn8uMjkckMTPfhqvB+gYg
No+P5U1HNHEADz4giTWxkzKm7D+fVQpP1ppmZGL9w0imxXPoCADp6PUXER3gjGIO
JQL5MTw1VpFPWtNqpHVYXf4h7rgif04TxiURDkX4siMFTEXTLOCymCtEIjM+2NCM
Wwtbt92plZIzUZuQ/TPSfIdNqD3HIl906/TYTnElf008OMvfQ6ReX7H/Ie+8KUBn
P/tFWRPzrQWqajJk3ZvhZzTmjh+jAQ0kQEM+0XNFCvHch8ayELi3z/RhzTXRYJ91
fRx35lgvy664+Ix9dOVWoaaTzToaAN4Agn2y21hbIHo28PMfkrGqHCI3U9/4dkGl
0hozW9UPEW0fgnXtZcWHAQrWcaV5bD+O8Uk/Hq0WeuLHgUasdtA/p+9J2jc0pLQX
U/18hxm6HxgnTzkz2DfJVbP12cfNYzptQROjq9AdTIjV3z025qGDyQR1YcoVw6kU
wMdftoiQ06dhLXutkUg6TJlIxzeJs1I3peDLtReEvdd1KIK72k3qfcpOWoD/HEh+
o3psAp1Ch0SEKKXnt1gvjQ6V/0HDF1BZ+A/B9+eG0eofk4BYpVEiwsglQPjRldvJ
mp0pZKdXOn/itdwqCplSQ+dZZXOI650O7exR+cXWfeSjWhsqpSqRqlt7pS+h9mgu
ktbgv6Lgk5uQPAFLpnEaRikv6kHIPw+8CNWDGnct3DU97HMUaYgis79RyyYSItFN
SVHu8vLoyZIVylMXcvO0oZN5S+5UoqtD3gGUh2L6TdQq+Dkjfsw+w62+pZKoXhNF
wBfxA4Xmk8Lph1nXXAiAo4saPV4Twv7qZKYL2fktiJJ4f5n/VvaZIqFngiWazGaE
/DLc0AEeXElVxaZSaTEa+ndKpKPuK4TuudVY27UUk/AicvI3yG/gLL9B+evkISGa
s+Khg4bwp4+jU1rqFk4U55vnj82EU97UZN4SmaTfcUwUKVo7hl5FaQSn7h6yVgTI
MGo2qtbuHFB3XVsmkVoWA7mEa+PaLGfCfNj8Gs/ILrWZirkTdFC5Pp5xGsJ2+syA
yIVjYW/Ow+IuKU+LMvpYOIhRLM0cXqTTnu7Z+bzCVb1UFD7DZFhyUbNJhzfqVtqT
B8Upo5N/6FFzWd5622tNvURsVZGwyrnAgZs+tJsc+h6Z345eEwQhpla8gbYjwZYf
ErMOI35OAdAq1dEoe7oxSH+yxKWKvn/dmQLzq9FxxidxHt+QLG1l7n3GSkGs6sWK
Ry3qj0fNKE0ei4cP69M5slPpapUg3y+CkkHtdXonkgPJRrTVIrwMTxK4HzPumFcO
uJW5mTK8WZFuR3BfbEPnP4uq1l2ZfUxTxqUQGrZ6zPZZLi1mKVbOoghlOx5RgkRL
9JiGOM8CJcfPsMhv7paGk2m3T0K7aP3DSEHjWq66Mc4rEmz1UWE7Ppfsrlj4Qrm/
zY9ah3p02HOac+bYeKWiMucGalp+ifjOtGNWjaBgsuN2Jifu0jdKa9NZrbezyhaa
zgNG33IFrFcTL4OgJhfCHPLpxpcnDMp5krBw+Cj276qNuLUbptyT9OM71M9yzfAK
HL8d++zw3ILrL/H6UzB4BcMAY8mt9oapWbr7hvSrvyW1T9LkpS4B1pGbG2vrEVHQ
qCPqW4jcVIFFPw+fn3TnSpiX2Ok4lndOwtOLDndYuPn2A+w3Nm8X8PcrbTwkV7V9
BA/Bcwe8tGlfN4aOGAHMQDItvAMiBxAPXOGwODas/+7wfB/NpNrD1taedp0WH6hs
tl45QlASN/0T642JMjdF23nOiVFVd4FJ+mkYw1xLkwFCSF6WvlcdM2D7vQoLLns6
JYrf57t/4iuJLzOEYIEouy/0fv3B5mT2wRskClHqcSbeuf4OHdNIvb/tfqFKjrfK
Ytgo84SAlbC0sKom9UmC4/KVO8aX3pBG31fgDz//7ckhoI7xc/7EKiwJ9LzeZ4+p
jc41DYP+N+s1/eqxniTN64KYfnTBMMFyAH1bnjEuRtmXDDf45q7U8ytl3rIvk/BL
+JE4nFV7DXdoAYgM69d/so1zaHw3AGAh3vJSHg+RqbzQ8C+nwAoj1/qRat/eJ4yA
hoSgUUtAJAd9f9k6qudaq+0AR2lu+MQyk+azDMjVYsZ9WVIBebp4Feck8M++HW8Y
k9qNpsk3Csj2BU3Byd0LAsmapXW9kWc98LA3sg8JGix8e6UWMMPcSsaA8yqMrahT
s6uiIW7LinrLsl+LWpG5CPM2pW7MSKR2PECWZyscsb/Nk/UwKfeAq3T+ooLrGVAK
oCy0HYmZxkEnFbbKSmrL7HJIbnzVA46wgMK+/zlx19DdGcKEmZIRLV2JjXXps1Zc
tRPJq/Ksa6UjSfH59ImM8lb/sB1Huj6YQm8tCmeIpMiZlt3G4O0ZaKp3NkRF4ewq
Ozv1gfzBLWVpYXjd4PeC/stwUlcBaDrTdvQxNLMuuSvSMknq5dmOL52Aty/fUkF7
9vXAUYt51GKMucFfdktoPg5JsKCgukqcSHFXVZdl/pslfBrXf5GeS05NOQHCHkr8
EWuZsnSiIR4m2Ekt+WyTqxEjnsgicHjwEs7MGXoLsDX2781kYmIl0K74EUU7RhTc
042B0EECoA1CQ1283+dyyxc/FYDDwbPVjUQRS0PPzFtFLdTdLvQ9uNg5+/mLzSwV
fKpyxFrxjobcEyXHwabYYzpI/O+t/HHJfFokJ6MYwT6EJllqaVLXeTLF8zm0sNVp
U2nWAxL4yn0LDfCm6LuaAA8uN/pgAEH1KGMZsPO3rvoH3t5qcWthcmuh+ZMd3mnc
YhZH/nY7yMKj2/rnOK471yHKu+Gq3yC5/oox96d5X7mP6dcC07nwAmJ1rGuThaGv
mKDPmO2TvnVsQkqRkaeLTBwFWciaLbF1FwQJcCr2afYpwhJbYOWJ2xmXt9jPCB4d
oWJHBSvssMvAml+PMqZxgw73cHdyBq97w7AAq50J4gVX43lY+bfRtXAasuzEQZJB
zOy1scASL/Er3m0RzphevdAvahuOjZqbFlEz30fQ8q0ThfAbArqTK91da7A4DRdE
ZzLvKY5bqNR+MlHtrFm/he7gG5PF8B6TgzS3gf6mPIWmSCC8bW+gzrVppYSSRTtd
wQlHd9G4O1XIHn3YtPGamvD3g7IgI5wgb8beKoM26CJsIsXGRAH855j8Wgr1yShl
PHUCtuW/Myh1CjGb3buODe2e3g7hoBGaDsGZTQjeHXsTEOT8NZC17tW2It5uy1Id
cPCNYy/KT+11sGxcK0YF6/ae3zOgk18l8+cLy+GllQxDSAQKDpElVI9p1FY7PxS+
TUMfnmIs4J23PABmH712k0fm/TdS19IxIMUE6zZxXQn5viWIqKcIkXCg2k9hsyiv
960wYcdrW6KPfQF4yBrpDiiC8Hg4itGgMtwIEdPBCXUDcoQWTwx15p5WSXnesTAe
1GwDSQOS5IePUldFOU0hE2/DIH30EnZuj5sfzVQUbr2GQP0pUf8g3ISMgMfH7QOD
B244ZunLilQW4No9Esi7GGW1f1QHcggWUFEeRD9sJkOcJRBr/zgMCMB4s3JgmOSp
v2nYIW1MNFQHtGfySD2N9yHgcfNuLZy2F7qCmh6HrqCCIWJ/8A3h9XHdp4ChoZgq
N1jqv7jRQ9mAtNF4Ijf2T2odZNZBFiPSuUL7dfJXVyzGDhQPsNVUCHR9KH8pq7MF
YGxDiHKYCI7vPM6zVmaffAZfeBx8Uk5fIMBe6hpsQD+b/Q0IGwUVuOddrJ3aXvWi
96N27hMDPm+GxNop/L11YaUexOWg5m6SIbVQ2RYmELVgGn+9exYAgaqDfv8EngkD
imrM2Zz39mYFt2EZspQnGwTInEyFVwCXm50sXFBDanhH6NAAC6yBBoXy2lHMzEYS
vI3/EJRMwr5Jc9D15ZJQoifohxrUuymMUHzMfrjuV54rrRHy8JbfWPit9oT0PKxn
sRQTGSm3Tl+VNXOhTVHn7Ual7unD4ljUoGYa2rrmDlZMyHSMruvWH5GJHN5JZQkD
3QbgSDbPqsUfvFIA36WRwoboTeJNEbTbK7lbNf1bMA99gJ659rr+ACe/Eewd8ugX
VyOlcI5Axvc/hPFqcXs4OsNbAHiUu3mx10YNJqqHxwRdoqxvcMJaQGgabAmnUtWk
nHOvfhK5ZBEiJAp67jvocOrc6B/qeiUnxvZMUzHSW8Yxk1IvzpPJK2BKRKor+vSt
dG9z6iOCf2uVvlauJBhzgAJP0eaBXJUBSmdHc71lW2Q7Hx8n3v3A+rhtFBa8ScI9
McF6/d721yInMQracKKWyIusGghIvkL4e9JutsskZAvijaH6T3KFyYNMQe2K3Q6t
e6wCthBZtKl6SXGuBvuqve/dcy6e11BFcw1fIubX52oDqXwl4y29xMWl1BOgEuog
wwx7G/wrEp9/Qa3E5or7yZ9oHcFoUH5h2vYIDRifiAgYaielVyEo10bLXXyi2QIx
LJppZ8vZSm56ERJfs96n/GV0ol8Qgu7l0Nt1lFSXbhTevKPGUo4OrPaMSkhOpjdc
33Of94Ulblp3yUN75n0oBXEvcuGS9OIVN2uxEbduEoNfAoy6wi0MKjH3w8SY4OZ8
LGdKV6+e3p7zozS7A4DdMGyb4g5Qu7k31VpMQLr8hebOP6xAnhoixNZSADOK+kOk
t3zWKknWI1A/dunsA4N3kpY7nRrxycRB7NB5W+d7HAFehRMxQyJCqfA0hfcPbjuT
6dkdYkvIXp7GbVv1Y08Qh3fpKEfLUyc0r01k/2SKkNMVVf47mc3AGRnShl62Cnkb
s0HTSMl8l8XbVwqIhHXTLPlYa16AKMnsnVsa50ZVGPMHDBHM0JchgewOXVamJ58/
v8ucq1MaPrrIz29PXoP8w6aKnkCwuEArx+O1pmkVD9C8gJ05JlWOn6zgxdd1nnD3
6Hq+TiV6xVtL0uh66ke55IARsjKXzo6FtJUE4ELgztpe9fjoxaqJkQhTFJTSack3
TIVUiVG7cN6Ovyt9Gf6/3bmNj/PVdJZqUAUGxyfXQrt4EkRA7DVR5njbiwpDFChH
zjMmXRpnhomin5Xqe4d85kOchLF8e4Nnwr06969vNOFNCCyewop6Zc/qQgm+Mv6+
XdQzS7aM6VUT48FGt7WhkVI1bn+vtaj0U8FlwlqLAAMKxORY2vaP79MzDnLHs3W+
V85edr6MGCeSl6aaRKUWyHLWwZ/fM2euu2vxmyFGlHWO5IL9q5FqxyhwCz+Qr4Bt
eULcEuCxAG6dMSRPPEgr90KPBkKQUx8/P6hmV0q1p4Bx+Dt79w4+zzZTWaqRdmj5
1XKW/rTu6hSxGIZ1L2ZONnrN30YWUlz3prhFalNhIS5THLoelIt1Oy65ZLswMYjS
51HZVr803bHbylOzKnb96oi6ORjRBjh5VZNCWOQ2erE0pKtjDCxCL+SR2MIm3FVK
nSyG9iPtJYFwBXu4G17uhwM7BlZeb7al9KWNzasMFH0UfzaUGMIOgF3/uGEyVimG
eLphPSdVfZ4vKS9YMhkOL82AYsjWdmtXVc2keKUucwo9X06dK3gByIBeinIA73v9
VtQ+v3HXkDC9S58+cMMR5boq+bgJzmKsav6UXpTTQ0rHcryaOmuam85ZPG8oEZvt
4+uf3afVll3sHUsqA2W/E7f99q410iX5qY/xwqlRwZZUl57npRrk8o3KMjogWxLe
52SeH0ge7rRUcDyqoYe2l2evcN9DzGmGuS6+VYd4HLmRv8v5K/2X/EQgQ4o3w1aA
LTuZ+ZuVo8aqrhhvPe+4vOFXYINK7q0kInjxYCFbDhDdsK4SyoqKxWU1auGpCDPu
1eqQAIAMmRCKecNKTlox2xQr4Wp7XFYHxjeJAJIz7C+ygzTVgLZl5ZHm9VtFrEOM
5fDt0jTC9TmdVDf7mFhSay1xC8ds8BpD9EYQSnib6rwkLzrYaAyuGaEw/VCr5Ceo
njlG9lV6Pnda4hu5koa7tBfho+mcPlIIrq1EPCt1gdtX9Uo6leIC9RSHasYCrQpJ
wCa6q53RxKkRRjSBmG/Xnjvvf6qqv961lV1yKG2/0heyTXmNLbp9/4dgbbl046gU
8WkHsk6+SCrbgscM82YE7UJQMjhwPRiGXvLR+4f0AYo8dqJvP06n0iaEykRbMCOF
Rdr+SxSlmGvodM6HsyQTehsOoUHXJv7wHjjg/8pL2j2fRQEWYQCKYOUwFgwacXk2
q17rRXLLHSpTGhLwTujWPpeyQ/G3/hd8Pcafk+Pmb1HBMF8GwBSjjvN1QNOr1EVw
TcRrN2W/bLBRjXmYkIiY8HmEBfYQNTGmyjU9tlnDUaWG6j0K8GkfdepzHbtcRur9
ppHq8tKNOArzHO09VBBosocCz6JNEputt7+4aeK5x0owEvJM6lcVUr9W4Fv1hTGQ
RW1Saqbr4cvq5FjLCkjJIkI1P4nlH44d5CgP1Jsw7E77JR97m7WTLmKcyyLNy8JA
Z2OMXIhWuIXaYhlrKTF/cwgJMjGg7sUpgV7B1pPSVe0YVTNBT/iTnU0CM0sMSMCx
A6o8lM+L92ckW6RVtjvgb/U5GlYn0JPG23KhO7K77J6IivHM9l3B4od61u4YJEY2
iVW4r41LAQBP3RiV+I4eosI/q78RnA1r4r/6TePUHz+c3NUshljXKqlhpRXzJrJV
xyDyrAbCQJYM7lCrYyOS0HZZswB9Y01IOPnmZ4QKsb0MFSnghZNO+eiC2HsymgNk
5qixCAWuTb5nc6ewn3cKjzhibvA/GJ+FP4Ku+WoNKkZpmRAmg5kxNXI6zNpJ2tJm
dweJDZgCRkZdkHBQCt9gbDhPUlz098Je0oROx77M9S0oWdWySINvtbPraR8IECaI
TYz8QZ90XfsujJvF5Z8NRnlywttC9bX75xMWRFj+fInapxWLdDAPApOmmlXDGAaK
4dOr6ib5EeL5GSzMF/n27rosk3jTF/0wL8GVqdpxRjEyq/0YOiOrsIk9XQXPNQBe
X0Hr1CTB1qPHpFrGLiUgyiL8gRODXEes7vf5oGDTedCusQ8ALhFjC+ZDa2poZtIz
qkFRFsu8HZbOogXQAByoqnxYSYsqK6lc/3VypXxdzNdqYU3jlD64PjwikRrF4DOO
u9BapDVwE/Tdb+HZbZBh8oHRaGth50/mqQ9danbwtkXz4aze8NcYlUBmJXwmGn/U
W58lgnXDjnbNQhRNB0tNwZujDli4V8Znb/MnCAblAfXlH0zTURPJqGYPDEfuLOf2
iF96/oZdG8wzMuZ2IOSo1DaaZk9FU295u8R/1yZYA3P3DZLxO8K+ZiFEaZkoUmM/
V+lWnSTXZyu0TGQaTZOEd/ypyMDWxN28Cs+irwuAS6P+9pDsy8bdfsAu12phieU+
1xe1JTTWcsqZfPVwB6g6tHfI5h7eeX3DMCrJ7XYLbPZmflXl+h35afReQFOOJ9SP
8Ho1+uAPhwU/r52OXVrTnCyv5EPGeEwZhp48eBJjZ9XQCGS4yy1yrbw/E0j5tjkR
Ny2R+d/+wZFRVTeEyBnoY27Zej+JS2gl1fOCcdFkk3GLX/P0Q6/Siz6ItDO6o/Lo
+AN1xe/+pna1mnzVKTHesoThVci1sf0irPYDIzzU95AACN4qvRWbF3b2fj3hD7di
EKRGVlDzUDsZnlWltosoTh7kqxiIdiyDDyU+vluUpIPnuuA+TW/9n62cwcCioj9W
cGHWMPO623ZG/E3nymyHUuPuFxfqgzoyH2lc+gVnFeVPCGYHfl4Eh+rQBlxk9Zg9
akuGsWE2XyqMGrtmN6rATMAhFafYD6g3Kf+etOPoOkmMdtFANYN1isEBpkTYC44k
JKej/ZfH5LZ6aNEXwuX2e+TED2Evh41QuWqizGqLTX2OXlJt+2JFrnNSrxhhHq5B
YuSA53xYssh1SasdoipdY8FW3k1XDk3jUfHv2ZEvVfyBw46JaeHhbhq080F8/ri3
ZM++8AgO/8fCIVygxOeYW33QQScI1LTYl4spG6TPztQuI3QegF0vfe49whA2l2oD
5hWFMSXRZUuocGtyOYlpFq4sieZC5WV2UUa7aMJie3llVPY66+PmD2+/kSYAFd6s
Uevzu/59G8Ft2ykjZxnDaU47kb73hnhJejS5L6ozA8O1rdvFtSMNh9W5AyJJdDTP
XRN++AtKU8kZlfMwBdN1JQgYruRGhqwk3pwsUEcDwc3eh+wlj/Fghq36cW0/zNq2
lcIm7eNP9dRdThaAyYAuOmwHjPjcYpHwn6glJLy8buZyy5714O+6Y0FLs6RxdTYp
3g6pHMPvhlIus9GfcNoiwOvlqsk7H/FwSvHZEv+kuhjUyR+nWImD3PfQd0tgZQca
sSJic4uwh/tEm4PgEnSkMggXIgqKbtG9gXj3EYOmLnQv8WP3/sz22ZTP6pbY7fEf
4EhuElyNCzUN6eozRoCPjAd+iCZcA1KIUUQs8lxezb9QLaVb4xxy/2BV/YFh/fKc
jTWxKWAgsdzseScphkSHHK2xd0WLqy5df02xuN3D8P336ESlyVRG+Zr5t3mI/yYO
bnVRj2o5CUjoF7TPjZZ7J9g5+L9o/iQompxaLnBPlSa6R6CNV2zUw63mENWEoHhH
tN0Nb7aU4ST6HO4n6qdexzkzN5U34LtqrdA7cWUE+YkH532wXA6q8dyhWg5OwU7F
6/HiOthbRsRPAMvKxtlKqkbXYX/EQjcbQEegpPIylASsDoeuCJA4fZ4E+15cQ3xX
1xTH4dekf+HjTrHc0m12AfAMCXvrHutbu9YnPMrreL9rm8xh1xHV7Jt1ZCmMVMb3
p4UwZLrJBElDhSWdlZ9tTzCxUQpQoWJ+ySGaNJizHjjG8+xjL1/Q5X9ChATzBJis
uCgeGMTORHor/Kg/UELIxjgReVOocNomkTVEg6Qzl+cZqDM9hSXcIrp4afITKpc4
5xk4ZrwWGslH7y8m002NCpodOgoWc7uzufPa505Yo9LW6xFtgQVLMMcHvy/bXy/e
UQD4Cp6v28M9wDdPjTZHXPqWGE6Z8rXuKE7xOiXeGDH2Yi9Rl6hDOAZXhweoj+Ck
zagFIbaJ5T+UdfK7ayF3Xvob/tjQA3rbbtoTmGBXRiinOdNNBAXEM2h0yymVg2gL
bQbYYrJXPNeHvRtoSJIfQeG3qXx4+WudFNPWlvgFWbckBZv7MOOcwbbzy6ZlEi2L
LEtTwSYo1lEvBjfqKK9zuMm1J9FksshCREBgidkT4/h5Xomqog40PUciDEWW99a3
3j00HC0PmzEAx+CEu0oU8nPj4Og8ZkKW7CiSHycmyWBZ4J+i2gBJocvzUkhsDCpi
Wa402fYWsmYqspu0QsLUKcYJcMZ2WTKPVGqGXtJrRzWIYn7UcyQAKSDaxaBiXUrY
pjJlw6LYsqT4Yj+HMWyIreQXWAAwxkJE/Dy8g0g/KeKMhon+GmD10k7d7770sKC+
C1/fqESOq5bBSm3BINXwwqEWi9E0XskgBn3jecjKoJS6T2mCEHqm3pyOJNzBRYSL
vFJaGx9ROW+x84TBGMjWR9foqEQqyTqLlqu6GNpOcDuQQZacyfIgr5YhHkfYGxKO
tkBJfYWks64MSirPWsAiy49rYnL1ebgh5Hay8HuYLR472uKhIZzSGCNhNziZxjR/
gdjZii8Xwt70ARrLCFE85cGp2h58bwtlDD3Ljc69JqFl6S0LUREshpveORlrtcY6
/Aw/bN+duKT4wD/rGKyH/lH/4tMjGAlkAdQN/+gYEdY3Ok3DPRIagEZtS+CunD5o
Q+TZAdLHx5OlbBxdQ+9B2l62LeVQGYjRYn+QJflP358Do6o6Asx2KcjbRhYIGRxh
C0CZG7Q8LJ8pGBTjJNnXzczzMtznsnEnyeVKBqW4/zyuv//ZCikOctABQVdIobaz
yzTaJZRPBe8YBWBWVJnDhRlM+0lyFWqFP9q76fMxVCvxMqwBM+njnuD7aQXqlB+d
OIJpfbhrTlC22zztwyuyhtk7qVB0Fyza+1Tb1KH4UMFYGhT4zY4634v3c5AjhseH
ujHuJXCbeJ7wG8WAc0SmIowucyssCJmXzHCe2sMi31h8A2HyfOCfPUKw5xYy0NEb
C0hUPXMqFcYMGiKLBl+wCy6vl7UKIdmvNz7FyTWJkHMnOnMrA9GeIUjxJCx4y5O3
KjLlUo9M3OzCdFLykwMZrkudIghBEIPwNKmIzM0TaYTQqwMDw5D0PVnvjZTP8ibt
zdKIYwz7rHU328Z1mWuYNu3O5kKFn87BHyA0hYwV47BadmF5V+FKY5KOvkPtJNCk
EaSTMe/o4w6Je6of5HUhZTih/0GhhHmRcRVmbflq/hHhZWuplL78kfRjC/oFmWmY
T2rfxbeTD756WCwWWHycvgek5XIZC1weHEK3sgkFaQZhC5o66cwiCs9LxT/85CVb
JWyoFsweBpRxx83/a3Ts1RKRHuWFqNxTNojESwgup0gsUPZ2MGwdZbXCTPlMZrKt
aG5+xLlxT57j+HKL4I2MmMaCeoo6VNMeZEKn/ocyE6YdM21ziiuJz8PfCbCHGUcG
qAf0mM4//lgr4oEHeJlwrBIBSq29L39+faVsKvVAfX1Hi8+QZiCMjFpEr0PHf7Hr
R0CVJPEd7uMpEay/K/mjaN7sxB747iBZUGEpKeTxMHOcJARPJ5MDZQq/3NYfl9+J
JnFvqVjOLS/TUvTgEUAfdkmbq6VOyxnhpo5s9Xvr+K+w7ZWqfSNEDzJ3vvD3nHNi
EsaTkCRIvo75zHID1QVG6p1UGmaf/ZOZV9LdXg2sROiLFJ1YdWGT19H7wznAnVn6
1L1x2+9W5e3yWw7jWCmvek+8htB1d5DDzYJDc4GE5ceWb0jlkFLX26RZ/Tp+Jhtz
vGiUhr+nc3Eoe1fb6mNyOKU9ZBlIT02BgIFR028+DaFXSk03LEdcd3Lz8vpmvT8Q
hs9OBqLSAKg7JQ4g1aazFHqTBJB+VTTc5q0C7TkwbidzL2OSh5mZz9+qF5xYMBMM
SOaI3Uq0q90yf+xEXpen0iah/snhtvEfc/wdidDrj0oTRWhY5/9Zl/Z8tZjLfYiB
P62t9qC175Tj+co3NgoVShM599ffhowxOz248U6oOg21KpAPj2DwCDdvT+jH3ntq
tjBcUxPY6uuNjT1U2pGYzdEe6gPa+mpEbjS8ttHqd9VNiYIuZkV+h3Q58fkysk3C
Tuz/g3CDOEGrfkoGfWRuXmU+7j0zepdyVBHH/ENVCZB6QgceFBBywdn+plrio7N/
2nQXR6gFdjvxWFGz8YVhRmTf7NQUmdkcSD0gYArfJup3yFGf/lG+Q1znMwTqwm1U
tjrh/W5lR/FhHi5/udIlk0ICewBpVdhw0WFmOads9rGdqc1blRloKTsh949skgJ9
Pthp9Rm27Ky1twBqBuk+ZrZ99K2Lg7ro78aMOUN5qw9ri7MUEvyAHqA77oQZkSVM
urCAHCfagJEIPWRp1Q6B7mgX8sPw4XL6O+HobXB/41smpRyXEw90Qc5roqsAhxAK
qzZQyqP9D2E4GEx5R5BzQ+FRsn2IcxSuotmdSIaMyx8Oqbe5rw5m08CgR6eXwQAV
VCQbU6bbe49q+pvhifYiZkYOdGyO+9/a2a79WVeQRNsOD/5lcqV3vvGs3ut7umtA
RGjTfBtQ9QQwH/rYFxvrxeYdLLIUOeRWkHS7W3eI12pVgexVnzISGHa5pXv4XBM7
nEU2HfUv4wzMaFFqqK00mopgSgWrhpRUOSwJoh6qYrx5k5mZ5W4qhskH3IrqENrN
mjv02hXWO2JG8sr4YH4uB1urUtfwdj5pfdqFj9COjLH9FgI2NEIP9y8AgDvbCFy/
N+xymvPwCW2Ok2pjFx7eU0Rt/62UNJGOqFfszJCjddSW1rZpnob6YC8QWsl0gnpt
HWmrzpGPByPBxVwIJdWFQkEL84OGbXvdlHcQepu7/qA+VsflN29XeD7jhyBQI+8g
7GDs9q/hr+n0J+gnppuPb+Vpiy4fhoiXmFUrQ79RjtUwTNbfzyK6j7PqpEVWilna
efhMcuxCxnGgv3hn8HGad9n76RoDQ3heUIyVrXymBGqydoipIFJbssFCD+M7j8zv
ZbkfY2CpcnffdQv1cl23f6V6La6bqhlPAKHtHM0dNQWBB6Kcbl3/S++hMbX9q0xD
FSJPefURnR1t/XycG+vk3FJnh5lLd44sPGNUiYo1HI6v0z4/Rbfg+6rIQuxX6l4k
eRq4LseyFJpKausPJXqp5SokGCJKyjjX15aOVy4f8BHpxC5V2hWVzZV/1SRfLyNU
vw/SsneVUH+T6dZl803m4ylA5+bApUN2JRFbOoUasGHVEXWNw51Xf+S2bv0nQQGO
QTlhfRltygt2leAKNuvX/TXVA1YtEFHswFJGZjMYGOw0ZecJN1gyoe7kUzVMevIg
hJWqZrgDCf9aNcY+4eO4/aHsIuHs2rQ42waIHqIucGsfK+t/hv+4irf0ph3mr4zG
ONUsVW/lh5Y1Rccb1aMODF34cpMUDOW+qbgHF4cl0iiFKc/Z5es3iWI20LIrsPFz
XgDMLH5jL5PKoxdDrv7i02I/khCUJlS1T3z+oFRUV6Oxz1154Hz52PnxxnzAB2LF
KxHkkdAk9Y1gWj+Xe3hDBsJC89EPNHOogkE7cH859oOjuW2aoRSdRykDanKobtGX
GJDiX2FR1N1h60/JzwiSo5awuneNKftKSMCfLmy1ERloWHZL3499ClXxojQA0gAt
qCTXz86plWwuaqajUFQ9YuRkEuC/NMyPBCZGYNMX0+gpoesQj1dGYXVM2lvRh8RS
oNWI60xFVDIZk3rinpQzKwjQGsNjVHcRb8zfAI+3CsPTPcQSO4fc9eIBYJXnUSuq
tbx/TH6WP1AtHsnuV82jqtvEGIHWvjJ2yTNH4nryIPY+03RSN6hOYkxbMPXwMx5Q
C69w4R2nibeSOlUnAg/haHkefPwWUSw7QzvGF2N5WCis0kXXJc4qrSYu7WkzS8qt
CfBzbpyzaIIlFu2WSvK90k3GRkjkUp16Ax0goSJLHi0VhVY9gApPAcXUc9iYAgCN
IJztjfZvSkLRUCr/WH6EHv7TTUuMryO961nuuIWJQah1iqAwZdXJgwj87wC9I22x
5SVivXhjFE29E68eOfUBAFp2UwR/BUQxHetie4w+BDB4vk0pZY7O9omWT1eLVZPL
WjFt53GBZutSL6oCIJ6l0vrF/dQN5exIMOOf9LzcJSaK7FtO/F7fugg92Aqz9jg3
bDPDLeqnC8zPDsYU6YXM5JEg/RK6xeAN+trjUBsJPnl7ja8FAS4JlLFsacHNRTYl
PLnyp2MyPXZXmOBg7szvh8rj4uya1xCUhYJdvm73xEFF8gQi+p2uJxGZTRlwk37n
N3oq/cWKkVhCb1Mnuj34h0GcOB7VEc00Z5kpdl+7lv4iTcDMLjXGW6Cd7ZvY+xHd
OYqZDEPf1cuyf6x5OntbeZfu5ZKxwnolviesB4SpSP3sLCGJX4rq/wBCpBhtVMQH
wowAPh/Rgkpj5zXksUGm9maK3rR30eOM0J+HqqsTx25z5jyGd8X9g2CR0j5b6WNN
hjIlBRB7ZBi7U37SwEA7v32Dce7OHKlfA12flv5pKmC37YNziHTd2YWHNAUM4IKR
Js4tc1+EvoyH3NWaoBI5bah6plQwse+/TWO+OdqICU18KPun19ImlHPWzDauI6C1
oQWDxi/KHRIJ0T21P4mGG91AwM9AE/8+R9st2hKPdh3MVPPqpVhYa6elXIU2Ul6B
jp2kmkAjaK5QcFiYBAPXjMib6hphLR6qeynYjvZRhGPUOa9grcPDXSv+EwDwfsD7
Bj/2aW/IsT1wTIoak+mrPFdZe/VWOgNeYiWi2v/KWCTnSaXHhmavdVdSh8WVs8cC
3bf7maR9w0ahmfuG2tR/pHYKUlCagZExl2VneC+TcVdO7RH5V0yjEBwDyPX34eqY
0Bs9xbEOdxESgMUao4o+tRIptDcpEWqc46JyUcQoKMUnhJnLcrdPPmlHnOHzgZpf
BaFooohrobnBY1j/rT/Qk7fN6P98jNm362IywjpZXEspOlqOnuI5HLn/Ouv/KF+/
KAcxOB6IhO0eruZXF4EsNwJVFgXh9N4TVuy3JjFS2LHthhRDj7ZZ+Zrx5VQW6W0Y
txVtJPsHFBu/3s/6T8mj81HAMZepinL5H1duFzZLtD15n2aXx5bxqusQ+JC0Kgvq
qz68IjyAhP50xKtCb7glPg0RXUJ5gjyqc0JYttl6V2oZGTgsxwewNS6PjhnTQmSw
kJ4xVo4Z4EjdYcMd2/grFnMldc03WYan7Jbe8XOmQyvRCz+mJywTUWuAENNq1wox
eS5a7MDFYOtc9NZHX3xMPYfBvW11JYxOkyZS+NUgB8d6/afra4f7he248A7Ug0/Y
aXK7q9VLfOKsiDrP6NkApiFaBx3YCBPCkWmqX5eU3bVN56D3Mjw+HtuesiI8cCx9
NCKF/733i8/C9AAUXWeXzj46DW6D0xRUJjhm4pU/oXXdTKSO2TAdXvNUVoyEN3oU
Cg4Z28zllrFD2KXUOBxd/1wLQlepnrMZC1yaQszGJphNNGKZdvu36qQgnVyRKQXN
70cvCGHZPV1WP6n+3PbOsh5cdHGXxf7sWEBpG8NBks54Lslxujc8GZhQ1OvMF2C8
CETzrXfNQFXTOFDWgaL4TPgb9jSv2vRvTXzLDbPVA6slEAOkZ06Rwo2WaNe2GjTJ
j5pLrcMV0wVALJ2bZT1xiLHnoPsaEJ2ldMP4Cg9Gvwk8st+zivHYo8Oz4cFnUwPp
3AlleeoRb8gEUB0EVcSDKGhnIUgxHvdR7f68hX4LrE879jj23EY6tWcXSYoolkRw
qaPLiPZzW/LcnTzVFl+hQSYzKdUpzvrgFGsXBfXwXIWdZlKIrDpne/Di7t3s+xUS
Mfwz3M4+HR6Oe7fW83MdMfIlNdf+tDbdk6sMtpBqH+uHBNHom6GgpbrmsY3JmEzZ
iYK6llhMC+Xf51AKXiBXWUQJI5mI5MzI88XJRpL/jxUaiLDi0WtvhhEQLH0YVWtv
df+56hQ/OYLGwd9haZl/SI7qf+EODlu+o2BjHwADNFDhuZocWaZyHPC9ChkCTYjz
YDXnhe3N+XRxY1HH3igVMJbwqCygOymrna/Timyl+S/oeQGSQQpcW6Jq+79BKpe6
QkV1g4hBOd70ar+yxJeVhm0Ge8YBKJIZORvEtWFRJCp+CJVBtHU5WKUHzVKxx+ww
RgGgalNQRMpQYnin04GPeld6UuUElmKnWqEG+yVOMjjUf9Zlh38gYcp+EdFyoCxK
ZVtLf8dWpbToOysLavw9t7M+GFrZNuKiFr2/pgMssTYgBaLaNqLykJuLS/WefVy3
ff/VpRRv+evfm8+cDgG0wiKH3EXrGVmZFhI9bGysMwm2YgpIqKCY23GApuclQuwM
gYwMwzBtpjykcPHCdtHe/3fClacOWOsS+YMcsEkBkHLorFbqladQN26NSTAJ8v9F
O8+tFXTgvSb8Wo6PuMAbSnLFD9zD/1cgdVVsOUI1J6/a8sc42U2Aa6/S3gJyxvAv
6B/5YVN/xdeVZhM3QDjTJkAFmMpSpZv8TW/5wqZwytZMAKdJH9Gp0CZ3q5NynMrv
AhYOVZBOyxhCq5+JgSmxXyIw0iZ3D29OjeSrNaZIYgqA39X2QBagGqGhITFw9LZs
ylWcgXoJkDtznDc4gtquMa6uEVxqGtaAx4NCCavHX2df2Oe0bzmdGQBkb8/fX2Ta
DsZSrxdSr/CFgxzwXn+HYLGmM6srCZFwBlAn3D9MhMeGoUCWbIx93/pNZeZLY985
sunYHxiAJOMjtUEPNX4SkWjw0xGrLLqHibh4U6MFsRd85mZhAC6dt2Ro2/qyFYJl
/pQ/lfIIsLI/KLS693EFFq+NKblTxk5txxBBWs2ufkN3YWYJwFKY7zuxsHuhoqO1
r4Q7y3vqTnxkAndzanrZOkNtDJXb8hc9syhxpODJODwmjaqg+mlBwRhVTh+gOgit
u1jf6ZcEXhWJu5V5ykNpm/D+7vg8VXS9eKONI0YMhKFMu9nshHwbMPPv+c6VA/Fu
XslhOXviVexf9DINH2GmpvZi8v3XXQ1vI5bqWTf1nvob3xHPvq24aV+CGE8Z+UdK
K88NXgVGN/tfq6aV3ovj8UAs1PgUNoNIbZKfzZ/buotwl9ZjtO48IVpGGoQH1Lef
GqOf+7PxD2lU/bE2TfNSRDt7SvgyEkKgLEzihj9Ajbu9vbrhcGfUfekbPoyuRhkB
0r9fwX1h04uIRlRlQxcxhX9tiCt1o3ZZgM30+5CLTGspDKp0ViZbakFzCPqGHEps
YbG19CkMg6WvXcHOn55WUm1rADHhG1y34d5v+gIq8tRjAuIYapyL+Lus8w0avjcT
DiOqd7ezDPgIIY+Crmhwj11GvJLxXnNhYj2uupGR4UtUmXPGpT8p1giXNUTjbbDm
AooiespbfYLI0DH6Cfke73f2I1GCUjDekUPBX+7m+oYmYtyeH7PRY6JlBrcTi2tL
dfQslIJQQbmmLQAxONuomun80oOmzhJwEPB4ZCa5RZQQvWM9fJfC5NxPkozbU1Py
hCnsCxr0WkKvkx7gfxoIrh5oCetDuOwMg7gzgLElTn864nIFQHvGs7yAKngDw7Nc
Vxx07M2sWN05ieoYikn5ZP8srbCLXDmuMk4dmre+MnGPXTqI4cjHeAlUzBlE7aHh
KjqFnFt0YUETA8oZ953XRfuGMVs9cN3j3F7iDTG7xqCCuW/12ttBiGQUUixJtpN0
Nn+qNpUJ7FarD8giW+3uEa4EyRW2QIe9WZOFDlnxPw6bLD7NCOsHaawKeSdZyzAb
uZIFBhy3RmWCvkB1O70n2krKG5O/6kW3TE6lnBI1xIFqHBqBnnLG8f3DW07zestD
LG0TTWs7XY/ALLGZ6XOY81CeUgYRwK+s91N8F2g4hqsTRRd4ob3Hcy5QAfwKledf
3SSQB4fwdkz3Myn/OPI9xQYaHofaUXVzxfx/j4Jg05AyxnGtEBVaxioBA0vRd1xB
JD0SjUXlJc+lpZWMPLRgIS2p4qrcU2n+nJN0X0JKjXuZPJJjwaqcYCBeM7gGUScm
8YYs2CaWyIC3EuB+0TfVymaRS6eUz90LpguwRuX9lRlA8iSA80Y6xUmYYBk3JbjU
9L4YJiLy0NfGpGmfuStPQGzcEqMkjnbSqkcCm1UbJcVH9v0IA3cAhssn+kzfBD7+
mzHdmZh2vtO/aE/2xDEVAfVUuFBDRG3X5EE9nb/CATM+y+hNCjTWMnxzeJg19Ruw
qusyl2wUv9zMOFnqDcZxlcamGqTmxdpHQCxkbWnF05S8BmX8kT+7XWCS/bW1OY0c
j0nwA5HyDonI4pSh/feugDHoTmxLDX6Xrm9gvppKGm9mrFvHAglS2JEatdKOHwxP
3WLI09FmHFCKNQ/Ct8mWwKAJ3mW4kZ22g9g43Y9YzzuT9LXF7kevhEuvBHJUhxfV
u+H51zScH20srFqnhqpxX54KPw2mAVUYD+QxDMlVlYJm83IHFzhlCtWDC4gvrybc
DrCQIkPDU+rGCWCrPH3UG2WkKulxOqorQcHsgp/Eiogwd9YOsVp9hJoCKLpuyjnl
/0cp42HOhNzIm4X5KMBMIiZBGuDuHtlESwJD7Fx8YXs5sXT2NP6ofSS0LwLBo4sV
8JoUqImpnl7RsQ0xfIS7koo58/SZqGawVj8iucl8b6QFUiB7aTfGXof3kYFKQHTc
+YOXWATobX5XGdKKCF9HwPoi5W88srzF3cJB42yjETqfBmncRC6mWwvSagyaEa7G
SJkE6AAi8AM1VPOLDbIO49HUe8KG9/LjrNCsTmMkyqSpC+4Ewu2CYdTx3WT4Dc0C
+USbgEmaCdDlld1KU16pF9e3KH+GlaSmRXa+xH5jVoNYeVJwx9VCHMaeE5+bVDv2
n2/DQ/iyU3wXBINmVVux1W2ElRKcGyxFtxpkmZKBAXuBzsAJIGGy3e52zGoZziLS
LA8jNFbccGpxsHUD+RerKwIC3m8Vl3J0UmcQJaL7X7xYnFm1hmLAVk42k4eWY/3Y
loX1+MUNmgLPjITd5+NKx170SfjUxL/U6qrPiK1W3T38X3ZbKxYSJW95rWFXFevs
EPJ3V2IdNVNLjCh9Ds0lpewv4W2pgoKZJxoTs0wLD0PfdyCIQ4PvQ4YXyt+XZAst
OgEuVUhY5Dshdg5/WJka4QFL+pLfE7+y+4bbRhrZOTbs+B0xGJy80Sg792yOyRhl
BwnOXkMfmATK9MjzBEkLAtJ4ncf1mH38PiQ6yamLhTbTPc45Qbns7gc76B4AX32m
n6duM/2aUT3ozzQqUUImV+sV80PCo6xlPL0bmVbx/mVzwM9aiH+ezys6rp0UD+ZT
iZ+RwXZgiI5EPowI3v/Srg4uaMFWyQfU1+jhcm0LjWFcJkIRZCC32v92LBwlJLcR
P5ZAGLpwHRF48UgL1Rs5fCXp/JyyrPaMDvSxHABQ5C+q/F+bqnWyINGK35h/pUcc
UNcAa1fcMj25dwSdYn3M33mn+UI+u9yHJxLlwLao0WLXDAxLpZ/QGhroeQzHiDJO
rfGyVu1JcIqXzqBhTF65K5xFbYn0uP5W5A3ZVRizcqylEeCexA6EDV2kpyaRbdyW
KxEZ9kWaOTMWAAYBf3RQZ7IgnPyty1vvzJVHDCzaIOM7ekgI6n/lHNIT769pOnDf
2spiEcrWz6Upp5tRGc20iGCFwpKNCWEF0w8h9v245QW/0LUE4Mj1JC9+HPieWn6s
DafyPh2sh6Yw9pypjF2sHFQLhQJiSkIMJW+CwTAxj5dVMQ6xBjSz4VedgNghQ3vI
+1rPbvgd7nOguLcpvjj4Wyt0kKkXadmOl4j5N7KCcBNb7sOJ9O2OIDUB6BOuL6Rq
pWwOV0q6G9FtbUIkeEY+MjevoJOB0/sO1TXubSwn/DYaZ8r6mfDhceDtxQnB5zoL
yfD+XlKOUzncu6Fu6SoqirQNsg3wKq+qdpLSd3RJVjRlVZzn7fb0CxnqZxqqA2UB
Duc+blnOc8OO2AY6AlL11ajPmnqCpKeM30GvYavUao5cKgsAW6ppLcS7mW8IDEIE
q63P/t28EqyVt9eBXGwNntwpkaCXQQ41HxGTY7liK5E93M4eV/vXeMRte90H0kNX
2hUg4FIIjVFO03llmbnFvPJYtXRp5pCHgDgae3NxUo5dfTsA1B6F+IafGOr4DrRJ
dWyDQbiiRGptYZWM0/6B0garw/CbZ7BQsyhdD9BnY8CExOUuBNHHWesstaC8LG3Q
bfIDDAGcsiSlISC6irzWM08/wBao6ybKht8IpZN0FOBgDQsPh8Z0c0vwbmW0Aq+B
zptQJ+e9985taaNySr+UujPUvoVClCAECZX2C7EQvTEaRcyY7O4kZKmv8TyxyYln
kCwE+x87Bht8wKmGTQKTVmtsDEcS83XYOsSn2j7n7VL50lGgNTe2urim73t97oPW
Ha1PTt1PH3qIgGF6krqxIkwLqTt1Ek2B/FSyggqfJlwZgyI+QvGmZm4uMcuUUQPB
x+CbXkJ6nzN0qvahfqgUA+7tx+ztMEbjxsMKvs+ygsgEQKaqIxcbTharZKNRDsyt
DDml7ceLsWa6isRySgVp2CvbEwNXV2od5drNhBx57hHQWEX+lMLdoMdkMKHCN4j4
3uRv3Q4X0AaV+VfHEie9XYW/VsbfNPBGZa1ulbLeUzRx9RgOaNyk2qLcQrHyEmLC
QFFwEd+hvxnj43GkDlWWqWQt/B3a4pAjo6mQb5AnPkaONExqPN9C/V5y6ffW7w07
MC/lfp5iPheDDuzE51uHHR8KpVRV+Ev8bpVrS4otMc6nVme4DTCfaEAfp0uGW5VX
YcViXHxwcafwGKGYFOE0RuUXqE99bW3ADS4LlnofOIgP1yqask8oJWTVHxZbH/Lm
YicvdQi2ZGjL795DH4B3Bn/gl4NWXTfb5OFXFfrw7hjY9wbTSEG7pGsGj2CzoDJG
mdJw6KXxk/a6kzjpZXQSoEJpzlCBOzc38ScRv4iaXCOP+7pHjq9KsohP9+ww1ceG
2AfT7Y6JmnM86O8EEYPQYhjdSatpGEttDveWw670lkSlbO6Xzb0rf/M/bC5zxV9Z
e/FYzTWIhWKtlqDI/QGvYKrxZs80Exj3+117Tv5O8h6C3iGKgTjFIj0eibgmtZHh
cWZI8+ZNcp09XOaWwfaNH2IAokJsZTUmcS2ha8HQVHyAMiHteDNmZZxWw73D4VVy
vqGgqnB/0jlz1xkoT3HAsttfqBY7PlviTdQk02MCyOE9CXKC2Mk++leD2BMxKhln
DZwYL02nYpTKG7tuPXfWSIcLX0jcQ30PnqJFnHUp9uNooztIU4rrz3EOw9hmMnop
vxnay6is2NkBGudGkog1b0hXI7FN/GPEXv8lRLPA4z3AvfL3XFdlMYGpMNSJZw9D
Vn6GNlr1XDVw8mCsP6lA3yaIhylpsVt6dGfMRgLOx/aUv7zK81tX68jEMw+9xuI5
+io0YiMbWh+50P7JHdJdqHfIoklghta7cLmqxP66ZeniUSeQhVed+dK3H4vERWcm
nG4hpNS1dwo8zoLiqDvXIftvvCrvT6jRzAMXlpsRB135pp0CXiDRU8Mcold/r9Ql
L+LH6wEi3d/vXPQBQSkYEroLmYA6Nh3zVIVv5gIiQuxgWdl15OuSoR2ZrqrGYejE
jquzVRmfWAZINmJv/11zTCQm8MnmrxOnCjNV3Ci1PHqG4I25WtTvt3SJALGz8BK0
xRiK6zM8UqKqjyiwyTm1Jl/gC8s2z3GPcto3UXpMeCKspQphxHLo1rsKLw8bi384
YM+NUf1Mu6RsFGvcvWe1zaPG7sfRUeHOuTGMTBWzt5Ks6WA5JviW0KPeuzeRaj1o
sEkeeOG1R1BWvgeOZTdUiFRxOra1AGAMFNzUgIvqYz33zTkCL21vHJlwN13W6OGa
6zHGnFyy5w5l4eyQY8anHXJJk6n71DOICWnDYGdZuPujAe5rOjZnNkwRfrToc059
bEnB4XT9u2X7C3uRY7ayR1SMd8HQnA4AyeLX0O/RE/QT/Dbw45iEojHvm7S75//g
zWFmg/JXdohjHl4RYz1UbKBTsvnEf1xeprSpWFhWZ+cenNrfp/Lm1FvR1Lr8obhR
J8FYp01l5MDRjnwNISbaH6Qj8jZVPy16+IIYDf/ipkX5p+NsJTLv5Yx4gUUybewn
nI0HntiFicJMyB531tj8g10/hB03qh4VAq5xaFY5OnWMQwKaj1XT2M60HYI7bpVH
2K0FGBZL9jvlkktTCyNzLf3FWnv403VLOng4QFG3r8NKa7h9qnGHuNt5t42gNI5u
yGY/lIputB0Lso7EvUhg1tRG7Gt08V/EpA2BCw5oFGT35+ohFokn9sDKv/2W9kuw
UukhUG8yqrsrjELVcAhSTplHwxXBaBpRfOgYUYAz4LLU5yS2A01ujaF3Cppgcgkc
pERjC618H3wRt8T1k0hZLsEJ1eeqHdjpo8vgivgBVm8LCqyOP3QXnvEC1KR0AOCJ
1ex8dxxeuGuQ2J2Ylup1bM9YSFznzsZHQgTrE24yfApeVRr2wVm6Belh5ViGu0YL
TKhtrZ1PUA2HlXMkNd8bHh21hN0YpSn2MiD42axYyd7NvHCGIko6Zmz6Oh8WDusL
XsoVQCfCbrTRHRwqOx5Bdv5eG8ceCuk+0NNzSfHRdWzFbzAT9uhqWaVPLjwSsxor
crNY72DXDOHEZ9RFLWh8LY+R72g0dc4rrgKOjDxSB5lW4G/WTF/vX/D2xQ5u2tKi
UXe90TlXiv+AB2xzuIiNIMUDtPcEn/6FlOanSwWj2BqN1xVqYbvzOvoUopaitb4h
X9uLi5nYyiocEK19rQGwq6MHoqn48lads6QauGPyTRYcz+3fNPuP+mSruxoq/g3I
yCgX09PES6ryhDw9hS2dfm9dCCRG8/J+tYp22t4CpaASSAuvh0i80sqpcMwF4t1B
buR/nL+/6KM4vuzUznXNQTT+0hXeRwCmRIox9IDrSGnbaVSDZe1hAEGhsRYmm9Cp
rZrvVfm/uu3KuXJq0hpBm+nB8DBSqLnwnmPX/ZkbC2geYNdobUDeqyftkOzL6ucs
6BlhZKA50fectPxKVENYNNmHuJ245AKMWqYeioCTls+Z+xg5292tMCb2nFAYzyAK
HfQpz4aZ2ITqI7U4ZCeYnb/gED8z8qSJm5XBdP1hikK0uTNwpfZvR4u/livOy6ms
3K5BQwr7WZMaHKKiSahspmEK+B2f71cFVzJM04w+lGaikbo+ZpkKUMJ5zrvC/8a6
litYFWgUi0yeuOOHcT6ctLmunGGTa2ADlKKCNUYSl/9B+hfHJGRg6AcnCEXkFdQw
g7p0bw2yeqRgBg41Ip7tBKYN/vk+k13nJSKdWgosWdD9Oa7AW3RQX7CdwgbdUokB
TEayZX8jIhL97TDPqeuvIkt+oTW7N36lRHaZlT1rVBNvAkLYcobSAWOfzIS95ph4
jHT5Sh0VDP5h7UIvp86Ph3n9AbKho2jYYIpVxOvO7yN76jaCAThrgB96ipmI0btt
ZH1IMYg+KpJdr53nkWtWou3blN8QZffWjvKf570G8ref/z83pVt+LbSKUQ1h0q3u
ksrQmkLLvZMnSG7oQzxp6kB0BRYsA7DGAfO0v/hlz2U4imSc+fPSy9R0g+qGceQp
BEmLQ+3dm15RGeUypJOM8vjNrBzltzDhrUjPwyysVkYm+jw1db5TMlIp+V3QoVpo
012vf5neS1suinyAOFeZNC4nb9JNZKbifRv9WLRat6i0sFKQNJMAv9TMEZMztyzc
zNP8ah0LzoCe0MGbWdK5G9kGfcnCdVeqlKDaZzJVps/XVLx3altxao1ppFdhzzEK
OOVXrQMK9llqua64Kyi2JWUPDGP2Es/sP+cZyiYEprpYPc1D7JTzch4EJbV1vfv+
NLquqUQ6yt8EVV84xwCkpvGuGvvLyUwXxCajLBa77YzcU3JmWa48MJBW9JZj6gVR
avup3uvwccJKyRH8S07v4gRrnSnRlA/L97oR8MX7Ii8AprTpGtclgMabbJ/DD+XK
PEeaNSFKmfO+6JPqD+uONAx9cG+rBwKDQoSwp1EuaYWYozThwMfk+Cq0OzkKahiI
mhBcPWz5nLamGzo/3Z9XVFxfd1VtKHcN3no3PGLbio6NtCrlHb4szKOagWLLKnTM
iOccknrdHBI0MVz4ja6WWr36ssqg5Ayh4MM2VPvYKa7K+DNxs6Xb0MT3Xm5ZbB5S
1PM5ZZGDo1WZFRPEwG8t6ZTeLRXF1JBTqkZFN2az1hSAG2x3WfkTPWaZDqvZN26h
9H+ssvnDj8bpyHSwseNyUxiYMsYvYk7APmb35pJfEXgfejT92cymmboQ2WgNQYZ2
nja+Mrlm1IhK2tg8ulpap06SvMTK7F0akUtlp48FQBa2L5euJv0gxY41yncXBO/3
EMQqr+Edn1ADOHtYHAg74GU7Hgjvi+pCjGCUqkROKXrAxL4m89PhnGgSauumZpST
Q7uTGchfPA9zdzMnDvQUsjG4gXYckL0D0gQP99++NjTF4Mnj9sIpvFVMeH92n4Qk
pDfESydvlZku4IcMyQvls7gUFH8F/+l5Noji0/PCqAOacxucg28VAwh/jQ2uS/S9
cnOZb8lz7BPvfstp0cKzjia8fg8yPQGVFQTC/GBDuP55e4ddZLCeFXjda0PpguPc
9DeV3z8I/OXUxvfY6Bj38ZQzqdIRHozId9JOhRbxnaPm7tMRHN7UjeJ59tPMfxPX
43rA4qjt56CAJbefOFjN16+rbMp6/T4kWBLkGluWlyLy7ItQ8xa4jYmA17QtzZUV
5CR5VAsZezBffZlpyj60k2thX1BUPyb0YokBi5RZ0GE0mLozfFCfsHMkxTB2fdWr
h1v61OnsKuAKy/+4xJEqI7nItAyUwbMfcx3OhV0Ro6UHhbhkGTS3G39zuwQwciwU
T/tC0ZMlDDfhC3SS7EveVnfjRNeaugau8Sef5QXCL2qrNJoeiyhrqhWmfshmFeWl
wNquo5JuwsyfJ8kiiBpYiyLXZvBZ3ebebtQ9P1HBRyXEeYRBwhizATqDsSh+mI9Y
VGZf/ruccjSvVX8IaIXkVe5HsLxZ6A2IqDpN5hkUkIEBXUqNJNNFh4HNtpk7RZOj
Ia1woOqjCEs7/jaCf1Okuv+xktSOUGcBU876M0wISHEa5+jyVI9ofesS/k75gjSf
3amWPZGBokXctuD65dVM/zgybgFbqPEQMCcRtCHcn1ejbXa2PkVzez4LZHByHdDJ
F6Mj/DDZSvOnZIHNF94Ui9YOy3Pw+7W6Pn6CMWtV3LrvGymVthqvBvyNf9dLNXN3
mm74SKzsboeIPAIzdC16svqu7hhEfJuDBv1MA/Dm4rWiNfZnjf102ssHyzOlcWHo
At/d6fnGXhJ+2RQbHs8kejH1TKK3pRT54M6qGawPrSDWOt9NSsu/6I/vgBNE8KQk
/yelIDw3TOYP6Z9nKOnPK/HQptmdpHkcL2zdXFXkdYGh3sShg1sb2TTILj8Hb9f7
9KCqEeN0wVegeCSGgcScYHIFJU9ojq/fUtkG4qaYMTHSYcc2Jevf8iV/e1P7lket
iY0fT5dqi+b0e/yXpF+cNnlAmaI7Nie2Q8GS7vKrEsVjKWY3tXnmldEeunQLkTvP
Pa7CyuRFPgJsi5AGUrIudLK40bO/WYHhFx8tL5mM0MAjPvJ5bb+fY354x2cCdPhW
5ctgjgwiWkSddpQnXLBOFl58Y1HYmij/K89iHZsb6ycVRzECTNbYw9py9nQUuI6M
xrbsfuO157ZeHFe+Mz8k8rl37+Z9PBa71j8NkhRXSHwxTDn3n2iGXVtOFGP30Lx4
ferg1UTMWlby5uImspb9qd4QfevYNNMsXe+cbKLdxB/wFMewWLtGC8g20UsnNBMP
ysCI8ozVeWeUmBZSsgJaBGvzBelVxKCFp0XZ25gv6diJSLQolR1+q8umW9aCTHDR
cByD3m4nCyGWJwkiAN95O1V/7E0Je2OCsJ0rvTNriEVepD9+GqHOzLlSk+je2Hx0
JNERvwBFiTwSaV8OtjIpqxTBvCcHkliDp7LBVCmdA8YRKd7rd1BJYTJAbBGax1L8
pW1+UMTDWgRaOs/q0hcNTslvIOpTTs4SaV3qOG+t3+OClPMH7DO9GpTzfxrry2eR
CiSjKOcUZ7h8AAfnYKCgQC84kno3ZctlozrPyLYdD+URLpjozHbsf8ECvATcc5gz
hZmCmbUE4eL82P5mAJko1L7/RfI+FS8BUzwUS/ZCDVhDJM7zWDd8ntgN0lXJBLTN
TMzFV8vVfldT8MD4sA4u3ITkFKNeVxFaoTt4OBiYRdZqmxqXMNR/LIUpfbriOuY3
9EpLrgKC/8VzZlIM4jeVsFbVWzj6BtADiuJHMO0ExNwMkWxk/v7rxW34Tst0BsN0
fThcbQ7/byek43xigYe7UvU333kAxwIZ/Oyw9P65jMTnyHTbknxZG/5zs9o8keLr
sbWkaOZGws0Z+8ocxpwIY68xkilSMAsa/ectez42sByZu/DRjMM4/yclXsgfvMaK
Vr7cALg5xUb9ahdbmh9fU1F96EgW5tZF61CLng3MieKa/gnxn3Uxgczy9EI6v1aX
xgHxU7zJ1hokeDwqoboqldJRx7zxySsPmTs3QRh5Xi2yA0onZ9de3MtmTc4Vda8W
9A4qWBa2ni/Xw6bim+6KzR8fU8abztiW+KQY614uwLqoqEUV8jtc6blMyWJBFKt3
49Enw9jUZ4bc+yAQTich9vlZAOP8jfx2Y3ECTJVezPcXsscnvTvegQhRE0Q5ZK8Q
rrtKwKOKoxoy1QilTa4oi+N17adqMr4mP6QuTd6RybCt+1xDLre+8YeevrzZAKns
TvreXihL4UpwvFxWXzNEQNTMf3fhyLmHSk0SYuxEHpaoxtaygQjyzdALp6phmlHD
aK/+n0KTHHviauYKTA2+lzhJ61wJYpHKmkhJGP29C9jkyUS3cTTZdEev+emv/9qT
+QRezkrKYamZv7+2OwncTBQj4cCWYJuboa+mQ9UTGlk621yXo0KXl6bO4Ty6NY/X
D/c862MYCsOOV+45hIDIobzEpdZzGNShMKRaRBL3vmk2XVS9sAyoGKZYJK/HUN5W
qtSAYSpMeGqe9ZPAaERHokZWAWh7tUUvg1pQu/wI3c4q0VLFN8elNJMJJGNpVdvQ
sQQr3Xc7i2bpa8iVS0jiUZCZ9BeZJcNaqvwPL++cAm/5h2wvfaYg4VeLP8KuqT8L
H7fQt0wltL43ebbVgbaX1WWHGfuB4yoNDjQZptpdL6syES3m2Ccitq9YgCKNxCef
pq3+ccR4k8FwrQZ6To/xcpBUOP7zuBgmL9lclgEUzu5AHl+nENDl97usWwQImCzV
dvYMC3ji8R22NZjwZt0PEiWWYQxAb1F2ZF6tb5lNjaf/HtWFhtKbC3EG3PMu1mmS
4DjMr5HMq8twCGmTLmg9h4k89xlYKYj52CFulzp4eQDPiyTu5mC82ucAVTd9Dr1e
aki7OFIpuaE0OfwZuCc1yTWJH+gKljKyEe0KVD8p95Jcv7OPvqHt8HjAIz7twEnf
aAk5X/CKlm90aLWb5O+IQTD2tIp3pRMB/zRKBJADrT0E4LQMiPKYvulYWzOPL3Wi
uVMIG9pFdqOSj/PiFLAPUYTxNncp6lw0oZW/IWqITe3wE1LraL2WF3aGHcLO+4cZ
QNOBY0eJttsXKbqrOmviloHcpw6q86mRDNSlv3IoYkWLVXGjqK6tOVcbthSmAbXX
BYSj8lDiRw/ShYMfLImB7+g70lfe6LE2g+OW0/AKitwi3xqt0cnsz5bYVt6rzeoA
t8C4l2Ce3i0qzR1+pO9uLUlCIU3GogRJJAaxqoumoCr4PasYAQe3nraOKSA8oCGh
S0Tf8YSoLHxkL7yJJs8hkBfnYg/1f6kzhxYqtiumCkE=
--pragma protect end_data_block
--pragma protect digest_block
a4kVkmxNzUPMr0I6KaZ0gXZ0gsI=
--pragma protect end_digest_block
--pragma protect end_protected
