`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UZm3X3zb6AGO+XvKvsx43RSnlRplCefs1kFWsiCoJZR911P0zwaMqsS/mYVPn9cd
FUgPyEtFlHQ7/JFESwOY9cj5EcHukpIkpjUxwttNsVZQOa087XWb1ctENn9jixV9
aE/0xGjTVc75wl7ilngC7xprDWAsmumjacuP8+cdUo8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10944)
WoBvZpBwDKZTuIPLuzUFW67ndJbM2frNeH5jY5XIcREDv7Vvv7WFNPkc2f0cdniN
me3sRzYLcTmx3Ann8caVH30qvdelYgiNs5LA7NC3/zKX7/n85QzQ0f7SsjN/OmLg
lvZFtd4dhcjuS0u2nPxWNueFmi2WMMIk2YLWHMFEFpIkwwYUuP0uqlS+7A8IdDD3
/WHGhmIgOnZb3lEhpvnoZQElXNN+YLGWQ6iUZxtg+u6zT4/DL1lj9oRcuF3Ab4R3
9BHP/SKEiPro7egEX5d/FgKx+6eh28ltaD+G8YqDJo481ZIlffBRSEVgfwnDi/n5
vzDm534IybXlhanptf1TagT00yc0dlELlnOFJAarIKBXQXSqZ2SKmOcbprhh+V5k
eHXjwQlVaVUP5El/xd23XWiNW6+77Ld+5oAoFQRSt42vu2dgFjnpbu6AIqW/Gbif
a8JQFR4baORAEM0JrH9BKl9IgHXDiL2iC0Vyo08cYbuSK0Z/pxg25KTEnP2EtLs2
6EcqBHb8oBosT7D96PQe2/CWoBKhhE3VoeYulz/dp3FH2kkzW0rmhJHCeB4G1QNf
dzE1FaJnnsivJC+v0170dB9HxVriwpq8/Uh4jRbQ9KvHhfXoz7j1HZ3avnONC0eU
luLD2kejtiC5gzKeTDezUeRTMJhVdGitWn2y8SC/YLaDfzGI4+GKxy8sjdTgiSiR
DAxPn9DYmJLgzHT7zjh2DZfY1Vrk9G5aHtlA42mXB+X4VDH0Yl4NWzOB27atF7cZ
jVAUtkkS22JS8ej4b6Bkcer6ZQuJiAzabyYsB1N9Y3QkaZlwCSR3dkIDUum479l0
pjnJiOvmgDxlMfaAkrNK2F8MDoaYJnfRs8wrbGZ+1e/9tA53FeEtzgnJY6l0wGis
uUn0jtiZ1ZkuPDUK2CdFSsgmR3DJjiR9oZcfafGGY85/tYwS+7f2TTCZH3C2iUaM
jSTUpTMeEirx6+8O2AhbWdKb+nJ9h8m9T3S+wmG0Zbn5m6rssQ6GAqGgy5bukZMl
Gm8cV4CMlMXPa4ZovhNbxwbnz+m9uEZ+vwqKmPzAlOSLZfEcKlAZLqhTZC3AvhPV
JYGlYdI1pSQGg0pqeaQjCl53cZ7ExS/tYG+OzQLxZtHUyK4eWUivvmyMelv4Yk/9
pdejDKUIx+vKE0abMsWGK90rz67rJtgbbd5OzorhZa3eW7VZATJ+2YT0kDexNVIj
fdud1T5gMJqexpqafR2o7xoIAnvkpWNP9NwzAklQ3/7npZ8whp4bKx2Gt3TrQGp7
b1bthAjnpBtkxCQs0uZaqH7OX3FecguKDZY2BsQyBCbRtdmDubFUhbbdQnynBCxT
kFaavsoVEkEgIl+AiyW5c++fQlZ4YyRmC4D8MK6MuEQEqx64p3rOlQmHFcTzGglO
Qq+M2MVmXqjwvAsLjfMuVOucuIWbL/NybI9shAGE/qazZe6GeygQKDNXk/0iXlrE
0aFXB07cwLbDHNujflwQPKnCg/DkWTMnsoq/fHD+r/obhI1+hceLNkYsNLsAhX8+
D00XQtSzaOwaCHkzqrW1boZD1Y5UOkHMBd8LAsTaYlPGmJ2sznQ+Ag6rcwJqsBsq
ww5ZGn0jOBktM9w8ckSlZShR3qe2oXM5+hpXqetcJMTwnPE7QKB2ofKxd4/guRJ+
UhTPO8VPIEoA7Dnne5rIaVnbn4QxWhi8OPkZSD7C+AkWuXBvwo53VrCAppT0pAcg
GmKdY2Eywa+3ZXruEH4nikOwTPa4COY6z8ZZc0KFQf3GROnTWZEkCf8vP1/OvYB/
UT6dSmvhC+bJPZlSFfZ1jWH+dAPUZTF1796xUGpi68x7iToyF2AyVD6RZDymHhqn
GAwRrT/+MA9IHEfuKjqC6DWzFPvAOzT1gIXuqiezsVJVrFA4oHkhdYX0JO2MHpRG
7A7xuvLRNnDrHpbuzU5NSC2ch1sytldn9kkPcMpoVZ17gnB+2Bvt7sOFR/XkITQ4
vHe0Afhs5xQ0Gl4FYG4pGPLzpc/U891zLJIJMtkj9s++K3893+Fkrr3hH/VKAKyo
CiMwILF7Q2I6gRxzRYo0bferEHAnmdMokGHTGGvukywTyr3XNn5+exCaOt9T+EOu
X1ZGTrgMNSki+3kO7qAYigFX6Gw5Pxwa7+ky+lxtm1cMgveX2keLPRHRPCDCui3G
OepRhc8eb0dc5PJa/l5U8iN0ZliypSFrgaO70T3hhcvckeq432w+HEHQLKpkKaT1
A45DrMSe89aR7oxn6G5TGqSXRzkEnMD5WwEuu61CS7HSSld66iQMOzzHZ5AUcQb1
eOAPNeyEXWY3S6CiE1OZ0xASj4wFn/zJtlS0zVdXXuTFsL8vk3nAt6W7J4xYXWuq
VWIEDdpOX5q44eacYeK02hUhUKI8nEeTLMPemS7HFuAwv07K8+7CJhH79fDstiGq
Gq9qKGU0IxHoAHZzoF0w03GuA6mHqYs7tAcFOwjytacuLKpxVio1G0pvbkB9tjmE
Vr5HT0oZPQRBDqBWku8W+p91s38h2dhg+Z4k0kLt8CUKYf5pYF2aYHubcCi00tCU
FALNeT9XbpLq/FVfLzMoRWtuvkJAiEtxN37W2277f41yh5JKyxynrz4cJmz8rokQ
HoxTKFh+u+sjMpV5xDOTSHlnsyg9Nr7TiWIssp0uDuIGPsTzKqFSurESAcrXdYSR
I7EbRMjl0MV8SYm4TI7MB74pPr1wNB1gOga1K5Lsd/C2aiErbqfSuKW+LFgDUeQf
8BdnsCtpO4+hhMiDe1OMise+os7Xj40vAab2HpDidf424HVFM5eMCLZ6W6RQ9DcF
op3Qtd15J2zouPdmCZCKCVa8U68UUpTZSxwsz6+4Qmb29YFRoKEw6TCtnjdtOtBy
mxOOrbE9Up1rt2EfqCX06i8bmNO8NBoDq0QHdp2diYQkOdELdUoG9Uw/dxxNQXYV
5iu5d8yLKrtWaq9aeTQpqUFtWZ5PeeY0VbkZ5qCyJkHBhVxdj1xFg9gojioCqRAy
H4VMtgPsEHOJYhSDdrvCHZkq5ahWQ7ESl7Epv+nLIQK3YKy/WcXfSofgJnQ1or1x
jm0xQcxM0WpUzCA5v5AAA72GT8Wh3wTJE/WBqq76Hw1P6ncLsnJ2o4dY9JhsOi4L
wO08Nu1ZKUe7NJABB+JT5Bw/DVrRtPTHE7RbmvnDsCc+bXMEaIju6NLej1HuAFQz
qKQWHn1VAeic8IB5j+wQ1D3Fh2KiV7Zharl2payX50NNhct3UDCXh2wt7viuM+ZT
OQfHSvuuw8NUxSNiu87RFJwspxIEN4HygW16G8hM3g0Ggq1OTvMPUKXTCLht02BF
ogW2dUHCnQEIT4RD8VnrIxtp8bp6Wup5Sh9cUcp8KgoeckefGU8sSZ8C+gXzM5xi
dhhL93nLVyQhOdVjuZAwt6z9axrgn1g15NvtZ1aIkkzYbHO7DW4ZYoqrMU681eHk
bsOWVia9S2BuI4GfQcae2z+GD2wqE3j9fmwhAW2CiZXjr+UM08T/NknTrrQzPYyu
tVqsgL48EVN1vnYAmfx9dkvHLaadEMKPg1X4dPilg8L9myJrooEivlv6wk4whNhY
hbOs2YGeTjk1cB46bl0KuzhgzFdvPaxfkRCGRKGtf4UrYiQFb4WFhTsGUqKdsos3
m8lEMfNeyI+sV/ayAu6Hbjbcgv13JT42/MooVfF4Wzko6LV+t1/eACkqW3aNue6f
YpmXH9rPd+sKGBpp8BBLQHy5+14jDw+ybL9et9Muk/fIBSRIL1dtUq1bgucIuPg3
3rpx8pddxsPbC34R0WlwdP7YqzFYL1CobrHzhjbrbsFqt3pwav3782BqnI+An0IS
2v656pwuJyk3b5i/P8BHHrxicYXop9tnrFKc0AF5QIXH77p4Mv6/LezDrv2wA9ZP
D2C4BE+eE6AGcgHahcKNplZQaLEpdhYOmdNsEBd1JhEBDi5qIrTHtU7N2AuESKKa
3QXYpzgYw8ayZG5KJ9Iq66npRLpn/eVkJ+f5O8nSYHPi5pRcUm7PN9DE/kqoFNNv
A5CquLKUHJDWVnhdD9U4V8RACrkZmkea67IF31c7Xz+AYLeNf7flMfKYz+KEhzqE
Ko72CFCQ6eynPRHh0HZtWH+o7t4DAMz7eEaTnZEoDGuWZmBiyMzKdK1C/I7CkynZ
M3m3rHGUKCpIs/5Ik5YTntH1jFN62n7aMsB0pcZuJI5Wpve1abMllx2CfINLu9zq
6PjzXjgO7wdfQ/uwPKgDB7ul/ax3IpjaE3n4pHYu0yZKioElJwrDS+f//EfiSV9m
Ef0l4OqGMRZn6E61dt75mhUaE+qXKQHGAI+dHi1UOnCozafKOArlwNDaeCNMA5HY
2OeFyJdhuArUBNtjgvlClg7hDhSVQj0pBeg7A7dzntszrHEFJ0/tMfwyYWceWjVs
PuDx6AU/MRPEZ18uY4vVocqiyn7Dm6c1eUsjQ7aGo8YszpPJU/I1rGWFZxmJ5tOt
7+tlynSTBbRXO2ejCJ+n1NkJGmV2mKhCWW4PJ+x4SPd0tV1+o9A4UQanoRPBgVOG
w1+vSkoTB5CtVh2PMeh3ieKlDI1K+Q/rLJIkZhzWTZ2WM7k4mx3LwSiMQ+EufIIT
nPO8Q/xGStpV3FrB7ngVvENDu7TA10jm00f/EYbbou88fuSgN1ymdp25EPU4qrWO
5ZR2JEcOiBbJiG6lTG+LZ83lhQsVuXUWsob2YgK467FiKkJ0ZxTXXRbicCs6kcob
V+koIYpbKhUyIwfhdceBP2P0zXV9p8KCPDE5o+bO6dSQ3j3F8/V/sntWPB2S4Fyv
tk9d/Nj4dJr/RpCwk0hYwXVBbPREUof7Auh2ZtFD7Vyj1Ur+6C2NbUqKOIKnaD+i
8AToz+fLhD0HR91m59I0JOHFs73Kq2W6esNWcUwPu2bK8hvXFlXS35j3KCuvIdG6
uUPzOBKVAIt0w6j7ut2SlE2atJH66J0DYllCDe9/SmI839gp1Fvuv2t296Y7jRWY
M2EGsa74eoTe0h64IFdK/wkoEf9cHoQq8W6GtI3mcDZVRoEQ6LawlPbvA6eRMqvm
C/4KYID4+k9M6oTRM9RX9svKtJvJxPxjkS0z6PA0s870jP3aL29Afxm5Nup89kHY
lhdvpuVFXeI/LxZCHREM3SzJ36gKM/ZYjOIqjCiAWccI1fN+K3yEwAcAAepqnYta
DwUDQQcKipkp7ax72cI9txkvNzlLDJQAZCZCLroCQ6NIWimb/SLRyesEMTb4tU4F
4oyikiGndNJb16UNjKGwhg8I0WsfaR1ROLqE7xJKRBhpgtqeJ9RNxSZpj4z3TuGl
CzX6tgupzL5wTC3XXNxFmvzl2xckUpFbegiUFS/5b4bJPr9f1gQFFXzuJIBmTmdt
hd4T7LjoYxOX9GyD0p+oX6R2zhXSpsm3Mce0Rjjd4vkn9usmCwwD/+A0L0vSwAMK
eu2p8hERf0GQQYf99LRBh43s7Wjn2kiFoiZIECrWgvIM9GMm4uybmJ5zMP+wzNlJ
gPbK7N5LPETsCl2Evi4X8vOdtm0VEQasQojFg0mM6/hbVypNIiuLYC6oXf3YkGro
TSgYH/jgzoZJytR/QQ0xhwxhUo1ykzUDsCy64zwHh5BOi7ypa00NSHs3SeI7UlxW
fy/uK56XowymKEfRhmErqLcE1SPziOwganWbdVVelcxSyuLiAFYFc/BGCYSPAdZq
HKHgywAV0sP4HgBtyRmb1JTLLVczc6eEKINZywkitV8HA1mCK+4IjWZyNpfeQ828
yGFCkrDI48GJzD7xSnF8FJWLHT+hgNz+k5eru2G3Wjxu/e9imsqtdkG0nLv/vi3U
+gEoaEbrMEVs5N2AXkEEWXs7WetFabifPptC8K6U/jFIIix3fg6+FyvAnbuFjM6b
zGLD2mw/vEeIVQsLa5rpISTSBoaXWdEDklEqrblXECB/rvpZXm1eMWBU95tbcmz8
SbkJzGzHKllienEBTQsufSE6bzHnMxxrjj97kSxmU7VloDYBBHVKRNbCQDovx219
crbiuuRh9tnlsz9TPjRbqdaoBCXfE4t4OPc0RZJkBezr39Ohvp1PNlE3nVt8kr3k
216P6qtL/oB2NaJX1gtFDOTDvV499p0eyMxD+3QCzP5fXLxfVkvbET75A+NxrWK+
eGD/YaUN3a2r4O7gHVRn7mm3oWuVKlRolQhNOhOCnPqXObjLrP+oMexEzIKSoMLz
jv3Pr81zAPXSLV4zQqjEStXbkZrL00A8K0jpJi/CkKybLKVX25mBChaODlqH7P9H
92Ku76AjcGlEerdI2L7CQgUjGAQrfJd1/rmCOlZfZ/NrDEDA7yc3T+fd1KVyMnuL
zgmga83/lbGVT+0MojROkHTwrirs+wGnkXdn+Hoa5j8ADFeVlsSypc/QQMS6jwq5
/0WenMaTbdSOBiceuVdLyNcBkqs00Dn8vZldhWhQQgHI8Co7PFgr7uKqMpLB9d6e
wunPmlJmJSIclbBdhwi3uETOS+YJKmiCyeSM9xOeM9EXwBlZQiGgdFoOx1wgZv0S
iYvBFrfasaWXqXA/YAXgkMAEHJ9m8xYaRcROiN9eeHSubYMQC0haQzT3QrTj3gGP
xDQGUm4hgJ+qVmxH7K0VL8lTTYAS77ylXIuczGAAf6St2NVcsNL99c8IlN5S/kAC
0KbsHbDfBOH0XiIZO+eHWTM3OwtNiPP/QyOZ+A/Ne13n9kJvN7AkwPNp0G341xOj
DbbHJ7ZfspUcZcJr/9F+IDv23hdwDIIiajJTOj7/yVT9/gGd/NaR2Oo/spI6z4Sn
wL7OSYZmRGOcWZpbgcheFDDn5hVORDbE0mAOYW9316PMXfw4MkpzGdaOi7MQLuTI
K6WNvZ/UfI0Zg9/1jJ4blLj2LknYbzmCe87jHpEcIZ+QGxcf+nQK2ONgzRCKQmBk
buvpPt1uaQVoCrBzL/NW+USLtUF8o2ZucuyKLfYhhdJ3saHrrDpNDghcssCcvWv0
J9wMtbTWvsmSiOTVeHw2xuU25jLTAbWYnNucL+vHkI326KWUyBwKjLsmh5G7HdpL
6+g7zA3/lnIA8bz+LraGXIyOq5oo7V0mv/DJ/0IUMtX1T9+uuyObxBhDTJA/VU7H
+2OuNZh+QutHY7+UTGpjUp8FYi+CHGXpwFKNY0m+j4aKVoEg1VHWNoSurscdtc3Z
mC1LkelEUTym7Z5oJEFZFjw9sL+4OMUcTFpO0Emc7XZs/wXJdU06ZvxzOD6Jaklx
3MpNpOtwHFVwgQ8Hf7ks6eU3fZcbLmkkWtgi8WzDVFuhHZKxuMX2jHd3h7ZihvEH
6tZTvcXvW/vpPXAj5cZjqUfDedvU9JvtJMT64e35XCCZdCm2MS6DEvbfCbZNFuke
qrxF0JECHiIV8VDaMOd3RzxcsWpugrGFf9ztMwZySeKvdDPuUqxiOHZp9De9Fmu9
Y+rKW39zit7kkUW9KtmR6ya1IIdMuTd6fHWUb3ox868aASyKeQ3zzT8d5S/a4u5u
9qmlREubgjLiBYNdiWm/gN4Q/IcEmq3Xecta4uR2DUOkr/t8rjcgxGXJNbtkvLtm
MwBeo7Oi/UDAC1Iw+S9aWIcvOe0gHr6R/cUHroBIfC17ztM0E/p/j21Uvno8lw0Q
T1rJ8xjr8vanRsHNbKAXH77nZs6xXb91NzOfX/KKqtzYnQXVGG6ESGNOwVvdPpvw
EUlZBkXx82UeTe1rAS0rdgGrGS513QZasQYKMCpVgWkjfJs/c/APQ3F77xsFhw7C
qOItFTFAXv1Fjyjp4Txt1WfQuGlP/FxIAN7BOTSXgqqr657UI/nZeiQXrAsHZ1th
CkPA7/0JfPcwnwRjmOyyc1DrK49FifT6xZYHART02QIHKay2X77p5Hm1SnlKsRVq
mm/mb1gQcxAVruIxIcOwON+7yQ5HZhPANYJWngBL4Nc3HyDgG1lwJf9921uLWBkc
8VXfyZOfpd9C5yOTbUt4ashI2C3XTHYWv0ktQwGIvwDw05hulQr+piItv7Zf2Exy
/IuqgmZOZJ1qpJKycM6vgF1GRkW7p/bzNd7vu0P4OUvFfDS5JKyLU5jhgK9DwBcK
II4mr2yniOFcrGOx4KBVAZRyIDPRwIQ4InxNdcBfpSYbjnUCU7cA8BgxLg/TbWyD
ZH/liPoGxRSBiqr2eek/FTpJe+7pkLKxuLWJd0xJqJpOrHU1PihvgI+A3KVq+0Q1
WHdx57bl6WXa2dxoZU2Dg4ITkk7yYjhPpTkk5PVCNDprWQwJGLD7j9EcrC684RjI
+YyLcmichw31g59FVs/oyealmY2bnBV2eOKm5QMUR99JDE2QQt+VH3eKOlVECKs2
ZBQvtz207LIH2VhZ8ec8pgCblRCp/H0d79CGBCR2DUDxqkQrLsEnuTqXGdIxkOU1
uMBnjqsOYpqmYJkYUakuAhgbwqb12USHj5Kkv4c+GtzQvgZthsCegewDzOeoizw8
DPmvfLtCMzrrnI7jKVyvDTKEZO7cJE8s+8ClwaCT3gljX7A+QiSPRIvRyWOV2ah5
zViQFpdIja7aU1ViZ6Iz1oByzz1bBcU3FQhkDpn+xwcBhboHyk+thX8KklF5g/eK
QfOToeYwdPZdVYIo1jbw6nnK089kNe5DDc1gCJAxa9hvTSWvFevesw7pStjluy6E
KIWyegGus5PPHTEw3dEltPAY7jHHK1PyreBcQGIxi5y+30cyurKigpQFvve8PlCa
WJe5IlUjmanUz73LfctX9SMocnFuTRApC1m98vneXo7aw2HHBiF92APQRXZOzSNC
39B7JFvu0WY4s5IkwwUUWSxnzdVcLNi2Khb1roh5211i3m8QdpIVnRmay1kCZJ6j
qDhCCTsLk+YCla7eloO3bYPP6ekTkjrHUn6XMXw2P/zRVvk+VgXf9vNKavZdTKAN
2HwV9INZzbhfN4SRPFJLmA7FQoU8uYdZyRyTT4KbrSnetg4fwSqPb44cipO2WMnx
uMMjpbtWM0KVGoW83Hr7kA3QF58fAkFGwb9qlasfoHWnyqlpdZwqJrlmcOLupS9o
ngEniplBQ1IrObR/vrYuHaIWsbyAtGvDU/dOkbYe09luLIsZJ/qswlFRkunUs//J
BoCKvZd0d0NTIeTxiQiGpVtlJdmFLJRN7avaExDByVH0nrc9ebL1uO/x2mJL27L5
E/8KFlq9/CwbR/92nVM+XXe8TsSdThAD/WuNxgjANeRoyymH5asg1xdRtJb4qQUq
ed2z9A6OerKO1AXehoE1xi13JLPDdsIb+9r9NFug4wbAufwTsy9sTxNlGiiZoz03
VUCtATffF93nq8J3ih6a+D4LR9Gsl9xi8WjJ4mGGuqRGfjEiYIW+u3GMigqXzQt4
PixZW1k8nNhejGVKHmuKj9AhxqumHPGDm3JFNTGRRoLAWEf734oVLS8mtwfXW8ry
SXyXZwcuZYR6ryfwex2slD0BtpBpzxsjHaGjpjqLJ/pOm5KhnzTJu9uLJL9hSIs6
Qc+7SJ1BLlMAiQhDWu3gxs8C1Te2tF0kdluUy17MYIILnhm5d18aOvE4PEDCFwpF
Zd/kPaLqgG4HTlrOg0s9WUl1vkaQm1830MNfC5Wxaxp7cj2pyktHiIU9iq3xzccA
JwlHIrnmLOXQ7MNprU0YOb5fFC54Kkk4JYj/Zkko51ANahlQP9p7uVM3FyMcw7UZ
82hda0RnI1Xvl5UNwr/MOxbDUXWWPsk2ie8VUr8JGpcrG5zyntkI6nx1QZlWapRh
jSdYFCAHRFurw/pfip7yKWxAh49VzSLnxjrXwuBlnDAbEKye5cq3g1VTP0ikXhUS
hCOIsGA+yYBlPNjJDwNoM0gEgm0ux6ljeyuR3g/mcqXS3wH5iS6JHqvp4rAXX3+a
HRjyRBgaiUV4oVH3ngMu2KS1/35vXrRO94BqWooxceKwme83FVULrP3gT2orA7OM
TOhq7IEvGnA1I6A0NFRcnBr+w0HcVjs6gGIGvdTQ2ZgRhi77yVoGIOEuMkpiF5aq
x0IZ5ZNB8jd/g5VOiuPlszLTK3PFy1j+nlVbdtCKeyodubk7gugACsnFqFOaUWV9
PNH7z7m14KqsvbZbfFW+f4Y5zmqYyigkeXlm3z8xPdMqzHBM2zHazOZHh5RgLcrr
deeN0Yp2Npob/kCgJDbi/J6w//QlmDO9RgIa2npiByUBbdUEJQKH0/t3JBM0HsOU
ONqFXlSSfXn/GURnNyu+XESY9bdw8dv6zReoSa9DtgkxIPlo/y8e8Wob/FO8bT1Y
RcHMfyTbx+7xVHL5m00/Q2zhNyMCEfsjOkFVCYj5sDiwwilt2bUFBMJFRl7HngdG
yHPoO/ySSMa+/ahS/xmEld1Jxnsr560Z2m/juOMiYlu6kEFi5xLqJRo7B4aRmMHI
rkIKB+KXWK+yoW3fhhvhsmRBywxoI21Fri/DEeuUsM2UaU+YbG6/ZkvFrcUA6Ha9
gp8G6MkTy+om/tqbF9vJq7LADeWHpPbGjuNzEf39bB/smolQ5+ENgZ2xzlyX6gZz
XMJV/V4ALIhHLrzkoCBCKGtHfl3Yq62f88eQw8CFchmy0CFId6s6YAj4qn79sApb
VfI82fqJarlVvMJQTMrHdvFu6rfCpVtZcswGfn19YDKyHddXmQuNHXpmpJnrzCfE
wto3IuEZRPwvxBgLlOG6RdrlqE4P0fkzJCbfegdfy0oBkm0wSNRszHfSVxUtwZft
fTTGbzpdYfh1B4Efz0hxcjRZhfSSsM6PhvKtqEyRPZZVY+ABbY2sk1wkUktqMDxl
lPaXrWdD39Inc3Yt6yp/5HR3w1jNfoq9ON47c7ebOzn4Gqer9GxfHEvdru67mzMV
eXs6zK0LmTUBpGmEPRrBqlcx58Z3YitSzixjBO/zJcPuFlAHn5eCU4yKSBhf8SwA
tEX2Tke+c/XqQUVGvoZ6Fa17n3Q8C9iMCujY3VmiqC44//DSU2YTCHOjVuWrplr8
rFhUk8Qjo3KIavgryUJ06WOBIVioxoLz6dotmPOJQcB+YdgijrLCN6aaAg1ChK/5
xAsdbO6/7eWvEsqEqRWhQ5jKRT8UNVCYdX3GSD8fyfCRgO1CJLgJ6A26pvyjO18E
zLn2NJKepM0Uvr5oh8cJrKiF6BEeYJVxvjE1G0FuqQLxxLwyhYqvCaYNWLoT3MCC
jkjHhFjjdXoF8AOTORwRz77GtQu1Gr5VqmzAsHOJsoYmjRixomrpRRnMIcJ1xjei
+BrrMqmQiySwpfgBsNdl1RnA6EE4oL3WXs0J+S4cwsoOoUApDBcBKdMfaOoeMl5I
i8BvMbwwgPX/KTMTyqfmo1R2SGcDjKS709FQ6Q7th86XiiZNnaR38WUs6wM7QXBe
8+G9r4KuPjCNEkysdo0Q/50y9ntKHxB2JV7stVxY5VgUv4GTeQYlrLVmAMybSl6b
0p2xSY5b8x2ARlfNTw8hTsfrpLTWFrLHiiW+1ujD5tSp8d2mvMyDfcq/phSxgZ7p
9Qbg2hHktTvOHnZNxAbXx2nVI5UUwLH5TAMB54KLFuQE3Fs+Clg1yMsZt8Fx91tO
CVzB6Jj665pnUxTiDrZtRw5pqBlaiafNXl4ayJc4JyxwwvtHNe9XCTDokJKOfiCA
b+Sc1xggqEALl6W4ox6MhKkOxJJ77yLUxUyGvbamQvFKVbD0/KWHTtxhe4RM3Hzx
Wjn0ayxw1zn+xsoeVQa/iCPo/wI5CusWM9AiglfmbYn0OXV3F/uPmhR8LCacQfHd
2HkLoX1+vTKQUKGjDtXxJ73SlXTYa6S6LN9IjXJoeXqzstz2xk4v8kHpkMxvPjlq
ORtgyosfb8tJYGXhMAZuswY87jT+UVgVkqQnaPn6v1hsFtHphWixoFwOElRPeQUt
wngLWPIkqlhgfg4LCvZ9vgS6ngHFmk/HdaL9TZt+2pt6X+ZqlneLRZegDRK8E7vV
bUKemjHRab8mVDn5Hham+Eu/7cbn7fNLzz3REmWMOKrWBcZn7j0i3/DpN9cvfl8j
SO3KbfIc6rCy0lnzL/HUSblvhtwwuNYhF6yl5la3d+T4MuS8BvcvewXkHyj2HJuE
qdFgczM2Bz0iUWLEQwkQfe/tIRN6KlHdrvXUQsTDRBYxGIbc5PJMSEmlSZ6yFf3i
hssg6j1ffr1twGlu4eKR4to11VpqMAcJveiWhjOxIDjlsvehNwEqW6ekLlSLO6nk
lEvVgzdF5ojOabYZ+lF8iyhZGxeOFHM9AKpsrv7ZgB3fXjT3R/MiqKizk1VCwwGS
7rlU0lBD1exr7+zhtPYkWRs24Q1N1Mj2C7u6JFblciqdth7Y9tjjl0STXJocKmQr
l35T5nWy9f9RcmIFy5bGcbOYlFk4GotkfLFI1q45av8GcbglDRGjyqcbZYK9rw7G
gpkMydggCHqf3c0VU8Ul3HKmnNDYP3UIik5ZgPoeFKwh+1MvI5rbl8IVytAz4u3L
0+ZW+ff3+RVr9MPWRtuvgd1+D/0Nbl54w+0h52FSnKFwK4Y23+UoIbU8oHY7/099
/CP99NHFxMDT38V8LNoe+eqIwp8vunjnRB3BJum0EeP8v/lwMYau3qk7fnEk3c6e
cY1Z3zAbRThSNrwo4ynideM+zyYDWiM3ON24KNm6ufP2/6KSz2tM02OQjEeqRiN2
AFIYswfB3h2+E1szd8Wpm8tnWIoXjd5V/iNes+QP5wSAV7dSErqofvdh7Dqv/Nqb
F8tKm6dfHvGbxKnM65Bbz6mUeo2BHob5fUnsuc2JLDKoJ2bmjzhWNhSW63Bzxa8s
W+RNr7Ueo/Nu8MZY+poEI+BwA9sl7PYutQqsJNCtsHxxsE5logRsamy02gf0IrZf
AFKwS4ion14R0WnVoILQpp4klwMZsDBfhnCh6izWOC6OHbZBVL9fJUsdzCVOtmZ/
pNMFx6daKWk532QIrhvHPmeLUG77+POGPfmgjJ7IoxpJk8R1+EHYi3BusmEO12/S
dxq5HUvCVIqgXdetfRSXYfaaQjlMY3mS+Dc0URGlZ5Edm9DqOchXbHMIws9D65Jg
AEISbm8dwKsm2MKQAPg/2xnHV6jcOBPmJC8wQ0DpQZP8TDvNmlqqAK8SIF0p/wKR
UBJvi4RaJ2RMYYb+HH2xmjle8vM8izyuXB6qEW8SRoHBCXKWXQs3WxB0+pf2F3pY
cvdheRWfMLni9DxxsGJj+ogF4UTSYWxGmT84uCSpsSGLAO1pzYCqVY9FAp8Sti0z
ebUVqk8peISkA0o0xuiASyWO9bP8GJCw/yGJ/MGrYlYWalR763EEhuk6OHLTjotB
hYNuqy7gPlUXHP/cFkU0Q4ysd6MkDFhmchZkxA1ge+YGgd0cn3NL3h+sWwGC8rJz
dxlXFhD86pIEZkCEUT9je1NXopUxAjoeGp8f8hp/lVpEbrh9swFAj7aebBP7t+qv
/x6waqW5qOAgNL5p0H/6FUey+aRF4xPk9lBaPgSeZv6f9jmxEYRbPW+YxJ8m0v9Y
E60nI4zV0wQgsGFv6nOdzZw/dxE5vk/Vgl8A/Cn6IjpIhsc5gunycnRE41YXOB6K
FNWgqw+L5Q6MDXpMsL/sebd3fGByT03V0enk4A7RWPu0K5P+lg4MVXV8UPDk5WRg
qJEGgxpQ5Tb2MnIookRwGfX/3ADoZ6zwkCxHsas+/SJNSuSiuZPAyTRYhZVsz1/5
O0HgmKq5kbQ0686bUUStq6eC0YXzQ0X28EACyc1bfkNOnjg/S3CupC/VSDgtnnw1
+LiNP8OmskFYPAwlmGE9BtxD7GdMUp4kx63gQJQPqwFDSyoJYQvlNpaiTmpbUmPJ
HhEhpUgAVlkuVYFGgl4BTfLR+8pFFt7IzUTe//OgtO8cZmoKREUAIiA8ov3Md6WB
B24/L66THHKdoPMTOOCjbki4M+thSs3NOG2oSxhVeScgAZ/eU7YaVS4ElOVMK7t2
h5G5Od8ERFHN+5ugWn2bT2h+JGiWBY4iCbyetjiaLVYkaoo2Y0upZfDpyehAz8mm
ByWXOi5+a7cpq6TDUvTtKiGY4hXfY5lJ0+mnp2tUg9BEZF500BC4+Y5ANUacIoeB
kmqdXGV/E9i2DlssWITua3+OdjzfS7lU3xDAyYmk1/MqdUGev0PLnLbRF3DyNjTS
Zwnqfv1TS/UNYgKcDgrHczer8Zs3sdG54EZ5fXWK0KSxsStxnON812LNhshcewj2
z4DI5UkcjUpu95ix05xPfbugIkuNlt+7IT951GV1k9ezH0mCqUEMUZGO1SeLYZ3e
XYYobaHGo6VHkusFLxFjzzFFFlxZEl+1/WYUJ/4MIOF9YnJAddjQFaJB4i1vHQ9W
THthEaEgDxU9WFFFZFQgaIMylSmaOIqlyzAbRhjvNtN/af+UZgwVc7XQx4p92c1A
wy6WxIWJDqeWJ8OweaTMDIwRlU41e6rfCAmAl6ApyVDrsxeCg+tNyAJHoZVze5sT
eV1RryBL1D2J4KWeeYD6YE92iQ8JgU/2ETynbNnmmdzpqplshSu+U5e1/zTBFwmx
icau4tPRmvvgCDJYLMyhTKrBvaXWpJEU2rTvYGsMv5V/DkRWjpyrI80miV+uTFd1
6F5yoPNTOLRuv+cPw9jd/xEivAvaozi3n2XH1aCT3nELpIc0skmzrxL6sslPppPY
`pragma protect end_protected
