-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
K64YAANp4CCts8S/MlLvCI16yCQdFEJEhOWBEqskwy4cUN1ne95K3RqQdVWkJv9U
k4wVe/0B7OuSUmrgMpAzO691BsOgog8T8g8O/MtYrhQlC8fQ+IEvjkSL57sSUcEC
eAGCCqzgiQA3Qvj8flpbGY7d9PrYQFvYzzfh0ftmtOQ=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 12078)

`protect DATA_BLOCK
iG+iWkic5Q4kWyRNcmzup+k/wjYuO0hev2AmSyEafZcD/qKjIXzOSEHLc3xk3QDx
/3WZZRErjkDUU6I5trkvERLhy2fsQfv+qDYAohKij1FIj6UZp/ajoiMKtzYPtuQe
/ZR53b7GMZIQNrtLGkf5nA8bTqpD5PQc5mfkD3WciWP0LdMsU4/b8gysRorM/AUc
TtdLvB8/+hRnMppzUYZOL44hkRo7CFkN2iuACzp/XNMK2mVs3cJRi45A7arE1nTI
CzO+y6ncTa2DSrUsCVoxeiG7nciLvH/Bqvtg+f30KaYk4H/5F/KrJ6pOLAPbJr45
waTrMxBWQ8xcz3ER0awdS0ytmvjxY2Yg69ypMrS1L/YxeWcqHJAzLcfWDDW/OCZl
Rf4GuETAOrLNToyh/WeItgMrCXDxpi6vQUXelz0Ojj1sXZVz27jVnNKAiyfQ+FlB
4Rr0jwmKBiOMnSCme/ocW9pXjXa49NttTemhb40Au99QsocR04a+v6xa2ULL8NY6
PV6N4IAMpybCcTsGL8H51vNotDyBXsBDE44cbeK7kMgymma7NaxL5aop07yfgSNR
6w2AYibi4GFnvJNt4MHhTrE5HIR7yjPZARW5LmWyoB8W4lviwpr8LncMQuHB6HIw
yhfF4gWZ4dA/ofLYgu2JXwkAn+/CStczQNtG87uA4uhcOOZ5TSxgaItqmMLk8juH
2w2BgJGMQkPPVQcI9WJS0Jxx76EFseH9mF1J3lE2GkrDFGMq1YpUl2Oqv+mJZf/6
gVXBR8jwSfQTCOG7Fr9sdTTXXzIZnAwvCwuuKKRzL/dhQlc5ndhnXqRm8ql9RmFh
qFEvkVOtqNqSQR6a0oj5d1is7UU6j9xzTGSqwUo9AT8fCJ+1gUiJAuln5ENWmgD7
zmegUTZe1l3HfhHRn2Myp6yfQvcl1vfbexowMWDYo8t3XuMZlKYL1xVmJOSSFzMd
X/EuYFd7/8vg3642JN/cFs8lk20rD3ayKxdgNzL4K60XFwYjioT6OlYZkTaZvHHJ
A2HJA9gqs8Xo6vorkbDbBsEiZ24HCaMYbtlhI/OWzVU+c5504kXNPdwiiz6QAtla
HMTrvnhL0s5sWtEjNWkLOyaSziiI12eFWyEdnD1kSMCopEusds7hsiaYozr1Gcky
iklfKYyGnK5eCq/gG8Wmhzk9dgjpbN0qB2CP4tuozJpphRv0ejwXNEWknEKsa6Ss
0QUyTRwJEpMSIa4XhRNQj9LB5Jqd+L17JhJo3MwgEPRxqthD17BPF1Z3sbNt+m//
WxHb/iWnt0w59XFimhgIm1mpG0W5lKwok7wdW4v/ABNMrEM+zap1Ac+IZiB4/4C1
myCCRj4dMVEQd+YzMgm3p1mUkYvzD2SpUOGnn/6pBC2f0N8JVZXN6Ed5vVedsPjs
z8O5ZclKDFZHQNg1wOi7+QQoj+JSaJYV2YoLNZsvw2jv56g1XqVGQOTYKyJoNxB4
8urnhrCLA1MXIMoSaQ+8HJuKlxMxNM61LK2XbRWqizGMN7F0JgYRR+ylwb4MwwIE
VMxjvmPkd00lTCBWsut4R4SYd+z5zuZi1N5sWMJruTqcMiEgYsIEkF6BtaUpZJBT
N0/TxTN61OV1SKfVyIOo+317td4AknsoUaCLwOtUlgfXemoLBX0wV4jDE1oWNmiC
f40dgxhMXemQiz7hRwBFxk7YdWJGg0nYmaZ+lmFDj3dXrjNQ/mkBepqADZunQUDk
2cTmMou0ZinQUvuX+97CmO2pg76CmupCLsk/D110dDDLD7wctF6+zbEg1Lnvcq+x
muFqvM8GWGGW3M0dE47OHaaPIt9iesBqJsCscuH3g5Yn3uHtiipyYBw3aFf5+Vgp
T9AshO1hwAlTFmSdl2hcXd7+c1L0mCQWn4jQgbouWbwVXiTPyNjJMcyu4i/C02tP
yGNKydjZfkpksfDCa52c1EKJwiL2nQiflgB6iL05JBoLPA64J6dNaav6t6d2nr5z
7CTwjshyYYsbt9guyDuC44ZA9u8WjbYiVJBKJglp78T6IfpgGFeCrKcR4evM+wXB
psnAV+dCmy24CMe67o7DycoanOMaRRnJFzwJqSooVCtsCtONibd17YIoYJ46/uUs
J6MjhXYReIiFOpkHiNe99ETI/zUl2BY6ktSGXdkWY7Ydx2YWWt+s9P/rWw/4o65h
1AXq378s4OaPsJS2H8QTH2m5h8TRxHsEmUDxge7Mlg1csgRKX1WcXEar2mgmXMQO
NMGbANIf64hGnJTa/mHBYVulZXKb6hujhqDFvRHlvhLN4V+aHlot+H93r8jGykva
xHmA45qFzR9gzJzO86GVIVIzn06QnDYeadTgen7g10OwjnOPsT8YzO5sZ5oPRDuF
FmH7cpMEkanjTQKx8k8AMu/Q/HfzJbcyb3p4JUcgrLvUxFZJjs4PKkxW8PpGkPjU
Y4yiuRrG6HbxJzajik1m2E5HtFOCjEpejPsgNdxRxXeLGnerO7PXZVQ1lzN4lko0
5lbTLxyd0CYcmzuOOssCb6QGdZrClJ0v2e9dyZylGM4sDNT9iUDk/ZiIuuVy/V8R
sOmqutp+nVJwPywYeuyNDVwLtISvU44Db8cZ1cs9nJqUKIS8EuRSKaehgOjrhTb4
GOVGsbAStlQRY0lM9Xv9tBKIPhZs3MdAUa8A0JqgGl1dnv1SIE5fuNGhdUvvC6hT
sY8yKgsicXwnHBpi6iwKsYswPrwqVn931fpzvUFrsoGVhyYe5CI4uFzj5dAKdT2s
6zoL42NyVWgZoAZpqqP+kTKsvdwjm7h/8jkINunc4HAo9+j5UzPO2Ft5lYVgI7PQ
/gJ5KbGv//2oP2VAH0mOhONThnpSqFH2uqVEMmAfmSrSSmG6CuNPZFwGpabG6RlR
4fyV0C6oDHogafYM5ZCaKV+Hoy+YTbppS0sSpI4T1xg66UZP7cXjvPqgN5Sa52XR
Z3IulKAPpC2kD9JQZ31xfegmVZUVpCI3eP1fTK+aStO210rlMarP5i4P92aciBPx
gUNasyBGPyYys5rYARdSSTTnMQezHEM27VCDQyjrKCGb1oWJ1kUsjcOw6nOscFcF
GT+aeXsSYdGazGn6sJBysohmYnsMFmtc6BUkaaDyqL1JTMYCdJgDDHah7r+GwIHs
Frhq0ACIYARn9q8/W9fgU2NfL8TZHhZky8q70UvgssDuy7MBzvElZOw5+1pCl7H/
dfqcqhl81zQsdZSj/sCTME55w8yH5NTM/CvhrgD5dNZjTNrGvMA4yCoGc0rKs0PR
gYAGwtvnDDnEWsGqHrNFWunBCNJCgD4wvn4MIHh0H+qWJCnXb57SHt6YwmG9lkmO
I+Zmdi2PuG0FUar2vV3BkGeoN9LrTVvDCUWkiRU2fv1p2sjsu7PAIY1fNtFH+W3t
Yr4o/86/zNMcwXKL3UlLUsxoW1eafOvmbt/DYLtNU0P30B/G2gdy1bl4nFbOpTKr
0x9F99VPlQ/gTm3IAXMxGsm7qTMoAVAmgGz8tAEjcuK7iZriq3NLFCYltvHWl+r5
JhPp/2Vo5n6Jo3uW6Qm03ybBZ//3hSt+7VEOZb1iDr5JB6Ej6Xz9mnUN4Kawh+FP
W3Qdwj6u22PTcB6k8JFuXkbaonkH9bYCN7IDrhD4fvzOWnF+KU+ZaYboKWLws3dY
hZofeQ+mUJdkrK8xKBonK70RCgbtnbgMzzLHg9jAE2B0Zz1doI6b85y36U+6CBXV
jw65NI83Im66KWSUlTGMx1c6IWfMugzjPsTHE2AsKx2P+x4a+RK2s9f2x0sklv3F
y7wUW3uZcDa75rm+uAQBAY31ZeNmia8ZMB2S00B9kKlCYiT9yLuDoXEoIVy0eZCw
7emxwyGnH0+Em6jhLS/p+kHuSG1KxRIZa2HjiCLetn/YaXj2/uHM/W2rjTkdFVNP
sONKNzM8L2lFenwjPorVMppbn4yu9VBsh8J6hvmZG39vboWKts+mOu5Tlydp2wF5
fS6DfL20YAIPka5RT7AZtvSWA7FRaqoq/nlhcfhyYCXPlEX2Iggh+EdlkRP+o8sB
eOjy5TSaj0Dh4b0A5ThjLhGSGqE4TSIKsq1uaBTlFORMFCDs0jtZ4c3JQpyzAy0x
JZMZhxY4ZnicH6mkUuHhaTCpVJUD10vjzN2m5DKYbQ0vlv5Z9qsYpmCajVrYPd9F
eR+90lBo0af8LqOZpmhALQBh+qd54aN/HyBXDILfvuGjd3uD1QkYt1DRK9/QBXqI
Iw+JqPHHSv1V8uZmOj1E/Rc7hshGRy4xgaQosO0B4e8oEx3ar+5kg/oJJLTV7GBk
Bt6s/eHrpZLDce2oNpEYM9rbboLa9vXMjztlSp8Su4bCicl5dmVJqbikIY3lNBW5
KFwrBHytbCAE6BFBlolywl0SFnB8y1qIdhZDw6TrV5vQgQPo+UrYxQmXTU+MaKH9
lnRE9RmpvLfQWgIB2gnzHe/BDBiQzrH8H9k6SBzOoQ9GrhoR9C5jBMDM062QIY4K
F10tYFIKTN3c3WyDxLgBPhwxsDAR63Mb3cdbWi2JaHdCBjG04WTzNwaRZt05Rz39
Xd1YMr0Kb27spVRnVynafSP2QEc9bRkbDp3vaAscnePbO1ods5/8g+hL/mUfbYfB
aM6ZhLr/ZH8cwYVSfCagAM8CzJ1HIZS3DJdJEukpFvhj0ZJiL1n92THEjUPG/59/
DhbHGKjxSZ9vmhrUPVfCFhnA9ZCTR2ILY7sU9t9gQ8W+XfG56DkYYp2IW3UVr8Id
yoQCiWaSO5UOc5GuGCO4TygiOr1VKzZUkWxlNsnSPx62ABZKSl0Pf8ApXFHPvkSs
utRgEYx6cOD5vrgGuElyFElVjk73BbLL0993vFyvLCpPOnrWiKhsZDq8bBUyiGf3
redfWBgNQUqyzKISuX5RFPhcbM6Mp21eK4ODmDLzV1kEtrWcNFXlUgDeXwcJtNt6
AtpidNq8ien+sUZUr2NysJt1bl/gJNp8XnUdBclJzxfV5U4eDxd2UyStVW00kW6R
gbcojA1evIlfsdO5RoJkUPLisvx3ZBZ7PJ+mpY0ZsP6d60GUJvB+5IBuPaK8XPJI
GL5FYs+Qjaq8RFHuZvIWU6lyUGpvka8Mf6l67fnlkVTdmtMbdkPyNNgTds/ZIUCh
6GHJMkWRnoKdDJcqxBrPWGIHAFNbh47qsd/Y0WMAsGIwUt0MrLMfgkSasZGL4lni
SONUCpYAY3PO9A9vgtxTqZxKYTJCvURprmptkQ7VZq1eeuZnx+P6m78IIwUXEhUr
r4C/Y+z8jR9J875bYJUFMLyns0m9ldQWe/gH+d/hW8qL4y3P2kYHjfb51Y8AJEau
S7SbB7YCGG5vLnjQhWaO1eXpv6zFNOPFJ3WpkOuPTuRNnflLqX65I0cfPT0pLDUt
lDwN6Db+y9bctgHLUZiPOq/2zQzoRL474IOxm/w+h0QldLXrW8LbB9ddmbnPMvlu
JoVGBOH/wtbXfpqAW+KbQdiPvwyC1mv4uoOcJ232dA1dqNjwPohV9O02flAPy/st
CsQRqntB9PqkSTaAhMhYQjNTdhjwHL3XdBgYojEJ3jhvGgDf8VfU5BcEAh57F/Ar
F60kZ04wxuaHhIWqjpxxp2mxKwEI8ScAoYiZF7x0NHdpNevVtTTYFFlFpk7s0irE
fqrrlM8W5o1w8AMDSpHCYkAcdtIv9ssy3rlGYrAbHCann79HaI11yBlLa4rEJe0X
DTL2/fU/Q516GwA2DKyJ1cXqGLMVJp3d/HRP1RRwY6X6/bMVaarS4lHmCwpSq7LO
EFnlAiLyS/Hb31Yug6Nog0BO3uZnhyMrKZV7Km6uC/6+z4RMBzm1H6qoo/Oq9iD0
ZG/8bI+0ZeAy7ra7ncFePzNCTOylF89hA8C5n1pZl11L61nBvjN5eaqItz8LSTZJ
6hPLiTTv5KX1iI/YMTYadaB6bWih3xrX2s2dKnKKcHNA29wZW2GbiJh/16CgE+2G
Tw8VpnlEaWPVsV5MqiMbJqV3CFg/JAx8PHZCUKpOQpw5PC+Rwm8IUEJ9RnFkKuVt
KyIIJbIPdw/Lj5mLstfm8Osqfia2U2qxYcS8sn1ohO/qP6eyODlTqHfJB/KZ2SPb
g+JdplrxQu3wDLIyZaUA9HAljBFdDzd+daYn5oHUM8sB3igUYcg9E3mxKAAntCAK
u1i2DOviuiNHHncOFG6FQtgOHxOmrOXbnyfbPDz+Vky419kPvYxIkvOkN/7MqXZt
2290v0BOgy5qZixEIneR6vr5FAtEdDUFQYNX9PCikJIXY/PMKIfDTObnDnWGRdqW
mW2qjjO/1wfB1Muxhww1ip0RVZHyLjGbrs1FuqJCRG+gvqHU3SIK5DuQvq2FaOXj
87wY2S7fjJwpzek3NUieQ38+016ubzsVE9zZyixCjgfuJQuTInCiOE4IRqG4VA7R
R/Ubfho2FFGsoURsKkKTIXxssC04g+gWog+IInexx4vy09iV1E4BmAnpYnDOUdn4
beBqzQ1ZQOb3/J5Sa/9/03M++ZqE6jBFmArcheb9uIgQMZvk8jnRmT6M72W2nmGl
zkMzzj5J8xwgNk2Kg2cJ3hVWX2+RfbvPxsH4Y4VnP6DOKHWx8BlTUtdO2S7zSZ82
wpouRnlwS0F8DkMn3K9+lQsDnjoWrzn4pepsQDYf90txQ9z/gp4k3hReurSTGHSV
lGWK4zGPxQX3sNlVTWXi061cFhM7bPiqM3UUNhyr7J/ooufae5QyogHnUZAiWFL+
dM/PcYJkuopmL1u6JwyV8oistagt/05UKkkMzbJ5xFUjZiX9LdjOSPqMZ37GcEYo
oedPB762sqGmZFZEQasxcm8Tmd/Vd28j53O0wU01WKndTf52WuFrJrQQq1yiV/EJ
GiPcapEUe+jHv8X+N6ngBeEixYI+QQJjADKN0V+v5ai4UamCCTWFuKJfv6c046YI
7TIlfzqYpzqUWMiid4RcGFUOm1WpnAv9dsx+XW8kCaVY4FCZ/eXjIiX556n8b3l6
I47qqe0Hi7xyIBE1wa3gJT4sTYTe/tHzXSiLKxnGcu+tfSpUuF9/hDXGXQMz9/6H
N1w98UfVmX43xn8DYolAXats2R2mSKulvgh1NQ1/acsPp1AQqNKpIwWNJvpesNiz
grD/jLS836XpjLMJs24OCZqj/SiMqzBQ1LVm8BxnC4UAJ/f1nxCFLHZZVGwdC/lZ
QIRGIrElfayIuQpqx2N/h/pZcnoAKsLjyHQulYRFy+zV8WN7jVc+11dacv2zQyjr
VXdMm4LxpAZEMYgSuUVmkHR0LGocny/K4izPzMa+gYd1xc6Zix5nfXpJu5gx3S0+
5nHSBhDrFQwFid8bz2/DNs5Rxk1rNCfpJoyoYuFIAmmZo+o+rBf2px6ctYHAP0Fs
Oz0N89shnxkbMSYzo2d42g1QC3o6BAh7EY11ZjuRvlE6rA4ESZf3b87WGuWXwMB2
xbor6G1OkMnq7OC7BelK/iBUIq71Viik9qkjdW3UfCKQRbd0JZGLgfe7BRcMl0nj
V5WYOpyihrCnI5UKX3ghJJ1pauHEvr093ge1M4Y8N9JL7IqYub4mQ+nURUV9SNYz
l1my2NdjQo6RIELpJZOVgeWGiASLJID9pRewTsdC9/ePfNoQ4cFilG5ZWMqAduOE
Ul1Ih6q+CoviLlxt3ocZgiChpcC8eSKsG0mlq6dRWfdZJG3WMGq8qMlysDoZgpup
pgCKYfSHaSLhVe89Rr74UMKO274ZH7fA7ZMy4Ipv4H0jzS2rNtGOaMv23KZiJwht
g4+WHh9HisasCWPpwqMRXt2mVRPIx+7YwV+iTJUo8kXCWKEy0Xb0DXh6uxA9O2mO
7SegixIDXw18fcGPgIO6Ig0YkhTjbWq8KrpXHNXEouZAMEt/IJDrBvcyUoyXV/NP
y9ybKdYFlOpKiGNWNWw2NU+3j6Tsm1ABvtH5I0nwDrLTcq6t0ZC04VB4eP2k7wxT
0vx01RWL+OTfn/oZFPQR2re1WNu9bwdjYldM6sBBhHICoeHFbveSMiDexvYklrIu
CFvWJ8VOaKPD5mSUcb5F5fnRfx85zw2l6oy0HcyVhlopKJUIX9ezr10/aOlB1juw
AbU04ZpOHN3lBrPhEg6yYYvqR0aqIeVvLUAnEw7SLAP7c8o+iG4F27eWbyojh2r6
0fYy+MJVJF6TViZeNmNFjc9PSbEGhJwm1xjX0Eve06EJQjTE0AYrXnOmYO3LbQXH
WQqi0sgGTTbs9XDAdisJCnS+n2Em1TVwYBw6L/QsBZEF5jwHGMKrzl6v/bjavgQQ
Pw8KPMmOU9Du/dhVC3Puwa96Yi7tpPIvQ8yJObvG1AtJIYIIqGf+ybEpWqHrSxH7
o1fW//t4a4M3bzNV6s/DG/4yphluvIFrptjzknnHA+6QqiNQXUi8nq6+djzpmBT4
v+V8uR+fRLdm4l57fKmm5H63WOTxY6f8piQJoox97qaV4VV08yFvXeZz7vr+HevX
XZFQWoRzaWoySFfdJrUFTSJaKZ0rGh3JRWSXeyFSLhsZXhh17gYJAJw7iOSmB+K/
lPRpYNGGX3NqEPQt4xvDBQ46oV9h4EZakNC3/eo3duSulRfcZruZl1jnngXRQZgw
I3YFW2GDy7vvw29qU+/exU1byhCZ2Vkc5MKC6ChRJlu5nukxTWfBee7/kUI90Nx2
aLFSENpNJG6XjxAr74SOkNdjnmt8w0p6tdmI6vKLcPXRZmzq3xdpP/AO/fqM5B0f
8Y8teGkLNJf1/CNwGM4aaOTJ88UvphKXFJbbKFcbLf/2p5+07fbe7e6f3YdQ8EiS
BKZJXVEYofp/i0sKzjgcoGoe6EG+pLTs/VbZvQ05AAmRd8E/Q5HuexRHIZg+WFZh
ibmgnNKYpqIojKHxN1uunRS33OVWB56CPdbtUL9w7931L2maw64GuolC7ZUo48m4
oC9Hn7f4Gp2YGyVRq54X9rXY8YUI7W7ZmCbGCzwaQ9X7hVYqON1VkfCKC0znP29x
YIJE2eH4s5YjvpoRnlcQn3wv8vu5PhDfSANZwWcXp0kw7HtVdQqT2tJmNNDvEXhg
QIFbO9lWm1xz5Rg1/ylgsnvY3lpqT8zIaugy89s8R+rlmXjcjece+Qv6AYuQm9qh
QMOLml30t+Sxtg0nTVJ2TvZoqiaF4ikJorrRSMAUjRnVGcxbQLecW0kvwExo0PBS
YtI2yB5ejD4SHqvoBGDXH7oiFGrUlBvrcyDE0XCWdwqee2f2BNC3IQah69xLIKua
WdtEYfIkPgzvpLmGZrT2jYse3WdpHgUyrYUI+U7elah4hmEAZZN04LqcKiQbp0E3
wWsUiVQBX3hPBKYJHgIpBRWrNBkrh2XxvyRmpb116npdMuYz2RxNJVl5YEJT/Mdy
ySWYbw0Yv4qt/blcJPE7xS3oq0MMuzmdsU+auMFqxHOZvo+LT0xc4cwEXhN3W9qa
xLPTIfMPwWh4KXvNtIT2JhxvnP7IY4MEXqhS8Jz/TyONJ9O0gQSX+mtLfaQKs4jC
QDSuDXEukDHGHUvJslokGCdKXHLlRGGxcNidRov7SUvhydPUjXcaohGmOPhYqZx0
g6dGJESrpf4JJUOl7JZcXD5zH/QgVtT+bUjgUqFc787C7TXhooKDv1tgd+SEVFdS
XG1zumfmkSnr9saqbz3cHTtrM4MoANYxEyyLcMaaUodL6PKebIx8NunEnIplmnFb
AyZM8MnZyvGv+e+11ciaIKofnAJQSZy424gv+RiAy88aOORsGyjQdEB6qlLe/rnO
HvzyuQ4Oel4ZV855RWTJ+mMxs5FlBB9RM9b5DQF/V8+OfqovKjt0nt7sERu96fpb
KXYEKRYK3waNObAvTqzeqbtkxsFawoMzQGXOKThhC7g4NRzfZiwf5UNSbsuWsBK9
4NTq7snUmwshi3dkWslfffc0hZh4muMiPBIVfSQjQuMMZeA3jcNNU5MGhDSFMD1Q
4shKNH+8u3z/s5ZpA/EJyMA2EFV8I8PIMV8c+p0/Q9M7PZY1vpgyOKQpDL8q9ddG
A42wQFYM8ZgQ88Tz7dfBYREG6EcHZ579UeV5QGYfVPpghkEB9PZKsQDnLrmSwx3U
T31mp5i68YwQG0Hr5sRuoCP6F61X1A+z9Hq5WFBz3bYku0vJrJ+uC0ZmuJXzAbMc
oLXMp8kFfvvU7xcQ8tsYXZuqXN0ZNE7U9m/dpNEwCZvGqppNX4Z0SHhIDquNWzcx
CzK+QJLaloTRjxMrckjDV+J03yXch59MufvSyi3r6gC68yfXKyvSoa0d5HFe5KR7
ko+SSOJN6vTC9IinDuprqR/7LunSnJb3gwAmdVT08y9IjxBBM0xABN5Qmpdj4Zhu
FSfLvT0g90pFfWOoWTFeyIZZryp5QuO6DfQeuqdcSNwkuVyD0E2YBwy9BXEjWyn8
nbnW8sUwUdR1zQtr0wx+KBSd/VBLRtGdKnKpnKnY7UKiOBcpIaoYQnbXmZowCeXl
gtvkmH8PJA2m1H6NxvW75965T0H5DimPGb7+f+y4HLC5SxmgCU62qW2jLuaxcEct
39WNAVZtDZFH/t1H+pWu/ZzsQySGZcjjNGwyaPSY2bCfGMnPUxIqyYuP+w/YZy+H
Oe+Z/70dwuOD+kjf9v7Rh9+Qe8HHqfV8hgoUZSrPFUxUiU4m5PjaaNiIQmpOr85j
he3m2sY9UasK4Z0eEMU6iBF41nDJqnl67q1VRKzQEcjUq6muU2MrylxP30Ju4iED
kNq3hzG0un+qgYkxy4w1N8w8pKJfhSwUDoqVUYEHsRy5WaJtXFpg4F9vxJ2uCPxG
9rwyyEFiuzmW/jTqrUwPf4BIno9jcjwq3RwuZIeO5IRWzPZYLoD7UuKCj5ZNXUDI
QUKPzY8dqxMBQDdw03dw9MMTslZaV87+XGNh/+9SSqvsAcFiKZVb9n6BzpCR7/1Y
jBlnxgr5fY8VzlKQFexcSc1Xk5wbV/umsEAIkalg/zunHNu2j+3l98bTtyn2bTUF
FYQKAfyN7iDm8xkJ8MxaZAVqFEVtB6xeCLRGJ6XFijuhGA3BwKZclC9i+jwNYDKR
2xr2PnnA8SYhhrLmTG5t6NL+cC0o3RVTvGEg1UhySq9ekw56fo6+MmmEeP1mCbR3
wwSkgmXjcysCOXnRhw7vdvgMGp5UHYuzTq808UwL/IEu9k6Xkj0AOhj/g1q7jIwV
ECfnC5dPk8wvCLLKuQtCMa5DPBQhKF4Tb8NYpra4N5QBxdxVrH++5kEZJ8FtV++2
kOeBIjVp6DxS5NzVL8LYd3bMAR2KQ3Ja9z/xm+UT584A1UKvXMgmeKpnkqUPUlDA
Y5vaRldIp6mL7PmYeX5F86n67jmgXOuh5OiSnD45uvxlbOr/8l66q8E6GeL+Dty5
Y8EbYKkFlZsoHBrLOyZN8ZOKuf1MudQt3t7VLVXjmR30YwKrAsPj7tJKvNEUDlTO
QqAVhvjkbwiezmONGNndsgbPqevmiWvw8UvEh9J3RkcS0BZPXb4fJqWCzeyRFyGr
nf2PaAlOfVHusUxZgBn8/KPzMqHfxjzgTFvIlpwiQPNffWo9RETXRQZUX/Jh51G8
ELdCpPT3U0PDnn6HMKfw6q/RoFtUr3T5FgeS7w6EeWu+SSJBOgVvE7cQPD/wFBNM
g1Aw4D2tOrcgMS1QZOYFzBmJVYFBXVcQnD6WHMXaJEAcWRmnBR3kRvKN6Z26uVp3
pWvb3HfKTS9u+cDsLWDalXx/9r5lP5Lbi5ESMRtDcUS0Fsj0wpM3KBMdzprHdzkb
OAlZKJV3bXyLwS8Y6oi61DrfiWEe0KFmonRX7hZZHGF1PhHztDwr1ePZNJsm5aFp
JbYfxzQ8bhDOD0ztCKjMPWov8tLB7VzbpmB5ZSjBgPEIDN/IFH7rP/n/YPvUCeZq
Oa9b5Ys8gje0jtYORoBTNmBszzmBixyb5HVRBFyDvCCZhS/ynzJBlRpHbcG0H0oC
dSkRu/7EMFg03KmemHbPVSJlY3A0tE0QTzYKupW4YweLO8QxVeyPxqo9/HWlXoOu
ncT5kwDGtC+Wn31af8SGlolNtBh/KEtJnLbBjSrxuU/h5U71bytwtiT+eKPiBS81
Ed2+dwKk/SBgFeJgvpV7w9PW5VLoACmFuuxvsCNNUt8eNmAhz6c1VyxBgDWszBJH
/GsDZgXIThiDjy5gCXj8MB9BRUqUikwuk8/YOrxk1wsmF+NtFIKT8Tn76Wr8ZLaY
bDyOAKWX3jI7hyQ9B/ykzfuT2oVOzW+WtATOtJPB8+5M4OBIYS36oW5TcZxmm/fc
Eztf3btz9i1j4aLvpPuG5j+O/izFvmHChdOqbEIbk12qRIGLGy+Njltfwjutjk81
hv5y033msa4Iveo1zw9HzgTKrSpiUtB1NbKsGjQOoMHlghEwEQQaWtUd3/e/5Qav
fHXaD1qiYyHfsv4ib/BeeH5UrHwp9A4UiT7vUopWxAozDG2K4VBcI7Z9PnVig+Gu
itZA9PU8aN+T5xsJZZh4QH0chbzMupJmtCnF0FTKtlRfopEEbAqT3eLSQFj4dBbH
EHftNSU2zHTfnO/sSWn1V8gix4RW8vKrlTmKFpJ3OgGD7wxvYCbNMnwbdV2X8w/5
ZshoaZfp2vXfxmNyEB+KaPqheklNxF1DZCiHIOWu4JZOxuvWg56QAqZVPLKjKm1B
IH2Z+zU/UJjFaybCE0fmNSuD9aoJSLJu5RQFDFaz42GtCo3ZNGBLSqwzIc6SuGYN
NezfXQS6N7/9WRRu+Suf+mEcNl5VzR+4u+6v0L43FyAYh9dESqn9OVhjaqTXclCG
uC8AlvDS5xgFa9zXhFcpttBrh5LUgmZ6dp3YpkKUTXDurytH3Ehr5r+YI+mcTg/x
NWrsoLCPHqpZyP+U5rgswhbCh/H900kI7mDjNnjRRNTNi4kv0cKWvQ0iHNhT/iyI
a613bQXp3emtTkoxIy+Pwd4kQdofef2ioh81s7FmyBQI0xc0PY4klEU2EWEfgyFi
d5e9qN7GiuhExIUsL5DaKeVjgHFsYXldSphE08ryt28KvhYP0AIxmoBIADpDrMRy
y4PQZKKx1vjQbsoVeff1dVCKAoynyYkqC8ZCpD9N+8rd47Ch8J43UOQ4p/DdHs35
f+WBKgzL/e1IVLIUKHhhsxbgKnzYmBSrtwN5GyiF9C88hJQKZeIyIxB2xujJZiIZ
h7lHM8vQiNSpS2CqyPZZXyk/ZE2sHNjK8s/6B6YlQCuZpTmVPWIT6rWn1M2Jcexx
3VMpRBCRYtbseCg/x5wQ5WkJiOxEM0m5DM8K0/O2Z5yYug7oFUYGolz7e1RcA882
RWc7EMf4YBgMSIJtBJf7zLxImi0QP87+EuBVO7o1LnwEJBs/tdnCUL2EjShux/rl
Xi5mXe3KX9jrYskjuN93GVzy6pmsHnWdA4wv4e1MiwNV3Y8vtjHYkyreui6HhuBS
1UVHUF+9pbUjeJg4j9OJD30wYzpyV6j3CEOcN7k5DTLy/U5wJJLAYfPg8jsoKU0Y
sf8u++82uOA3Hn3LuV6MLmR8uzoWWtI9D0shntz8nhuIl9xuBoT8IcQfYD6jk0gg
s0lBV63NX/56xltLTHe5M3Sx79wh4nnmTcW8wHMsfCU3eGxiEFGVQVlYOmqMgrsK
QVn0xBRbasdLAthHEt9YGCrpTbyeKlZURVe33jK6Gxo5GtoTKgluFmI/Vi1QWnVy
DGY/HiCv0ngJlLCt1SlYpV9vvhCHOSQHDrxek/OHTYCI3FtObNezOGi3R25oS6bQ
slxlQeKNSR6rkEtdk0uFNCSN6Xk5qVx59P7oeY1vRK/vNr8QRZHXn9m0L3QZXBvk
WranXa4a8K5eCB6KK2+K7In9Ff+99DUk4OOXbflEqUvGjXMZEvyX8YkIGUT2gJGY
5Zx2H8vjK2A3fkxCn9xI9aq7PMO10zjAZrPT9CDdFV3qiY/VFuL96AkOyrJrt/Gp
vwmWTh0qfBejmzEJBbLtv4GWSwRhPSNaKuH+RYCZ5UKRHP/jCmj1NsoYlQ+gq59f
u+9l0zf7aay0KzRJzxp4K18zOuJCNYiRV42ksWiDOSoP56GRcNysj+tUCqIJkMFG
tYiRd9pLmPXsGsRT9mo9g0XepCIIbOW9oMGi1IRducT2vr03ha5VabWQfbm7oGFZ
GmEwnbytEJwhgN5Q6jaM3GMxNFryKE9eYI2c/nUQwdNvKDwDY64xm/gHvq4GFytT
70AmByWgH/v/F57nB3od6NvxMUhsByojP4FDg5PRB2W9BVqalsGr6Xe0VRRhn3XC
ufP/sIL1APgP/yW7jn/F9jKXq6w+9Yx+hEs72kyh/5G2Oq3pgTJeEDvh0w2/cynR
UanWxgKiwZ4GSclSTV4gsE1Zeo8dJQfsReN56PJz+QTyDozAtG6mHK/+3jnVgJgA
ramg1drMaKjX5j5jKRwnoswT+A58olWLr2/7Za6+Zdrwt9rfuS6XEr/tPZINx/kF
Bfh4vMiA+JCqQdVRTnm5fs9MG4YlYGkTy79bR/wFvER3heGzvgm0MOsuBh4mVmsu
XMXbWI65r+wBuXU2dZ1Ev9fC7DVD0uxqLLPJzsznXK3ZbOzM+1Gf/4dmNNlJT6R0
XT0FmmJRGGQahmXVjvNI44ZRPvX++RyJ/VwRy9ug2NGLdxcp+GM70AFw8vVXiXSa
Vh423E86uLwyL/EaJkxfUtXxf/x43V8D8UpCA9ieJ5XcRXrqtI7RxBz+xwzE/4m2
I8Bm3hkLaICywgbTjYZzWRV8bp4kkFHXadc+u5oOEcMJvjBXPlIPthbUWSyC4tl9
2tkQU2pcoBiBq9BdALUw80B1S6/sfQj7V+U8tqRk8xVVozRbtMuPBjb6yq362TeV
2c83gXlYRb1ZU36URT7sWFe1iEqLyabdqAZ3DlDEAttFrQ5TEpi4IzPGskZoZqGg
P9ZLxtHQp2lL3YH3/c3y/yWWvawlPJUZvIe9uKg7HEcdyw921nXNm/exVH78Y52S
vu5EowZrMoTK0IGekA0TQ5OWRURGFKk1TVF1iEx2pWCR6H9zz1Gyi9NIrTbOpSC/
NxjPNlbjfqGA+Bbmq5I8T9vo2XvE/mTWaWCWapwP8ZiWM91pOUBnrrTTlyADOwTX
Icry4oXt+yzo3TVRSEH+Htvt2n5IoYxVGMtI/TNpC7Lp8ZR74cz//ixvTOBV0JcR
5pMGrwkOk2obOnO/EhxMHIa+DehSfiDtxc6/Z3qr87/W2vEup4TKng9V5JoKo6Yv
um10np104xI5mB+D+IsEynZAuXkjYWg5BtN9VRH+JpcpKr6Ufq3dlAu97IZyKmJv
h3XjMlMRJp5uc1lX8mxSDz4Nea5TjTbRDYuo3OeK5oxEHrEdfyZJF076/HUqYo/x
9ghXC/KV4lbyWBsUR87T/dnjBAFvADCTximomkIeR+I6L1/Lxj055QFNCXyFeWeU
/Tb6t3LdUrNVnhL0qqjENIYVrzEf7S72iAPqa9RoF3vWhHUWgQK3U0qRHWwR1Dgx
F+W3zpFJXCLYu0ciwBr3LsY0GrJ6VOkLUq93qBUbk+74EprcwVZABOumfKBl2Exh
Y4IJQnfrLbwJ2kHrFfKrvmkWPOKhw/y8Jfa8IZXRfZmEZ9NOhFEpmR2VaCd7d5mf
fTtlloASuS+nbwbxweike7xGD6G0piZNR+3HI4EaJvaqiA4aKChmmaaMobqAjRol
Ce3yobBT/KFjrCKuYONFe63+kkNdAELIUrLmf1uc8SY66k0yUiip7Ik33Xrlc0xn
7fVzjUVYggsXHhx6WeEUDCOYWqDpAyVDNCh0z+swQhT5pxgzqB/524EcVlVajth4
49bzPYKJjp062CF3ui/wV9hTRcK8QuYCIdph9qEJJseafuT6S3MSGd9o/yhEfZ/h
IpmnWm2vdbDiAmuv4Vur46AI6W8iEB80TprUx3J7COcUaF+R300s+0VzFGgJcOX3
0wYgg1Ce3slnZiTF0jzdPdKvwwtlnlDr7fqlG1TzTouiyToFFlTRQ6CDwGkfhE5c
J/YKM7wIeYn6bGiNvwY5T8F5hjzhxphEDKIz8sqo0dzU0HzR0l0xB5X9E20571Vx
jG66LL2Ra9licUgijQ5OfXHm1RA6Oxk95xbjkc7HTUfMpbzSNcC8jAIwPZg+J01t
FzY6Dwz60tJM5Hp+Hv1AqWnSjXf5RqlWXTIdSrKeNHlAdTOl8K05NIqKd95hCEwA
`protect END_PROTECTED