-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
--pragma protect begin_protected
--pragma protect encrypt_agent="NCPROTECT"
--pragma protect encrypt_agent_info="Encrypted using API"
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
--pragma protect key_method=RSA
--pragma protect key_block
IT2TQFjQ+iTFoTDkmFdX4V8KO4iWR1WYChyEEgVicZok00Ke52ECbjo/BAZFoFzI
oeald3SS5s+mnSoSN0HNN37ubdisLUYu3UTgkAgA7xfphyS/VSO7IhbpMudCeCYv
1PDpe1C0AB4AxAZb0+X4Vca2LSlQkWgqkh6rLYFCAtejklZhIbx/hfe9YVznSJDP
5Ef62nMNyPZSTMEXOZReE/IoXJhQzkw+Yyv0bBWWXQegEzPl/m/imtDGNgMofSi7
+aq/+kbHLSCnYBwoIFcU1rtcYitpOsn4sr/WRbz2SQzGp8vPAW6M0NtYRYUOishR
kc2LFmaYvuj/XGh47a6ibQ==
--pragma protect end_key_block
--pragma protect digest_block
HIRoA61VA+Euvfzo5GzZkTwszEI=
--pragma protect end_digest_block
--pragma protect data_block
hnQ3My45GQKhWbxCy/epUX7BdWZQiGSZbnHHRO9/V3V6qLguJzt0FbF5Idlkp250
LSM4xwksaV0FpZ7v3z4f8eP9pn6UuS0RDL1b/K3D93HPG6siUo9CJ6fsHHsuIdWX
aPpcHrf6BvDj8Ak/08phyosFWycNPUA3zjt7Cl+KWTyYMS7Qc7pUJaFQ2/XNJlLX
sAT5QVbPiQnPk89z1bdsxJPjzRVfrD5Uapp2Lb8+V9YrQMGsqxgo2aub6ad5yY0T
ugfBBXQj1abE5qCUtvXqcl/lPykdHHfkGVF5cUoC0P+t4D9NTv3Kn2bZCGSa3EEO
/SEWTD0joIDmZhF4R+fYJhwJihnjHwIFkeq3GlkgrkKKpAufmAzuLjo6qualtU1z
fNG86ARsVnnjzvyvK2PXSVDE61EIp51g6hOD1Xig3dqMTQ0bV74GjK+atJ6gNWLK
74lwtCxkkO9y8lovVOJq++/i0AkqX/LqGNRb6CJ/5OLvSHmoe/Z1h3L9Oq1Bz0jd
imj9H6+RVA5525VwKMw4y6qU+nGkkzruU3HB0NlYa5cZ5qCd5DCP1xEuerKjur22
l0yXKgnsOaoSlQQpIzAtsgGsMreNXC4H06HkRwnq4Dr61TyFoPCP17DtQEdg7nuu
2WVCGaW5JbIAfSxHnwzgEma3YXRQ+DeeY6LYKk0UHaWiBXz3E5efjJ0DJxGyOSTL
zQBk0ACmGsbfy+J60lj5oLFaeNW81eEjOhddJ4WbyyZid6eIoJAZrC4tId/+g5qR
Dy0kLndmA+4DBki3cQR9we4AEFxwPNZy/gcDcOAnQPWV5YiCyf8y28humNuymsAC
98ciJoGMAGCAEPNOSvqQkrXDtscqSIL2NrGdDlTtLxdCYfW3ZyV9Dr6/5xHwJd+m
ligWxWbERqAHP6eFoaqL/r+LbUClNfI+SUhn2eBPK/n0EPDEOTFdJB0w8gIOCxBS
mEFhkOhmOSWABNj/JktKr+/wj4Ny//ESEfdUq6W5sG+N675OvWKqgXFIBwD6pOnK
7KNGANLAyeCM782WL5FYmqJiWmh2OBgp0oInrruOyZRaFh0dJJNmExYNokH3seCX
3nxOGLv+TxwYZRAtNjZ/kSF6ADTu2pkPD5X8cO+GjoHrWoEjSnsJOSbZMZ3N2ENz
GPRADPqhTc9VK+5iX2R71tcHlozHXFqNgTfb3AGeVNKGTE8srgqyo/NW9V8fl3AT
Oq02m97XWxQ8uBUD/CDoiAvAgra6trlemBnWINhfQm3AoTttvae5Op8reK2jTD1R
YHx9f0BqgfXpLaKWIFaD/GXFVpfNFMW8HTnVy1G5ao9q0VoEvH8V/SIcbv2mdSwo
vI8bAgJynHZmEirRB5B0bkE5rcaKB9gTGSrJefB1oy/c17fI3UC2C1j5kPD2ZP7D
VC1Euu9LV5OPhDYMm0uzcYUe9X+e2dBC3+nGkG+8IeypTvyVNUyY+xJsy7sHWtWg
0RM9zHybXTwqunTkb5eHS8J1PZPj91LATXNhkO7sHxgP5ypDfr4fHtBQOc61RyEZ
eOeizVbAuM53vCtYhMcwMHTkRFXFWCAxWpOneurziV4+9IYUMU2VSZMbu01pGpoN
gJJ70Qr5GC1heFrWS5owr4BdmTe0KxQoaxxnc9eX0Q3mF6Wt2JzQHOhkRqSwYg3l
J1B8GTmYSIiTLvXf6hJqR1BF4w8T/MWIghtotZHqIGw7gc7c+5rfKVz6Y5PbXpGd
k8LHm4g9Q0YkBWcBR6mgDLQbEq3OUZuSWgKDQWP3wKhu4JuP4055UkFMYbLcKNk+
/Lx/IItgUh8cbbDnrarT3eEzLcB6SAlRQJ7TsXkU6FZ992wFbMJcCHGNZmdwj7ud
voWEblOx3lRfkVFsCdlGIwr16NKimENCGstdJARn7axkL4klflDjJq9OiEN5Ikwh
SQ181Up5d7XvOledxhycDKt1b/VRKJRBtN/o1HfyKrDU+po0gesG/XpjnOZ26eR6
cEVfDtr9qDLDVHzzmm29L5Pjxf5tKGEg0hHe3RQN1zn8Y2yzj7jEQdPk+Sxv+sZN
r0/o4m6ZtKqyOVboJ2+hnNFDa1WqmaK4ThUVA0Hh64Enk19jSGFfX1GzWV0o3hCK
O4FOQTJNHCHQ6Q7xQID1DASkIl8eAJQ0To48lyZxM4BCZHXTEvyI6MOCNHcH5fNa
CI6CwQ/Zmkpqry4GNrk9F3FVhMxE7UwkmB0wzy9T1NjGK4kJD45O9Mjifvfzpzsb
Pi1cnPY2FjM7R/ZhyLkaTzO+YSeMtwkTrGXx+0KDHgfxbzqAXOUd7Q5Bj4kgi/I2
FHsh9gmUj1z2Ff9WR98Q2rprASqRlesuSoaiWpIfyX9XqFWPqb7TLZ35XZ8fIp4K
Q+EarYxuXHdY18pq0AI1QL71dquri40zJeJce0j8BXGU0hPxLHS2ifdnPXas0KQr
Mx7Wr5xc9o58ekVO38s9CBRnDXUzPBG7HNOd074Ab6p0dKvH49AZjAEBRSdQjYbw
ZkPra6yr+FXpJdDTqQ9ezP0GKqy9degzgs/PByix0HaU41LWKkQaenXATgnfPpSn
+bWiNAGam7AjzsksLSKA30XgKGK4+H0Zvc6+YrcQgeTWFm3SOkGxvDJtX2c9JEjr
SuRR5quNo+b/YUeuVJZCosYki+kPBjbs9R4GFylel3PGTrUfyCeTdwqL1ypV5rEl
A9g0YewP6sQEfJfJj2Rj8LsAPZlQB2Rfy5+7DjQPFyBvUOQ5IgwBm34N+KJtJL9D
pbRuh6Iu7IQGmkN79JpG2+olwk06SvZ3Z+GkGcl8gHzR4VF9kFYapbKFWBWmVNHZ
Xjtb1C7VHsl5VwdW382LqVIZT2F81nch4jBh3Ca0BXO2hdIKmTszLTbpuJ3/cBdN
obNIOBeZgrJAyTzIlrDcCb1EqE3uiFmFWrQH9WUMDZXaYd7lOcVzLCZRpesEvFZ0
ZVCpVKvDYlnk5hYyUkVpgtAe2Q94VEgXHgqhlTk4i8y8Vz0il0Bo2vKDpaitU5yU
aAhdE8Nf4mYCiGN37lJ7spzi3e/5dX/ARZ2aH2S0/C/+GfBnwLb+cBFV7rjs0Ia7
MKosMCVoQ2u15x8Ri6/1UaezifCGPFnowGDGiz/vV/isscZ0s46Wsa5M6w4wuO4E
S3oFIzIUw9NcnH1HbxHh+lahfWUj8GIxMoU4JiY9RrLsAFpazig/2m6wi65LL3Nf
abhdKt3KXY3RXu1nqQ/H0hBJINDSKKgPBepCHmdEOuhXJzWPpffOGkJO9XdKMYr9
dFDRW/4VpnAZj9k8AZc9SwF0o9qoj7yGlO0DSdlivWOsoOMbsLBve774t1UMKaEg
SeLDztz/yCHYn4iKc+PXAlFi/Q4P0ifR3IRz1JeKyy5vtQd7EROo8kiJsAaTpc2q
XoOErjZMb2ph8x/vy66ujpVmtm1bo/hYsq5l61N6gJU6NyU7AlVkholgSCDy1eBw
zkO3q8iineNoQQLt8R+lHTbBSaYPt55ctCIbleWXvGvJccpqALd0EHdrFgEe+XWf
A80o1wuEH+bqgO8Ntpo1Gv7B6YvbhLXlIPMpHrz5tZKcDKU4VKXmOdwRLypLXwfi
3S9y0qrtIjyHf06U1f+tFd+BWHLDq0uyE4Bij2twlMZvOmRyZEkYrMlI7UbupbU4
+AompI/biFtHccA18X7Cut23u1rLXefGE/OZEa/Zt9QsbEN60pWPRxCk4zbIhG6B
Yq6utiY2WkWD0g3aupi1BFcvPXDdWu1oSjzMb5ivvtYWbnckLGk/o/SbOKw2TTbt
ZGBYYDYzYib602YnOqBjNxpDuZQDQb96QuIhMbzbwBwL9ExQeAqxvDTdVg1h+ZaV
ka4F6sMbKMEcJYeXrddUgXbBSpxpczqr8+i4rI/16RYbjL5rmccMj8FYRzh4qm78
/qxNn9KXlpK41BkPWeVJXhAgRelIav+DQPN4YZjRdX+JsaykL7ESKupIkhZt70jZ
JMGzcIl94GVBepGtngv1s2s0cac26rQaXfLJO82jTQXmfzj4H29Pj1e1kzGP2SCj
s25wgfucC+d/KdJtrTCODex04eO2wF5gBlH0ND0rT++pajEJzfhBneWME98siEGS
J8b5kPBVecOK40NfW6tlx1D7dj9e7ALily+U8du0wD5gkMk+yP41atj8xGMcUE9m
Kteko1c3zwJg9lz7iQ+M2whAQA4TgNY9d8B8k5hbG2QP0E4/Hxa59ZD4LFelrXoC
zFuR7muo33Qd6jdGkMEk/gt3Q13qirAyYmIa3IUPp2rGvzNSh61+witd6f24sgae
pg+BTUJfMkPUSZ8hQL0NlyDvTELl0gwG0NKUrciOssRSjaUrikMkrTnYmexevtok
YMS98W54SPV+ENLR2tYB3kiLNFoJL3dPbCB6AgKF88zzmU6AKZUWe+prleM6rVEz
ZPjyFoqgtmHLQcJUEhfcCQ0MFUVCcnA+3P4a3HCsPGNERz+4+kVMfq3De+jALhWg
O+oM4DYZ8GI9Y13ppTkNI+MsBaGOI4pQWLNvnstu/0cZF8yfGwn1Z+Cq2jxRTa1j
Bo3x8Xv6oeLG7g2TsbIgl5i9PCt2t9YA7hzZSxjEWR2RKhZTRRpU2eltsBEMNCCX
rn9dOqVet83OFtN1u6ndkaTVVVn8jWisbcrDvYFG/BBldbqitIUO7E9RM6fakjTo
vsluvor9N0J0m8HB7xRpY2gj5JxB/NhjS9WeoWkgYJKNqm36PEve/hk/knK7zn/f
XCzkVCIDcoyfLxrpHMtWjaX+VM1rS9vSSOuleJCUk3DT73H0ujeYm7tUGTW4RmMo
TK2AEtqAmxEGIUjpslShpiY9jTtei7Zjz4yg/m2Oa+eBnC91YnKn9+QwCAGtQAcg
m+ZWhQhvXDLyIfPHMNgaC8js7uqescYCnmZCL3KD/hHnPwk2l9VKLEj6SbxMXrj2
2oHrcann0PN0IFo+aTKhWyRa/fPflMTyY4pUORZlhzyO1r4LF2GTF9M1VsSAIK4Z
bEqRDR36EReCCOWnUq3T2ALAyXl400GoVg9+msBhcV2s6MbussGL67K48zVdpywj
PH4i7O1iJ+4pyuXbpCoQ1f3qeFZROjppJDS2DjFvAq9JEbMgOzOcu/xhGdyUmKpg
gTBi1emrbH1ACAZFtPTy8AQTa73WE+IeuM4Ce8R1vgklpdHYACOq7zgbtyDcDAS2
s1YG8eJXh9mVQSIoFv1sivhAqbybbsNurxNzIKpQSGtbPcn8aemZlue1orPA20YB
65hRnh+o8DbdgKJuWTeDjf69glvP9h6CeARYUk3jvWZ7h4Wqgp/P/haNTDTOMxKt
4KtNtkW7KXGb7f0yHYO38J8DrVfIFOhUDMcTRPKwsqSCTpOgjMsGr/GVtZtBcIeh
sX/thtJOd26bdzgXkOnqm1akgYjcZ2Oky/9AAoZYG7vsXaZWDoelwZwHzID0SlzP
3cikqMbmY7giHTjVeeXSW/6vqqM+IZzNQ445DZR/adlFo69QbwxT+Vh9OWfrMuIM
3h8qpbQueMVglbxAWrUKxy71lyh3dUQfH+heExba7fSyqqqQAQBAk+4ClVhwL1UX
k76+YghwU07U9Upq9/x3IxiCFdjkMVo+A+zl3MKUUKS2TledE01urP7ci9O5AsAt
AZfRv5wWtMGlZfJBm1/jkkLQe7HbAnzlnaUzBBu4LwDUNFFy6mgKzypZolHYtkJL
nwXqcPs1uqbnTZN29njtLpQRtTbZ2e3dLpA4p2ZNe9J4w0ex5lYFC7U6R8rKuvA/
AWx/vVpqoRAIMHNtVBsSUnPumYJXgO7bLH5PdvHeGiHntSHq/DOX9fzAvmz2T9rb
o2kPes/F5Sdr2czTGUShx3f7GhihxNABTxhRunG7IeypUAEE0c8s21y+DrmGZHTh
VM0N84b6lVBkioHVFZUz7ULGScss+Rp9gSNbBv3naanWhivH8bIwc0t7PaG22BAr
6Mp5oGZqHVp6JYGC/47Rrh8NJLD5p3GEG4mdaidd1HFk2S5EqZEvabQkDOnnlV/x
JBaKtilzkSBggYzYZpLG805AdexGUFkv4xd9rnh9+qfTLnLwQd510cLs5fN4fbCz
MhY7dNeu7IoR/7bi9dP1oLiyRMRqTuLUKtpGbxG4gluDaiBOOrcFYsZ0eH1TFQaa
PSx8JJr15GO6U1Ys8iKso5ceSyQvZ3kbpiRPztKKs4NNNGBu9XC3+egs3NaPCrR7
Nd28ao6M0SeBtJqniX8BzHs76IEHND8YAKfKrtsb8i9mzaRT1/1ztFNj9P6kZfEK
7bfByJCNs3DyT/GymufHDCCOUhTHbsa+ldmR0eDOWnvZ2QOJzMFWa+22TELHYhC9
d9zukf2B1Vugc52hHSGgB2l2InmL9GGF+TDPBly0W/UI1FP/7CFL02Hrku/TMUSh
dEwwQJXa2ZHHZJ6odbInulXwPomtD0ytoYrmXK04yKcwMrhUEay+3i1KnZ0QgspX
cndqU19Z7UY0sJmoyeMlqw19fflgM7N07lxUysjEIcvwXe7wXE8LXaEqg2Y43IiS
LxiHwfLiJQzpB0ZQvWSsKnClfrcAmyBwjE1mtQqufFUWlfOtCH10kW6uRYivwsk4
deEqUAYA4f9qUcTvNIrRAFKP8lLp8/IE+B3SYO8hNyRUFvCK8SuekLhkdmZDKYJU
8hoJ7SrdDKqW+I1a8qCbCy2+o3Oh/JxCEctCVCel0mbQiVXOa7RHhuhi3dpB4Tdo
LsTWu3k04q+sm86iIdN1MMPYo6Jw43xXKbWDGhVYZpdsLgW+EcAImQIpzSVxztBt
cf3kBbhNY2rfoERvzftHW5MPDhTPnl95lR1YXe5Vl3v1Af39tNmZAFE3KMasgmJ3
Wku8UiscGAuR0bxyNaF2yEWc0BVtnZPweP+DjPT5XAYGPx1a/PZwkSl2mXNL+z/q
fgWsWWHvXCpOos0Z+rNocvqwk/jOgb7c1KLjniFD1DCgV1joe4xeiiIrgAxYRHD8
kBXvQyqcuVRgYnesOKzbanKozfu3HKIQn4p37VOWfV443JCG/yQ2E5DEkOnhcadi
rLLeiVEPfxURKHIWmNpK6LuWuwkfpGPhlPdtMEDVN2GulIA+oD70074KjEHQ4Igb
JQADOYZGAns2h7AAvmtIa3X7ToVYIX4sCMYt6KwVuGwPoSps3HePGtprlMG41Y/b
/j1COh6/ahf80g3poeDa2eqY48swPSBVF46rTbdddCPsJOKQYUsGAr3+a7T/J8xc
gms6X+8LYa74X8RyjqUQufx+Tx+dLmO5EybOTkJuxwISIx0W5G5YsW2sr1zSoL+e
aPF++yfmO3K54B0g3Tl5rAuUuWSnIPPMb/p9fS/aPnn06QJ6wqlrF2zGKB+EIUQJ
D4ndboAyUvk9kKv7W4uRwiuj/mspZimhQclM0h2GkyUc37wVdLCOcAu1gdUMJHgx
onUEyxuzXy1iOvCrUJGvz39shk1/e2Y2p2d6ok5R0TxV6X3dUWPcLYzwAoXAbvwN
69adC6UFGu81JSzsdsya3s80MEcfio+RXQSM/RIzhZ2IpGHL/W9CLw1ST2y6v8go
ikkBgJ+OL/erxTl9NITizzydjZSoQ1uQFZKNx/SrL5dBK+q1G/XASB8y8/1S1QR8
i8JLZACeIX/SG95BxHtFKcY9yXp41CeDQZbPz5GXm6kYdFlIS88dpJRK7kyveAzz
T0yOJKgZKJGADmUxfjIq1EJJKw0tC0Un5Qy0qrEJwCEidL/KH6jcqVCum1w+i8/p
7lPViy0iOw6CzjQ2PdN4U1Y36+7bIjc2B2fzNe8Qikhi/lhaz0fSTG335N7YojTm
dY499Di6VT8TNKdQmwdA6RqQ1M8sTw/6gTn/EI7Lc96UMeJfdiHYHMToToxfgkCv
HYU6PUl+BOu6vCY5UsLjo57SPzY2j43ZpnLSbpL1Pj5lPYe87x7ffy25U5+QC90s
4JhiQyT+ONr3ZkV1WXubdrrqFKT3QjyddskaXmb1Mr/pkZoq2tZyrwI3k4jA2wh/
ZzCvJZcEnMMl0gdKJd2u9JioM3HW4c5jj6f6IN3eAKM+lMXtgkaQ66aViKekb6cs
xguzExU8OYMfsIo4BViHI3ug+9tWpsg4EhAN+x8dfsoL13da3W+NeQBqM9n2te8w
1r6iXwWnIMP9Si9qL5l/OKQZxHG54zzl8NgyogLsGYXHN4CkEC2UCwT0rBpBRYI/
5WGFlqCXWgnHojQk4LIQ9otip6Ln/gvrAdiyy8rlDXn6I18oZ5TFNWaDl+lxIwIN
XHSyvGVqp5d9zkT+TVkEwmzDzkFHpirJ4UlQn8Ndgfl88GW6sHltHpdad/KWNV+Q
5ylmIR+GzIikl8nyDkohUJgf6fsfVyutP4I4sjtc36RFYV4C355nm2tLYDS4fXLp
5hlM/9xQYwHyVHanA3vX6aRhEsmikFwx5czPCeDPLIJIvsYzPlh9wi0WBp//WN+E
5B6MIRsvKa4CBZl/+sZlltUalRoMQN4E75J00LEr9Ay4ps7JmfBeNQb6sucb/EXO
EIaOmpYeBHi+3Y+orMay+MmiS5hoyhB8P+0+JgFRbdTE/N7mo20JTCR7DdCL17AB
N3FLILoRbn4gWc2GbVKBdtSrHjRbx4v4+0uL9/ouEbyG/O+83dENdGFr1El+QY9B
yTeHhcn5ndYVYKK0Z0xVmmFKbMheAfZvQ6H834bIX4Qk6dwLrzxk8GJORFuweMOV
XHYvkOo5eq1v8NpgCvKKO+burS/3VPCdU8jwEXM5yWNoaoKcjr0II0RAo7bIbMOa
M5v/mveSYKzU0sfJXlKUF2x65DEUpRb2Abv0aEgS+bFaKlx7kmvw9Rt3/B2JIhT3
J3obaP/KxodUGfMshYucT1Kq74v/j3QHMzCZTrLUcNtIy8SpHzk4IVSqOK4iRKrD
C7L6t6ay4BBJmCDg7IxbS6GOeYDGtIT0U+VKyaJgHhxabeVGBXsvH9lbb6dta0Nq
GkhrKGkueXINMQseXEtZ7O/DZ9bOOceQqIwHGcfSLIWK1cYiWd7MtSbLfT7GZIUu
ZM5D1WgZK9j3HhoHP7lSbGUt4L1hr2VJlJKujmfJ4PevFSuXEhhzV7ZyF4h+P8Xc
tcFEsr20bIBDNTWtFIZ6Ww/iZANHt+VATqu6JW2dxW2ZCfVnL0R09Jd1BHxUpS82
FCdHzdhlnEtCjI4MEeyFd/AqxerMnkHTwKO8TbHz6ZtqqbbaHcWzXgfUXc/bfNSt
duUBRr8rzKNIY/27FFsbmtRuhjbQlXAsuOuUGTSbfzuC+bmKbw4YS7s249H5h+xi
HgAylfTT8NwosbiCjRwKAo+2nIk9kzmq69Unxa/2MFG1MN2VxAqhrMmOx8IyVgny
UQBXKMnKUne4zNxMyXLIGpOlIh3Y0fahnhnLHjA4aZ6Oeo1erA5utw6LdQHHTwyJ
RJQ+7nTb2iAAY1ffGP9r9UIW15xIFnObLU4E6NdGl/fxZBrbVxB7JH7+nhnMtE0o
W5Wwet998Lle/j3T1yd90nx2XRwa5YWiBu58xFW7jXbYCHOS4Wm02bVdPYUmQ4yd
jophX3aMGRA5EpyaQ8CfGdPjtI1bYErNCs+20qw4bJHHMeK8tv582Mv/WW9FtM4U
ELTZnSFEiHnspE/tdLUTZ+BbQnlPdNJbf88heJzdoZnJ1cL1k4X/Ha2vpefosgVJ
erUKDPkWIpDyZEgJgEbGCHwS3UHuLx0p0WFRDnphzqftkHqtk8tB+pJys2fky5tR
Xr/8iF0wMMNhrUqX6izJgfKLrwv5Gz6ez+OdZjD6E8FXRl44FfuRbwOfA7mT5r4Q
F5w3jyjRHmLLFaClSC25c/OAP0L3EVK9OfbWi8cwcYwyMOG3O7ySBSP253ayReQ4
20g/UlvSoeLvJ4haaOfvDfhpAcCb19xfy2l4F8zxsu+MZZv6JWJ7Qw7Nwu8CwCY+
BJ6PCAlEGQMEO30nIGxLVhHSzpdta21AEqIdeuubdPjSIbT7Y6Sd+sdeWB3Yqr/q
aqYSij6I5bjJi3CiCuq953ewR1rvsZa4IRKXHsL+UdHO+o/XpRisA3SWtWDnnQr+
wCHnoBmTDzzSm+BX2hG9pf6ydz/g/BGF2tMyFoz1CBTSCOgG3ZHxWj/S1GkdAa+B
JpRW4eBu9TwSb2Pr6aKYl4qINmzh5/UdZh+eNyzNkvljZ8WtLwGZKPWMARWbDzMe
TN1J74FO7reVzWFKX88anNhYIJMZ6phWIOqXpdZPpb/ie5f8+clrf2ipeo38Qium
+KvHo1Pfobg9JvOgnkDfOLbkbClYGToH16M3x+OHBoushum7xdKQ+jF8Zpxd+THz
OiRwA1FqW550VfC4cgFDMOwRsX7RWAQ1A64QTiVMhpOdkVsX2c2wwtsS8Jlae3tk
m5c7E4Q6quxtSnvqPF0FG6CxWOa+h21linWzWG66d45vOdWzoa2MUJ2dhDU1vfDl
tESD3A+zdxBHIFdleojdgAkGJIg/vEF0+5SjrywOvUXrvyowmU7O8retj07A33ZP
oQQtFbnn5WrrSjXiN3XpGxzyWyYYNr0ArOaIFXytN3BV3l28xX1dO3jFBh4K6Qq8
ckHBnh4ejlmYCSl4kiKV6ciPyPzgRldjHo7XIe0Qu3rTHDcdupIM6ldIUDIF+AWe
+2HgU+lyx9Q2v4RNgkrerMQqKwnryVR4NSZ1x3wHqkCwpY3LQjIU3zVnsBWhlG/3
Q4ZpsxB0vTQYzrRQKBGhO8PdYbohCt8cghPCvDrBcqW4S9glCwUNNwlPeKShq46O
ebbNYO4G8kkEmD7saA2i+Dw81KLgyKlFuYB7T3GOah8LoFyxrF4oMsaTouuTDC9j
ilBzHauq63GNouU4L3P4H9vce3g6FOkBE7gGQDj6Fqc15R67ypJyEItXKhYYk5ul
syDTpL0cacn61x1uTOUDEEqQ8N8tGqg5FpgmSskfnO+dLfhtIt+7YKcZec0cvyOo
gSUJDm+ifFUbaEfKDLGH660EMaGoMm2uvFe6NizkgRaLPVL8kNJnXKgrN5UP+YBS
3jRvGvRc9Nr1mnyd/4GQYcH8UpB279jq4ZC5zCto3/Wxu9Nql2H5QSD7MRr8Jirb
DdE8TgCwIuGcBg4iAntlltFy9nqL65CzVUf8cGOHieSx6A0k7PKTXGGC8FdrfBEO
GQg6GQFClzs//Q71fuCixB7XvKiWk1w+zUzca7Qnr+ZGZlrzLFOz1rxZLjpaxg8d
la7+ZMWC7/3I6PSMd8NFd4k1mBEkBJste3PyiRlCRismOcTl12z/rbY87LsWuVbo
oUpAOQMq8IYfU4nuJJ6Gn0ID/vHe9j+08HxfgVAn0aN7TS/U76PbU/Fbh93ZH+ex
fwhgNoX5rRJcIzc+BIL7dTgdbvXpR3NY4Jk6SimY0t7N+CQqW5C1VEeOcSxopKLX
lKPVla/7zpYEC4Xba4+Ygqa61ijwm4d/Vi5PBjGkWzgVHvuj1JIr/yQnHUmp+U0b
stWGsKMOWXAz2xq+VFGc8RQLwRwlaw8d3GqzX7L03H+0pBML0I24deq1aPZtwYvH
IC+QDeQwApJmgQyBPRhecIYaMhXx+m1ETtjif2LF0Q3amUJO7l02dljhqpvkemg6
O/gRvFU8ioLPc2Hns+6KyZyvrroFE3e/v9rMoZXDFhHzZluAP1mjo4Zz6ct9oHOi
2iRBab5noQyZEuDs7GuPIVFyy4BeMc9Qy8jW0/EeBz3jqXF18WEKzjdSQrvoBG1/
LJ1KxJ8cmJhQkYmAeZ/T0AKh6/W54WXG1WDrpVqd0ZA7lKNQl0jJ6GXVdI47w07m
GcL+3cA+eG6HdB5atcTGvUoePIF+OURKQfk7bnPv3IHSIPxOmMwfRGQavMIk9nDz
xuTWdx7L2a0yn2DdC4jK06khW4WtAnoI1ChNNU58lBhQROCHGClxcRqcyNRawkzq
oE8t9IeqEquzOautvQYXUay/iAz4lqAg1jlRXXEDqxleuA9+DKLQvCxDQLEqxWxr
n12V2B46XWCvf+gkWQKRepROzvssz8Sbq8FLVeyC/JN3M7euE5N4lb7Sej7ZFRAu
tIh8elECsgG38daFjequpWQl3f2z9giWYlrH6LP5PAjTgfk8z8GB4+EJON/jzIAC
NfsfUHS+mMKztoMYnzlH7RaP5U2RUPALSF9n0NQ5EuVoqwtrkZXQF27G+VewzZN+
/C17bIM+s9wrI+bZDHtTuXw1gnHUnn76CYOq2EUqOvEPzAoy4hebyC+sL4/AQBkE
y78G0QGPcfnYVmANJWgVCk3skt13TxZA96xfIK0ky8x4eu3w6oPyVfwGnnyUWTJh
mqSLh5+17SAmd3PnEJ1i4kuRzTCBK7DJOAvD2yKxgL8GilDwxIfsmM4Oa4herhCe
c1Ov6rVKuOPCY2e8txMS08TQF222lgTWJ/0Jlv7uNb/F5hhognms3qtydIO4/zVS
1DI6xwwro1CmUvpp1fEgrp+H58hAV4/b8e5sv0DO5Enluc4kTlTreTYBMUAb2MzX
CjfWx9W8Zt/QtR3kpgBPJfkA9kdtn2MKTkVvjXuDHiZOHCphZxLeR5A/NdoI1VPl
0XIvohV5D1S5s6TEdpdu9XRg5yrgP5c7o3eC1bZ7p8NK3aMOclhnbc8pDtte9nR0
wHudEGa2DZeoItlfthhfywDIML1+PU7NGKVF7jVdgwMHWxXsRR6UwDfhz/wvmaRh
oP7aSwFwpTAqW7CQc1BVbqU4ZnO9VTKuATagm6orLphFicIPXSK7SkGSsuoIjJOD
xs3EOlVDmm2gnEnCeO0pnWyBsT01kkE2AtemRZCHWTNVkLc8bh/vdG+tqvFhQqpj
OhF2tGkFHl4ZZQLuhLzln/kkjJroh5RohTsDDIbKSUAmj7je905cZcDD9LgaYvmL
b+pX2ZEwdZw8cE21+fL/vBbdTk9Ta10Lr3xAF2mTiMQJil6UdOzXSfDV9i2p9r/8
H9WibRKNOSMZsW3EqwPbphQRDYfe3UA9sVtfkFghGCNke3motkWpsGdPDs3xYaeY
gdAC6Rl3rhzwHLVb+++oDX1UMhaGz4KSL1iPP67WzXci4N7ENNoIKoakjqcNQpz7
6xA2zVq+vwJhjiBR3vc4mlKHgkI/eU9C5QXS5YFi18pXiJNHOc7eVTGHSg85SLQw
UDCOjHLzIoZ5YIAnb3vYwMDkBH8y2chwv0KhAzQfImpB6ALnsfWx/pWAZm9gKwqv
zFf5uryjWEpDYaoyFMZ+I55wu9q9BkVZ1idvvzi9GojuYGt8vPG2z/Uf6keBh7iS
KCSUG5xJ87Ol7wNFGt/I5EapTURaUM4gWgW5cgtDC6djTCx0LF8gETQwXFL7Zw1E
F+mzp0W+3n8CYpZqm2AWAlrFWpOOXJisXgijpZHbw5LTdkjsfx1TQveBoKmpt9pX
zNmwEO4kAl4pYrx1V/9qngHSne3joAJWnx4hnC+fmUiJ1+zhfJ+bPc0yBxug0JbP
Zc+6r5oSEe9JIdyvWZTpnegYBuqoQUCIFk9OyYR0e+YzdTsNV3Z29vc9R86vKiQw
9cJTj8CGeeO9wC6tUuwkNzHskeqA+uPRFVmNx+2ISThAZuDUTv+333fI3C6TFWoF
NVNQEnfLD5j54T5gEs+GVKVi7YOr+yxL0lSBuVHyJRtYxP/ew+E6qRY6UfQFGoVl
UEyy0p1OkOKBCe7egUVYpZZjyKkklRLWWg69yP539dRAfaWwia5L1oLQA7s/FKlO
nEKFWv4eHbuqRnZlVu1gJ2L5qt3B7iQ0SHEpI20jakLapyYu7lSyAprpQmRuj63q
d1CvJgsBzV+YFoy4KbxjK/rLODEFJp3SpPSuENfGSqD7PA0piElPztxUM50GpTUp
+hLBTCwThULD2aBeuEzaQ6KX6VqBh/hXTE/23mrBiSS+EyrG0vpU1EH44O8JREjS
TqhaAraWVCVeeik+LFPbAcxH15NzCj0+rI2uHV0FgB88qoJ34bLV0Fj75RYQZBiq
bcFUk1e7OcUVTe2UV69drWUILv4YDi4ZtWj8AWa1dU2mxiQ1kYmq5kX5NqTbkDcW
bT7yXlnucRJKluNbCYT/w2ds3c0Pntb6kGh4xf9zsLzyde0aM+Q0xOyhRZbN+C5x
lSir7P1TBhf7m2bTKRzxd8sWUfNnQZIbtmw9wUFHd6QaX/f9beMYZR0NP9TnyJXK
SgX5QBLsQzLXg2kFenzSxjgqGlY6k/Ro9zfot0QndQn5ctyLajgLIKSoePBuyKWl
Lb5Y4rIRDySuTpy773d41vd6buyR/L5gDFA8pPjl4zs8Gwvf5MSMcttWrpFzuNpH
wW+jjq7WEnsEE72IfEKLVgCqpeLKhvv0gksUfeG71ornTOboGJlj0j7htwLvQqPS
29CyHJa4HSmLOKnURpM/BphYgWvC7mvC8i1Ftx3xUyR607PETuSPMj/3We7Fjjm1
ZTzvyKTPMRmdelpS7XOj3VVIpEo7NazXSQzols9EFKwpoH8j4hNsovBxDiSD40Wo
nhZJiXAEH895ScqnVitJ9nDf9uGxMOQIQaWrjtK7wbFAmTGpEU1VD4HQRuiyaTpH
99NrxK619Pm8c6zcmt3fSLYag1LYa5sBBIWL585T6CnhxBtZvqAVNyIs4mskbEiC
XA02aZfeY259BAzL/EC27lIiWRPbhvlp6ZikBqoWnCtwDoK1GbJPXQIUZrDwP1gu
YkCd7UiIxMX+JcssjedTINkCVOaKZeAdpvC+d4VpUU7ellIASWC/sChx379/Ugvh
tCPxAtquGsQzAW2c+uxOMI3QMJ8Q7Dvfmm7Ovu0XkUJdZB8r1Jp4fP9BWg3AzRJQ
+F+EYBzl5Pj3paeB6XdtJ/xg0bTOEl6fJD1KbLVcaU3fANIGFb0apQ8yrKIP+M2U
Ng4TlGylnqylrLGb4S6oWK/bMQISxWhZoXD4TgBG4XG3t3szp7kdbB0olbW65kq8
7MVwzsZD6xBb3SKUlvCC5N1hwNZ5wNPVqIf0XAeAdYpmvyf1f1OAHiGjWJcm85q6
or1x2O7OT7c4n7Usx1Mm+LLqzPIC0u/KJdtM6rmT/xPfVCZ2xZfG622rXljA3E/6
X3Vy0M9n2IO11N1wfwtcyPD833P2aeJy58V2HbDlYDXwNdeNjche05l4/ZVDNzW6
6Pn8zS9R7pjIKTnh0p7VkS2JGZ9R/emd3WDM/G2ZO/D2adixiK4+2BQcrv+WJmMi
VUV8POIcQGOAsDNSDin1SXAdHA+nq+MVXaqBy+RSa9P7RK6mGTbqwOGSEWi7Zw17
UEOj/29IlnQvrhklwZ5BkyVDsG3GzWkVQS39lp7pzmMw3iSB1Z8yeD1ZTxPV9Kcs
E3+y4tdm6nt+OSspCQugONuBOE0+SyKwfIyiOjwZ/Ivtixwpi9gsd4lBs5rGcXo9
LoXZQdZtEF2vSuiEnh3HteZNKe3eWanMoEOYPXaZKVj820Hfui7MN1YlruxHAN6N
xJNfA/5edC169s5er0uWYdjAiygXvDjBvsNsx7E07h5YJzSSdS5lPa2Pbif6s5Ft
31tVfc4vnZkNO46v4xcFYXcl/IbV4DM1dZtQjCBXRMnu7wzwq/P7xaHYlYQ2PlGa
egogva2sZydzr46HkEgJ6C+wNpsgGDadN3WrWlHc1UaBBUHHOZxkFgQXr8TgXKSr
h+FviBUADi47tWyT3uvDCiEQ1u+vZ7qkoKXvWdEnBt2sC8emKN8qLnw/nCQPZU6c
lSghDDvDNoCqbgtaYEolodtybhftbFdzA/L1LtnP9/iTZfLeBfnXMGdKBfQJ8VYL
CS6LEFmoWFQ/NLHEqOsZNn2Wrp7XI107wzzKSRw8S99+hqyi6b+t4z1V1giAP+3O
2QEWTAo8Mt/1f7yo6Q7/19BBOPz+PdsbP5yWtZe5WChlE7WXBSPqyqoKB1K/WshE
XaSExa1QCEB/QLcddg5ucJTNjyvOjz73dKVVimx+BhXGwyL5P7NAXflbUn5Dv9wn
VHAMRlN4cV7vSm6S+mDBVgSiCfLvCDSqE44K6+3kUauLlCWkgxKdL5+h02xHPxP7
kdkIuiyFDinHd39BfvyNBFT8DjIV1zn7S+1RWkspKU12hvGf6EtQ/tuwHdteFWT7
lyrZUuoapwRvaAd3PXTqhGjD3ohuIb2kY9URSBZTF5bcMXq6KMkICXg0L4cMl+oT
cbLyKeN4B0Oef3lG5NA5jdbSjS1STgeOD9S+m4nMxTsRoDU3DaFDd6QBZKsbexYr
7Lnyt01dM9FMD1lv0Znbm7ToMz7o6+57qXT6UkxUAeIjqVwPGAwteOS19wCI2ptJ
zP9P/JNjo5tVX9UmSOnXvjahG9eVjsoeSTrCYpDuC3iGU6squPBiizhj+leaXhqM
83kbUAC/lbmTgfSp7T8I9ZIteEiPxHOKONUYcL1OgN2N7xH0l15exo2SHh9+eTDb
Fs6LmwqBEriLlybo0kjSHXm9kKlrr8muBKEk0h7PviAlZgCy0VPnj8f0P6dBkhlj
2xKzKEAUO2/ZfyD3MYxDfk45HKzNLJkIVnc07hy9P8eN5S3eyBa+ctm0eJwshQef
0RsldM4z28aPibmliDFeN52v3BpS5RPjAuSfjsCG15TFUCbDDKXdjUMk6iBU3LOV
qYwrCDr+d5yAEVIlTUybm2r6tDLLb+bkLZHJRUCJCUIszelfBmkPdaU6NNK3A7uI
vapaTiHyTj7uESLPNjzpkPo5DRGlqz8y6d28qoyp/NUvu2Cg+zp0bkFNOalPk56P
Y/SQ23pU4XWDDF0CkJ8xmUcxqXkuR7sN2vZ2HXnCA4U3n52D/iyb6gfYTDOM9sDC
OJgRqPqDkZbAGh/cErXyXM8mmisirUhvUj+HIW5Jdk1815h9JnM58PZM/le0r0Pn
G651vWQQ5/bqFBTLwpEf6Qs6PjkvyhjO/uIkc62UTZVzqIXP5gMVC/5PeyEK03hD
hxV81EdSOHi2JCcth9rYrULeo5viHClEg1/u2QWkpexBGKd0j36X8MAkHUQXgzGB
9hD5m+job5YpGRV6Bvxh7Kt0944WZTB6fdXpLtsgeuE9c64p2XldbvyU8Mz4CBCh
0m8UE1+kSpP/EEr/XwWYUpSXlkVg2SR5E+0K51T5tjX1SA1NQWPPmJx/+8IsDOyR
3Uaen3G79ClOXaVjT9ExLrEMrPW2YfCUSHNxB40seLSlejMuuMGZ1tGj8E9pnysM
bWkiKcQopmq4iLtQZDQlZZ9ykDqvldKw+JPPqvRIqWGomm+cn+NTnCoSfVreMWcL
vA2VeeHygythI6YpbpGBUUIb0+Zt0QpuuiELc9zHkpoJ98ZCto0mGRk1CJIrB5Nz
I6QMSelvBkMtn0noGYpvM/Usd0H1VFfAarjtkppT8oLcSipAGyJARdKt+KZBxDuA
Zsw8jNtlvp0Kp//vd21wP02bdkV1k0fqOk1gZVXPxdPFsu41Axms/pPpd3Pv4aRV
L2yAeXVUObet/jmHtoD1jb56utAK01e2H3Mb75fbh7g4XlQCYyQKtGnsBUI46VON
e2fb08FFtXiWVPBYIH5nTH7Wv4FNelPkapAdVQhKjUb2RAamyjJRi74+87tb/Cyf
vcvcnvOTx2pqgaQZ07TTB+GeLjx+raKSbIxPvUR2rR3w2B/fW9E6Yllk6dZT1bwg
LQtKNoFyriMN4sW5GKKnBEhmvzE4BUd5HCrvMC2BzP1iry2PRYtiPRQ/TACMzQbi
cxF7fqam9aqm4iM0iCtFqVTzN+4xxpi7G0sBwTl4jJlw4n2IEHhXu4RoEyflPEhO
0JLeP58Lmop0MK2T3plCIJoIxBhWYtoZ1I8/xWpbzGkVenjaLCSm0hW2/x1VAKlh
HBvqRHXd2spyt+cN2KlZpda/w/x43Xc5ZgPOIh20fiFKsuqOMbeYVRVrfcRiHlBS
ZFRW2D3wf+yC+DBeEQ6JAzXlTCkSaV2Jbb6vWAgBiXRreKL/MRkmCQlVdxj1ax7+
7N8kucQ8OzncwWGwZN9TFB+4yvI9lsfrdXVldzatXVHpvclcnHJZVD+cow+vsw4B
SYKUMG/d205aLj8Q6KpnpAHo5nVfvOCll0qRaX3tlEOcNaw5iUYyERUW5IhOQ2S1
w8YLqr7k1I7BrbChd+VyZnxecZgU84o0hXE+35qIJqZPE92yyq3c/T8Ws7pUHjjG
UKW/5FexbU/ODC6Mf/W+yQSpMvJg/5YNGyHsogOtF0/HAWIGtXsNYx+fc8yXgSMa
Xlu/cTYBHAvmNEc77QUHR0qdACEWVA6DrQZvCVkvXlJTJawGnQ5JOfhDMf3yP+Qu
4+kvJxu9ZEQknAPJsi8NpHcClGOijyQAdDes9gXxBycJbg2zESFTW5x09WZNWQLJ
N2PHn3zB6jwnGtRwluTRo/wQ9M+9iLrMRWrOq90TS2UKvje8sr11Iwfip6sXiuH8
lUJTHPUHDUXvLlt8dMFaMCbvccdI7ffuXLP+JHHRdiakwQ+QMb50m0n15aIjoxWB
7hELC0eiUSxvio76ccheWXaKwlkylBGvghyLmRv3iaHXDP/qTz0SLubVRbsAHqKc
Vzg5g9HyckymD4EUd2iAWqiEZwJdwxqw85QnSGQyii5jGACsLWl8rlf3+h9JAl/h
6gxF89cQ3aEImtPDdT1JN8Pyha0pcoeebEQ7VLQqZfcv/UGTgSGhoXF2tVSBT1tj
XGs1/85QlfaE+AA/i6vbLErJVL17suGBKMH9P0l3zAnLw5oSTDD/BoAXOtZh3ElT
iDYJqo6HNlNqL5jQseT2QtFaOtZIwHFc/QSe9sW6jU3sJVvyGPAwV8nJkB4ADrIc
mqLJ66pl7IokIPvNemEUhZJBduKsBqpN/Sg90CxDxpDpc06DLkUk4k0VnNSVnjgw
41bTtY1qGZh7wSGCNmuVDv89VlF+XhIxpCZdabeT3bpcG3/QEO4AEjSbS+N2yv10
xrefDq1hXNwuTxueiMzqBXskIExTCV0gW8EMKhWQZU+0aMIUjVOYsRyuvZdRWaEc
Xk4A3zJ5/rzS2nBxP4zvCsUjBU+85VBQTHdgMctUiPPEAm7IXfazkXwJTtaO721o
gc4uAMMQRf5BfsshQM23+a0Meq3RU84FV9qVLQ0FDrDmRZ3/y9ADtbI7zZDIO+HA
yX5me3+pN9Bj4GXKFkGjnaylMQyu+v6/9J5/NLJZ/HuHBt6lx/WAMYOGcwIYMmfC
khKP5L1S9bucIu29Ipgnq+CYNFixb7RNL6XL1BJkPEhKmRvqy/JkohA44OzX231K
XmlVqShZr6YxsFog6MZjsj45PBdg7mexCBCKXzUFnh7KhIRLwK938GCiV4dXeyr7
oRAxhpglrcjqsqjd3f2KDaSJqdyImU1q5fE4SlmsZVGFdM0GybRGPOFzyZB2r+YT
xSQey8FG432AgxY2I551rVXnGu8k0Iz2/tAVe89x/HtfGBXlFXNvIe+y5Nd7gPRt
xcb9gmzX9KCiFw3sCFOD+tAkvJyCLnHCiYnQhaVfi4dX7N3MOEprrwfwpZpie16n
6trcP3QP40R5Erff72LDXlPWKw3C2yhf95umeB9Xd0IPMMV/I2TOiPxu2ItI1Tct
kN5/YaWPLftEnpbEtnAVAgZhJKl7ugYbsJXM8gS3gWVapI0EjQ+xBpw/+25Q9LFa
wH8bM+dY5hxiaqSJKAPxMZ1b5qBVe7pd9Xj79iLJ7pVe6oP3ll6iP6vfQF4V8wiP
ZdnPHyimjjttdQCW2Xcjgs8JmWhTLDr1tx4ePsRc4+443C6rcy81B61+vKhUdzhQ
redWGxswLcPRZeFdT7oqoAmjvkVglWAe//r4/ZldcnMMy9Dvvp2w+kvTP0MEyD3m
RxE40kstG9kKH/8oVklzr2e6RRcF9JtKSEKqIDuHtynYwp9FF1iu63GIMkmmuaXu
zrOb5NdUCxzGRQlMoNUK0uSsrOcu31UQebSXz7txjRIhkmBmgPAYoznGyWMVi7PL
t2tr774fgr0r0AFwqFOmE0f2q32gNK4uZUh9hpCuSHLsziIgmABJEy+vvu1SWMPv
M6ZpqdguW1R8sB+E8YASGqkZaOq69ZgB3tP6rjtUy2mh3JwXfYkk7AbAbj2zaAtk
4OxyCkuiVL9z5AUj47Sv3CHYcXG6C+KOtMn3R6Cmb6MlaXxNGl8T4Alv1P+Gz1bs
HO31EVhj1TeOKaJJQVnnXYQjTjD9VJYs4HlRzB9cdVWGi/rdi/aJRp79INrAE003
cZ6eWFhEMMAAA0e927uZdC07J+/GoZwquZrn5kPcTrSgbVPdAqSDKpKSFUTc0sy0
3Fe8Fv1FCp0Se+aIwkwn31lg2bNF357wfqOQ7dZWLQhjG2EgQlYM1dMgckZZx+6t
oIw01FMYV5xxJHi0iu4xfafW5hNpugVgqo+v8AGZghfxxZS7+ENPYXALfD54kO6j
X/Dguge/AkOhhjEuP32A5uRfcrIGXVUTYft31r8UzNYYyBfDVPPLzi7xuiBmz25g
pfr7UFdUc4tNOXkua45sIQM6MkELue6B1QHRURtyIoJNvmD9RkuXLLOQrRKXVo8O
iH2Vwc2eqn0ed8STem6yXDtfqTrFMtaBafSBV8oUPguPqeFOlLI3oETGeAjbeQvm
x8GD+X0rBlplh6/MIuuzvvlOmr+f2HvZ5hhhbydxwzfpitTgme2crFr4hHO85/yf
FBxLWn3vH4BOwgtFDBOSzUv6w/VcbYUNC1FzXA1hCL/zpdsxA7ZvAxsA7X3IO2Kh
wPZKMtrr4ntn5pxZl9/+vA8GqAf5RMRrcuUofbCIm1cd+i6rHkiEJlpIYET5zBbL
MplZxgH9+SPYjJXa8x21Y/YkoSszgJKlASENXHf6y8j6ru0aQi7LU8xP9q6xhE1A
YZfeTGjqPCcaGvMwqNhrBwhiud6S1i9PZkMETgoIG2oaKdnLsUTn87BZBFVd9dz9
n+daign4JvG/Ld3FLYbuibn68jglcdYFh9NZMMpJjPY6DsChW1WMfPYmiw1DDpVt
AGgKJWWzN7MODNlyQusu9fUHDjRX6ULlI28Gkw++fgqZ3mGbuLaGeJXwu+DE5hcC
YyQmVeocs8UAha+0MnYWu7Uxw8kioX5csmESSjOPcpnq3/eGI3BKOxTFFaliVyfg
0n55hW5YZpOQTWq7q/EHoTfWmrg6ORqffAR2ap8EAAJPJwVmt0diezu64fKgAJvY
zlrg7Y7dPrnbv70/+oxE1OEZO4XFQw7ecyTQ6pDwOxHqwTp6PIstYGtMviw4ZG8w
0zU8bbzzhTb3SG+J2bRBXbJiuMjDnaJWDbRY2fvElwpeYUvYcZIWtFluW5PH/IGA
NYGIVwSaFpyuvlvT/xBZzvESMxFmM9da3fkF9ecetqlxNCDPt7TJBgoiRfz8qmfh
O4T9wOlu7KtWX58n/5TKz/dA8Hyikwj5d/P0t8KL62MNBoZBR48Bv3P8rCcxbdjo
sO58lnx/TKrHDfFCMg873COvTccqz6zKtyutEKZ9QnjNJdrVq9dXeSaDcXlJvg/e
qe9sK7/UVcIcDbeG/lwwZoBuJXjRFEYuQACmpTKiREAtF/l3GPRVZL8GYjfeegfW
eclljo74vVjnZx/NphWAGuIP7LO068ZaK3O61bxhVE/bFT8A3OZkBjlRLHbIMXfl
eu/cqDBkL71KG5alL3qV1Jh0l33lki/vdPfAE42KjSi6/AQOJfp2upeSiPlmDX2A
iqtZJXSax/c4t5nd6LjAspyevjSGj6cFnZu8GGriZaQOWHO5DmpkwCVYDgqxfSvL
5HuIixzW+9QEYTP5k/6Zcw9qShFA9uzpmS/6vGcpMgGyvr6T9V6DNF0+nI4UKLCU
NtasBNkqtNiBsbGZVoXItymyRI+EQsE0u1VCn4NamMyIuPegbHKj+ecitILX1djg
tUJMxo3I5fNOLXJUI+q1cho9TB0X3YYHEh2N/rq/WGd90EvYoNVLiybI1LTJbZ5d
kGbZuc84SY2uQQFZ+Gb/Ne9qH2/GPeejF5vbyaK94wIwIomSfGt4yzUJHniLjm53
uXaCx+pbzLwaRpeRedJ6vcb8SLFPz6kY5lTiKP1EnUngWu7b5JhqWUpZr4nnboPX
n9dbV6asjlg2JubW6u5pYi0fXSkrN3KIrDoxjf8ZSr/wnwjXw6n4vRP5mZtmB0if
HftKCgHpj/qd9fk4TEQPEOhW8YyScrtSbLytzGW45p9kOHlmQk2IlJAMwR1pX2TL
bv/WNkxPc5ethzoAoVDy6sIMAWPKlBxnWKuAn5cCmNYigaRX1GMge7mCQkpwr9B7
/hDSjNc1mTpGqVk9ffhC7BNN6JwkM0p87qFyrZuIRBUu3JgVFTLz6webx2oA5+Og
WbHs2t6zsK4HUuX81bs9zfFsB5AEwQ44/AvFZaiOBX8QqEljOr5TEwIgifvVqkUP
Dd7eKC4lc1g73+BYA2t82cdURibStiSXim3VBC9/q69g0yWLgTkMI5ZgD+ZAX29C
XBvHp+Wfu8BmQeL/Gs0L1xfLg13FJ9qyEcaq/6uscyEsZFnLYhC99YWvL6jgO0yc
GAhfGmTjE5AMRF8CZyoYpTnt5iJfh9Olk8FZ7izTt5aDHehKO84e+86rmzuMCC16
QDtWUwVilnbRkpfjpdC3NWyuGw/kaMWWnkyiYZvucfqrgWp2k7+7RcbzR1SPzBEo
MQ4Mg2n3Q9Z98v8dGKC5kcBATsmS5K+wT++cQ90LxD8Xq6mz2z9v/XQkjRf7/3xc
ODohdDmM8Gcun5ftV6Mv9RXfN6PgmFhgqNTpf4yTrhHax9vGMDe3W4MFeq+xK2K8
OUK2tGI5ngFKZ/DbORvPeYUP3KZmh2azA8q4VByNhY7HzH/ZacJshxX2KbYravfB
SmLnZLmYi1D7AbQvZH7efl/wGgclqjOKTxvsi5wMWOYjvaYVODjs/7tjQ3+Wl7CZ
gmD86xUcDQMBYlB4W6ncEoEwOSlNreLm98Ewbn/XdVIQmqgkEHNVp++3qBdl7aie
OyAfRKbkG6CP+S2LgSP4MAQJOnSVizgS5UEAt3KlJyrNAqqzUPaaIJ135rzJxtry
AFYe36fJ9lOLzyPlx0q4NLWGvCx7GpS0i9eJQMHPI/bZCB24WP0FrFmPP+LPIx2j
x7Djd0E2UoUqXm3oEk5kxenkAjNArwxxDKy4xhhOPgJwtnJkXgggOvP4SuNKB2j+
fkm7nI9y9X1T42KPaWw6pKL6lUdQwpZQ0PRUiP9zukpLUeLAhQnDES9qQaetViDh
b5/9rjAbxbZya07p1QCNOxMKdaliYHevx8qfYCZkZq+0YnQqN2rS1uX7lWCOoxy1
/l+rVL4+DqMMXYp5/Uf2d7m4WENvxQjakvsNmzuAICJRx6L3oHXdcJqkz3x8+pjF
+EdBLALmCoNRNH7tESFl31l7dH1l+1VLLe5gisqyWFkIn14cU0Sq/dDJVN9XuYrg
CztAjeqY0aOQS/nic6ypylO1GgeolqVjUcAv/OI8OML2m7UqEj5vpgopIdgNNK0U
u/h2QMJE2ysNt/ZVMtdJiW74BGJaLeYJ844vfdfH56fpxNhnmFbGhKRmzGWCWwyq
PXmrwULOBKC3epJWldgmdtT/3NEYJqeXuz1qcrVyaioqZW3h6CX4tD8xE7YSAbUO
thia4rmWsPqv/oERRecTk4VlmlAK0pcl02JAr/dTJWyMWH5dHC2di+A6K2v8mtqC
ps0A/L1lVwYyrc7wegCNPt4ZbimHZ1xgtBfFyX6ULHEPbdIxkcMQFRlwD0FEQQio
PDNJeQQw8obB696mlJB4IzpuPdjCgwt8fUBwqZ2qbHa85BZL3EHuQvlFPvoU3Srb
1AwfFg0iFc9YsJg9fyCdSWDxjhMKcD9I7gXsm6t7ed2pJeG783JtqsVs6Cr+cKpF
/Mb+xeabKsx9tENfhDNvd+grlCMmbIK99HJ0eKotLd6XSSY24R63A0077rMya9SI
L/ieJAIR4PTE7Ie8pBLtBRNoe+5I9oqCqURzW1bH6VZKOokcgnJYZ7NLraDkK9yP
vOOK7ntNvbtQM/PFpQl4rmpnzbidLa2k0kQL2vgoMoCjq3XZVAfaBBAVFUMsvSk1
qluCvrnQrVhwZ7GCSX4gU3bCQ+r2B2sKi77EQX2zPLlDL9JgGtOKbVQQLv+tVAzf
ma7nBDmoC0EeU6bdq7mZ3t2U4IUMK0Osxvs9j1hmWC4giBuyImsQHl+nemcuzxWx
Tsae/U5znIAs2NRzn0x9yNGEE96nqe13PNq7wlG3ZI/zeH4gcC7BSr3swH9Nm0wh
SL9Gv6K1BU0DCJS1qIgIFL0iMtG1UyfIGEBNkPjxQoVeUXETvlEG0svgPBr2EQ/E
zThTHgLwJW8TpJtdHaTbRhIXYkQ0ZEXwZ3uCxYyqXSpO/js09XjPc3QnxKfjYiGS
u+c3NayKFoQa9N/q8vxhMK/n+NK1adS+F9gYs1LW7m9W7w2cJoyEPDGmwn3EKGrp
5W7/1cZC16BG32msvWq8zBV442qbwjD60bDWGYqYPe8MV0s6xUzrj5+3WxWMxDid
jbnN4MQvDxpV7AKUPXt/ChqVGBIddWYveXmWArkhwFUKRB/J9oka8C97/Q86JidE
0uaS5K2oych10XTUWINv22UC5pQBXwMCQ5FXRtQ4Oh0HyKFrh4/tcS4IPdjUhbXv
GlHnDF/AFvep5TC2aE0fODu4+JLnG4fWAhVIVhgINfS1C6JhkGS7Osw2NpyIPAds
LHrsxUOhQkwAJQo3jpnVK3grjDkhdSffeGCI5igVdyusk15Wdk3VCOuYD3p5W/gm
VC+FZaBO928k3bKBmWVGUYu8l2cF0BugjFp6iJGN5QrjVq+nwnTB/CPnkyXTvu2V
rWE5pdauXaYS0j4sv2D6oZxPHWA93hPCrdL0OMoKdxKMWMkQtaB8l5QMToP+kq5v
eXZknQwOksFqCe5PMnJm+EmmdrIJjOEYGnsxUNJW+K+qYqTToixbR6epue+AjMk6
q7cKRyEX0DeZ8jZjMil09c1Z6WHdpYKsYfFxPV7YtDu+vsmWp6NWGIdwrV4grVMM
rs8l3YvFbxeqLbDQHUOWTL2dlrUSn+QN39/jz3MnGgPAB+11SYg12yW2MIyig2Dt
XSBMIm/8wW2lqALChc/a58tKeYkTCDZW/oXxAqtKI/pXs3Coe3Z3iAlPJCYmKYEt
3BmtqF3fNkEnw9V2rLWbN4vcFKd0ZQLGlUAwg3wjaZKRaH1D1/f0fWbDTm2TySVm
GvZx20j/NSR9WOWbajQwhedpsWB5nDQQ77jDO5lg2SrL45S2G8kP8dglcQff1VAM
E75dBNkpGPYXhoGVWiFf517zQEAI1oTJyeprJuOHa9jNO+WN4ibaBSGwy4DkrXqc
d8Cyr0DftrW9wfO83S9s+QVFtlaTlbk1kYup0w9+IB16egxWPq7lcm+DHM164Z51
Tw4aBgA7ujRihwkvh3sDpU59yaqIpb7lSiGb0wZ7b6dJhp5X03Jl/w+M9PhvFdX5
FGAhK2arUn2XjarvnI61SYnFyHmqdbOIjG1cCO4staktOi1EFcL9jFi8uKPbGpLi
/Hu7pJyidUF5pYUdItTFD8g2JBqhZDD/XkJkZr76dBkBHfAJWSeZn1dQHQKGkybk
99ul2dXZuwUovCInp2X4JYgHcwtWlY4lEtmNHdBQgTPYe9hY/6numUH0BweDoP7g
HQ9pf8aiNaBJsorkER61cof8MuzYmFifcPSUe2AWL/1Zf5U9IGIwEsoEvfTv9J2E
hnADCZHuHqj17hHsDi22pfuzZMUomdongl/tjVZjaZ87MVrkO6FBg+mDw/6rg5yl
M/7tJOXZaYi0jzFLqxTI9NTDSZdzETp0AZJ7qrM4FnFRnJMF3zUQ+PC30zaNuEYW
HRdW+7yU0sk6TOXH4qZOe3jCVh0gCfowVz3Y++U/BHrt8kOEhDWgM+hrjlzsoXy7
KTSZ+ft7sjryE64XXDs0AOr5vCbX1c1UvyM4N40BG2JGlbG7P2zES0AGbS5bkr+/
EXHdgOntl9y0BMq8m55aG38DoxftLFx1b1VqC85LhyfgoqTz29u9Tj3bA4JWCCuw
wGfNyHu2ZLosB9RWrPbKhytK0EgaKIUhGuJxkMU6ZPhHbw2fNnWTesTHDJyp5Vz3
sCVcgUEamu0JIEg7H46A1o6Hhliwm6D+XQe0bFiVdjIvXpoFsR/XlWlv3S5XkK9c
y2Lpo3DOvgsJtdqiwGHDLNzdIYhneFdFZgMc1nFraJRh8RV7ZxhP1IAAwu+oq/bJ
1H+CoohdFR4VpktINCnDjyRH4tziFEeSnAKH99GQCo/cERMapSwfdusgWyls2vfQ
hguozwLIF8e2NCN8oVO2ofwmFDjn3oGZnqitp/BFuDYWUc7wXZBv/B8Xk4auTqmI
qtgs2I09rf0Vv+x8FM4CTQZN1Y1Va15pruVH8Grta30f/PlOEQP9yA5RISye5Lh3
O1NJ4XfLMndkPvExmUByCbt3rM4pLFZWgs//tKmCUcxAMji7y3ibchf2XHw3dmy/
kUeQO6aaPOENfrd75PgXzLL99CuVSG7boJBwKH+Eoavt2nAGM85aVhe2G6R8Xg+Q
iZ9RHReL8jrg0Xd3EmgDmxqtTa4a3v/WYgv/1Ndt8+QVS23aWYLf+waL2GYXsXrz
/gHPMHQIrNrtsqakkXwMd9Xb1syTDQkjKaLBhzRvOIt02IBWGpaEor+S8CPVNt2d
c3Mod1Yba8sxqs4vpmPJRKxb5k1tYVNohNT3Wx+SMrYaOMxiR+kwIKCFLiQQzrAV
BNNxq/KIDSNim3+5p0FE9B4gJbWM7sK9Bvj2RJ7/OizeSWXVeQ7/uiEpnefBm9i5
VgSlakFnx5usOo/8KrUUJJXkyM3VE4ilszNiSh3ile6bkbf7KDvTVH+sv8JaPjNQ
WywKoHscjQ7V4kHnG/mXkAJEi2ds14EWLVRwxH4wCig11jucBo30YpHqPnHIlRsG
mv71UZe3ea46b+au185MSl05FJj6SaM920hWWwybhhbr8yolHAdTkAfW7jUf8uFO
+gjOtlBHvntU80P7m7kH0LLAFNthy1cxGixscPQQxDMnFg4iduf6jH558k8t0Aq1
Nxte6jjfET3R/601PUbLfn9OiZNbUxWgQkwiE9wYbZIWBDR8H6lZiwCVi8TaeH/Z
zDt0W8JIPzEs3Jb/voAvzgzZi47h4Eh5DVh0rUdruHnwfrVArKFi2ba/L2u+WIRu
RpThC+xaFRM1VJOpZltFoo5ogeWnjgimOVm8fpvBQWyXbpvrjsOsk0HkxgY2PziP
2o5g/vMMd0Z5ZpscdPCQXRTz7nZKPJ+QV6g1TlAvXmDrA86X25TTdYprS9nMnHDN
pdpjQIOdrJnGyhhFayAcqFoE+8ojpi9GzsksXqrxD3kRKfCUFUWtD3y5l7Zca4gY
Wu9joaKh79qdP723NOBQjmPENK+YbtidlRfDSjJx/qGOlvvf0yt/ouBtRuyaHOA/
cdrKONkV7W3KITzvK8yERZV+sSvd4psjpvhzwT6GyDhccZ9Nwo8m/K5kU4GexOJz
c9br4GQT3zr/mvRNMCgQV8SYwbbiK42CQu2d2Q+jRuAnPh9niDozvA/EVBZE2KvE
OAZo2bYkgBJ9OFcAkiQkYoVmVv498RYR79teXIesKqne17gES6Zqo6Kf2jxgOYpj
H5RA/0ehCrYjt4WlTCxwKkkC+q8iXgMFGtNZKPB1pvyCE+hdIY9dXxUx6Vntjh9k
AWCCIrU03gj9lnlCfsJ2SDYDGB4+/D3BT6vNG2AcfVoaVYvb97Lxp64CZllrQ6Yu
vo4dDjLMvB1UH40eB1jIzy27eDmrsnvc+7ETJOVb4sye8NqVH4rQwXxdOpMBZfQn
+ys5DLRVCOrF54FVUvI2g3GcWmVNB89+9QlQ5ez/LZDhpUnc8mslVadNNBeygl7U
b5BgLF3jmf4l7GxAmvBm4lI4GjfEATcm79lWVfWsEnHYzmqqk1vPqm1ZAkl/1ke+
YDG9tl5xyGIDiZystDiJ1RnSm1CFHK+PkHEZrVXDbyw7l5z7slEpF2vO8js/W+xn
e6dLGPKhcF5OL1u2JnNWIlAripKaRWXQpVy04ViQX3bj/d2EdM+DhzvsGyv0XAn5
hmM6r0qMYFIYTxDaP4Gxof+c47sNgdNZFypyo9Ke146+0sLCMOICpB9ronrUfYsH
/UqAMr3wG+pkUJvokW9u9oA+bLOmrQ0aSIUhjwqqUQDCNAZcxXLhzM2Idf7hpVS9
FtR506YZ4hEh7hOOcUUzOrgk8Drt1d8k79x+Ywo8NeGLXGnjkMJ04mSSexAZW3AN
CeFM/oeS4pFaHziKyVgvw0soCBPCOnPX+51HDLYSKpXTzuUr8Fblq9xK6AmwSEJ3
TTgjlSaGg3NNyX0FqWObUEm2qswQtngnJG6KFYdENF/7zLW+2ckJmrQSTbaL8PKv
nF4ger3oj7IeazuOGBHg8YakT4c8XeCnBU5oBlleJk1m9qHp/O/32Xpd9+3ugDH6
CjlSAlQFvMQLoC5DtEQbXvW8MLTQ/t+6nq0viX9fP7pLoroHBGQmu6TAmVGqLO/J
wV9Gx4LOvDBjdl+/7/7TlPxGPYMLrWLNiACgp0E27fdGNgIlOQIb2xRKc12D1hZ7
7yYPBX73GkOVGOQbRACRXZUX7Y5qIjYjzcaHXpDqfQPqQYBeAtgXEJvrFuliyn6o
CS7yQZmYkidKctiOgoLVtC9zGyOZeNWoVdxHdzSlCh9H/wsjUCMxaXxC0HY16nPm
hfpYDhycz57v5GZBHHR3yMxgk/cVsxGZ2YX6S1FlcfCX+t5AEjhPFsTylS+H0XY7
D6b5z74ZFPBRhpbtSVbmhrHEoVii0xETUtTxizalf402FDGTW2pcY/Ks5OlYax9t
PP2o/cgqRh7v+WRw5tQdod6DMBm70iqnoMH19wVjKaJ7wXW2N9GOwJnate7/CQJX
crx+FMuyr03jfRINubUV0MYG8UnqHYt+WwST3ZwsuiL06L1gGDLWWO6/eFqMa/6H
G99/pWYOoNrOMaBtbaPpLwrpoZgoiAt4E1nc+SMnixr0djsYU+XchSDwqGqK+fsK
yAZXkXljAB4EcEdfDe0wmbDkY6rK37TBG1kCtLhJ8Oee/rXL274VIYMFPnmdEecH
iZCNv5O2Ctl3LtzAwxBOOyYw5ibCCD87jlp7UpGNZ5Dy6Uf2zzVccubia5ybsnZT
RqomzPD9svI6/5vCoBBdTKhNSdhbTIlrg87qBqpgKfTDrBS91XEiXyrFn5HZmc2I
2T+tlJ/T3lzJTKTr8ey2S5sGTc+RnAEf1izo4proMl2saK3aIQ6U1VN1jTF97Ylz
O71xqUIxwLXkzIsrIHXehD/QTj8w15R+cSYedOJx46DlPUwS511iCGjvEUF+YYHY
FDDflyiwVn7rFvSV0axZHNKbYUdudXiSNinBU3WoW80+hGdbd/oPhxxiZS6f00qN
C90Fl2AdatqcJin830OQWCcfn1z5H0yGCbjbDOCPhAp6ZOwxtB2vPaa4vNuUxqNb
Npg19R6W/ffDP3VbgUUv6GF4XQJFvTyG6tF+JSy7ZRxJWmKzTBKG+ax/W+o333Gb
wSIshJX/wgQLVXIlV3FtIoPW4zBhS/MXOqZm79VY40bRWnFaTUR3P0xBOlmmtb8T
9WHq99QH6VD9nANRrMjnNxktD86iBDZ8pw2GDJz/cFl4bCNmb+yaaFtp687i8XsJ
vOY3ufqVJx/sy9jcYjQZ7RkrhKegJNbAz06Nvgr2jsic0agcpHFIax0qpVwzzShX
CISYMEnF745ghA6pI7aySYU4E1xmMRYn6KqH1tvzlmaFg145LsDMawctNVjaZXUc
+FTyFyaZBQsMrgxzfVBSBWejV3cPDZIYXF4avbrYRAIm9lEQpTJ3PfiUMVaLTsOl
9HkJmQ873voK4Qb5Wi8JyVUL02Ldx7NGxr3848VntpVvZXmSdxWoEM4OmkNjMG8b
cK6DU+lLBcmEPH7CWhT6+sqLavXnZ1Tc94psrHSn7sSZno/myKnZ9kOnt1Vlzoqf
qzYBt0YS+BZk3rRDp9XGG3YbP3med+4rMEL0hurywGHdmz/+FkbQKNNXMhebFt3V
OnEje/w7M7j+pejI1qCPFzWYtuGIltYddS8hTfmkqJroH9eHEqVXPJYvEDbvVU5n
6aFMDUVuIcrD6bMRwNJioC15f5Y9QGkOBJuODv5iosh/woqCm9iOIfcOjC4bDTU8
nnq/GsLtWXKgHuBtyNPhbILmSyRnG11rcrHtVQOxQvF1cBdRAsLs6Ygxnk5Z3s+3
hkhkiplhhCIhzfNgbx+P4HP6NvsND3Gc7A7AecSlplUQ6c/SKPNDiHepkA7LDx5W
BpzrZLkHl/cctVzya1P85BayC+UamuqPjRGUwBeG/Prus2VuUOdfOb30BDgmGaJT
+7yTHcH2EJ3i2/IneG2Gfqze9XKbApTR/TPtjVvlVQ0Gr4Q2TAi/k/rBO7G9YSfc
tXPkE9CmDeFO/ybHBoN2rLnJFZK3F7ZF4JbVbVCsrB0f1SFaOnecpIB5myx8WkaS
TAbEcJOeJNbqJs09viV8+H4GfXxsFSGCE3aCgRjQO6CNG59pw7z5PD/RBbZ4CImC
Iopmh2cBpO+CFG+Z81odZaF86RV2Bdx+2qlkMaWG0hVudzCdYOKkvq+jCkeQfn/c
bGMmCjBcWD2kdxPvVmLGi6lMRuYxjdX8GWagwIH2sEh388R8gKd31tQPDu9YaNMO
1nQQLLUCo3KmkJ9TNU770Ie9uS13XxE+5YThUlrH+kOKANgfqsszWQeW6pxmDr3R
C1JnClJ7WTiW/E/vJ0+8LG58zxSvb8EXoNNNzSWX5Lf1XMwuWXy3MblHERnq3ixa
PmnfGhyAVT8cwsKohxb7A7VhSb8TTVjrZLaPZExKMkXR5Gjp2oKNfNQ43Go+0e93
jxb2WTzG93nTB16XIMuNoVFT8OtQjW9MgwCJw4/8B8897y6iFpj77cHDWO7pC/bO
tQJaD+UC51Glj+dfqGRCrmfylFlUk5/lMn76EQ/XQZHTQxDJ32MI4lUdo7HiREH4
68vcDiL8Grt/lLsic/DL1x/oK2/W+x9DoVvfblo1dfVGi/AuNlJ3sp2n6t85j+Gt
TA4KS+oQtNwPDEWVKaj6i7z2q/I/3sUfrViesU735tgx1rUWxqjRz9rY6aEqzZTs
+k5/0IJLE+/cCJNszNvJ+iDEukzf6QhDKmeGEVUwdhJ7qdjdy9X48rl7iKyJeUld
Iyurk2/lQUW/XuJQ9PTAJTWoadL61M82bcSSNLBYjUWyuVIB1wiPgPoKYrl4brj+
I4bzxoIpcDcDb74tgWarXT16j9Iy1VFfR7XA+aI+euOyamVRzgcSAMGQBlU593wm
sng/kiB6mAfMfWUXfwG4A/YZ8lpFPjlug/XRJtvk0BNpNwlLC/9HOs93/Z/WwChq
fMHhgl9ffhIx8G2D65VOjlYvjVNoXTJafOWz1MB/4HMtAJOIaSkGxTNmRQOu+dYH
EV6Yk2nm38GHfCAGWNjc7qbuxr4NtfMaOqDORIwXZ37hbNgxXqYlIHdF9rRLDQ9o
07IYyUm+dd7Tntck8liNtf/F/TCg3/XupsZtWWY8ha5C3IR8wmSfy415GpSG8b5A
HtZOirgTjRUSgPmFjquDeuvl5a563Oh2sgDBCxM07Yh17ZIk8XzJlT/wpTMsnHUz
fEUzHQtet/ZayJxY/S+hoO0k/XMfEuJrsFM4mwAU6goXFvWjDveSV02fzXn1fOoq
7aghGwzfwc+sEMB79ucCF7y4udC4pa2MF/9ZGPRuryoMeeie3LDjpUcIUFuRXFeV
4TiA4xD/cPvRUdKQXwcERE2RFGmGLp5t7BKSQxDqiC89OkSOW0CZ3NR4d18DXU8f
NtIeqpQgQojMenL8XjLLJDZTyU+2OVGYwrwfQkQtZ1hKX07rEgdJBy+lwwKsbYwm
wJtCYhUxmYdKae60fzYaaWOcfOSK8OsEbutQueyAPPAyu2k9r+ZNpPZ8ZQHpPwi6
CSmZ4+eGkjURqbWhu+1Qt5FydbsqVuXX3U+g+ohKUavHjJnosrBS0xvmJKqis2BV
BszxxO7LfildDzFvYqFVtKAQjw9ZwWhY4Frx5cjvBIxypK44G9jzO3TNc+pjpDwS
8A2Bhnik1eRyR8RI/hHKqgmFLMKqfRz8T9Bw4HNr3WBNEP4aybARUXZbj4vOWfs6
sOoxs49gxT+P2fLofgJD4N32bkbAHO+9SqRQoR4ad2WWDmtYMCtbipA4lw9FvF4n
176A9trOhwvlSUC1gCrCkJayGkif72/QCCvGQCz/+Ac9ynaDBsKWb+KAZWIUXBwf
VrS5r6MT9RC34f+iwkm7RhDVV3BnrpUKb8B4WRJ8a7/usEDmVjoH2cgrEfG7Sblf
Pb3LKd19lebmmZdvrMh4Y3Z9GgUps7s4FiLYJL83W2BpT0xAN4NbwPsbXiR3usV+
7sEYMi5mBc+wBgfpf3JPbtX7Sg6MXlE57QYIzB/IpUfM3U+LyfVrBXZc59LIchrh
Mu6ByKzfs1nvMrpxNqPVMaBtEMQ+rE5kgxtiGAY1sio73ZBpc0XiyjR8PRFQCbir
PMz/K46HUkiKGlyIExv9TYUo6/lKr4gweptxrJl0w3j26zizNJRNDdSzcLGHhlxM
XsL/fBHY7UEAtr20Dj0sUbLWj4KUm7SIXrarlQHOY1PK32P8qdZxhUrO4dVZneAX
q6nVgmyB/SBqV1+QzV6IbBDOzuAScZrxflVcmk9b5a4oXHk7+CfWPEmSIXUo7e0N
Dc/QPQsrc+irG+HZ2CT8qt203dyc0+C2botsFuD65CxwoVbASXwp+a1V8OtnvhV7
Y/CPJs/X04O5jFTP/KiPDsQgR6i1yRajRdcuC97objedN9gUKVeFXhhFktJFmcOC
sq+ziveiD0ci8qUwWXaJt9OKGyIuJlkp2aUpaLksCKRlPkB80oAxZpGXh/2PNlHg
xdNfFjVTvBAnxDjv/Qj4S2ajPArcZQmIvYHClhgMveEznPttsWSXWcq1Ns6LR+8S
A90yr6EvYCqB5NfGfIWpQBkYgjyuneb2PjuGkXRokj0s4E9NGNQlNe//nhuONtGs
95BjA0jkptr968LC+6a+PaEcPfMalw0cQPVvAPRRBPvzu0ZQHLQ5Lqr9apA0rvmR
jCKIHCISyxSp/H+xVc5qJx3q3pTKYP8zUwTUzS8RD2Zr8JaKXAexwEdYX41Zivk2
FdALdYXXmXxyy92qlIH9Fl0W8rln3dk4gV/+e5BOF01YV/hVvpO2vDOptWSAZ6VI
ozENyUG7/rLnc/Ty0ylLAl9wjTd1iWisw45GqOwSYo9utDjCHZatddWJqbDM7Kku
EF/BkjYCrPOU/nQWuRWQvMvWXwq8JmQnMaq28WCeXMZ62Bk652CLSsHpEPYC3xhs
Y99oYI1y/YWT0ulFvd2tmLnA9cZbCGrcNaeGpHcGx4LtarBlNeay7s0BpmW2C8kO
81yH4Ibl61Ylr0eKug0vqFXmC1Qoz9jODUz93uy9eWlEcNM3UoBImGlv2RFYURSo
utG1f/27O00DZXT2U+5Eo8oxNUTcoKF87fjqbnJmfusA+IHKT9zSRRPjO9AYhxIm
smQCqDpKMJDj5Cae7DD4OQbt1GH5NtELtP18tIShnJUtaV+1E5/kUSIkxy5DRjyj
hOpxDjn7n5+Hj1pEp+T/k1HycagKw6iLeM9qjkAD82p6dt/LfXD4OBZhu08Z037t
Oz0+m5Eln28Sg9puUbbK2ynBG+BaPKPpTGVDdt+OzC2bR+pbuX+Dv+c+EVAnoN2c
40YFJOG6dTh6uzbmzSEfWEjS6i0T+38JvIiFm87gfPGG4f8d7/3RrZ/D3wx58UND
XpiUMzhCk2D4A/RHy6k+Z8ooBT1AcioUqQjSF6DsTwS+xuKBIfBBXvqek+AOnJnI
feCsbo1y+PBa047R+f8N0Ew2gVHxwBmgZ6GEhydfqeOoO7kFHPQusTEME68R52tj
kc0hA3Fe2l8gtpF0Y2IqIJ1S88W29Ty6S/wbRciKVezF0/l4FzdbW1S2Sp38NJw5
xvUtAXI7OfVx5xugGoVpBeI0rEvG2Gr/hMoGRnFUizW8pvn77BIcDOUDeyVHiCyY
WHbZWtWo9Xx6s0G3z2RBhNe3dKCxS/Segg1bNsCR1eEOsns6Je5C/S8sIQsn5irI
lk+BN/LJYK4MKsZZbIBBDOQNHT7m2W5OLzeVZ1rveQOs2znXlHb/MBEoK5+n5gRe
7EJs0Y1EkUC9rPVwRwCVGMA+WzfmHgWMYSlaJ7CkWgZAQyFT8TIagiboO3j6YvII
MjEF0bdkivOiF7K60LzZTM8C68Pepl2ySHggADf/mFJL5xJQ8MfW3mm+SJ7W9lTV
iLqPCTYvdnKTAHDVw5Bf+OyA87cV0ny+6+SMHMZgi2mVq2tRtgQnJkKFMhnnqoUe
Sy/2HZSlp49u+ZS5LHL/KmXVFYVeo4hBH6wQBgwSlYgY8F8EuxNA4Rx9P3oenvzc
6dTEjsUhw4YPlO0mlnoYedXtFSXvRcu+/z1QkTxdCrfnuTsJUuQS4GBUdORTIGBm
cZuR0S4B0Y6Osyj4KIru4GTq8WJk3C4NxE5ullwhSrFfq+Ua8eE4JckypN0oy+hv
yphaVH3bzQkACZSQ1IRey2ilJQ1gT1Ht87E1hiG3Rt9oTUvlWxVYy88g6WIRZ16k
J3nrea+gFPs4Di95rYKMX5RVtijS7dBQhZBHLRP5VqjCZHlwPfr3n3ukOjR5YAO1
K5kxSQ6OF0mT++QoMzRxsAEoVtgA4bYav28kmwVypI2bBWbEpN58DyQSNg+DnzDV
6L4ZjDIJ594qBm7cUYk1ZzJ9MmcOLETEUbQUiOEQOOrWcZB7F+UGLEa+SnQCXqpv
BDjhHJzX/UhSiba2MmSN+VlyUPbDw0GAR4oeIJ2/b1C/FDUhdI8igR8KXU7RMkX2
TvAvS7CVWmaos0S3UznIXZSiiaz1UTl4Iz9JGfdE21z0IchfQbMFHrhD0akVInKf
ZU1HGAcG7ONDOBHYHjUDc3LFigVhDM5TJAraJZUpaaiJQ6hZ4vXN+b45W9Xfm4zJ
A8Plph+UALwpKiHAvQZX7v+gh/OGpPW8yrJOtu3qrSh5kuh+c/7/im9tJTCF5EKP
/7Jk3beBFGg/rk/FtyyEm8jBqZaaYFFCWCKhO8F6dlLd3Q8V5Cpg12Kssy/clnqH
Bcfg+ulH6sOFgI7arEvFmuXJyYwbxTU/DOQgRMOOlg/7T3f6IqiBXgtYtYsg9DIe
0n/C8RzGoOW/s7FGNkUIzC44ksu73CI4Zc/7yQSlCQhidbF7aX+U0IDrqzwaf80a
l8HPUdrWwhZ/nmeY0+2f/XReqLWnyyV7lJ5HV21hDNWvuCo3jXcyPxCadqNZNJHo
4hZkpUwKpS/E0blMhXxj+Ft85FW1hQRjY711IBCMQoqxst4vSjpOuhXvBC8y/AOM
JaTi9vJqxAx1PFzwi+/ZNO/TBxU+boE+5x5lJlGi0XR5LK72pTn2Fls/YcG66bGJ
Q1lenLA5wp2uTVD9/2DnbJRT64CMGEXcUCni2XRAjl5+Ao01j/fP00D2uRZjGi8/
aH4fwS/7znA+ddSTvruSP5alHmGy7G/pSA9qmjCZ+cd24X7g8c12x+EBz16zAl2x
z71Ce4EN67vF1RnZMPSVOhAhpnzlQN7CA7F0877u0Volpcf/DzRXpTAIXpKHc9Gl
ZyymXb2rrmmi7XDWIxTN5ONibKMi86ifs4O/9k/N2KR+Yuwn1EtW/Paa5zSx72Bl
2p6GVUPFTCiAijkr7hTOpJm3LX+Oj90RUIlZtRkoIRQubBqIQGM4FXZu+YNfkzT+
xW0cnSv6JL1/fanHbu8Z4ZyX3QhhaKjVhWqaDX9UCxXeJnFlnxDd9lP+qHBR5tVo
KMcQKeoB1l2EtII3es7/zbkjUMBPU3YiAhta8IzxqqsSk5KXWRkVdMkuXOgo/VmC
yMhEyLJ07nTdP38m8aVRARg7JKM63UFSfh7/744hzK4S9BZrfsQHqkVYwxnLiu+5
K3P47l2O5scnJwKyFcUKoESd9AoMOQyCrUp15Ikw19RwB55kqeEBDanWKkn/Qzul
N3KEXnkLuPlMaVfksg/Gp1gLQTNxWQIitXoTINxG0RFN0srRB4W8tDn3lTBnqD9J
EmJV4K+5ZDoVnxPREWDrgnU9CcaCvhN5MXZpf0uOiCqqbnhYNjTyqCkNMSq49/ZD
O9dUmBVRd+HXEL4iozezXYW/BwBtIjBbE+qqLJ4tHZPUR4WG13yFHohJU9Jc4BYm
FHwZXlvTR8hhb+qzOgBn0l9/1J5VSmvyE7jSxOxz414DrBoW+Ik6fKmJz44s6b5a
WqO+9CleECaEdad0bobWh78y+zjGr8ORTbg8VfWIjEpHIBBdldqdnrrqD/kcq1NY
yKMLbrSG3aM8iEdBzXWw4TGioC1V5mZtEekAV/pSuOg6+wh0+gzdWLgNhzMJoI0f
RMRnUK7lZMPfoPJ3pGReBa9HdWmejUihDqB5UpA+HtyCpuBx9KH0VMOHRngWTsXq
ECRLhB2lWsVfOFKJdXKeiybJKWQUN+WjgISKv0O+Mhk1gJlGUSvVcBosvEr1oeA7
KRtRuxR7khdHMzoLaa9paL1mRfnOIoStQjdkphvkTQk1CQHc8+mkWe7CyxMOZfpJ
da4mcYYTGtqDuCDasZTE4gkId7gX5hgyRWcOOvZVefD3kjUKBStOqDIKqc+FK/S8
kkxbpNcqHP/nXjhobmlrRaj8haKWhmNz8yANb9+daAFNeq6I4uZs5jeXbeCuskMq
9zJSvW/+5ZexEDjg5gpQwfsZw9khrGhAdgsTynvFQhWTER+DCmJ9PGQK7vRHUTtF
uGDa1/+vSs9iMpiP3GIIlaPWLt+/wc4n3tSv7MeJLI2TRAWobup14Aook2YNlN+6
tl7MYB/FFkiy5RlWaqN+SzMJ9ZtzcKxYf+6Wm6eRuIixjE9mO5dCud8ICdxUo5nW
v5oUZTjRuoOjMMoE7uY0DmwA2g3Ek6e88+2Q03x8E6wCg2aySAGhiT3JfxTk8dCn
tx4XZLh8K7wjkSEc3ZYyqAq20DHpJNNytrv0IVpi9ZX/Rw+7eVtOngv4zTkEzxOV
7et0K4E1dpcE5lwTNcvb0D1i9NV3V9Vr6T/GBPXBgneCBtzmrWDJcR5B7cgz1bsm
AsKNXFf8Qv7knMLX2EkARU5RBwU/2RqX2k1C3C6Lzs9kkwm6ROP00E6CDmV9KC1L
4Z0PV0lFAHmBAd8kkf8ZU8/izr/7dLjnVrcO7I9soYaxggMHHuUfk3QlQgy3zElE
s4POTe2o64YpuP/01VIUd+p/7IP4qWlgJSDH1LOLQWwuLwniWG7uW/JQmwRIdgwC
zrmhb4/sXQV3cP+Y3CiANMp4INS+H4Th3XROxDQtP65ZTVH9UOZxhET/ZG8ZwZob
J2irJ7KuovjnptG/zBBLJhPVb4lW28hDggFEJKU0WjInpa5xdizM5wCD9iunloVt
+Ajcw0OLuBYYG+vIVXly8bxWou7gMZBCIKcTDkCFYYJuGxEQon6WY9LMP7OA+kRT
ui0c8WTIa6Gcs/69TTfU22tHDecAcKsb8f9ESQRbko1RIHdpUNNENldkOJ/V7Z5N
eydgAENLtFhRcy2k+2l3yxVP20lfCruwd0Avp02wF7g07fETPnmCFNXAOvCqGXcl
KTbBT8CgwfZxKZWQ+oGZ6i2Nvev8AiFJcYN3Cg7csPjVhlDnUQRqUye9x19YGqaC
xUSWTrgapPm6d2rfqs6ibxi6BP06Fw6b2q1xh/U7rwi7rPpCZIJ+uuVrcYZW2Hx7
bn2b7JGdtnOuaxbmW0rIGBIpv23fnpzukD1N4hQW9zSqpaa6tlXJH1AtdJk863Vl
9jgxho9SnWj7w2nUhDU5WYIT4X+LVYVUdw/fg6PYiRPzkNHgUfbHkaHpEa/fSy9A
7yIFOLRHvEv9wPw3aNY71t0rhty8JFoa4YfgWJSrPVZ1vfNjsi1c+pd7mws9BFlj
jsIh355bep2cQIp7g7Wuvag0fNCBYFhgXJ+mkz3csxbM+ZU05nTwdYovvLkAXseR
KCHXq8j2nEE+nd3O+mw44SE9EIUC6ufqmgmUdB+G96PIr4YVTWfAvijqNRi0fgyb
DCRrXqJ1dZYjeFALfVXJtGtLsySHK1ND4J1sgVkr0ctUsWL7wYRZAcbjYb3bJQjl
CaQYa3YaUFY2nhKVyUVTcFVimbVDZcVcQBvjDXHKvZKclTyZrZzO7w8ifLvGum+4
hmzmnAphTdgkkLyuvuIbptqRJWMTy9ILuDgi0gwjXd5zQF2pTYn64FJBDd6xBRg1
5LO2aMwgSiH2G9MZrt48hD0yLACEFtKBenlHx3su3kq3+w/l7tfx296NPpjRIhUp
QcIPEYUyKu6pTkUzeBguqxZzlNbqEMT+MC8WDcRS5+RaqhvHu6LnB1BnjaKSI8Fk
BcDlpkR37c5dtouQylhoJjcZanscuE35OAYBJThc8GKMv1kZh8u6b6X2C1Axax6C
Vj/ERiZhxHknvx++AmPz/0x26Qbk4VIuwGLBpiILJSNI8ftcH48T6jQpeU70Pfgy
fOFD6fBvl4qu+E3r0HGvfHcjM/F+vhv/fmLG5DNc0Uxig+/xms7nGEvr0HQRQ+3M
G8IG3ijeCVdYDnxm3e6+2rmfalfe7YNylL+Z2V5JlkJD5yoaWHNcXarK+G4+1le/
6aHPk9SfXYWl9mlRxZD65K9vdpgcvniDpMlAvXG2CuPsqxkdBXPuil/sn9tUFAmO
M/rzK46TJryvYhFcNfD2QK7LAEPyaj999TPwDDlDwno8gMKP9iS05xaxZPFBjSNi
qL/WxbKWRAyUwJgBcQxbXRdqwoRsX9u0Sjk9MDkIutcUBFcBORndpWW4ZAYoxtZ9
XVnw9BjqKivnZVnR5jnr2KsEMbl8iGQ2rgiMcYVtl5BQNil1HKc8yDL7BoH1HQKI
fCQBN+oRwuVfJxiNy2HfQLT7A6tHNhAeUdBmjpGZ+zDVRznoFbvYYIvcUqfYTXmn
LypNfJxOME8WWqRvVPNeNnrLHVKFrgOpEcCpe28oLdf2Wn0vDC8nO24ifoewoWDV
7N3yTmd/OP/T93DWIU1xd+6AHfMygVYldmDsLQm2nnOKa7TIbejeWXOyf3qmqDsY
QaZZarDFQqUCjHnK1z+o7y/Px22HyhXd6MTPltX3cYBOFqTv/iSRCt/CEoVPzU03
7Gphlr8aGRMi2ovghH/gdKDff6qejD3N0NHX46ymaqV3hUfOo6oLRXPPWceiZbNz
KW9VkvoGKbTtThULh+0M1lkOHkmwCO9SH6th4vEVgUw5pGGLhvWKBjE5qnp6MQeQ
kGtJ/vaJFYWe9GeL0uiYVOC0yJ9h6QQj5Vj4zOXBw4cc67FCoJLjr8kEuvUYgIkU
c+EPkjToUmGHjSAwHrcFJhviuN49+Y7jMEmJLCGRIF2XhNwtSPK4Wv7EzZEZ8YNU
hHXKNAat6GzYDY8PHMPWgWaCINbv2MtWM9BWkDsXQjBujb3aWBupz4ECx1CFCrsp
qItjFcOViWKKuE1BzXsfa4Nwc4Jw6uimyOPu4lYsvPpJnNi2pPUi8jftz9Jq9k2p
vUV/2TBxRJe5GGS5pVc9akcihnqKqRWet5oSLhmvW+4qR/Rry9IJljuPVJxoS6o4
IrVgLuGT+rL114tQC6g9/aHViWezNR5J8wFFeGwOaTIuSO8TLPuJfUwCC20RbVvb
/J8YZRlua88188u3Y/EpqZJxibCr8d80gN8Hnamq1vmDEaVDn58HB807XHaC+pYY
SmHT1CrNAfJj9BtXY9VgA+aUooI29sVrFQPOBbnsd6U69iSIeOedCNDqvxMVwmyt
/a07wOyw55CpR64J1mne67/n4+uV4g5NB/qCit0VHD8bp6JAyMLwE4qBK4B2IbSb
7b9st0eUXf++LOVeTx0IK2JPOj8X+N1eqKq0D94yEE0KEZBvFoP7lk5qkMtykAXA
4IrE/Pr1RXIR8dUWWRsNSHelkCX1cxLk4jDGS3cWKwdeV3UfiRVh1NlnyOd1EDZg
A1YV7GQEtBKGVdLrHm0RxWzwepPOx6DvBHwF8U6dnCg3E0XKrxg4md887GZqDDrl
haB3I60203KeUiL8fmjewtbLTjiBcBDpxg/YJo5v165ZxWYwkbtZmdZeVHkH/DwX
Ue1Gp+5sIQ2TjcZpz1c162u56NKUyCN3h8hRQWctV/GsescslsLi56ZjWuI1hM75
fMVOd1bJbpvcMNyVM6I/PwDMKUfFKrU6Qw3vcitk4mgtia7h0nAM6IG79noy3Wuy
/H5OAZmKu70HZ2h+Y4ohyIMvaZSIkj+fcFdRp739rvM/TezGzlvf7kp3HtR9ynWw
k69h+j5abvikius7QqAyyvPa+ZBS5cREjvk5RRLPsWv6NvsgZ4N25QM6Olk1IlaM
52KjeDDjD7Vm4WdfC6medcXgiT5rx0jVd1NC+qySWHFuB5FC9eaiem2EIiVa31RE
KYkimLRaOnlIYonTg2AvHWj+07ogOLEXiHZIo+Vh+gvJ+dhYi/8KB9jf8U6NQdTV
M0R6wKmYe6C/TRtsZzjyho89N7iFNTTQxaomxTqqzF+n8WMJweaVwl5/oFuEIM9M
to7lznw0Jd6JdJbkUCIn7WcIUOcKOevk+R7o+oYnD0iPmDfq/2qbNZ5dIXtE0Pyy
30fXTYT7P+uHpqVhI7ViDxJgt2sraVVP3CapqydBDFv8zcZeHU1LpWiUWFtRJ4fC
88Q2n5O6LsDO/ZGAOX+zHVVLqLJO7TgYK2JVCEaqeOtDB4CHqqcrfWpPdzk97gdS
uZ1/E4Z34rCFxtVolNvc/bPzy/UHRjRGFHDltkO5sQtG3E26nR6VfAOWNLlK3jFx
2sIqi5Asyq0AomHPf9ecZ7xK4axsESWVEM3GnmbLlbVUJnM/pxosK2M4O/rNaNfR
xxVFAiuNb2fL68xA8bmMKpE+T3v05vQZkOoKIfITzsThkyeiHp1tFFQ7cRS/4W9j
3c088vvoVuXMg9plCqBSe2cjCxp/b9vxY7bfuRl3HLjEpBYRHLDbMoTc+5dlLWSx
imz5ITTITE1EOQUJbXNqshLEdnnvK2pwyqdvpaO9eG10K07XMWPO/kOlHc5XILrn
a2VhEOhPjR6MxH7mCfrq+VXnlzywev7awzvKgIZ8V6bxS5DPHCALWl8KpcAEiN/P
JLxa+8eYChFOUkMm+Wc+cVk0j3NPfJKw63be/V7sKm2fPiTRQwsmoy0SWW1XH31o
1ax2njb4BUzqqvurdnuKtCLUuUDCMSqfXhP+oW8dRLftEPkR6d1xcYHCVXYxO9fu
X3RkDCqjyb10riWeBJ7rBOO5/TzW83Bq69WZf+ymnY5kl2zmHOUtaF6cuz2K+jWN
ksqUwZRQgXB0vljtn3tyIdhS+9n71r036goJbJSOSk36Oc0BLGCtKDjLZUH2fAsc
VankQ2CYYLQn7XvM0AUEYGtrOPZ3JbY+sH8tOXEBK9TizQBgNe72uXKCEzVDHn79
v2ttk0L2Gl3GbO0yBd2Nbyg4XpsXKoKriF3Xwf9bGIgvC1kTF2GbFVSzp5gcyIo1
SB78bm+fMuYX6kVMt6yX5msMbdjg2EwqSuLU0QQbqQoet8LhnRlPRRpX1DDFE9VO
aKV9O5b8r2Jr6cW/Kz3gT99UwxUW3XNgw9nehqWydwN6lli1o2JqfZ2AMv0dA7X6
erzOAZSV1iuW7nFCbzwoa0JV4pLVEMNPencSMhbdHgWek6k26ThrSgMzGZy3oOJs
pJkzq9YYKZhQ/Yl7rKUfYEyyrTA5XXFzA3m02nJ6ClrBuT97hqgfusCdGhaz+Zyp
CL2kox8rwJ5hPKyqu/MDwUgQlEdBanUHK07mWsTX3arMaEN1IaIZyuRETeF0UKPl
k2fzjcmNtUxHD2OXBBsoxsyPGWR3fYyWY1LLJ72i0mgktGfWivAxeOtJ45f2VXVI
m1sqin5R4ddJkRVDr+kum1jk0QenqRyzZ+kS0JAY5d9M0G/1YvHHEGK/C1Gf8UQS
R0ExQCZkU24N4cEpEQsSZrz4PpJZPAzG4YFf/5Cd8oAhAUw051lt0B/TjeB5vEnl
PRDq6dJg3KBgBdelxo+XT0bzxfULfA5OBTh7AyKJTGigtIOBQUPEgoQhBa3gzKMC
w3p/KbyHYUT7RXqb9Ht7gnodKVjGDx2H/K1zcPASNKQPvbBJjBSSlo6uUTDWkrpk
4Rrm63Ge21wkL4WXjkEzM5kXa4vNP9LNFSXL/6Z4MYmCueb4H92gvmgiORay2ylZ
wDz4HbzCtPtCJ/JbOTiNG5AXjZGh/WDUksVbWXdYiPzMFM2CH4WZuKL1e3G/O79z
fx4CA6xQ7JqGNJyW/0gwOFr9g5LKKxCG0WFwlv/eA7ujOGIZCyUg4+NAjVmQhmnf
gyNl+l/y/1rrlyaHeIa5Tty+CpAPJ8/NQYoglVhHR+mDGZFUfq6WmVz4eSVsAf4M
qU6IV4VbXRLW/mF4nQg9N7uF67jMAjYKYHmp5qKPZZNJlBaNlCXA89OFqin8lGMf
VE40rlCjtQuGKvEPL70eD6S5ExBojcochBHTIIhqqbDKOR1I13BqC2cR0/SVY8Xf
TaUpjEDGDIUaCNt5hQjBJVV3UDfN7Z0nJSIt9QGDQe6Qvkd3dMaSICy4OWD3dlaD
W8nZ7oC+2tPhML886CkpuTmH3K8lSCQeohyOb0/pO8TR33YuxKbxs3dLYyYz6kaf
AGYEhLdawH3p+yctvH4fRfPa2cCaP8rkv1OYiHAnIMNn0a9XpKl89D+O/4kp7BRk
5nbDzsYy7ssG33rZU9hydCdm8hgdp3ymSxgxW/f3V7ynqqznIim6SfEuvGder+Oi
0naqrws4njHA1CekNBJ2Ir86jozZ9DEi88vgTBQrjs6+xvVAAgy5yv1ClTGakVs0
pyi0E/gyZGOWdqQQ0UHFFLzITY9E85ZDnWPr6XvQnaRSacgjEC8bnOgNxe717lFx
12wCwgRfLwzLW5A2Ek6KD3NTkk7ZVk4Lfg/7gyiFW2oI5Au9kj7uvi/KBdr8e50q
Rh7W0t82HltsbR/qZ5uLCyeg8uUKvcjwoyW7Rf4CXx+kWv0NX9qBO4T9qnLoXpEW
Jq4JHoIHRnBG82kYZzB6QILHBjCK/0zh96XtT1fdgWFh7bBgnmiUixlS1oXolgPG
KjbGFqJHxh/V98faEGg7Ou/HRDE9SKmVUpE5P2s7eE/pkr92Rk3eF1ZplKPEru9d
BSbPw1jWnRVtzjCtExVjz0z2oAthEg/LB7l9gQ+LaP+g2PtrUVeb+vpYnOF9+IvT
uZ0s+9ICruXSyL+u1JhZQSJI6q2yfxoV+8VpqImiFB7UCa4XJgw39mFQHaL4Qjl2
w8nm4hRPYzhVTXzgQk1WG8VJnxQwZT54iVulhsEofQ4INhz3rTn/EJIBlX+BQ4l+
YLWKARKLOaPK/zA2yUGCVODOrVgQGNbnwn6wB907Fk+LCkaBfjfeQuI421LGgj1n
G+wjj9OpIyOkErVqSZ+8eba6U1fKhL/vm7BYvGyQ6bEbnFrhexMlefNEMe4fErqo
6x7W+9sUoVxnb9Z7uEp3kV91F0mMxfcQBELEt+jUHogakeO380gXOdC9hQL554O+
X1L8ugRSpPrPJnhV1ejps0zXQTpxjmcAuKhenhT/Rc2AFDU6WRuWYNRq5T+USu0n
3Ax8VUTE/L2q6d122HuHTS5p6Z+nYpUP7xT6+3Aqr39eZsLm/LWKNil325iio9BW
gknGoOOGB/aWSDtlCB3he0j3parKTeZfl11Z5vxsFZw/ngmEChlTbmnVhVvLjKuq
aOikCeDuDCibDLuazmNOIcLcc1sEe0Lh84C7YUAlTXyvnrBVR4G4ae9af182xOgT
lHGIgP7KpUpbAN79r5JkhkyWag/lM9d3BNwLLZsgET9LN5lZHzjpoBo8rODyP6tV
bVJkgdVD5Apha7MQfRiK4+tV1IB1UH4vrEm+ZVEoUUf9dKFs5oQwjyxWQq6/3PGc
6Lt1isTYNFgxLaxy3nFsJa38kVrnJVera5tX1CEjWFI8JdIZJqK0f3ezc7XMA3sR
ZFO+XhsHuvDKQoxZywn7jR/9HfWyYNU7R1F7Kg8udaau5UTlK3Sn+SJ3g+h/Q1FM
gEnZQzaA5rCttEHzuhLajvta9FdJGGkOb0wBN2hQZsLzlv2Fu32LAdlIwBPVcw3s
62A3pyVf2uSnOLNlg5RFSaBiG9yXDCwPXB9zTe3PCe48XAaDYtcGjSuTv7o9y5Sx
7t+ahWb78C1QnPgLxAMN8cYdryGeSBeFbIOYjKf0bt9omus1TN9Rk7UBKDHdqCw0
GDYA1xpIDb58bmqALWiv11PADsVI24vBrHk3WgI12muKRhRr0FWs6i17IUxCVp91
bqg5DodfBvW9yo2a1Pwha7J34Jdgsc3Xt4xgMahRYBPpefH7OMnWs3a4Ems4Nsp4
0CTHRI7BMSt8CALVqRD/M/O95ms+4uLNcbz4tF+2U9LcXiUsstjO8q90ezygKE4E
bcjSYCySaD21gE+4yhJOzNkrMiQqkqds+6M01Gv1TuKh0K6FedJrtB3HZ+2bw24z
/RFkgZVyq8js7MGSEVnr7e3V0XivvLrlPH09uadyPakXiqdrEfFgsICMRAZ4ERfi
DJIUD67VFGgw77NAQOUeWZ+vkir4gJpJQcG3h2BN8xw0XO5J7ppRoJaVjfLZGeyo
WvxibzREemtl1f3AVtn+wLLoRhiHsQZoRc/MHG6vMGNxkE3xfBPig4smf/1Ouidg
Fzj89nEBvFUU+TA3NQ3z8tj+3ZTYoEnS3jh1hGS0z+NU+Y7Cwd9CWVwloUKfZHTE
fRatWWnbKX0pd+CbxpCAc51p9vZ+eM8hpYlODcT2LrVda2xH6cho0v4esE0XM3Hr
RX1JYcDR3Akk9NIWG7k1KnWevHUkM0/YLG6ChGMzOiQZ4eFHC/hNFonoRkfU+4ZT
3zPGImPS+vy1SSMZ9KGClb/ol2W32J8tTlV50tK4xAoEDr9SBzgZM0BCuvcf7n91
YvtXPQ5WaG7gBubVppTb19n0VuSRVHnyspUhZ/S4UR7oqcTF8q24e5j+3Y1ri93E
BSq3MVU93mJ6V+DWuX0Kp8ZivQRBGZi7b82ckpp53O58erM7P6Q9+U2K7AGww07P
LgBHibDu6lVt8HoXX10weJ1/LSArr1S6Trho/0Cmpt/A4Exj6urKpBhtnSAeP0Ll
vnISlcaVtbZviK2ZEoudt7yldh95zuu86krrwJvWcQxuZWijivIJLOcSZvoTKqFH
jpHkgo0MUgSOS8hkpCSbikTc/kIrIcQwOVq7+irmjM8g2DHNg+DYmi5QezcieLGT
wsN3d84ZqYlRU/AWLHmNmne3KaQgsR4INcyoBWgP4AUX6rFBs2klDzfHUNTI5xTr
/h86eScsfC/D5EfU+ccaP49V6XVgn5LzOqyWDuQDemfu3tw4IQFLkS9fd/hAfMO6
oLOcqo9IPngUkIL44yWyLilRmRRRd/zczs685lyf8IV2Dts7rKzJhCUSJ3SAdErv
kl/YjlEuNJqmScfBD+3FkxF5jvulaHsqDEHAxJuOMXULZpmtGZEoT8pAd8Jfjz47
UdjbkWAObJb0SXqngL3nDyjyUxgVyFSY2SivZoaK3jE1khmPDDfx/IfZ2I2kfKsB
YqcGOLqvivk8kH+blTQLg4iq0FQdUVHFU5dB/Dn+z5Ykxio0g4AbixybL18JCNWO
YB6TRAZ0FLHGtLItxZE2Aln3wh37rQHMdJH03H0RCk1ojENXoq1KsIRB+dAsFC41
A2OhIO/Po/EAYimg6syKI9pOOvTTKEGAacYMx9UExVeXrFpCMhTuTBwl1rziRYez
G4r75DFQA/t0fNfEe78PUWxezev/HPsh02bdSKS5Pk9Gg0zKabZ7fKKhOW2zLwLG
Vp6sli/tIpw3K+70Qo3jUHrkV+r/QjI1l9NomfC8Ac983im1N1xqzDmYVdrgi4yg
KRzmTFiWyDJhwOltJ7ZLzglyBhpDDpBhmZQ69n0MqFWLHEuSPIGB+jdnm2kAgsXn
MKpR3cLrBsvBHSLOJ3CF+GhrzYBWeBfnm05GXHDrbYK9Wk27hUY9GJwj9diVVNZl
twl4KRdId50zvz6ydOaDWkRh1VWYemIFVVMKPaKt9k19u4EZ1g46JTPDgVGkT5Bg
oANS05Q5wICclBoUkbhbmxnwVwpDG8prBLPxPXyHJ2fd6hoS/+Zkj29uPBGqUTlN
L/qZ/s4fl26XVRfUbVQl3MMh/K9AuHzlKB8+CRmMHiK+I82xNlzX21tH0+32yanz
W3IRYo0QF2Ado4OdFcy8BzRYkavlc51XovftfXaRKvgLCo0h2EHf4f3j9cAikSZO
exYWjW1igFLNhwO2KWZzl89UdoQPgLaGDH2QwuoApZ0cLKgfXFGfAEWHkeFJoPqB
lMK7/N+00qDUEXs1BF1TBzHQy1ovxv0/cExEUo7rvO/1EZCFvbL1sjTzgyKlWTGv
vDr8roldOpUA+utuZVjMkAcKsyXnO56rVLix1BCCVvSxDg3rRCH9Z+XVJvBTiwPi
PS7aYO3SNs5YyATENg5npZL064WJwgQg9SrJOMIAXYEzdIX+v3H//IWQe+qUqk9m
A8B60RXltxLBvM6LKXKNalg3ZQ9upBfFrmpmFHz83u7m8Qj7O/Sp2cdD/XANsHGc
cNyR3pyif1E2uaGiXLgGguCUy9HMrt9P6haBS181sfPKzJjvMRnEUIHE0pC1mmoI
2DDY4vBEj3EzGeq5qzJ9P324q/tMRRa1VmGU7sMNuAqv+itZT/GHh9uor8HD+3Fz
aehvhF9cmvtPMxtm4q/rwAS2sslXro1Q7ebiFMqf44lctfhOaANe44Kj+5eYG02V
G3bybGnHeKBQKzMjSvZvLZ0VRZI63BVcdTQxDNE5hFuCALWDP1mslGdcPitICbcj
H00EIZlYbVIEPpFhhxLKAKvC9YQSMe5h3Vim+jmpr/H4LRgNAgs0O+U7Ud3yMedk
4LnpfyCAHNdQhb6a+d0ZpDLxWHvY1CBzVb2XYwURbeC6zdWyQCS2IREikKxPuev8
1Bv4/5lG2DUHm4cJW7tmZd/zJA6l/Q+4ly8rb6jEk8xE4VErNa3+0e6kPegR3RJz
etw5V8QKS4ObmeCW7aL0nacORHob9bU1KtNnn4t6QjQG5NZ0QotJbHH2lu+vUVTi
YN81zHfIXeEQgbXjJt/JwIkAczXwjaRXjvUl5jpuBjn//ArpA3bY+KqYFhzBEYvp
tkwTfbK/yd8KuCi44rKksGj/fzRsEuHiE9n1OSE120Kd+lGoZyCGySDlsjfSQkK0
1OycT56T/Xfp2UgZ7xgQdYRl3hh4XsAIptuQsG/BUKYZwmen1h1PX8yKI4kK2HVa
DQD3DPZdTG4JpbXAmwFZzQX8XtytBmDRZYSFFr5rm1GLfMdzZXA0wtkCaKzPaiW6
6YkSv1HBSZy4QnGGNXUHC6uKJ9krS2VNsbvy0BNhlJCsHsDO/MWHLRYiKtY+lWVl
R+yVfgiGa3h65mf+4qX84Eik3YYGlkQMpLdMcPS8DxAgBQN7YY1v4fALScUW3PWU
FCyhJHcGsKGVQXvOPL31DYYqfnhRphL2fF6e94mG3AjLDF2TEB6y9kKNe+BnugIt
+TTgTbVx+Tua/3EqicQamPwWVbPFCe6w4jpDRVwTekMPr7NVQ3X9kGj7PYzz/os2
+0XCWFILNsxUTTks5fDKX6BX9Yo/e20dPBLoBVUKXfAKkt1ZSssH0xYvv0DbC1bc
46HA2YDdmGO6ifKIqj4EtrsgOj/ow8AvRqeJOQbVI7X/+JiCdSjYTjn7KGvSMpz/
pi1sAFcfb+Wu2/I0qWpYcuC12bopIMkGz3GKmqZEW/NbTwFHHEAEcMF0l0Y2yvqC
13OBJXUTWIjF1CO1e62drUflPBUb8OyY6nTU8j59439BiKNAEEOGnXAKtyBnFozc
2wIlFSxpZa1AG+FR6oQoRT6CVuWB4B90/zrs4/Y5XZyV8okcCSy+/lTLsDJeVNtQ
7H2NJkiYpi3CfU8P8HoL5B21ltp3GJjgYoFkSFen9uPJ9QXnNR+t9zWKSZ/C17pV
bAio2RD/mCNsuImIKB3MAckhBsdkhstx070on/E6YNWnbJ4DXrXfsVxVzERm+0gq
0vjEaZzN0P0DWiie2CahEZaaB9gM6ainc98lkP6xrEDQCLpr5bLV06hcpDVYAyRn
gaifLdLu8ZQ8aQTLIe3jRRnXP9vanfE3ZVABqlf/ynZ5n7qK8wQSjoQPLt4zjeXy
WNCuiBeJQ0/bpDHaWKDVR7MnPaM1RVoI8LVVG52NACy6pHMoOHMqC5mERrtwk0zA
AK+An33vSlt/rGyaxVEKWLBtEidbNCQUBO8yDAjk7aV2u+NumNf5nUYP1+nHbhMH
JdgBFAerpJcnv/lkzHAnmgc1eZclGcodqkX7WP8iLFv24KtOpes3N+rE9bn6/NfP
c8CWd3Ga4/FIExLt5zUqVBllmXa4zW/HUUT4AFhwvB5lrHlQeO+NvJZv09Af/dEm
Jj4NgOKZZ48AMBWELur7P8GAPMFbMThIGG8kmqxjPc/FAClhP1K8J08z+i9t0Oa3
aiJM08B0IYvoF8aocY2hp+NX4l7di5U3xjzRsfvHFBWFJLHel2k3PcOQgsE213oU
RPw5HfmTMr/1XcENTnCbQm+r4Q2SQPd6MbyGkcA3rcH8ef2elFJ/c4YhGDvKbSWH
R45wWA+UalHrgOgtxADO8eC7BoKAp5jd7BpBoDkZ2JgRzGRhiB1BOQk1QTnR5va5
8KT8w6/Gq2s4BMkw95oTu5khYBEFdcSlQGoDeWodm09cQo0T2KGVHyJJ03WKS+S6
I9iKxzSMIpb/j9/QeyEpWPsokC0i5mJqBDhUcD/S8QaoK3EKVKpsCxmKhFK60va8
+mPxpTzRUGGdRZHdi+yvQaMrNJ5m20n3lvFTrEdUAJfHpHpg8Lneqvz8JqK0s9iy
USx6pn1DZo1m7BLNwGGobsH1hsKgswQIxWh+A6n0yaKOvj7uhcXVo1sK2xLQNFko
d0QXKEVgcXv9aFLkh8FDM8ijb6b7lhORzKTFUcRZo/2PZbJU77jfjVRoVPT0K3+1
wwfcJz+NB2Ul1gAuEfCRgila8woTQ6n2f7vlH4hIiKOlOUDNDkVy/SzL11mGmkCE
yV6Qy5rpMfAyoXpGPGyw4EqSklfibrtxEgDQVsE9e76q+d1QzRbhQoJdVT7tQwz3
cjoeydezav2LUbV+p9KKHg7Xf59YCxK3CQ/UMzqOJkrrqVYrJ6ub7ijV4ry3frk0
lonoTyEDX1WDfY/2q1r7MF4hcEI+HXQIBUWra2bqjGmEKwpeKzI4xS/5oHMgdQqm
pqMYtxl6eKFm+tUbPDDO65eLy9qSrcdl/loY79CybtSlwtvlZc/L5TC2prs8IhKb
/ve4sP40QeS2b0KaRgWTbzOun9m1pFAZ+mFD36p0KXv0o3GXvFxXDTnT8RRY6lKP
cAXGj0yoNOruQPbOA+RFO4v/0BeqVrIqUiFrPWBrcfmTU2SCD59QSprQpKGHNu3t
pTmE/os0NMlrZaPNgnNcvw3gaG8NRs1Y8kNSAclATchKz07TgYYKKaqkzrzOhPkq
8ooZ+/8ACLT66tngbAme5OOte8l6D42HhH59p1IYcQ3hHz1VqE6d3eFobrJehlS1
E89s7qvIymUOqKwMmsPVChbXgcAWXaKBANptopnYldm0avyKOpA/7CqVSph7Kq08
0N7SiiVg4UmBTF+bGbg5Uhdfk61IixgmiUzlQ+XaAoGJm2QQBaV3tLEM+1BbrVj5
lOSvhAOlJdTjljeklD94WpKYZ+Nr//AsFE/Ngw9ur2CWZ8WSIAjdEtvkAvt6wgcl
Q3smLisTURNcAA81sAZ7mc94W50W6SnQVttZUZQCLhFKmcx4jGwgYHTtZDjOLTrX
a8e72sFnUJkjtmnIk5SEem6/hJuXtbF0ULuJXDIOGIIUQG6NZTPnzSN05aONPPVh
PnDfuG+Bh2K3SW6rpF/OPOi6D/sLTsPSqdCaFUBSzdEXx38oMxMT8D306nN+WFg7
0vwMvdAr3LRrzpUqy2OGYcPj1ykXnmcJFvRRHs6KYhnEcgCD963Le959JIn1bKgR
+zTmMaTl3DxOteNblYocrdF+vnNyxwqOy7laJ7fimE35OT013KYA/46s09xPLqKp
GnK4xZYw8Gu/e1GbZiZ+tUfXVR4Go2JLD0hUClLdG4FSvvViF5TMbmJIysBTlP4D
3N8V8AX5+AEB3GodEMhNeZxoVxz+qRmyLeS5lmf7H3F+j6sEotCOp1u4hhrQmE1l
KXgexsZak+rkxk9NPM8OcSwfAyypaPSRNF6crIz2LuW31sPhMcmiYxm50Vlwo91Q
+UqQXL18FyB9gUWsr2ueti4qLZxfVgCxiTfhhplvLRInd5VnAB9AMyoPjUo34Phe
jhgB7ktI5wYl7/eVqW3aI7xTzDPZjVECkWo189MqzY8WXssL0zXuKsj0EMX2avDJ
11LCAn3mYFz2Rz5xdXhzmJxjE4zr2ajTHObr9GrksZxuLjkaex80+N5obvJkqH/T
cjoRyp3W48sXbtocyPE1lJh00sfKK/gZocaGZElJ01t1oFs9fEzrRLkbzg/RD+9r
lR81By+Au/ztlWT64MDOqtLXz5dzHB0yaq3JB4CuNTabrk8nNh/ISTgiiGieG3Ie
YHWrODCUX/otEfY7TPgD5ApT9J0kgurrbSfZbGHPZu5zVbQOx1Cw3wdzXlt9Obb+
H/20gND62AeNO9uc0lPUjUU+BSUsvVFiM9sYlfo/jqq5Jx6y+QCsSdEzDTu1Ajbt
rI6Xbd6HQSZw1Eq/qdrv5ecOY8OK/jjLrbcnT2yXbw/wdko7nLmbVv1qvvAst/6l
hYY1wlWGu14waSnTi5AGG0qdkTs46DYKHHeBa9ca+xa3JuE8TWG9niLTjG1YolZJ
gd+jVnhWyqsYyAPuF6ehDBaSte8vcJuY/3NtlmtWbmo+vEUkb8EndW0N1pL6NTSb
yrg43sNmtrpCWeIpeYQQuw38KxncEfrs/2MJBrpztWlnI4CFe967D7O06Xyl+SCB
zSFcdpfX5GVRaWNAOX9xfLfTokOPRt/7hy2nEAdQeqXfydqQKkV55mRqz7ZvA3JH
rklf+UzPaOMagJ2lQ5yoe7gosQkxCgtYVJ4VhLcJ68iKi1LQWAQAaI3xQc/VnwRc
JnNk7c3wDWOS0u/EaBZHzqgeImtmZD4kh9GfRg7SEzQcIKlCV7cAkS1CewsHK7LY
4ghW6UaGWkBkHBqfcbHSwdhXCealmb270oHWBlbBMgLJQfXgL54xAT+px+axbDgN
4FISUTezqOBMXc/uuyhFnUmdtxb7vrG21dlzjTjQr52KJq4VGt0V/Q9bDfEtEJeH
2oDKJPaBZ8wBCVZRFLuZhQvnCuY6n+RfQ/rU8UHoWhKFjR2NNN7XeYJPHfGflSFY
NM2/lbZ7RYW0Ce+qJsYwVKh2ZrL8n1tBID2MjdWSwGS2TUgBelkO6gbSraZl5wEH
lIPySI9Rr/S5Yjze56TkEA36Jycn/y4K5vqqU6wrgzFG0MQALJmoWL4hdW554Alh
DuAa7n1wiYEwy7Vyveh6zhwq04rujyy/crPv9A7ltZBmt0QIo3e6924CgxYcaWqb
8t4sWvWd2YSmy1ijmU1uJJ7X8Q/ORvnnBMamHht2iZL4i/+TKy3pTDmf3ziiS8c/
1gmVPM/ZulcRI2RFFFtFt4sIRzE3igZ18hUFU9gMn80qioah9dlADxH2ToqOeYYQ
hSiXuXchF8tdLaeEhypE13rCx8Xpf3gqyDVOhOhdhupkRJAgSY/lLaCR4hoZUHWc
mSKkCnK8y4G/2650RSqFFuIZb2PLAAl0v/c07nqlTUX7v0MxZiVQyWa055JDLDjI
UUsCF63zlZVz5EH00Q91pxJN0yYFqx3e8IjhDe+tMOKaQV/w2FWiy9DJhyxNg5d/
ndebv7LKlWMU6ftFhtdikXGQvWlsOr2j9s+5Wuvb9aIGEkB6qu08U29or3jSs3Km
fP5nGHrWZStKPRVguxEqvkvoo2BTGIQLsb9AXmzS/NOmuC0+cwx+56SZbZeXmpsT
oIrXCct6afdQUxI3muYfn2fvTY9IROd4mYhR47svO2YxCjN295Km48Vhwplqs6bh
xxtvM8luNIlHZO8573Lvg61+NA5jIGLc0MvZeIoB5fUuSJZdq+cY6CI2q9od4nDK
vs+fRyE09aEweiSVJbx2jLryydkQQdGDNJnACkGTtRtVOiaQ0FJl/x3/n6gFKiql
i9HukXf6QsC+KcxFUOEUZ7+rb1AvXETAqiSZc4skCP6GRlRuP4md8XSsqLGx97N9
HSmbjS4d9lX1oXBfP5Oqv/YOP05HqBfn940VoTihgj5449CG/Qx7R3W4+wj8UJoh
AGanE5VVxU3yeY3MtsAXVedrjBiwF/+dshuEOSkZwALTfE6c5M81EieQQ10jC/w/
oFDg1hW/xbEvThbIpZobp5a1wugxF/K4krdVZEtXB6KgS7cWBRydIRH43/lbnI9R
jD/LLvxxwqr3JFYL8NCiuwiecVasfOSHltuBRrfMo/e4Dk/s2zYRY+pbdg+t5l5L
RrnMFiLyH9h6qk0o6HZWxLJ3HW3vfeAm07Y0WBaOR0xTz+nDeL+adIzoDBLPov4m
sRJCxxR16/sDobdmD3MZkMcx0TWv1/0+SBPKP1Qimf1xn4KXnj3ckWbvGhbCUXEz
pp/wqwPuaQUBiDfJoHzq1AsW+8vqtowLWJTzGj1hb6w3zrpNbNwpOKYTgPgLttAn
PF1VsVTgHanTxb1wTj4PoU97eRqrpSMb5sRj1odkO9xmBLx4BnAfaoO7nmyaxbs7
rAh6XtCpYh8RLdSqnZx8DZmn942VEZYPNJ1D/G3vAE+rR/sTsMKemNKwMnii/BwD
46/vviMbdybN5Q+ilQ4Xpq4Q5rK8Ujh1tis+BpojCv/LEAJ37z+2Ns4vm5x1WhIn
qpKXEGUwM9Hp3hG+0pEGBY1o8rRIMqYZpUuKNoDxt7tcIaa+6iRHD7HzD+ZFwC20
dEZmqJtVW3XI8RdgYNLxokBxe5O+17B5ZBUSfjbMfuNbeofF3W5XsAATu7CHD/Jh
6/wtfRfwDrABNhmsyFXV5DfYfALsP3yaPwgmo0TM1It6QC6h4O+aJYWuykd3bYam
2gYTrZUYK7QeUZ1eV6iEgeQjAUfGhy14d0eTrm7RvnXkUJJIyg2jsFyKpJKoNnMh
xJFvDwXLamY4nJxlX5TrdnVXiLkxqccyLN7rZ1qsC5Gdul13Mc+hb9wFCriWyuWa
0CYNypWkYpVzxEkU22tjVzEszgoQ/YcvI8EPRSMIVvDAWteylCQqtlBajpVpwt4c
EqylynJSGHfSCNJxM77vNGTGgwY1Wc/UF4BePN43Q8m44lWyDZbORrpWR+NZsJmN
zP9asBCU3K5N70chejwcAo9xG8AUvyQivuNTRGSy1GF0D2u8g35E8hVCuXBOigbH
JN3c+R4/ON9yXHq8MICCspFGYgoU9bZMa2Zomk/4TO8Z5QGOISErmAqzcO5bjvtz
J+jtvoQqBgpOQE+6Hc4OoNIH5A5sIJw5fymo/0bmL2rY33dEJ5LTXuC93QZGB9/G
2bjWdK1TIQPLBId0ZEgDDshK+dkYHhnE815diDnX4dhNKHwgxV2MJJmJy4ut6q5q
mmkvowtkm+YrIahyia99gFsoyVJy/WUQC5qZ1RYZbj+WU80KDNxFwOrNZbtIvIHf
vfivqRSj/UawYzEq4OjfH7CQom0wRdeiWQxcOmsUpaOPQgUP1D/pVbwubHsq/zpC
cB28QVvSdh4HNmRTZGapm/1DqH/YG1OS9AH+9p8Lx2mjCtucwHXyK76htR2w973j
JoQlYsrwWsJAzZFG0ekxmgCUucMc3GyvrvjY9QMCpO31frgPCyIDnkbDPg1S5W8R
JUiEMKHQ9bssT1bhO5q+hmRkaITtCdJl3PkGFzSU07/KxuRQSGz6QUnqNihEnk4b
0szdFY5RKAAfEdseYCAoFDTjKUmm7JtuttM1R4vQ/pLLtEzd/IFoQOeH2KayMiBw
0M3xaGZlcW+CkESCMehZ+Otp8d/FacfO+FKRRz25mUSpeGdZMABLEcR3Xjc15vvn
f18/ex63nA6Ktm79wCjKbRXt/espEF5dGckvD9auoZ0iQi3epSKwjfaJWJv0Pydk
nwuS4Do4BGzI/EIJlbUa0N1PCCz1rMPbZYUCfgIv3gElklbvn912lsJjXFrdUWdW
ZJaXbZV30Z01cHJn7grMAnBQC5pU8BoMHJxsLguvNBc+9BoZ2byohmyO0DsilYF2
GphzbukZ3w1HvybIZOWUMTcC8d4cBVwSxLpG5X3fQghaB/XA9aUfvcmQd8O2Hxt0
MBQTcNu9plQxHg3NpvX72xoRgI4mpfTqk9jdP990ORXiYJS8NoCivBLErbHGuuMi
IkYLTreQhiH8REctCV6M5+lP8ji9cWpjNAc3eKN86QDcQesYm3HzD5AVEi2x9zyL
tPY+wQO5INk4BIR2w87U39lhxGwC22H6BH4pPKP+mVHjPR/aT8cOTuXzQW5mJA3o
6NfxA17vXadtycamZcwsTu34SNeId91Hn7jsTatyYqHwtO8qpC4HfebDB5nJSf3k
XKZsGRnUB2tN9wuWg0bpyn4x9/I9y8k1YHii3sInK0zc7PXo4LeGUqUmQ+d/k4My
vpqeNGRcbWPicpo1P3U9ki+dNtQ+9G/EleaYTRaB/Z4g19eKkTCKWjr9Zjljf0K3
5jR9L7ZUNW+0cx1uQWWF16QnMrKwxSsN+s4AGCD0BlwcnoBjUD1/+EYuyxD+bPtD
L60KsdFktK4e1Q4tqb5MQMxfqpKqI6tIvaiLXsR7116jlXjzdBg3X6X2tHFO8CgZ
N7ZHUv6CE7Hbyyi4ILerrq3N3HPxbwjiRSHbZWD5TTFMfJ32nvbTP0b2jW0Urpsv
WWoOebofXyH0ORJJRkPhXyJBlyFVw4Hn0Z+UmJEN24JM/7JCzJ19E6jiR9vRv6JD
0jGFDRqeOpN3MBLxahOpNEc/xTzJsH9MiqngqdXSoWCheoQK2Zxfy9Kk3sjxN2Yo
yEBwl9L2F1PYtlnXggiSfPeXuyaykiMw0cDSRwDaaeJ9vbiwigNHAJ/hWWrMJSfp
1ioUaTbQCgn0SoGPNMUfK33YD6GSLh4weNbZJ0/8J5OGivr3y973Tenkt3ZCT5kW
cG3f4hRm8XU6iklfne/zENYnj18iXIEL4OoWXY9bRfAcLPsv/mxUQUthZGHNG8c9
j4QmYYCuAUKOaNc8FYPOoWnyEU54AUxgMIp8/xXSh6Q9MTep+TfNCytGTQK/Ap+P
zsqM6i6O4HuM7LH7JdTFbpTk0c3DjNfjlv1fBhoCLiNJoFxjlDJOgBdmLtpS8Pll
uzyglMTfmOgXz0x2qri3Utocxle4b2oUsYp5SxCYvxb6VVzN1o2ggmGZ83LQmtjM
izH0nGgHCCPgmLQcDjgR5RfNmB5JRgU0PCw1J7lp0mWjNlcrLzrphA0SCpKDtBvj
Iq5+W5YR/deJ2JWq2mAPKl6FUOkhUpXskXtmZySYhXESVSCwHkj6K71+adiNAT8k
nub8AgsWWAURshI/1uZw0nm5W1dTt/q1d9g9gpx2W+PJ189QdfEq2J6LhXtJ/qMe
nV2e6lz9de36nTBkNYQLXgbdNS+rqZB/rE9/JQcNfIMazbzPQTYoAFaJTNCj5KHy
851veIfEOItNouL6jlUh9H6Cum2tqBEd34HsbWl7mfPF5aul4Wo+r9Br06nNC71k
BDmOIQjEX6eWaXJ0l2UKcZxLi3Ok9ClaGZnzK9rqHMJvftZQweGVvnHUt+dg55uB
V2MLbxQCVPSXIsLIbu4Nly7olitSweuwXuci4NryKNubm3tYxPUK7M1NU3MzPhnG
T3nUirLcn2F4a1/Ee65ILtS/HMPvjzeg8hpH6ZiyGbNhQAVdCWDB+Y06HEt63a2G
MbB+iZ9v6yGojhsKplnNi2kDMp5upVJ2xNHkeKMu5iePMjoiHVUwkJczyWHb/SDK
xolH3U12g4wND57MG1zT0JpLG/cqHuWV+BslPDBVChm66STadnFLRe3ImG4BOT7X
xF8WZ+iIihm8Ghb6jTIMF8sz9Qnklpe5PMoHymJq4KR30KcxEyX+pVdpV1i7QGC8
CUlM48sp0cw4FaO44VKVmnWWOOhK3BR/j6IG9/cb0ZZ6QW0jh+cZ8zl6lr8/w5HQ
+QG1Ms1FVlj7QQSYhqtWSuuST4fAFHPwwz/qgVSl5eV6erkk9kfXNXSwTN8w1eii
gla7irQsqLXgADBo9UmrD1PnG1udPSeJi4VF9n108wycxKAl+6Rq8SmLpyEPBrqE
sr0BQxIS2vdiDSIrMZea3T5t5u60m+DVaZOdvUJ/Fxz6FiOQxzCmxOqRAMot6qeV
cqQRtLLvFe88+mLDyMUd/v/nCYCr/cGq5YbtUZF/z6Lqp2AJlRUWLAC0FyE++P0k
mYIaefI5aw/C87osx/LJLtj+B2g1l4N7EUXbm+bci0jy5d/Ax5FWWurYlM+GvgiX
0rd/87u1XNcu7GRHlvEIdrLSNjRuQSYTRah3HFdUFDMHk7Er5eYpBQcev5pmPP42
fqidgpAC3hZKfUEZjEf4RaRVIV/ZlEu4UdmX/TRGdD8VXPiSdFAm2nJwtRdg39Ih
Qs96obySo8ZmfE7dlvq3a7A0VGtuF55VkS2f3L7pH47CfJTJGjUDPVpRqlHLeBxV
R91Bi/q3nvRVnmMJO8xA15iYkuL7QjFtvkbaGQ6cZdyq1T7vsxQIbpo2/nBuTk+s
GECWoeFrcPVnNo3xLOzz8lnIacTZOGaHtX4FYq54BDzptqnhDVHmms8zM+mVNhQX
puW15WhhB/qrjX91CGBZake6Lfn27LP44oxge4Q0HoYm1NtVFavKdxksf0wDZtnN
hd+dn3qxWxsFBz3dh6px5gPyWI0MRq0AIhbWSFl/54nqlm7NKpwKn2PJIivu0G+o
YVkSGKQY+akOi/rTyRvfluCfyjuutXDvsNuuAVbb9zNxQBp62cOM4hz/y2UJ0Fop
vMN5NfexDyvRvogZOqeEJ64s6Vr+ej0kuW8lL/xUjR6Xoh58ohOs8D17F4EnInXI
tFeT8cWJ4n1GrA4yVlv1aTlr7dRbu98vqKZloBo4TSyQvqeiI4JorrVQZUeufnEp
GQ23t+Y3pTzILcUSk4yIOWssUwLupAs3p+bHpfV2K+xGKwvQpICAaav6xYhqN33f
sQWkYS2wZU/GonCPccFVhFBEg55VsvVOegLuGRC/zf4YXs2MPEYgoW8fjWmckcdk
6dnN4UFdV3D8OyKavGga2+kDz53XK6DP8oEXkIpV/8T34t2h4nAoR+eKJwRJqkRn
EpMOiqgV2XRgxyx3LScFD4fHjthnnPqvE5+PodiMu+QOKTdkGRXHTiWn++dlU9qm
olY3mBd4zbwOns4A0noFaT0GX60YgXRg7Sa3GZPzLAp4ROAgNa7kmCCJqV3gxV4D
z5NZADXm+m1KnF5VruhWwlhSwmi9CPLujq4PP+4Atqeql5HFiQz7MOZTdaHZ2jzr
Ji1nWT6kDPZJpFsTX8eNNOVjHxHemRUfISDVXYUeSAuotRIOSgUpQvcFEL+92ZjU
rsXvhDDo1ATsoi9j6zXSGBqKpcQQjmSktcRsZZXi5e9xjgk5uY8Q7U3Quc4trqjP
aDA+zAaUChUhpj8lTUIDEM7fAW1GO2mF2I2m8J0ztu84G5QMOozBUZKrQJW41cNT
A0UKohrNorkxBib6r1AW7Ji+uugYFEPuWkTXnWXeHvACqxX/wGGoEgcXr8By+ruZ
0I+ik7bptQhfL/rtPIXZTD3FJDtI5HR4d0jcmB8P7GDPGL/ttdwBYwJQBAtrSuFd
Ufv94W0Lpb9a8CCc2G9H/pZ34m5XcBUURWV5QqKVHbVp/wBCKQGXU+1ZlTIbu7/F
inl5xLEXGbvQq1dpyeo/cnEldcLh1BlbqqouKL1JJTRR2FOe9AjqyabGiRe9XXjN
15pnenU05PA8SRIepEa9v+DjPg994UsVyB85DGFmTnWm3cBHdAORnP16F9pxlbKC
eByQ4TQOp9Jg90h6qxmtmSVvTVw9ZtRr9TK7Sd+jKhLSLcuCmnaXhD8RKYnwRDj6
x9lX0uxcMNT2UkMR888QAJBrgWHraBpH+FIUcpJGHNfjHdQk0fsecCpXIB8TZoM1
ek8fO39Gx4lBfMLxzJcvHd/bTGYAIUWmmDl9yvYrwnI5L9EumfqR7xQOJEdLTnQ5
2gLF21cX0BHEk5KLlMmVHmyE7m0Pgg7s2ODRbN43Rwvh+xhjpxODBtGCa1vfu3mg
OGQwh1hExPau6Nw1HzDt1u11kRVRMbgLaH7LcJOW3SiaOLHKayxGONccRDjaUT9b
PWfDPbRuuGr6WGJ+snRfNYVBTGxrIAtpYPJi6/fbMMiVSJd+6RC5LMBO2gYHUvpR
l2GSC8iq2MlkbmEEAR24bgLZylUxrfqfRmfIhqOAcS//hghHwtakaW0Gj4kQLAPL
debkBFbUD/17tplSPEEmDzKBXlk8P5lJ2OgB+2G7o8sdzs8Nschio1gSmdz8lSah
E1GcDHgeZm4e8hX9ycoPOKwJQUegB4RK1/Qm0AJijibGblEc9YUHEcSr3RjbMReH
ceyrwnSMKqC8TNskr3LMSdM36DOveDrchoq3uOPBDAk/zXEq5pS7yzHuoJmWI0pr
dT9/5OUsieoAGwZ6WX5bGHE+HM0KUBV/LvM6VjZ5kevp6OE6xrS2IBHbPTC277VX
Kw04TIenOxS9XusN8WVkp2TeQ+p5Ot9OJJ2YNKW5XMz99LW1//uFuSDK7lOOJ6hi
cchtAL1X4wiKm8TnEPY7WS8zVHmCT0bvMVkndMP9X3/BzLVM/pj2MTsnw83gShEg
fvprQkBsHcmwwLTkIAtfIwLOiWME+Cnouh1XLbRexrX1MT5C2pNfpFQHatrqpT0Z
guno+WPMkFurqsyYGBplesmYxhepODRF94TG5pLd13rJPZ5PNPuEura69lPAHciD
Lhh9DDt2OEwR9YRubPDMU9Y82YKM/NVkF+d1EEusXVJv14J5LOuVhZtofu9KwwQi
lIxcLl3pGSDXXAJI6XxtkeB34UPNyTP9MubLBVutLq5rwc9OsxoGVvp2Co1d9QZv
Of+waFuNbHeMB0rllPumwF1Ppdmx7Vxu0dRGCtjgu2Mwx+ZbFasMCPTcQsXe8hUz
NaTefxpiRtu6BbIxqDAfeTAG0jGFKdNCFjXYL/9ZoJ4sehTKY3ZF1Qnyi+WTHo/G
UCRfaRJmMVuvLZDKk2vMhny54VOzjxyClPCUzDSVo3FzDA3b3kJpM4yrginPLIL/
52M8ELF4EJzEdJb6cvfk98DcQQYK72kKtP3u4c3xTHuKgoBAJLC3xDPXZe3MhZGR
gMDes6eWzhwsKl/A5qiuoDAOBZS/hMLNwzMj3zYF77mkOIezTLoK0W1FRvME2WXO
o0cEN4fBCZKY6RM4wVB+ByGZc3yYs5UQlnBUKJs+KgJKLE8+WNwD8ZriDuGgZj65
PJxeTsuuwbWcJd1Y7C8BznCyxVFFhjgXBXNeWfyoSWWP3FFGqJLzhSQb8NsAVNqY
GhOacaz0am6yPF/V5A6/CAq5CQBb+6S6GCDNFT3D3leqURAZBBwam5FDKBYSXkwq
EWMZKvMxL6/tibbiHdRI+g+AzWrhXsUjaSbK4Yi+Dlg4KWfVryHgGVP1F0Sx/bIq
AOE+PMJM1m/gIdqSSvgaN/D7KaCI07S2pDLOTRkekza3n6nR8wv7qvYHc5wJxbnE
Cvkm5A6EOBVOZz+TOlYjK++kj3iQGdkOoHvHXuXH/6R3i/s4qgwpvJwb0tWTpWeL
lmgiEJDwvdH3/r14BnC0/EIiKozJAw+2rlYqUF1TSrpG2rVjWRZNGkPNEa9rCM37
7acZ2uAyBSfD9PEU4qifLnwGUtr1Hij43XjDBqTAxzeujrNTNPKs5ZLiBWy7EKkv
qaJjXD1LEFu83XgvwBdvrjAG9+t7JhuHSy6B+BGSZKc44Hc2pDiPYwEYoRm1SE8j
Zk3UCiXIt0ub3FRCaE/ozXxNjA7DhVw1xN9OZJvwp+0Tl5q2oMgOIqa0am3rLNRW
wYuDPBeUfGzV5Gzy3y1OeL2wcAr6moQLsmpvu9MKyKGnE6AAJui7hgaHBHdZygSD
ZobnjuC62KFbLIEil1YPKajffzR+mmoUrIy0shvovyichlMAlUPhXbgggz/8QD1Y
KK3qbuSCu5lL6Uy6us36uUN37KsCMiBmtewhrZqxbPyHMo2rQwv8e9MNjHbCPNPR
n3QT3xDqH1ym5SQIFvU6VzjhqcevB9ca/Pv9VhpaDr6u4a64RVzxEt+BqE/qPnfw
KpKe3wlmaxNIoP587X0h2piiztXgos9CBC/uckNgH3eYkd58OAAm5Sl0Kdbxq4TT
lOJjGOMYBa8nlrVl2VrnrCw87cf1HBwVGuK5Y6pr4Gn/LGyRZ4DwpsvWUIyuA6II
VjtWvXsr2YGsNmotHOm1qD9hdkwN2wVR+pz7lPB0F6R10S/3jCQeuMcuUb5CSboV
wNHP7d+VXHEGtaaB9NxXlR3KOJAQUG+u5Dmn7hNnLQM7JFb0hElGv5/DLPx+0R4G
h5zsqgSMCoa9jHYlm0nVG5ATuCLCv+jGyMerRmwge/o00zaYXR4VjVqtVV0XWcHX
dS5VtYSDHJCKhT87cCs1Vqm2M0sVBNBilGCod8jBzwNDCHAlVlEZdz9a3kmwCTAA
XqCf+ONuUmtsfbMiKT0y/sS2pw7ZQs/s2nejQBkdOSO8l2ehMJjsuc+zIIZdjiQx
mq3pBONToQyeDadt9T/+K6Rqxg0+lbrInbIynnxJaWh7HJRW2n8l06OMDOBT97bB
kHVSqn2NhCRW92Z3iw7cQIFxjNpaPNu7pBm7j00xnMU3o/CUgSj05fvEXwHr1GUj
zeu79UGR6pwsbdhmvApgETVbYNETxKtvd8QnEl0VgTtaD0FVtQcuSp6rIoteFNo9
aGNmwGn31HeoWGgQ6Y8fo/HCSvmCIEpMbIoJFtNLhXZZpb6SQrDbsIE0RYsRngHd
QQCfuZx4uI2w6KQiKjbyfEBI9cRCbKo4wOWamavNJtAaQEcqNCqgNSItDgfqmV4m
sGj9EXYDjJe+QfwkY13ap+4r/bzAEpALcJgqlf8igE3fIq6+V+tRoa1OOZXEHMcP
PRuoBZ3ScCGPCtFyNXXg66MP5k9ivGXaENFVkR3uOWx8UOA4+8h43kBPKkumYGim
ofD2LkIWnGLGK9DyNx+F/QgS6eK29UTm34/wYmSUMIhWd47DF8ETmgG50NATw52J
a3UxO4vKSMoSncTaf/IuAqwDQdoLn4XPipytV0+ydFPyGv4rlGFMPV6ORtn8tksg
pA3Xqod3g/Ztq/DBz+RoGnfQA/WoSVOvaQoByM+R4XibUoMyzWKle8IyVpDW2TD3
uuiCUk07jSaB4lP5ZmVV+zC8JZNr/Y1cBE+WGw/HHqJM+cgXidekxclsELJcQm3Q
moSJYbQPnspykJ3/EWOyfHczjszos7pTCwsp6/W7VBhpl/tW2NYPzWB2YMv0q/Xr
Qe7n3SiG9UYSRn217KLCK+ExObRtlEJ3CHwRsxdB5oJJ20c1tT3TwLxigWhrnbJF
1nB2rtE9UzT9VbEkXbsiVCNX4vS/S9KFx6FM8A1+qOsEwJ0QKoaaQzotQYHVkT8P
iA3S3evnAnfulG8U7t5ZOaYMnCfCWTiF1w8MfiMq0chlHn29Z5REVWve4Tf/ZHd1
k8YJWNzyx5BirmEkVKxRBqZEzSLFMB4wkzB9J+7E3KyonfzWARgB4v1C73KQEom5
wvKLhQPSykn+bUgB0HXluoYrsabkcdiNbk9oxaiw88njnE2mgTpkL9AQeZKqhYhJ
0nVeVYuVmT2Xo3U1RjOFAF6GZtHh6H+njFRFiMvafslXdtLUe0bV6V1OiMd45VQV
oVmi7KcVr72S7eTu/GYwsRLNrLAjPs8bu7Pl0X6VtGWF2UaoM9KvLuW1QCqB5cAU
6A6hl83panMUH62zxArLjs4svAb2z8Ef25oelDDkuCjMxFuy3Tow5/AfsueChdrD
PouPQfJVbkJlfBgObXAxqvWVr6QF8mEh1o8CRk12uutGx9PK5pcuEjqHUnWpKx2h
7nKhxcs3pU+h5NAV3NUaIpoKZzgCUIWGVPevMUKk9bCcSK/d7+q5Um/3jgli1gtZ
/anAzq26fl3Ehy4JIVytoCqvFtKurQwswBtC12wvpoO2wrqfmecRsFiNbWJI/kCi
veZa+eFsucDJjNkJPa1iOmBgYNfcDgtdDF8mn5KxUN0YL2j2RyAlms5FEkxXEGDJ
V+MfTuQy+wIylZxiN2krJPP0EIG/cV7PI+LMrJXZ8UkwqaJhUrCFlA5M+hMjaRi4
3vabf3qTgENmsqdlsqarwCm304Bt5WR1hJ9J/HA5LUlVBvrj1LByIch4ouQ28gEp
NULRSC/NODmN/zQCNv60DBFmBhAS8cFKwj67MoaiLPH+6ms0rVUnNu3FxR6ZgOOx
pDK2mpGKSE2+RxCW6lY8whGvA55rkKPgXKM0HMt+u5We8aDkFdIUPW7PDbRDqACJ
+eBGDixIJkv2AQjFunCJdQvNo53Twr6uKzOaKmTIUq734qwVARyXgVElnTpjamdg
MSK0KjCZGuEWAev/2MFFD8/9jzCraR7X2aaJvPNsET8+3pUbisSoBZS6pd8fypPO
m/PyiL9RCdvAkCXeBgsGnAcfq3r76Eh/zohoT2SSJF/77/6IygHpmWLB2CY7af9V
Z9JfVSlQnmoXQNQNNlrFZWtE3xSJc6OCfhGXX1bt8XHY/GD4TabVeA17u1JMew7M
9MNM+r8xHol0pcHjJOyd0S/4Xs86poBr3nEQoYzqRMomnYIc0n/y2qN2YqcUUOMX
ZX8L5uMoan5VuPRwzN1L9u0c99bGHBR2p75R38AvWdr/D2i12/6wjHay2zIGDChU
mzb9FIZFwsxEfLyzshg9B6H9Behbc6sixm2IY/K2MOsOK8vfJOPbxqb1LzXfRZZf
nfTrjiSbHl1LjdCGDG9C8Kk9rC55WpQ0sSYvmlhArNYkLMRBkiknTlAvChfTGT/A
JkavSkFkkOQsuh9P1hutXyQSuC8DumWTleMfgVnIrDh24JvEleG6/WXfvYtmosle
UklPzts1so0ePDTvoeNBQp/LX7UumVB2bQ7WI6oXw//wZKmaM4E15qEGvTfk1UJB
Al38tIX0rlE1rV3vM52UinlubK0JOGKAuV6zAd70aSHWpLCnDp1X/pjVYEpfThtC
jXVIuhr2LpKLghNC8U/5dLQsyrRTXYq44EwPK7tmnbmJph0tUNOQD/Li4oFN0vUr
LH8ee4701v9hHJQ1iItwsWTcLgN82B7p0ZNMkkZ/VFSYt7mD4uOtnrEJUD+OUuq2
vm1mW8XM2URYJgNSc5dV1Fsf+hJNCxzmj6jBHhGlIgX23MwoYW+9H+F6vc1rViNB
EL1w8nPiroqTo8WTuX/tTDb0RUfnzLW3WVoZsIgnAwdlLilNWqZxrYevVpvwVJbP
mWYAonWXAJBSXyr70I+F3fO4RDjgNBy3iePZYhxmnEtkSASXUOgCN2uuBthVs1ky
SpDmvSQ3JnTbKfk++Zq3U14V8F2wulcqyKjt1/QCxEzBSgH/KHriwhApJWZGt3LY
SBfZIRaeRAg6+ZWuM/xkFMm5WwLmoVNV3OzvVuwrs9xJ8uHq0bW0xqPa6LAVMY8b
B7CQHQf7QWvTPWXu/Vuvv0tZdqCtAyCc4y21bdNje1eG+FUJFEehGeNSb0A+bwLu
bKv1SoGwYlqlLUQc/Zs0tg58NrZnO3hToi9ddsS1ag2mTiUmKdL59WVZmAiDK1oE
o7e2ntjhlCzMPfpPAJVh5UcW5vyv/DXYuz5xsUC1QrgtCFxphCF0hY/tdxowJ2/n
1DjvVG95V5Ixpp6b9y/9w0vlpjauSxJtT/VgcfZ3Q2iWLPGNYmF6EbwINxwctgtl
I0rijjqLbJo+E3m2gyb7f3NaXQsOY+zyE+nn9cTLSmeCwQA/bIX+BcaTbbLK4GNt
o5zEFpUExE7W6FEfz34l211jDM+vIXyBa0M/T7EPIbefnEr+n2aocCgiStG3nPIL
MtbYdQmZCXlx8sdFp65Y7Amqv0QsYkyn1mzIrKhBf61NBBspxiVzdjbrEIWwjUBw
Co/AENAl6BuU36h6hxTveYeESLndeZf8q9Qw7jHLkCuue7z6VfPnibJYKUaQPT9e
PErGcfS3AHiP5svnZOF4iQ4zRFq9mRZpxWr2hHve1ROrsP2hYrg1V848WM64APGA
wOtj5oa5t95pKuZTsjZ1bYTm+5Q3ILTZVvp7OGa+OsIrQMHzaYpk8JxKD4PzQfGi
lLQvuuTpPqJWDtXcQxU4f0jH7sKjuwwVhJuXYoJJigJooWsGoL6cRvlyH3TOKeJS
RCYiT7I7bIgx+t+zNtGCw3kKRHxiWqc+ov48F7e9U2p2pk7Gtl+Xwmhpv+sYF6Rg
rkzuCScNKRvcaBOzq3R4VP2pxLWeCpa2jNokA1vtA9kM4dYXYVvyfTkM6FewnZuq
nJalmMU0o3T43WL088z/zE8GdunVgcdBwz5S8Z9VDVJ0z1lqNVrhgCybrfZS9Y/S
4TDDekzsT801yb6R9HVBHfnhpbur76pwnO+z0SGyt7HAyBfc0uBbEsQ/gWSYPh2j
7Z5oX4APHIIdsLFeSHybzYQGGY0XVS0ljZax7S36nrnKKWjvTBXhcUnNGHzfOw89
Z2Kwp9n4nOTyNbRynmaTerDhq9NSp2R1PoemeinKUZq7DBvyLlJlJu+rxwtGMglI
LVcztkTBLPy7R4MUxlWJd8FsGWQ6kd0yChTlFTBBuBJOA40o1aeqH4cmcoD4T/yP
U9xApTdMhwyCpwa6tFxh2Va3B8ywY+m1ERgVCcSvMi0aTV9A1zH2CU8QuuP6stuk
vhDEh/w2X7g8XPyj/M+DnKyipjK9qEa1x6/6mQin9CM1ZV9coWXNWuLFKZ51FaYF
KqtSYMv7s8cSwsEGg7j+xevVvY26CDZoyD299zKVS7bZpmi5RXqIjoNFT12je27U
6vy7f1pfF+wKGNd2yCxFt5YQe3QdK2/Vv6/l9+7TUlv+/qApUGqsX2xSpGL+n2jO
NQoYitHb7ZaQOrEgEr/Avt6mt6twXkJLFRMj00M78MEGy0HzKXoF9pF1n6cfhgEh
xVXiRKd5WQ4yXhF6Ck4ECm1OZXgUQmpI1CVLEtVDpZmmqpZQ7FDMKCbkEjr1H8af
CY91Z8xRFaHBsN0gPgXMk1ewn5gNOcDm1eVAyB1w2xUl/DROM96uq2CHq2keVerF
auBi6gYfmyIZcRAeBUKDhXFCVt0C1ua+bVjwVaDamgNaNcOMGh2kVxfMbx5Qgh0S
M6rVQ4UgzmkRUJ6X4HEGMKN2jnc9QrTmFGY4Kqo00nD7jlM6B17v3E41rU0I3yBs
JStswqwruz+JGzwLwfME4+fnccO6tQCsMl425dCT5qw+1DmvWckNov9QAGQWcORm
TbOx/+iwGaM8ghuEZq6UVJEnjmpr7rv4y8DRV14xJxJguoZMly/HF2Z5M2/fQ51g
hVWaAewCbZfj7rf3VwwZp2TLxaToM3XIdP7bK0zSz1LzBhuocQ/M4oanfPRPWjRB
m6Ti7NVeGJSUFtYIIoneeYaNYV4Dz9eEoWNsWU4ks7wvrs5CbaRS6AxbDVyWrGFM
sKrCJAluiEuzwgxe4kvB3LqVJQs9IaZXU52pZjLMvNlifiqI2MuvXfBhEsOdJmhx
feMKYfd5KhWmx7Sc42aJcUJiayDURR+FCoeLOMcseNDcBfrA915CnZFf6yBe+y9a
3DVyQcrXw4A8bkg9HpXrbd3956TIOvmQpAkn4OiuqQMWItse5PlZNAl/ubsUIAL2
6KtEK+TaGZKBsp60uEC6pTMb21Yikk0NJzE/exmahnJNNPF5gxEV7LoWMFAC7xrd
I/bSz9w4W/cTQuLlZHlaFDtbW/gVvJMFq+a8XS3hFYf4DS8sY25ryMKjTCjShQj6
DkmJjzyufIoefJM9pmiYxZJwkZfsKKn9XDQp2hOACNE+0KBkuBz3Y5bsDMt/2TS/
1GM/CWADCp5x4h4hns16owCRLtoZI0KyjLn1akSKCPkM4PUQr2yIOXzVX1l9gRm5
IhCD8IbQ2/E5yh5j0rYKN+P2iKZhkuOPIzqO22riTLKX/f66YUIRXD3UP+6tuBG4
761atjvqZ9WWUrCuWOs6xJFufVPwku6tulEszSEjGYqfDaSnHba+BAnzFzC8yrKB
0Q++TbBmW+WkSdGNYqM2+HNz9C67Pcolol9yFFy0CZj5PamPKgXTereZpFMJ9t+N
73DcAQ5o+Eiqfp0VCMUFOqDKITTAQ+LuQuFSzUrzf+6eUZlVLIT65xBcA5Sic6Cz
FWT5GVyT1V+ZSTEQ2uWDHwre8VgBRaCV1aoEYg/mP1AbxIPTxhEStpjUyfw79CDt
SCRg4a/4i+WW4FNL2/DnwFKp561R0MbJGZn3AMFl2Ei4kVocltWxUKTyD/iDfNA6
PTyBgpc6MjtDnZf+fG+7kjLdd2M7mbkPnNQ4mVlDoo6xQVsfpQZpZskL6SxIDEfH
/wJRCftHsD7mPDCVLXA2vQSJKxv3+tE08HExgTYzwkDIweqx+X92bXxXKJyKOWBr
VfiyWvYSIS2PUzBiKkzUZdQe86/9O2G5rmHRg6V+DNQlq8E8rNPdnx3pcmPxiwWE
imJXkv5jyCgbk+4TVP4rGnlXZ6PXF/AXOTm/3eu0zgCaBfS1ehD4HlycbDVTnXd5
tscdT5AwHnmzvMlJKzXzE0nwMJoxr6Jbo4+0xoy7QruQNBt5Nrs3tvQIFNiiVCsY
IWmU7aRDm2VAmGhL1Rnv5llWAXv1Fiv+7ZSq338XBbtiADRk38RI9QB5DylNOyf0
JzQLm29LBi81ToSXXCivzQy49zjKlM5vQ2J+LfSCU/76kNXQfJvqu5W9T9qtEIeG
EZzo5Sieb86n8uQ3sXm4SzT9RhGWpC3VM7ufbCU9HFxITB+WlgK9zBORjBWva7yA
Vd3UyNQ2F2/6MVJq8rN0IBy3xZsapitWYY+HKziB41+uC2uyXpipsgAoj0+HRkVu
xij3sKhJvW87DJxG79UklNh2kGlv31DUyaqSLAaUejpkGU58wMw0n7H3rvMdh4+x
tbS0TdadO0FwYp7HyEVc8X7+/awHH5+R3KAY45+9rx73F77tWVJhWzhOxXdZBgnt
3OZI8EeduDgLcCUqVlpRG8Lx8eSUEdjNZEJAuKXw+0A3XqtWfZ655cx5q4by7sdP
OwX+B7RjvJlsm59ppem0GHPbe30EsmpDFM5LhIBYX78vOMVL4X1Wbj4P/6VUpOpS
gPb67PzFBiJGfAWjKJSC5Mexy5GqMFOGlpboqM8SiQFbCwXnXUwTjmitLTp6a1S5
sLs4oO8c9FyIRGuZ63xbb7nxlrsnAscY0Lwp6i7ERdmxkjC9yGxJxlp9ken8TYaR
SUbV5EhqqVdqXGDL3KsCCuqau/oJhoA1AE8yrnHrU4dpKfRx/uRpAr/q7aRpLuQl
e57EBgNpMfdPMPWwO/sLhamDE6fT3SwX76e8ynb/6O9V6BjNI/EwU07Jc3X5UmR9
Mf4faxwi+WY/c5M0DicKxpNO2Cpxe+/FY6cpuGcAmcn+G0w6Uoqa5o9WpqxPXUyV
iXMWZIgLljCZPMliZtWPbknDWtOg8ckNjRwlTRn24WuPRlFrLBG3LuMpTq/rvKkY
KQRNTFT0wAVDAl8mMhRn2fPNdUehl3dnZSE5CZ64N9qBe+SrWo3ZgWNDWv8k1weR
EdYc8nO5Rk8qxQNdzEw6+ToVAamEOTX/aqOawj25idQ++5l/Wz65LUH0aNKwhZaQ
Q/1UNn6ABXQOJCdNDxdO3+DSCnzBrul+xmj0qzgRNAmA+Bxp0npzVWZuqAeVmQ5w
fHpA3TVRmsgY6NmoyYttHrDxlOnTjo1YFfUH89NM/GEGspLoEwNuYUrbZYUgZfy/
dFqdtsJPJi0RVh0p6cCAniBjLXkaLUUkg/0Ezpliv4xR/OmLqr++CSy0DNmxUNsE
tbMSR4CmcKH5neWmLfI2OLA5IjkefNLjxEYbdcjaYR0L7BmA0UUSxkOAyBpLh+/v
Q94mr/AoYWgao/llRAkDha8KhQ1SK1XrlRDloHlZIjfXRqltnzIDt6DjjDX2QGOz
Ld+2QKd/9kxTFdmmyKxqB81DWRVw3PnxA7jhO1WTWuNvS5m6lHfcGgRUf5vjVzQ8
sy5C8BDReG17pZbQ2ElUh4c+JbNGJEEQKB/l/xgiUtwEaTRQf+zHemLBTWEbiKEt
nsF6zhQLojNZeQ7gRRS1ZkfkPsPk8r8BvRpyT4Mrs5qvO68cR+MbrBXehCpper34
Yhgsffx6rYsHaqq2REnp0HzttSmb8t2yJHXnZslVjfbzRaerCiV5inVhq3kjQFny
VgoZHVo1Y6tS8RPbLm8oa3oNwh5+FnVnmEVJXB+dLRsBcmpMY/IragvhfqAnfdAa
tKM+6g8xwlH9hFd+hsGL3unfPZSZ6+aLIYDOPgexRo4sCxG2LPK08BjJCkN+ghfp
83dZbo8hG3J/2xibCIz4agSJveFfVhJzULTEnZnwjin6zaJFLCdpjwnN4iL+ku83
bVil+qLfgnqAxaxfdY3Tbs3tdl86xUrI50ijtyfALAG/gcBMHCrHqqUjcIusiRan
80PH7pOp/tD+GtCEJTLonfai2FykRnE0wx9B2EiJKTgYpCd9pudX+RAQmoqqnNjv
p28g4G2cgfjt67wE8gjCu+CXcdwQjnXDdEnzwKEHa9LdEdauzXs6cEZeBkQHQio2
SFghd4dArTV3H2ofQgyFnQvTmG2ONCHoimVfM4Ji4nptB3gccGLuft6CTxxqNerK
X2ZHJYyPD5gRSWfogDxtMHReG0r7/rbNGTDxbOZeDZwuDcoMBZM3IXyWO5DnndeC
i45qBCxt3Si+F6THB3bl3sm09rAXs2zkLAYFmOkUAwmE22fYXT6YFegueLHphGJd
DaZVf3f6LyZAqDuaIQbBDOd8qLkpXqy+CqTDimpFxU6EPAWTL6M4FMILWmMR7nmK
lVxzVkp/GjhAAaNkpSE2dnnLJE9SankKh5NHd3IqMIrLl3qvlE90ikNi61Vs+rfr
2PBIZ7VoPIUDeivaapZoC7VxC9hEhgR9GD8tO8w12IRafjfhiuVk1uQfzQg1kD9E
cQFrn6aJKCZtz9y9OZQZAnvcOFGRQHOMCPcly2Y+BkFmLCAlgN8Mjr86IjC8hNyK
+Z7WRl4jxbuQxlvRLvw/fAlfPxYhxU3y0HGT8fcU7bzwopoaRgXibX8peAYdOpo6
a/cgkNCaPODDrHuDsIG7E9cDuL8b+bUmK5r9NLPoV5kA8XqPkbx1SfDdFgNfX3wa
M0egyFhRqkaeQFCEa2PKiR0uo1dN5aOpN5r/sZ7jYTCYN3aEQ9xLmMmrJaiOIS/F
8nn03lqBaQM1zCK4X8xSnMMLj3oB+5RxAAFnWlZkIGQL6YGsktTIk6UQspx2rnZ0
KMYPqQmoP2i2HM16RXjHOffeutR+nNRd4UpQW1CRNiBmMF6H/8Tq2eGYeuhahxvS
4m70842wNVfpjTxcQ+rpdge30q/S/2GHUCWWMuWFX00tAawFZ7RIWX0OUAgOmr3Z
YBnJplCndo3A3tnRM/SGB9rDgKiq9a0mE6HzYHPA8bKM+sAvfmWr36OW0xGY74Ki
XiqHspcMMJtOg7tj1eO0ydfWTy/X6spo+UcOJWxrf3xQnX5ALPUzjMpAeItrwbML
Hp32pdCA7NcExk5TI0G1TMGPAB8EDtyYnYYeWlrCyZjNhKkUZgLlXaux2ZHyTTm8
IRuJK4cAAQ/8Y25YH2axrAlDVDWjYK/pqXuW37XEVW8CnKK0dAws8eVk1Ct/dShL
Wxw74/ffqpEsMXsHZ2Mz0DvG24vpfQR4tOWgZ2TRhmBAqbS7SwrbDdBtxqVMEJQm
Pet/uxXln1pyoWuoTX6LI+pIxIXqbTYwy3po4AMkQSFErU2jn+Rac7nxUzxIXSVS
OxBDgMPOtJ21/2dOBByicSyA3d/JIZ/qUYMbSkWejNLRFVUXzImqqgLke51wsyhm
vuI4C15GwQ7U7AUcB6D6DqIwv/QxW7jCeMjKlWA2fpG/uN7yiqBIDRhcZ6Pu6Lhu
qkVmYi6qycq0dr6ESB2S3mvtUDeKYgvuJ0cnfWEEFR14japRDUREV8yEzIEmi3vq
wl3qQ72HcIKRtLbYBiA0dQRbllKH27oZZRczLQnzSyniOC5HSur3K8LYSnrvCA2D
haFyGXx+eD8DgyvLQxlkQ7F7ip4wiV7w7DfEtTLGhSgM6aUg4X0k7KLK3j7ROEYg
B5oSowKScqUMXKfYS2eO4Hx24yk5Wm2uI5l2/30vUQeeKPoH83R6b5x1alRQ6HWJ
arBInQbJDKW1E2i9bxhxJkIR8PQp+qjq4x/6pDw45fbwmtcEmXBI6AwLDB7RR7rR
2ode489NUXdnNO9zIx/gN0U9qLvECNVJn2OzzlAMpQe1SwoUQ6fZj4cE8/RysyuZ
eduB6l9SCAVMJgkbeo3bQDR7UfvX3eJXwyyOzs19SRVl5BAsAJTy3DH622YTAxPv
g+lgipvh563M6cRXXW8rWLxBObeDn1qv5UbI7X3I9W5x2vJ/+kEoby013M6QIBPh
JWGT7LtloC7Zzd/MmLGdxI837I3lK2INyQ3d01ysA1lneZx6g3oD4hp4cBTVGMQG
uC1TKHIpgzLrVY1Y7kC1lCGamWqCtDejIYUqWCY/Dn/Ea6IQIOUP5edVyxyNuLId
wk2Lcsqrey6foyicOIxG0Tw1QwXIpSUYD3DMrEzbk3SHV5qYXgxbIf1Tx4Ws+WIO
n67wWaV2GmgNpGmPWHsxcRUhqqpYogmLOV/GTu6oIvfTD8Pljt4xekpgcwpMbm/8
VfMvxnxn6rD6p1NKjfBmes+NCz1PVsZTn/7ObnmrbZfHodZk6z/ENfY9pUADc6uY
8J6RfZ6TLaVwQAhwQHjKmnmGjAr2DC/vnVy4Wj2T860RZpJnCTOP8Form6ZQET9A
lr/jUDbF8EW/ArJ2FIFwUO7uDaNIJEUEZezNGo6X039ba5FpnBSBEZ5cLFTWnR77
O+A9hseHwOG5xdNfZDLl9qxl6GbF+TC1HcmBHMUNrX36OzfrBUJQpJQqIRk/oJsx
OpMsOW4CfpcSsdeE6/x0qDpwsfq+lIaiK+jE2hFNBUVwKDLsGsFFgLnrCJm0P/uH
MUmrEe7bVd31mQVx/xNMAyzrbAnz+1YMktoAhrR9tr+sJZGF2hqX/tYoRYqVmf52
FQJEtEeWwEiB1QCEX7bICRGWhtYfgFYU87I1iiCwYpQZ9XtCUVAAP6whB4j0YLbq
0YMLU6IbgDvfVKRfiSNxcJ6vrNS9QMWzgerRG+o4HlgqyxDjjfvt+gazXnu/9mVU
IylqATKNUCZBzTO5JAp+C6O+bWMaFi6UBvg4QDBamCpuHpACYe0ldtY+qfC2ziYx
y2hxT0iYH8BnEzf5CDnHt2Gxbm6LMEqYbEUVVdQsIYSCjnvZ8S26kyzaIGGpcWwP
XBQ7xyLVU1iBv4fOVL6Z6WooPjeE6Q8SRUY7bqd9dSa1sLRNRKawkFj3FQ76+H7z
lsTuokO29dL0i1VH3YMlFZ4V3icPf6A5M2OwOiIOLbquV8lh66Vuw2b1H4wawnOW
QZ6lnareLu9i3wPCMdZ2VwI6esyLEcLSn/aCybuoS4lVomhpOcmJhYpxaA+eItwb
J3Z+S3v62N2nMOepilsHWjGJaYfOi/G97wASPjN7CgX/mfYmGB2DjqJq+eSXSnDG
zMaJy6RVY69oJ4w/IFkSqk84mVMZkdiOOP1bdFoJZCnrcBgemz130dvNLkdnMqgQ
BqN25DvFoYvKHqNv6saSKkCqRWcNG9E69jGr5Pi2YE8mrNb2ksor0MwxmeLyJj36
837BpK1ltHphBwSqT5aozxKTVwQHcnJVr4WR76lG9QmnT+CUxgZuNnFr8BoNWjfQ
GeSZdGCHY0KscadCtDAO+3kyw78x6JPuI26K/ckJWveeiQ6FeJhoAxIm7vXzKV/p
Q3y2+SEhuxEYg9vZpckfZk5HAVNezTKKeWQogrm7cBAMoTvVCZ58XVyBpOxsOvJ3
J2NIsVx7VNGUuaMr2/+COgy6ihPgQ9+i8nVIROLaQVK/ufStqdAstWRdH9DeJ0eF
2kNxq5Mp3Nb9Rj6FXWXBZl8XRrhQxgihpyR6LkMAOs4wuObd0+4CzVRCqnNbBrtu
3UpnKhBHDcD3nKPDWh2/10djS0IVXJwnSpoMPfkPk+5hAG5c+nO8EVv3lUcICJvU
XPCNlsA+nhzmVEVEAfIqWqu9TgfDVsJzn8g+guy8fH+h8r2bnmi+85nT8Ecbkr6j
Hlh+dcRakDI9Gz2cFXVZbvufuNTlTqnJxTY1qyvwQkHfsm5hP7hddKXBS1rSWVRW
bf+jf9SkrZ/2N4BFs+2zS4v+RQjhHVqO7kzBtzoS2z/DUugmYKrsHsSg+0kHXTn5
rCdiqYDssiUycNOqGXzdYcmQvYRTS9iyo3p/68tkwAmzgNrQ6hECWUaqDtRMXGgZ
nivxxCduf/PAfpXCAciOOFkVxn6KVOPUqF0ISiBUjbchQNKs+q9Wfd4cLR5s/uWV
xT02+7RCrHCfh8LuQhAX91SzvAOjdlnEWOK7nZLjOTBWXFhO2Hv55W0wKVFa6OW1
b8VihZ0XxhW/SJHrmorB4DahkFM3AkOr5ZVQq6Z5NsOrpUNbgaDFXVRawZrttphe
OzPwFcBYXVB6X2pGSb/7WNcRC+MB8TlXpgtsedAESceX1Y3XTvmsT2CZqVeSi8Ts
54MI21KCz9+uuq1+4v5+JgIDvV5EcIxZI7zXPPgLcPn4Kfth/bSjfKv8Rzi5ZHSO
kg8SUjOzN0GtQZYXKx+OROCRDItYlKXmjYsYUadQnoOB7rJKpEwSj3UEoHmHRdTE
ZvS4lh3QhpqHJXfHtF0eJBl51sVADDPJuDmJ19zXBekTGcpC8dbN+DCQLoGMRGEl
NvX0pHssqPH3DVjXnrpqtnLM6y4voYqR65fbutdWsE/23Vytt4eonPj4wGUsABzA
N+mTFhaEro0ydwLXAorDJ/y0or7jMqH6Z9Fwy9229s2Z/OVXB0aeEoPY4aDCELmQ
VvE3l9TFAW40HT3Kl/gKdxZFK4rR+/1tCdjCSIvdrVh+27aEMR7B2a7aprnq9BkG
3ftNHaCT0+X4R1416GwfF8Ch+7bhlEZwq0ul6K64XaskoQwUFunugmGgeylVpe6L
rsDbIlU03lLp4RHgn8Cl+ObsEySIW3tTPlcUcfyXXDyfbgE5/Sfz13yQsPbI3xNR
U81R7Ad6rjSV06Awa0eQNTRpTxSWl9ub9Tpdo+YG896vGLgtDr3LgOYdxkNPjvjI
silsX1WGS5rM5p81nXGXTR2FbsgO9btzLBWiZaC4qgmhxxy5JZPw7d4ZT7YkDkoH
kwYdY9hn+ZszV1EKmaTCh9lQAKOxF4dk0AcNjKgFteh1WL9gL8MA4V6X9J8fusIO
qumWZwcgwFdS5KBEQC6ztFDq8wfPmENS0tGs2/NtLL2j0ukQ4ia9zlKiZ9XL3bxf
xa2EBGTlxNoJb48Twmsq8MZiFOdFs4PYg5Opl0J0dMMKkQf5kr0gmdAIN+MtRfhr
yFLcEIkX4Ealoevhv29S2qHsbaZ4zvLlzoKnLp8TjV0NzVKpGaNQQ5dtXbLMneok
paJhlhUVrtxnvNUjUOKiqEOUxu6n9f47aysw/D6l96gHX8MtuVEKKvut1ItIMQdu
u/1XH1iMAmxZOvCXmhySAgURoHoK/3OoS9RZJAqr2C82ExoLqaYhxIs9RVyK8JmM
NlmK0HC1DSQoUVv5FiTFaKVlleY58RKmrc1CFnMRliwj5c3mzHRA129vazfgeQn9
clr/pfINvqmS2AYjr90yQLnB+ROll9cspExHv28TXmuoqmXQwK7zBHK84ypDCaZ3
r9yAEwSpP8AJLFaCcTYuioqJHY+0ZRpuuvTX+llBTHgrARtVXIqT64OQxGjkv7o+
2zqLQQFGM0mVBnZxWJ42nG99qDiYRpEFL6I5hNh6ITRDJO8KP/Zisn2hnliGKwvf
suSy5WzsLE56GRTEaHKBennJyiuZJAlofNetkLKGnTx0N4vgf/qNOML6IM/hA5T0
kWei0IpuTcQbINO7Y2o1EZpyn020FGgUWKkYx+aD04GTDdxhXZXRZsXQFh3VB9Ae
6jvxOjIcEsi0qPZ70PiVlahnCfKE+Ew0UIr/BZf9iHdQx0qq4meBzc2tl6gTUySr
xoQWNV6JN6ZYp2plSnSKmHR4PLiKKMZZ3Pz+s4hw3xJK2G36MKk5r4Yr23lPyxLB
UIi9fuPA4Jnc1bx4VC0QIRJssKPcPH87U4MMHg5YFHKiJKj43RHCLikAuRyJf9S9
EulCw68jLb9pzsXqez5H/JW/2PA8kt1FLFcHGz4i/2rr1BjJKMuf1AX+yE8VMuCZ
rbW6p4BnYahF+OYeW+lK//crugr3VpaYx1zh1WjNA+TSWFIsQpo91zYpKIdsQhxh
BaUpoEQNMdYIYRccF/XCIDXWiI/6pil33jpvSzTuk8LitEB0OsnhgbJo28JzwVo1
9D0HClQYGmNbTpn+9iDlZGgARHsoJ51I4I1wdhTIkzAfAVScCcdqh6eZxm80JZ3Y
U0SzKXdlQe6T6Kr3EjMwQQPT+R1XDBMWw3STBkfpqEWCpEx0wxcWy1H2TTCqyFkA
T5NhopBOFtXuIrPkCSt1UBHCrjGe+faN+FV6LQx/+62KXdlyP8pcuwFsZCS/9ENz
BbC+gTBFrGwuGQa1nqXjVN6U3iAumPZ1m8DjJgowMK2w4wY9daqwvzWIAmZglK1M
pJFfcE6nw+zvD3e6S0/zMCwuyApjfNmLIU7vdxEAJwPHNEE1ouMAGmS3ZqKs0wWT
A2vBGIHtMMHFxEVL0IzWgYz1fyJYANXsaVw5vs6D3wcdEysqOO1NW4wl6R32wd5n
gO2aJUkMr2kdxAhVgclLe1FEmj9yhcK5z8btaRn7DE/ETsFVUIG6Jt4Tm6Iq9CdC
Atl7Ud+qsqk9pnH/y9rYUUi61RYl/KztMCmNOMKH1iVpDh+uNglDjVoYxvdYanAO
S5aG1Squ50OMWorm3B/wpCkUD1xNYfUdYtyiZbC6PivBMo/3JRYn/EA5B0osMsbP
aj6LGLXY3PI5f+O+aaR5OjZqAvSydcpTn/+CvuIuFUcjiJUoZPxbeN6+SCr94Bpy
lmWCoQwuCuZwLrSERWSHP5qokMgcc2kMJT+JnO7KxgsVjuzqhGv4K1ikq6u6JAXO
h0KohrIXhc32THeYuuJL6KMzG8irq5bJYV/Bf13kc8xM32S2cQhJIRO3SPnfHEGT
Pez0+KgzqKFL9lXqFoD37XTr++XL4jtvCnxsE5ZxecbmKRg/LtsQu46I+ND/cfU8
hXSXmE61CbadxmNZXrFuatwa/RrBob32I0mC3pd5LDp6V82Aj7iFUDhZa+oCFz14
qHbFLx5Hi2DfLhxoE/MiyDHbCWlgOLy8ZmlABmWLUAvr6PQJMeABBGmXbXyAa0/i
9eysaU8gbCE/fxDoruLW+EsZLehrI9DYxm+OeuxvhR7W2elV4hwGe9K/67s8dT2N
D7/U526YzNRnRwKF8muA9Ko8wKUXebAp9iPPRJAlCIc+CmGtqr57D69nH8zZLxHt
svFA+4MDy0Hta6uuUcSDMu45r8kUPhIvYrH7A5GMG4AeejQEB+qqA5z0RpWE+dxM
j46AMkKsWG2e37Jj4mgX1QWjgr1JzrK3s88QV/2A7Gtz5cutsIPuSsWaIFQF5UDa
bdY3iS0uqTZYDiCYOqPtrttYH7c4ZWzI5VdRsSLC5ITa9qWDxA6ceVAfZvLbz2PR
LyhAZ1pDaI6DXWJAq+6z1RMhFIVo444n6mKfnto0/XqoazlEjC7D2/1xzpf4OX+S
SYCELgZnEJ1G+9kkE4IgltsPvzZPm19YV1/8Nfd+CpP/UW/XfXrxh3QTTMQH4331
vAmqkxZ8UX5GxzdclXhq6QcoOuOKDHNHcu1cdU3FztJMbEIrD9WjYmTZ2DxdOjMb
56vfJlbF6fea2Sf9pdWGhSKfI64Z/W3ulxb7ow3h2YUSOmuY6V/Zkk54M9iwv7ex
1UBHWLmZCGGuzYi9zaI4huu1ny0dEWpBCRF8mOHem6nIh7/2/faOUH6LJkN9ih7e
NQeV0PD4b/+xEoEsWPSa2oH0IAVM4zxnRsXwoeOwN2gNPgBYoSIG5w6t1NxXmPd4
DHnWZu/eIX9nf6P18/eWswKiP53xlpjfjw5vYkKpE/hUufFh1fp5uZf/m7sNE36Y
OvrctVojeodmppcxEIczIsByc3drx7hlHDmQlDQ/OGidxsyTD6Of5eCMrkphK0Jv
y8f9vw+ZbBOGllluUtlposL+S/5GGpC+XB+OCi/cGTbGT+YrhmM2TaD8MENSFsQ1
5orxVqWEFTKA7KE5lvLPvzRJc3SYxg8AffBm0SdidBdwEyXkYgZ8hImzJnootc1A
FZwKntolt+JJYfF/1HrrFwndBmWBeygoMBqTfmPhhbmHeVmx+bC/6VItUTgfco0K
ZauW4EgazPNlCSKlSUmwJmu1H4tmldvU800D/uRdDu1sB4d7ZN0R8arCmC8fg/FJ
IOdMr/6DLgOxG10y3Jweu1JQeOS4SD8cTQQCKcmOOmbcm6Ws7/9B9tvD1/0EODjl
aWgCriY2S2qkL5RD1IoLK92c5e617M7t7Hlxi0cYDXSw/vCvfD7SqnRD8V47sFMU
3Jve1Z8mC65/+DbW1qeB3TJQU4nD5LWi+fY2aoRGOu4331KKz4I4GbJeSgoB0PgH
yKfYTBKXMTSH/CgB7QiDvjHMSNwt22RBRujNhxzSTsWGJ0yqrmF6CGPEWLvWKb58
huS3udaxDd6Hk0BsSuXMael4xB4reJiMqvAoYG4prVgkdl9rIPKMaz9jqpk4ZFvm
aRlO/70lhb2JDtM3pzQgy0cUAM2zJgUDbm6g0sTClBBTqoswvR18avYK58kGKOWz
4eo/AO4zmdeDnAaht94BFCuziwSwEiVSNCdS9haWYTdMlIWg/tiiYbLLrCdj1Wc6
IDa2k/ZfUsjf/iaJao3OBgxfSo1IRtcKhVDEZlvysZDdIBPH9a5cXWNX/nSFq9Fr
lgTwllbhcMZ4nnltAwwVUybhAl+xUy5JVoPAtrOv9aWu85MAkmwZPNZKl9I31z+K
SJkLHRGKsfUf5pKcnAg/qsk0U0gyrO2kH0v5L3GbiihMF01XXN3YkDj773fedxIW
Um3LGWjthYbb1u3j3QgOua8NPNdKDz3ta/q0Kji2kn/jkkL1wW8bc4g3lR1iDBWJ
lL/kHPYt72mNoiAsX3E6F57Ok3ovVgdgxwRBH+qX6YfEXWMV0JOpJRil75kPpHI/
AsW/pCR9Ng/1C4mA5ppHo1WFc3z4I6qSb+efTwUFBymtFQixTSxyQ1h6Y9a/fxRL
aB7QZictfHR9VVI9stTLFYvRxORfEJcqDMVY5PWBry6qG9zxaq8fXvNXX7Mow3zN
g6fCVYVGZdfCKdZkwZwpaK3r5CGfaHIMCMMBCHNUnbZLUep1gowsLVzD39mcij60
Bp8OfMZJQI/tu7rcPlT+vKzt2c+oFEFnOtY7o/AwmxEz1dBDfVT+egVN4zjxm/k3
26hRxQsnVvtMl+iP7r3XvzSCeWIjn74yonR3vcYswoWWyO9bd4LrF0/zIYGT2gA/
Sk7C8pj2CC1Z3teh3stt+JVekw5EcqlusTnmMtAcIXHvUgm0BOkcqouZOVsvsgg5
C24kYGPCdtLj20+yjVXdUPeHZYXRGYnc+ufHgz83Vyc/ydpXc4tR0m9U10bXoF8o
6EREYz0aXwfukOY1iZTBaN92+Mp9IKtbUSdS6qHr3O+BJzGFpLngPYQ8hY2qn/W2
IyCuY8cGNPxXwRMQULsgmePzOvutlk5Pe7nFLCo2PkLpfET6cBcvKwWPOD+OUEJK
6a2MFfdXbo3CQYfHKZHkYjPaGp6KIBDnty1Xs2D6b06qwVjvk9hg6f5BNo5D+2xP
nPFp09Z/DOoj6BJfSFtEs7WyZ5PBxP2tEciXsuF3S4dMdxGYAyYz01WKVEJ3BT4Y
ubl5GPXueB8AFQZEvG0bP+2uNOUOLfQm0pAxuEgIfdWnlippNHhWqL42HXS5d3B8
Mc4WlymrlwxbDX0mRU2NigG5ygea5wjAMn3rQ3I1ZSs+kOYthb4U6+rbtUuYJfzl
hr3fqt2PmvsghYmhMaA5Y7CmzFiUam4TQx3KHUKaqwS1EZJdZgwl0B9TfP9ZABCn
HoOyLwyceLQsMUDnAdqqueW4WP0PQ6jc7COC8cJkRsIrOfIG2jcZcjeM17mtMYdV
bs8yBX85KSzFOOjfNVRN6KWVpShaqh1FczMS23yCu78bWpLHJ/8S9MZ/ERhQTKt/
qMh/kGVYT/tHJR+bYA1np1hppeDZoojmVWI+A5sWsNdb5ZaXC3W7TRb6KYgF2kZh
xOpzrd0Fn8hVL6Tjql6DVlB0AyGQRGEn4kSlpPl3vmGePAfq+c7KYIlb/lcrPh75
/jwKNnKxsR8uXukmfj63vc0BcSBK4be6zjE5E04L0kFzZzPNc2gjGuIR9ps7Z3em
yaPlHks+gDffiRjiyzM5J2oEszZRBp8T64ocLR32LJ2rO3csr6NBavA3j92iqzvA
NIqc3D6kjnokhA6bBFnxE8LcxxlIS6BCFtMLzgNkP2IYRTwSyH9T7NBzrnLZt8bw
WfATw46FAiApw/XngAWPwxeZDsDI3C+vcHC8SZPVAmQEURYDOVCJ61/jWg/Wu/0w
PnuZKjTcf7roslRvPS8CcEw3/oOWmUEQz/Ll3Y0A0H2/ULNCfRvSWRKUn1KT29mE
RzGLLQbDeihfDLLXPFoKfpCvWbwBpgA0GofblmrYM7TV/mLHm6WbUD8rZPq3Cv4I
dEav0k7ikMkD0OzSmdL6O7Jn4vtUGnROAnv5fh/3MWPhbvCWIQ2o/DlHTSvNW80N
vd7gQEiO+XS/vi2X0CrazuNb094F6QEoL5NIYnRo3y89MRog5Zz7lPxVB03B1wks
ApaTZSHyJ4CrJvqY69s4Tuyn+AQI0I1HxvuIYet84VDNrJdiokFSAOlmJvupneuY
xv3mQCX2S+Id3HMIk+KNcOAS69BUSeUQboLsi+xva+0lSZ5wCrRYlGpjyQZ3Ao0r
q8gZR8FFkg7ySEa/sETkBt//fOETkT7neQrimWWYIutwvm23l7ktY3dKtj1lbRuq
s6sV12GMeUAP544j6haYkiy32ZDNY+IUkuuvoCVkPjPLemF+2xGWU6/eFPo6Ggyk
x/Qe19nVQtwsgtTKxDLjsC9XOcrvOJ5sNRewC4uFZp/mPOJjHzEGsr9ByVNSiGfA
b0SwVlKQch+J5UaEmhjZybXkt9ovd8pG7rzmuoeZncLD6bYcTTulJbhk2SElGJw3
0iJxpfGgBD6VuXHSaxFTphscgbVu60oujxuvFxizjJyRwNR+yibutraQy2b8ldM8
tK7TJu/lJCMZg/omvye56Q9j8GHLD5jVjOnAiszVEY3mTeR/UCh1/VRU+n3IpVIL
NrhX/6KJLtwZuAzjrueft4g2q0gO//1ZMP8HWnVDZMmT5meUY6oxmpMZGayAdT6n
Mc3vrsxLlF+9rTdp1OhxketbzlAzaKoGsGeekUg1PllKcvrab+bN7wFwd9gzYsOL
D4Qlevakw/YrTSuKztWg8HhsDu+PKAYnJQK5ubgnzmjbB0MvEKT7eLVGZEpAzPdm
fA4O7oKoWI0J60ZrwFZpwTJamZt8t0KsquRxNDc9NQ4WJPCIstJ3lY/SsS4+e2Ca
Yy9HP8iWg8vTigsjJtxNid9OveN1JBFJfc6MmnHj5c0eTtw5sTL5NrWlgmxc05qU
CQpGuCUVCuAvCRJUMpmFOPqjnzxNCiKETWksXyJmgg5xQcr/anmihnQ5/ozQk8Sk
w9sPgi6CZJ68pQf7Oc9nTmCf1Empe7but2jX4tm+8Td9FrIdCj2jC9HnKpo2TOYf
TpohIFdwIIGMcUIRwiUO/an0S6tyKy13ZXCQPcgGMx1HVTuwcLnb+c8RrdGTfi4v
x8U3xI1Ig10Ll3auxVBEwG7Xvt/WmCBMsbVXrAtC4E0sXDVON3VXNYsrt7Bv/+CS
u9FgfbZvIOXSzWRo3AQypnlmQlqGBms/KUhdarVaNYax25nzbVvykZwvFQmb0RU/
geP2Y20Wj6n1mrsk9KlzphrSlYoTeTi2xWf3FA4I0h5oI6WffJmcrNLxiDTzUcQf
EmlhxjK98rajOGy2FT97tDvmsGrBOAw+9tNPOitseJHu5cvqmoeDCGxF/pjRuF3Y
nN02K2mfOJ6SNvNvs5bvelxOKEzHHYoKPGab8xoluAmXcLcb3OK/TxcFAWnRp0bx
n5RaR+Eioq3XxRrHcuhYtqBhZBhblA86LPEgLimatboty/0jT+m3jxK+98lGnYH0
y6SEAuGdx0BBhB7KM+NXaMkL8n4sLeCCPyUFNJjfQSPppwSQBhIAqnkCXI2gO4HO
dyoDb6Le74prswcTMCl8YvAC7eWEzIgv8ry/1SVeoGQ28FBW8NNXhKxbK46p1iOD
R7dxuzzpgTlhAadMNP8x3A515ii2ZUf83xbG8qIKNr3QJeDY0sd0HyreDKDY7J3+
GpXvXQi/4AKg7uR1GZBP8liXiK9ibNt3Az407ZuHtdukGdOEOZSWOubMahBZOMrW
e7nSs/Ze6GbsPOWObf3tAzMSeI2LDjzTAjn0jIso7kLDQKiRQYQ+0umV7xLwFYVK
E2Ie+FdRUwW3fkzed49LpPNRMbrWfZ3fXnkm2LxS7AC3sy2LguSCl+/v9H3dIo0S
BCANIbV4vhPjdSKAHIJdofkRXQ6TVlN/H9uM+Qg3lKb1zVYD3VADqxpmPaao/Pug
HSqT1VLjZKgQ2RKU4vf4zuptoDrGRlwxLs+o/SLwtRc9TxGTwvcZ4rS5qOPDvQF8
4CnUL2y0Hj08XbOmaWQ1flKx2vsfRbhqwCi67MGuKTFoDJBJ9ypXgf+iphHm50mx
7sEF6Zx0N1js9CO5Li7QQFcl0w1yI9UdYsXgKfipXsCQnBWrq0u5Za+dFSH5Zr5x
nvwaVWlTBwP8jOAd3kR+tqbfZMxcvCbjT0VmQNL5McE7B5bzCZkaODma9/mji2Er
FyJPC6yO31+XDeM3ZmU8ldnMOqAJhp7kWHlvAFpWW5P3K2doQlH9CpvkG7Ho70c2
ovOovnPCN5yoFdMnoUUzuQ9+Qa+SEMKjuMQ9n0pcPBHXZsgeQPGxA1IqkuzHQzk0
UIQ6ZASfYIn2KDmFQcIW8beMA9MHTNhzx96fJVdnD3uN4lK+Ere7xkTvsrmHWs/f
KmqUai6kE4m502N1Crxubhzi8k9ieHDR06kJnHVcsEvlgKmZzczsTnMUqlAN06lw
NymH+lPXh+YyjUHemr4djy+R59DZGM9PqC/+X/dJQy25Ulfr1Voxm1yu5rRXQD4W
BHfyu+c0R1HQXRJMaawJq94z34NOUga8FVSTPRtgtyR7tGjPaD8IIQwrNU6VlyDk
QHAahl4cP9Yl4hnPZFs7RxGnZQ+Vfb/uAbQ3YCae0qU52snc7M0d4bQ+EVdutNM+
/f7xVVrc1L5marSKlkZ4EG4BISd+1bbSE4oukELxp/oy+8NcKtXtxOC4xUaJxEH8
nZ8rk5wbsMYdX3wD4BqnQzz351YtiGblsL+wvnoWOp8L4UfGKL64L9heAC/VBP88
A63z2kyHUFBzCALIoTdvaeXAmGJMdqdE+lbgPqktFagSXE1b+xKkf1FhVyBgdGou
s1k94FdN4DrFnrpdgWxBpey5PAWj5DIhd/DfwBJwo5tS9EKs7+nGbfIaWL6nKl9f
DHcI5u3z6qLPll1BU+HOsHRis4nk5UZH8BiHFkoASCu2uq8V8LLOaETIDhnTyFWN
SWv+sl+TWMBzgo8mTOgem93n6KHR3wC0jolIjCt7FccPI949iRvdqt22d6cdy3bq
I0mWS81DGzgwFkBNOIinyWICdsqP2SyI0iMmkf2Iw1ZImRASDVK30/ohx9AORzTE
tG7HV1xvsKkivrLNHUoqTS/33xPAs6RaKL0MdozMxFPrnKNn607bxiD9i4psTR3t
Gn7QbaoZvCDXYD/76jGj5pY8oB+IKpJ0TNS0fiSgru0rsH81Ir5iJCs2E0Pj9sXL
QtlXH5RyqwCfY9tMQJnLZVgHPl6PITTgQRyMVQWPJsmy5eMzuzETJcCptsKcLNPe
02d6olxdkyLtslD26XfOqdWsGjGKN9pJEFLpaa0zqCIxP1kM6bzQybFjtol+zpDg
afOhDHsLtsC/mz5exx1JbXYIyyAcey9nmg0/6gx03A45jycDu8he1P6O4GqzyXpJ
pjdJaZVozwZZs2+TqnwqoIs2HxTQKd5yihYS1bFo89gVUX9LPgZ+QlQ3xCnJcw9f
uBVeDGxAmhwtNdsejlJ7gNhSqQZjob3ib9VQ7FWofIyBBUCBm4JBC5fgZkgmyMl4
PL2M1kkEF43SmNjtsD3alFcvwr0kQx6ASlFHy1IZE6fwWrEOOTQyd6/fYtdoSMOA
iI45+0p4n5MzLY0fZUlsql9MJwQEgPQmQf0/CkfTcHzODkd5lz/px/gztWcLfQQM
WmEzSdbGrHTDA6fjd0zz+wz5L44gvw7LWqnBT355l9ADpb0MIDt553JvBJnh1TvY
/vhj3NBXtOFuDIm/NXq7xigMVxr/V3nQ4pTWcGVkdPMzK8AKZqiZledjRcmkinsd
8j3AsUSMK5eH2zROweAMEla+duvbIdiA/6L89YVO4+zOrHhM4foUQsWbyQ3BDY10
lusD33uEzmpVDqKtXqNZVJT3j3lfuEO0xAO3xGvZ2ecJgz8n4g0Tx7EKsSkV8zt4
AVkRxYaSfYIyKK+X39yEOzChkQ0ozBhsTKQAq8SLm63ih2ZUM2IsLR3bUUc0NDE/
3GavIDeY2/m5Ar/qvR9lD7Mnxb+PY9pbV2i3IhVj6SxOab0K0v62MnxuOV4uNWr0
b6a5Ak1i/GLeIA/fg43QGptdO8Wx8dLmgFICnmZ19lJHCAy9GoAaF6aIo0l2Xf27
2SySWXbiNjYOWsNOeN2woFjhjHcAob9Ny4yyH7BXHbY84kNh7GWs9y8y1OL2MaPi
pkpjxET1FSb4LVIhdIrAskuCXWC5sQQXCOOrNYYGuwBj/YNVz8fr7/NGDOp2FBzr
ikuXmTYx3/WAao9uEMDLtMvap5FdIaD5/IC3zQyl4TFjmxZK/W2eqwIMY3tZ/A9L
p5pbzIQcQmJf2TV8gE/bMbZUMDE1gLELtE1a5A6vQzJ84Kjveno0AkZqhd3mL92H
xv4Xnky5cOVDx5TtMnWpRKyDoAwupAOg0DLE1lJkMoo2trPyljyKY4jkGuk7uMGb
m3Z8mMPvUit3vjAPP1yC5E5muUnirF5/UeFLzo+5QS+9cQk4B7tYIdvqd1UCZwB6
uG89dy8WKm8vhsZC/FkB8xWqjT0UVAhot8AiN+QdoMUcHAsFT3gsBT0YzlWOVtQI
JG86n2G/xLNamVPGqtCJgoCv0dkWEYAjBXAYcPTHZfSTpgUVQS6BJnDEfQpaoguY
q7JSRM0cCEBZQwl52wW7SE4rIrHpQSvHHCzKSxjnGhRtVMCvOjBMq1tkZBl7sFVQ
uyOwK9sHOwAemmwjr9/C42SJR6ZQmaHoD0bQbapfqeHElC/PFSx6YlfDrSavLiwY
RnJomKeiJv7brdsybi95mdwL/Kv+qCFu2xbEKTuS1ZX7vFcOosY0mDFvad+qI1Qi
02RFYURsOUc2mgR4SYPfifde5eDQTUoI07byrWf5RHkoPnwRr7sttw85PMb1tGrH
w/oOu9P+AJJp+c/0BVKCjXuIdoslNq/P5eQouWQZyhmWirCqKNVDWqn4UVH/Wht6
OmDr8s0F8m5cvo/Wm4N3Ce0oql2NdXj/oIHQctkRBad0LR8r1WltDy1ySv039utt
7Z69y2dsh6hlkojuzNlOG4AOYJRQ7Dio14w8DyRfj6acz6fLmpf82nBXtFRwPt9l
dc53gas7bDvGPUbN2DeY3XNXuYMc+DUX4evoXHp/+GM/VodKRiZsUqTIJjiTYTc4
1ISH07MTh7s22bZwjbE2KJZtgjGPLCzt+NsMCgMjP4JSD5L7OjNPeYWxa3/XPdN7
CFod/UrOLcvkYo/341iuSgWQ4Z84+as3YKekZ3jEeKvuonZJ1PqFNClFu2FYRR6t
2HtC06KmODzhFc1eB2sJyABTV9/lxE/GSHo/ddAwWvkfGTK9olMePEGaMwAbYz6J
cLWYfW+aQ7f0waYWVxEYR/ld5V9aTsppEUg0eqFZUjeWY9kCA2j0Rm2pjjIc/aIU
JHkzXOJ7VhVhH/LTXXUq7EAJY78aq5W73B1WlC73GwhKkBpK4mJo0z3oVBOc0JD3
T0mSuZAel1rSdlugHVRgrXuQU1+bQIABeRft1SufVXdmW6TyKMxZJZUya+YUVvme
gocZuj7/AVMkj5V6UjezT6TaXQ3t7H+UYI9Uu47QSpSK7dQPeNsSE4gT9LCRr2qD
wL6wFzyC7yNVpqDHk+WylJ9EBWKrB34oKtYDZMacgvj46Ro/zM5B54E+XXlE6E93
Wy+zAPHRfzShT0jgiUF99/cmZjz95v/bAukLA5fn5eOPqOI7HgOxVIO/OJNw82o5
lTIpwdjZfj2XqBVpc68xcHgG6yepPFVyo9EqhiSs7r5tKPBuLvit7YPQot5WsGVg
qxgdg2+ceALZkSAJl2xNsE6vZ3T0LXdXCeKIPDoS4r1FvMxQRsCCheprot/iAbJO
i4lMGV47AeayUU3SxFP6ER6fBEWMxcJlUAJfoMxnJNBaTR9X+Qv/DxVMOJmTIzQ1
WNa5/2aBwgUuRcV+EMegbTj9OLU1vJAA9OvGFg7V9TOxb3Gpl4vrldoOK7eiHDw6
NNjaPQOxm6JuZ23HE/5qAM0S9pKmxxJ0WTRS5hjZKqJtuUwQ0VqyjWi3DAeJg3/5
QFCm5ob6tX6U00K77+IHg/RgirhvSPyQ1Zx5hCw+qDBPbaBCzeNgg1j4cGjJjLZW
j5NWrEJMEyQf59hPkolPfowwuZySaKIxA6YfRrvhJmhGjiH5HBhhL3a2yg7AGdbR
UR2X19uc8w9FPmlmiLm8Da0CJ1Rp4GS+RLSkMaQKsHLJhWodmPAEzgs6PmtORGkB
wcGKvBASzZS1iyswrYxfu9Dry/bXdWeMHZ0bAJ62XXDphUg5YwRXQzywoFhrd5+z
KqTdFymHQru6zXS6sKtcNLL4Zharit45iJ4mkMbg9Aa7rKhiNkyG2EJ3xwYyQdpy
vLL1bIKEOlDz5eWTFYdnu7ODpeqEQ5prNsy9BAPP3W2UxM/7HGjDX5Pv0EsZhdFJ
1l1wJtJb5/TtQThqfMBUQ6ljIY1TNlqrGtMxuj5mEFgsH1vvWdLjiZKwbUhteOqz
hQz0oXiq79N6UpGcVnTH+MzbSCZTtcO7pAMyZTOfGyNerDpABImZfgrG1XLPvrr7
c7rBqyYGlTfV2pjVzSHHHWwWfZ+bDrXT/a4y4Vys/iWtQSI6oMKPUNsBWiKbkqge
avv12iTh467IxGoPKHS2//QO9oF7tX0iI/8Pe9KqfaloZ4346E/5CBd96s/1zlFi
WpfL2DAGgZjpvWWvyptj8p/G+1OpVLkwnV1ANgjGmIZfVYZFzHIpIvjh7mkB3Q57
8tsakAXe2AhyYD2cCQ8awcMC9vi4bEp38Joc6HudQEhQ5jhbmnf+r+0o5nuPEnhs
AC7aa+SCNnn+UJgqDcBxpd0OcZrCzp9lQroPO83yXiHJGOrUT4dzpYboeAfiIihe
0MH5BarYRmcYifgnG4nMGChJJiyo2ZM9x/aBQrVwp8/JSha0xOMQHwjStlaJ06Xm
7zVewH9eMiFqWw8RqdOyT/W5BnLsYdzksaSgb6lCGI4q2U0Ujywz0RwKVhz9vbee
ovnX4rp5MT9xonLnndunRhDpFB5ZBy7p6nMev9/rhD5hqslHmV4SrR5tsmUkJD0A
BCCyDTS7UL7gltCA3sZNmlQxt+8ag81KSfZqT6bzwSByUB4Njy/RJftIMHQlGqSE
W262jMi3+hMEhftj2scYtJfsXYHL7xgnF2kO9EdaQQuXGhtYskP4BT4o3dDUsq5f
cM4B3FT2mxniOaRoGnfPN2uJjFflhhA2mY75ZF9dHa1AgS0nnjHACQouk1bx2Q24
D87mvJCNlLIfjG5G5neXa8epbMWrVWWt0Yku9ku5d2aUGwCva2Db5fWGM95jiHCv
Kt2w4xfCJ6IfYJiwFHqeC9ArRWe+Dlibrr5s+SfVEUiOpihefd4cc/IVqOND+lW+
sP8E9wpqEBSY0N2EjmZ53wQ/EBRsgEQnkNaXJj0RDDXLD8IBWZV2/PFjRo2SVhGU
Gr3wUeV6t4Aw3m5FqtM0rjEwm/wpgwrA2EMfmQOhNlIbkSr9Htw/RuAgojPgRYua
+sr3Ya7zUqWm1W+xca5RszMu375j/tNSBahpFgdSK7roOmTyqS3xqBYuxUxcJ8Gd
/qBKUU7o2rGvt8tdKEjJqS4C+HFQ/nR8OKnmGxkcB1X1sHq0+L7W6IAl7g7DQ9yv
+pstTLijVYhnQkfaI5oV3YqB2pXz4z/u5exBbGaHXYDh0YUH3xRkzK+ztTZfXGwN
GahTj5pBMp4POs2IbHX2PFiHXKXbgSieoJdbDSIEEDrdL9Xf9K/NxqLJMci68sqa
c75L7KtlvfnU5kpRuPXf141a4IsHr9lpOUavc6E9prN7I/+pUPqAcWv3nRWtCFc/
Js3oOCsIUTOaS2bzZg8BtYvwgOHpgGBtK8mw2kiMrQvEnG1F51warPfMuP8rXq8e
M+M0Xe13/Gkhe9xSQmLWcamg9fZ3YjxvVLK+6jGmfSHi+191X5w/zem2Gi1envHP
XCZXHR6brT8JcF2XRuJtiGMBybBTv0y+V7G94MjCFxSKZbCSd6rBhnVfqDK+BSY7
r+dSO9xwKJ8S26cz5DkERtvfN+Wv8edBW9Zq7SW7pagXHvf4/VjuH6WbMx7sR7fQ
jBKqjOIm1YdtURo6MWnfb/mqclGARQgSZMrd7AYx9+yFXrDUI+idxKGkxrMltsUV
W4KnXBcldZ9x6UpkWlqZML2L0PeqBpcfIyTeGLZ1rcAku1LzQrUjOevACCkV80p7
QLOt/rHUmsrdJuNZDh5dblL2K1sYMqXfy09ka8rX0+PIO1hYVdpEwI/AbxXBHZLz
dKwrWzQo1oQDncvvMH+2ecV5Pdh4mQCZlVMZ7Jmu52wIP/2sW0oThYksohjbqZWP
2QhECn+z5m5zJ8xfv/X66xtP1l2aDebyRgONyDOl3fN5xJWPBwmwzvrPstD6veWY
TuBWAJQbRtG+tEiyVxN2NCNAGUxc77Yxi81S2RT3mshY/qMSIqvWFejT3Z/R74gp
fiMU6yTvK3sUS/wavovWXsb5BtNiGzvtq5HjM2/qFIxJBT5fxOY4Wevb7/fl9tfL
DB7sOE4UN6h4Ng2IEdU/LAEI6H3zlLvgRm9INGirLQmZdKHZ+qILo+fI8WnsM762
EsPZE6KEYACGVlYHyacJNY/gpd7IW1ChLU3PlKo3k4Jmv/jCPnS7I61uggggA7Q5
qF7EYNR4/paEJ4hZimwga9TWEZBHx2eLo3c3/3yypBVj9HZZTePYBrrX0IbQwp5y
HoA6dRrYL5D8cQMKX1oPXCUJS2zSxfqGde3Zgcab62dRvOnRp5AYDTG5GMV8HT3/
n/I8bmQ4N84JbxA37E2PZ9wvfwWbt4q1xPx2Fhjr0cxe0J3+sNJg/jSGiMCY7PDd
hG27Z0fJ/aIg1N0HrdvCPOfbULcR3hTEMdPmfWAvuR39txEqWwkHNgVv4h3h8Bl/
aPWOe7P9zvA61vTK34kfWpg3HhVuZnB7EWkt7WePEwGPvVGxLOiHuyV2GIx4ywqJ
fP9JHNnAg7wRRNeWmQxId9oPZnT6EemrDCw4wPIyTkhZeaYbQ+hiRQPBaRsQqK1y
EcNyCPNg7T+r3dLShjlusBxC/Sum+9DqQz0D9spk64oFrX/yk/4jQ0EqKt7gciHf
7A5bqiI6BTqNrjb4do1HDs1euMWsHGBEmwgAVrWbIxh5TrQy9NkOmUI75a7LdwOR
WqHcmFdg+ZEKoNWXKJuYNxDPvwfjUh7jLlEJdEPzKK7blrz6Syogk4GJuggYE3OP
kGI5H9iQCfZHNgS7sj+8DXk1LxP/NcysDVYxyVQy6mY9AhnMHcUh6Ciwn08lcwSh
a74zTbggn2dbG7kaSXHr82926PXhLoJuzRA9z4ZsxcFvjiGub6PDUF9+cu2HFgdW
av1RpIl93maADuz1gZbLh4QHmy4FIgbSqGYJzlwBKPHJr6hixdsj6QeuWtYqwsjO
nV+ytQH+nnQk8stli4blvbspQFutGlWDMR/lX0t7K6xR+5AM6G/MNzXyPexizjDs
8WkjBX14Kb68cox3aMiQl519JG2BqELYM2poXuaTvBTjULFa7xV1p3cmPyXxFap1
0sYCdoYz4DtkPinYfmCLN/qYnTO5lRHSKTRYvue4i6sAM186Ax/qlrIL/qqIYEhY
rKQK/b/s8nmxQgE0/CVJqBpvUCp+ZfyYw69SNUEk6xKe150k7jmH2AxZcV5/hc9w
4A3AmlYNSPbENSUOnBvKpz3wZLWj1Tna2HRGLG8NEPt3RWseM0if7YcDKhHolkgg
flq6of6XmwdgUTq3Fgp5JQCTexOvry8VXB4QIgJq7vtCh5LO/VCWmLplrKI2GsVW
LcVnTUHiBlt9c8bXYpEUUInhCHdhUslJaMNrt0YRPR7I2I3Iu4YA64ipoQm/HI5l
UrCe16ECEsjLdn24XEYkEjpqxceyK/3Vf6bijvb6xdSgBWQGYeAlRyLlooUTr7Aq
U/CzoigANZ7IQFsps5NuTn+jFSRJt6783xGXDTwodV+JylgKNDWRGQzq0UN21LMV
BBUaU+1dch6b2O+rDzdAKc26m+00M/mP9z0iUPXuPPtIPrm9rhImmTxqTP2Q/yq+
Kwrh/xhnpAPlKts8TvU0c2qxxrs0SHofSboAQXWOzGfOo2bWm7Go7tgzqMqUH4sy
vgRVJyi/SbM0LN95t7LqWyhAVbwf836GWCWWEWUN81ISVmzIYOZwNk71z4rbTu/z
BNnIq4nPuktjWCEEuqDaCdhj2wl2/kES6Wwd3ZzCl9cybF6g0QMGA1yFZNznSuAB
WlRJEI3m9+mQEr7zFDxmEa7M5AA3uA8rlwyX3hvC/cPiWxTBRSmazGMYjQiG28hn
GsPf0L1MMLiiDFhLsZfI7PxudeszL9qipGhi3HV2SVtSMSsrFGur/eUGFwXbFNGi
IrzfkTyfRQ3HiuETq+824fG9pn+WRZDjP1AJxR3COestWTAX1QqxKua1Fa2lDUST
QHvCTWS6eVU4UDcHU3WQinob14/WsVYJkIaelBO5rR//QLXLCNSJdkOSmmKo2g7b
DqBDi7VnxvBUfa7f2D6b/CXxXSEdSU3CHazOhl/iWF6+J1JnNeE+aXo0qb14DzSZ
nvZhTbJLRNpFTs9jj1srRs4WUSR0lu8kR4tbeyAioQOcCY07/SthpTfzGxASIfd/
0GwfyyFjkYrsV/KJwLjOITADVmhYgapiTruwP/UINSEU1nd9w/pHFE2ziP9pGHyi
0TBGQPkWGCEC/DyTTKd62jY9POJm8YmnEtDVMtXA0J9edsgQ43CNs4u9Bg0CI4cf
lFqJLAFyrtKLRvkgUlj3Am545wr6YYY2sd0TA+1zvJxYMpcDhe4bamn97cUAH4aY
6sOXTmgmJX4xmXv4xhtaA8lLUJFINOFZSaf1zEf7M/zT/LyvPAnh8AofCzcbl2s2
rRIXWq4DYJ7OYBiI2SbSkL3QGECD9ZGObvreroxsAE5t/IxOYarVmKOJ/ZSm8TB5
8E1QARD3GTY25RIo/JnlAWLCrQf1b2LjbvGbAXhl2/YLkx2xmyt3D22vJRDDV+8b
5Z8CeqLdwcm0OM6KHdNoQUH1CSrZ07RyuF68RUEKkGbRRxmy7SAw7RX/lljadwYV
iM4X9s/e2wvroEdqxePD9BCb/pf9G4eInylSWZS/GIqbY4vzvHTgIW+xQaxmB1UL
RzsozIqQqlXPZwerWtDhv4V/bM1qSPILlTxGncubqTvbZxfsIGanfA/n7IL1OFIT
O5w4oFwwVQTXg5/wmqol2HWfr2CByQxv3MhdTaopYQzVYL0TlYkeP4+zqpqpbbrZ
ls2QxzVToqq1qKIQHFJqsChNQco/en06pJHhjyGVNI2Bw50EzI4/dZhRmTqt3qob
luVSmRkXfClXLiHUUSlU4HU3z0RSByUWZ+OmWrKs+PwN5Pwdg4I1c7igHSnXFevs
D+iE3lP+JK+v9oMv95B65ecol7vvLYpwYW4ww2nvZqjT8oOURvR+ExG+ubkpqSRI
wkQcNruyc9SKchEwyq3MkUUG7yMehwxGWrNQD0FlW/O251MTDO2LlUP8M5ohNPG4
vBzdxk2Vb76nRyhf3KMvEAmqGhWhUNTrUZl69QkoCu5LbDQ/CXzWTJayw8RecWgE
x8MMpzhFskm4yNKWPksfwrhAiESIiyBcuBek1wnAIk64ERPykOlNrZFN4CC8rEUp
3BgHWMmqozMQhvlaCNP5xz+5Zs49HaWr+XEcmx1UsigmWraubXQfAoVBj8d0BsrO
m/59VlHe0GYgJZkzcltcb2wv0E5jIYneDikWmBw7BWSSpq491E6RNXm75HxWuhOU
MNl4seVSYtBQ4sHCBLWxdMDBoI6JJyoPuJP73xXghXZVLTYp4P7FurjF7GR6Ckko
nVj0F7J+1SEUmNzfdrKRBcp3I9e3HgpMZzE9gok8uhtBbUF9nlS5hRJ1J9bHpoWq
85HPDFdN157Ag6a7Ds6J014t3EYvMdNaKhgNmDYGJ+6MIXdfwdgHndk7gNQ7HeBm
rvgqIzj/50Nn2ArfQHvWLFls4AdDdDubSoBcMJ334FxiwSrENttj68AjHmz0k6py
GRMQyGjUrx1nig9ZrrrKRHadq6WwFWvK9reG/fOrOY5wNNscfg6NcQaK8szQp88Y
Lc226Vs8DBGvcI2MnraAyKhqAC8v8ZjDS9MYdxuWDbBIoyw8kTsiNE3Us+iIotHj
ta62bWYc5hkBua/qUg5tKxNiLGyZ7+yehmi86szQzjxeq/0ndQGoq0Pz7036vZg4
pSmvINphu7qfCi7t5Tu55wfi3Acl5lKF1rYLUrFx5e4CbFifmRj4a/soefex415D
n2HduOV2w0kdQ0MieLnFcRUVSXUagNoZO+qeswzkogCc9SwoTX1wKyx6S8x8vSpM
J/R0nKkJXiaiZ0MxxA3FMqKGkKwWpG4IapfS1aScXFwoSlP37tMl0q/jNy8AIvjn
Sq3tn9AnUoWexojkGFGTDs9kM2OCV0KxD73yoFFczT3UESgl029Hv/Jg/2RFcH+/
aSbZPSIPRUx4vtvoW7nTxUZaAqg4c+Aq7DbIrYQJJvJPLJ5ZMwcHcUJ/HYBeHtzQ
Swu6O44E7prpPMOCXGKxLjGAfLivYiUmFVhCDiPU0kHhTF0iYpiVA9+iBhIAASLZ
4MFqw+LQU1X4XT+z2iparXc/Vs33NfLih7o8L0MjzqXXArxPEzYez15Sxpz94Hh4
y8pHcRje8F8QFanoMu/2EPjau8bWwScRT7F83kVQhBiJ/mTshWppHl9j94lQrtti
oP5z+hIpsWYlmTCbWftIGBK7mSGrZwru6MmHpaVDUXlhLP4ae8FHsZhNSi8zWRVm
HX/n2Bwk5NoObnOD2w5KH60YxbrBBW/YrIPMb5Z85NxAeKvalz4UxEGidkv+9Fij
mxkuHNdP0NkPLh0b+l9rDGjw95SuZ+lZmL2ASkicE86jILHSQfEmwMDVjOMggfLi
Ka1vWwliBpXCnhrejgtzJI2Fi8I21ITev5FXGEi4r2/4c4w8Nrhq8PVXAcwRjm4d
/wYgmn8p9wJsMewUD1chqOjXKM5uK3Z2+XXFRlHLBnhH9z2b4m9fQpmfNL+UjPME
LEKfgMT6oNlM7tRiS9Bqz/TFxgPcQZ1L/APFsIQIjTRcA9wBnA6IKN55HKA2isXC
YpPcwXU4O5tjVMHHKCwh0lL5eIKXlNspxKhrcycL/YiD8DB0NZ6CB76hpsp4Rk+D
B+VOB0EAOreUduwMV7PTaopFkNMfokH3hstFKdZC3uJXD0mhrwUt8KgDaWE1gQMd
vU5DfRWFNoRCDhQOq0oaZM5CvN6ytXlRL646cqQlQsFNhK36i0ZIBJgQdAoqGSk7
cCmZWdjE15hal1h12QZ0ivSih2pXja1K2n9dhHWRudLTNULexv9bqqMNnArZ6Ff7
VRjCMPOpYmDruVctlkMKbYyQcuyXDOW7V9zxG3uMOZkJDsiCsyKdQVvSC2ul22tS
dX7ICQOOTeZVLOjCmsL5mCKmgX/rwQ7g06aeKIfp7lhKYh+y3HvuHLZL4ojCiYSn
hPO9eOsCDMinolMH1cdBgYA0WKcaJXSNx2bJwZm+AjBhrebBTRc6iYPDzryn0c7w
hA1vj3uAPIaLet5MZfu6KffIzRnlwHjVwggKf7y0yCQVNc2cWbjkbK6uQ0vJm8uE
yCAvzVcM4SWFj9C0molM/1hqXGoF/wjVFDXAEkHpKmTkFLU6mAbCUHxXlsTR/Gyf
B0yesmDfpbpVn2Va8vye5srIPR6BR0dc+1ZdihytFwsUL+lYMLyryC50TzN0gr2Y
FYzgWsucbdyBpyYVxOmC9jHYX2UyASLFHl1Vqjtj4pI3KyZ/Rq+YoCfQYqR9vdkh
lTaAcmHtVDTu/E7DxVc4LncjC4xWSoSZHwvnhSsOLSWdq0Xagtitt037ore9ywmj
/z+dv2tpGPhg1mADpTr3AVmzSVO0/UcJkk8iOBmy+QK4Jrhom6CRuuf21JNVdykw
FQazDc7mjQvKLzP8E6ji6tBKVC9+NRyo/VlROZoC0vxgEAlDflY8J2rrNGGNFZxB
dllkyOIUbcFmB9j+z8e3vlACfkkNhnYjvo8gAQV9aAc7+9GIrMHjmsv+TufFOsAe
WqVv0+4wX92jO3bJmfKHShOCrYDNDCyz1ipsE+8VmKtmzpPaD02b4xKPOoSE6Zu6
qdG+9rV2qnM0Grr+SVPy/fRdxjiiwMgz4PF+7SOwlyD74kZnQPGpqE73FhP73SCU
aY11fgSQBN/Z+IPc5XUeBSyP2sArWWasRKrSRHSdrbO5Rbz4fmQtxHTnosgyi/py
yvTeCNwVCaXqPp/CVaT9mJGCmVlu8Tm+mqQ0HdqEIPGdOTY5M/4tl8IuiQ9FXf0v
O9CmUoXK7xCAleVSVHkczIQbcSRymnBLi4zRsGdfuvQv4+Mc9o4jyn6FTCS0YbJU
nYiHRKAIMQfeCdANTimGbQMh3qjsWh6hd4n6H7yC0Z2lgdFNU5td54Lei2WK8oSa
bfv3XWVjhjGRVr6o2MUU5kzSJSidllD5eJFc+mmr1TRPTtCqcBcfANdKmTghks0w
zL0lLIpQDTVqAM7oD11V2HE1UyXGDsy1KUFTbLGm3MVPZV18e27QWRbNRlaCtr2N
0dCc+w261yPt1zEajj4zxU1WPcWrGhQMusuPOMrtN4lCiqk8aa1tqqwt8giiSVRf
1KGRxwk0FCmbbWzEtclTdRoTQCTgd/bw1V+eq28KgyXTRADNUMrtdRLnaTtaE0j3
ZE/otX4/Vpd8wsH1BOH1Cr5X8KJPFH/Wv/EqrmDYONZmw3scxgQVsrgIRgkSYs6I
FP3OcNRHaQoVpMDk+R7JzpYLWY6XvtEYPoGgxNJUVsbMoyBMAotk7j4W42JB9quJ
kETRIwmGRrrPqr443ph3y5SxjLN9dEiylV2YUua7HcmQvJQaid5lCyQNB8hDHsoI
/pct948KHRU9bzsgdX7igCcZZ3pKJtxhrs++wCsuDvcvcAB1hYtwfQwbR9+sd+M+
DulnQ0tC408teC6nhLBr+Ew4NnOP3BwJl05fdtHOROx7pcLZ2FajYrs5dBlXmO5O
Ge5EiOxS72dQgTHNBtrJDhKv6euOch12UxH+nK4kHq1KyqOEC/lA8/8GhjXYBDQp
J9bsAmCeJRebHuVp1Jngwitscb1zqD+HlsnW6LAJvRpcrWxPpjb1PKAqnFPlBbsF
Qdy/IsK3X2ZXiHI6nPlwQoiGvYMzEeJCRfS3ivlg8I6Bo+Ej5I9+vPuXYigKfKgh
TLwlUGG5PiTEhqdq2kqQ9m3cw7upSppvcYNGdKCF//fOjgTNZOPDRkxpVywtpaS9
ylVdvRsxySIzk/7hLL4IUyJ1wYTG7K2IwT4ba6nb8kHCUUPjGi0aRVrgCdiw6Rot
hgFqB+dUWHlZyo/GH0xqYM53GEPICYmRNuJ/ilGEFhCjXiRLGSMzFE2L2A0u6+AM
ewi/yhMHvkTQlDXU6+bxp/55q1T7qPgIlBD+IWU2hai5htbYEJKGou/QL8NMJN+P
94Ov33WpSHdbz8qFZfG7KQ2thG6Me/5yifQkVhQ6GhmzXW5FRtP0Hlyo9lH439oy
5nOvWs3rJNgDY71olQV7oUYh3dE+NyHNxbYbJvs+JNotkrMmdalkuBg0++xLQLO1
/tECv+njbbSbK/rffk+gAJpFqGV8MQOHi5HDpDqZpVBew5z6/nI7LoPgXXopG3Lf
S5J8/vLBNa547tPF/P70dyFhKHR2FDFqiA+UqLaGNyXnH47s6ttEXLsokvNPxOf0
4EPJ6+6WWqoJuszZcme7M9I1sLyoJYidTpPYIoEgLVWcPPrZ4qDgIjbu4pjb+ky9
ofYW5DD/VSTVEHD7ee0RBe+ZpchJ0koB0hU/ETvtzTI/NjtaiTf7nzsKunQxy6LI
6Wit1YIpCSwu9H8+zYvShRYkNWVEXklBUXYgXxdkUeht8EkPWXUnG64iLcLoGXCu
NM0YqDsIT9Hm9sI9EIUn0greIqEq+UDjyxdcw9RA7neBM1KfrYn06dPigiJi5Dq1
bZ5O88WutFKDHnB0sI0GNL8eRId5/vCZCncEhvs6bdM2cLQV2U2LUHxN374vUREQ
fN5Ba9Q/No5j5BMgrBxxx5VUc5TeOYySgJIktOAP6hIgoH7FZhLujkmWwH1lyl+7
+CFR77Dc6xUSD8fIMvUwiK7ExBCQ89/gg1PJxj5YhzbD+Te3zKk6vDHkSoOp3osq
dN8Cb2F3PdS+h+D3MwENmygXrLGQAyyuvR38ongYaBWW4qb5RmERTFABLA22HGl1
md0G7uwSy6W2ASz3yAM1wlEn18t0QOCjPunbXNCdA3f4VYsXwuISLvV8snr7/2BL
F1ZVkNyhSfjegewnG/mJ8qmvE/PmBUz2Nxoc8pJS4B53dvjB+DanO0wJcUX9YQkR
tMApFFDGL/RHxd5vS47pSpqZPcv9KrNUKT/00D0b10QXCh8RERW1vJnVls0p/ufE
1KAjjSH2J7RSRn3FKu63f9tXLVBdzRFYf9GVVjZlQORouWmu51xZX4PabhQuikvf
umUYaTj3W5QQq+w+iSbhBoWz9hrwW+LvTdOEIcXu56Ge+f9hCML1uBgyGN/AhnGm
CjvIzGYDjxnPd49WIcqqXJACAq3XeP8tLG1GxpXHoJ77cxfP1NcKG5zZCPmEOWgH
XWode3NOwetSQpw2yqkfWj9NE0TYk7nA0n1iyecYfTXU46mYQhq7o2G80Cqe+HsG
M+Ydsmtheu8QzrwgpQES4b1VGpZeBT4KV8a81mUWnRs12oxtcGVCCmInoN4KDVkO
Rvgl7QdV5sMOP/9u/n/3AeyaSvtC+OygeK0X05gGh2YlUKHgXXUQMuGSoGhBYuzz
RCrFHveplWiIhUdVzwSRO9BJfGnywbcl+3w49hKZa0sPZWxskmldhshsHwBKTWB3
nd5ZiOwXK1tzg/Ty1byg3+y8gUbWiznYT5z79BIFCLiTTL3zufmLzEXSlPE9ZfCl
0YFQYoG8CbZV6/vl4atIh71COA7aLf7E35/KbjzzQiO7YA40VFrT9Jpe+uQTD90N
ASoT8mGwDYX1hY381yI8GdVHqV8CzgbjDoYi0MNdYjq2xSl9ROiEhJ5MVMYZIFaY
r2Z/OWRsIlstrgRF0g48TC3agn4VPA+epMVAKYona9j2Ye4/V+76gVQFvUo4HAkL
a4IZZ/m1T+nbeLnu8NwwuS8S/ZB/GKTL36p0biD3m6N/jw6ErnUC2nTyGR6Qnjlr
0e/+o/mR0rRLBG2taAlsMYxUfV0Ql9UL5p2cHKaK8yeIwiC9LcreHbzDTd4s6vL9
qK7ECA0/baAndTrdO7l9RaD6+3mY6WnlTO6y41E9CVvqpFMhQNmJjVYg5fD3aSVY
LbV2vHACdsZ9xRUPfEv8fJuqrLIDTcna/jxOrKmiEtyf4dNt6sUIBE246LNpbct7
v+/NmDjm55x4W923V6wLu93WIO0xgJYjsEZv5Vesu7EXGytMMyGgR+d4yN3OXj/U
YhdiyE5xgNqSdVsAlw0mMpxJTzebbwhtWS7N8LCLFoS4Ywo27w4jM3rCj102CXIE
9Iub6kI8JVzz7DVkl+aUY2JF/MsWcPvsnI+YYKcHWTNDkNZVTNMGCjxlN5/tDk62
Lxmzqp7uWRg8R0w8v4pYM29wuWtBylbGLSgwoqZuqojMsgx3fcfkeF3vN3SsNo3v
4ig+VkIoX8AcTJoioLYWU9aG/pdAf71LMYQIIzNfLfLV0oEo02pgwUmG1XV72jMp
MiDSYPg7PAuA4fqBv/ubCp1JnoNOWJ5OyJPJ1yRUmT+R1FMCgA2+gQLGTby+5l6p
e2/pgs6ehRRClg3rv4pWqGUEnrsZJzRv77WKiigvKuIyv16Drdi+Qh+5/rf8Qe8q
qS0whv0AU6AliwAjOTAIjNH37zYMW+TeHYLQZdNEU5AcxviYsIgO5nYWFfElUEHq
fZfK1S5Qt5miL+qlujdBeWUcwMpXQLMmMgavrAwCFdqEBgKzlvNb5YKJ8dNX/IdP
Dhp/S5NshDJ1RdkEKdsYiJfqzB+vABigbxo3MZtYh0Ul7ZPhbvy7ozG+nVK6eiqg
tf62nhUF6RZjunCRlZk0oijzCrZG7ccZjpGMhFsobFCO3j7Wokyiuz+IJcolxy1V
e1m7M2JDY7BtHOnW7X/ZqSL84Ctsz991ng0kbp3soVPup7r1VA3EnQFdmg458EWN
M8d+Y/obaNt9dIsvrArBYGfwgboXXHJJEQ4a2A3r3z4eNv5DfMk0CENN7Uj56QDw
YRm3VCox+6ZPLc7sznoZrJCWxI9JZruv73TWvCUEZ3nKmGYxEBgByWLK8zncDLOa
v/pwPg8sOpbFIIH1fVTs1jivpCfurzGI3JVYPGz334OBsfS04NinjqYQxpkGdl6m
2F3ZCSIc+KxafYEfAYcE0l63/Z4lWOZAqoTzfr6uV6kTpj6DgdDgmGFE87/6SzKy
BDdyIVrMFovHMfGNeqSo+jxKObPId8jBZHUSZGI3n30ZJlaQ1dcuqYWZVXdzYcwD
UQ4w5lYE09o2fxuVTrjT38Lb5Yyl2p7d4lWiPq/tZkmGfeXBUWr8e32hXuhn/6iL
u9edlprFB+k7glTdU851Dji2F9965STURXjW+XFSIRVyTCTzQiMP5SIwOxwBlKhE
Z1X9Nk6uPjO7tOZLs53CM4d+D+VM7BXNOWgwKDJZrxAZSpPEVBYhkvsRSXE7nYsq
jnsRy7LLfMmrcbOSKIMF4bHOjlZlynqzH1AR0zP6LGgMUOv3IFrz59BoZHAWtBIh
vFmoDKExOjglEWmGP8RWplvT1CNWWiFdjtU7ZjU1CUdtxXd+h303ML/rQ64Ee3IP
xTetk+azymwNtUVFmH7mO3DeVNhXaPm0Yxn01t0qS4FWBaVZM6l94IcQEkQRbOuz
KwuuHK8Lp9RQDhETFomxuXBs29BTQs3I9TEKEAyQ8r8wz6u66fePfIqV611XxYNc
qNkFmi755sbNITmnoaV/qfZG0rVsHr7Ba+1FeH32vrv/WfgMB5WlswJhAXhbg6k3
Greb1XKQDbm4XsuB9AanSAc8IfRypfMoijicDT9jbWyXT9F8OMRiWR2GH/WZeIGh
L/nLgzEfcDn/jIKJN7ClhBJthnYqa0iAdpQn9TwT/KZlrLxxAP8dnCNzAH05MRaj
a2vq2Sk9zsYNux8KrHbZdA7lvx0FhterZaQHG7RXS9879AZvIWlv/a6SDjUm9Wxe
4urfSeRTVSz6n8Vz6s3HQlZgP4203P720Y8VbnWxqkm9b7wEPSoJPf6aJuXbyXzD
pQnWnF4IOPN2+aCKc80X2iT2M+eU272sxccp0uJ53UjhM3Pg7ZdLW7fpT9WOn/hc
DYJKek3t7O1HXlwD6tjsXYj+MunMntR33bFM/iShC6ZxK0AgOjsF0miUU00mWJ8i
tP0XGYZI8ftga6jKYVhvXg10h50ZthDGHW4PHJZygYY64Mby7nLN5jV6NOJZX1FN
fWCRmMao2n7rEEk6SIwaMB36F1gV1pEmCIXQAvv/Ieok3KEsSg4MSNKZkok2Gxrs
YWO5Bzw2GjEqLnMTq+ppdc4iY8vDjZPqCFLFIqg8LBjWnEuWNNXIXVVIjEfJ6e6w
VN4D1qx+AwKHlZR8xVpnZ/3579DwUJBehObxP7/ZD1CHDno+ni8mf0TkyZI0kfcJ
RNZfHzKMBowabWVr9QjSSpgoTviSoLwqww72kPhUFnGh7G6Wik6R4RuFTCtz6UDf
ehjHUsdGatBZ5c24Od53X5Wt4CY6Pg/zpRO5xsp6PPPtpw6qdvjYzqWF8na+Bbfv
jm2qitaet2oS8tFWnkq8faAPr+E3V5S/UsaKdfHPgHFB3rJgjEt4EtBuHQ0Uo/LI
AK9DmWRXsJ+BVgaI80s3HpONWobEonn96l+a3OaZJFdANXtXVC14uB4i144eFqB1
8Bkc4HhAhUNcLU7i9NS/p9qAiFVSrRM53+eEdWuXh/lqHdzVPIS98ZVWKc7pVy4w
EYNIaSlH7Wjizdv+noreWNV/z+L0if7lQf0w+aO0XulrVmIr1VOBbnjQsAadg25D
e/Dxe3TTOMS+vlkm/0gA2EJFW5zCUts0SsI7CHjVa1hh7uX/i2bYs3TCp2UmMsma
dMhtxsWJOTx0MO57QOvs//5GVFFfnvqCOSDqL3fxnCY86xY7wUfY3oyZwb5FFS7j
UaI7bYf7jswe0E1lQMcZ+1XHlnzRwVuK9/jXuYdNhWfKuz83SI2htvJ44erytCvr
uihDabVqJKyKdgTMoaUiCMbjJncVQ+zx9IiACxlcuuoDUH9h060UOMO8sfgOQw+q
isu+VWtdskbYJzHloezKO2mjipWVGCK7DvAuyRhUJcR1cqrNpWo1/cva9HKAg87Y
uV5FXm2irj6/3gK00xTZDwfvQb6iwBSNclfpJvzQN0KrHBBldWkhgH8aEBPcR/ZX
qC5SDFyL1AY5+4YAy15B85ZTtWUEF3q3RfWecZXyfjCWouBUQaL/XFvTbuEeFfXo
G/9WgemDhyTFfoF+KLpBUOLr5JPqe3A1wjogEM1U24l+U2gvgcMGhytR5FSAeP3G
sLHgvL4b/g7nrg3pCBrVtySOPBOjZe+nPCCBsKY/32FgcB1n9XveGgz210ZfMC4s
1hyDOzqL71CRzLNH2A0RK7Rlfa5YJS3CUPMLlhGKdhw8td0Ys9GB+QDBYoURLCMY
gCK1E7bOb2p/ku0CcwnMPqGgm+rAyR0TT6i2KLfqlkXC0/mXJZ9bdveQH+mt67d5
DjC5BIesQo+mwICoO++jx6+5nXah0NxKBDrrfDfw1mhThpV7Wl8yUiUlkGGk23ty
qje8Ow0WLNmxl9OUSHQW0NMatsKD9nl/nDKr4Oe1jS+JuYhJv2xnC4vwIFgh8Fpm
XAJK0vy6CGwSultDAjOE2Km0SygyJPsYcw39kuGzuUoGYtlWInHMEyN6tWWzxNXT
XRyrM/WdKKkGsxcC3EerE/X6FmLnGBEidnVTu6m6oMn8xMA6LdLrcBGwas3yUn0u
UC08FItBdF9S5S1NJcBoOFzrNwdzKc7ylSAEawD2higGOTyfi/jBBNMZbmt6lIgH
MtKiElp6M3g8jGlzRbvLH8e++a/czUhGuCBlkddUtfBP4BO04AhzkS7NOmIMezZj
3D9oKhAhDRi09Xad+RYivgKrdIKdNFejqzfEmCMjJIOBosjc5ToWkjKGDds9dLk7
JKACSp276ktqx6uStSzuEFAh6yYAn1R/RdqD4dPKjCm17XVQ5urBsIrO7DIDWtHO
LSEHbGXvh13FLkcHluy37z8FlhJDJkjIcQdXAGVRHhQYOzCnCN239ZxrNezgviKV
LdoAxVMMbHVo0eOMrZKMZR4Rzuoqr2MGP8rI4vRbqSOXQ/gtEnKHFL6yjGUrDlaE
jRR0Yp73w+gQTo2gc1KKNTO/7MezBqzkmZ/vOIxjUoUy42Gt0XoKwVBQysIW6oo2
iZih9f5AweBWslMW+fY4Vyp3MK9MM5t0a0OzU0H2QwzQZ+wahI5DOdjsaS/RGUfG
MLIBU9q3lyF0YQF1dPbp4pP93+X8oxJRI1QR6D5UPyPyh0I/ZTS6zxz0XXAVoqrr
9KL1KFwzlg/MQFhxPxvo8RZttFJSu0CN3pihHB9ScXUBMQfzxdYeOFklIFkNnYGG
DJaK389CkA86dvIeEDCf+tfGLFS9Wc88KBniPAaJZE5mRV+4pRIjnIjUSimkWqPM
3dR7CKykX8RAnSLjBbv+N+UKorijrQ2netHmor7WyKQHxoWflzSePs4uxxjiCb+S
Aj+/eubXyHY4cSDEpPKLIjbqqYvtwjrBt2qsbRnLUPxqsXWJ581tBz8WcXqOcmd3
FuV11/9Nkp5egyf2SgblweDvkOz5wnVNwBaBW4cVxbGtwITqj3vWma21yodnOikD
3ghYQ/ODxySNox1iAApedhVAPg80PwcviDmD7YWdosM4Tj8ZVRffGJ6ehNq5HMzM
jDTeSU8DQ9/v0d/nbRTN5ty1zt4XG2kUuxxbwHm9ZVXg+2AU8hqgzBNVItjijFWj
9nbcGQ5kpPo+f7riZGQMKbAMrtorwQL3NJG8nbsY2dqvd+bR9fIVqElKMNLdBoud
zEgrs1gH78cLCZBisLn1Iiz935eDK+iG4VPSB3saYzEcCnxDZ5FYR8OV3zj4EwRr
7nBk1/5vp6AnLaieJ0vOIo4sgh1mZQ1OGG3Y/+wbMdSZgl/bWBTPmFb4HY9+tGPL
5uLNcwum4SJgMXDCPWu4fD2+hnXfunv24piZwsuzZ7qoATndKRHCuaK5ZyCwSWtp
Na9cPDQkQBjkn+1DGTyTstqcxGgZgLFsyM+UpFKBH+rxRVaUIz8pta6d1LmdQm4y
CcMIZmu6U+mcNpYk7N5DUTP0kodBCEvyJGZvZ8AYkF0QqIpVZAeYq2VY6yX6MoQe
Oo4suAKJjAc8zCeVZRJtFsQ6lgVpLu2wOhf4HdMggK0ww4cGAF2Z2J/yTnGQRB9+
68/hM5E5UFg6uaQ22iJku8NSnOBWRSfvDZOPuL41muAHv+qhu5pgzh8zfSComZUQ
l2kGoLrzb2TJ+OJxN+YiGDOIv/IXtzkbMPZ2qlJD8yY8p01nj0D01QjsSd0Y4Vlk
8i6Dl9M1I0mqyJUdv5NR0al7TZHaUNLLHZGi9TGAxF+7ZOBakjF/JXFmDp7PqY4A
mHMjTPn2ziRbLvIFlX2x4q4d8Bezjl++nsoG4s69tfyA4n2VZ6IE2bKcy7WPj+K1
PsJzAf1Us4a5fSmSzbKrLiMbYzGEJLCxKOy/IXRq9J38h7YHHGwvWfrFGRNaffcz
n7irxRsoLrn9NuEfo2wJdQeaRynS3ue4PiZHRI1bibHwbH+U42kIRvXTWN7peNDE
+HIrlwq1DQUjG9F/D5CvEvG4g/05DQSe5zQoRaLV5uQemhCTpnENKW5hy0NdvsBZ
77yscIvS6hWdRjFVlXYCONanioUgDRR/HB+lGkcWUIU6g+p1W+ALIrPg/wts147/
Zseb+x4fNuCqG201PDM2kIhQacHgBaUO2VxUOIsVbnkDQE3MtC6Hs7+GekDUGTKT
Atu7gHAdNC/KWhcwteWe89ayjJXBT5wKaOaqL+YNd4geFNSrjKvxFd3jX055xkl2
hHgaWHHRnD0QSKxnuY1fVoT6UcvZitOcVm8m5xGSbYuwQ+MMXQIuG7T2yPiZxlEW
fBohEvk0YvxDbmB+gs6j2puCHOTsp7MemW6QVQk+NjagD5IyaUzDs1oEYDLsd2mH
DTmywMe/IpPN7KRF9snFe6GKgRVDl4LY95AWbu8myXLx/o72rStP7D3nrJcbxLrj
OxTM3fntXuEkErFpzQSBq4pSHx1BHEeGcZ5g1ZrNAteTrZ27IJCHLwQ+UR6KhbIP
aCJxEQF7E/P8/bHH8mUXg/j1CxEu1bwY0BgLW9aF4I7czRlPfzQeOKN0ZClCB2to
ihbDrDNOgAm8KR6cVMewJrBQ6iHqAtg4xopHL7N9uDur9Jg2X1aGYInQB+GzHCtH
pvtJx8axPRRKuL7jCauUr/hQbqhy1MIK/4UtmGo1gnLSHLFwrvgguObW/ZOzQH/I
9vD4hrBNo3yrw/JbrHtw11d/zNFAFkrET0M2GGQO+Tx7ElgbhMgS5/uF6C9kr7/E
z0qVUkOVNXvoYN+L3lZAQGdiboIH+0sZ8U1U8eFJTiURs4wBklseoZoRBMP6hL7C
gtYeBf6THPRtK8wP2HvVzlzZ3EPxwNh12QPH6L9i2PInfJxvFpeUTZ/Lhxct6kF9
xlP/TZT7x4vZ1ehprp51BC6fvuVFGx7hGW2rTreq3lZZDUxN3jidhwB/fYq22UHY
PCk5RJbeaiAuWr58tQOVn7PVY64aQGVMFtc4gH5OKPA9vOOkxvIsjBVhJ6RQ/gcV
vvr/h4KdXIWzluDm6DA6+SEeZeaWhMmXrYalfw13nAMwdWfuA8opwHLvzTAQhQw7
fRCOLauELXS1eNJeP9rO6e/XdZBB1w7fZYI3GtPLcKyfY/rUxPBR/9ifdWz6uNSp
cujsY3EIVEirFTlcHqC/6IyTWWdsxUmvoA1QpHvSxeyWZElZ9oICxcFjkLtw3F6r
pGOuTpPCShzZFfycinm6y0Cf4A69fawmigsFE7BGattCCT7JG/+TbhCThkiwGY6O
Iicb17SZHwKfkE4DPx9RV4RT/lCkSE/Ya3I9Td6GCnk7u7XGkLKZr+52Ttzi/NH0
WiVyYaVXU4g+o5T6Ndun1mFMpZjAW1eaWRxvmUhnubYugT4qrVet5uECEqHC1PmQ
s1OAT0cpdJQi1mIQ0uH6FvAqDEDFb+l+2SipIw3NXhHRQvjEOydyPxJpUusA+A9N
i0Alqr1rFojM66QVdC0pO30hoWwrTYtp3YkfAzACHCVBcEf9pScdVxOaNOaOnU6G
YZaG1V8/JvwJtqi/CP0dXUUyyWNCGR6vJpktZDVlHaoQ3wcud1ENA0hWRn4LocaL
vd1xG9c/4WGCt2ykkQSnlyf2rQ5GgA7a2D75WL68QmuBADpTTg2HJycr6Qr5nj/n
K9lWglRQEQKBiPYt2xyIMmFvn18rUlGqnz2ulIXYlT/989iyaBf7FVKWb3Oee0oe
Bs4pWkhQehDOOj+qasFo6p8llXHjcWPtE1kUPni4u0/RsXrt/4PrzmB78pwWemlY
dDdVda1iPWAK3NNt19WRFhI/ALTxGNPC9+g4yWIkqM8lBqN+2yl6gQIHsPopBGlt
XjdtRB3SdokSZvQNefgT+2AIJF2POiQom1AtPevAGwtnkTKvXOFDAtasLhmHnVrF
GDmmzQXUofDZQODUOnLY+pQqFZV4Kh1WKpkN4x+0JcnXy6GQSJRq+JsgHQXZW6fl
VypLddVg3Ga9mxZ5EGrUxB7qwRM/H9pBt863A9nGx645ZRgAK7UTZ0APOp8Nfl6j
RAWH4XFyo0KGGYOUDUjZWCew2Wr1j6BY1Fbnbaa0rsTveeBwPn2ElAgG55oX3Kb6
3E5Oj9N0u6om83jK3ue3Ao1sURidm8ZlpboW2BgR20AUZbyEy10ejBhjfAL58G9u
NnkclW9SXAqRX2RL2UlUtK94cw4hWw+qk+UvVaq0S2239caQAzWv4i+MemnLf33P
G8bfOaMubxucySx0eekK8+DsY/gbGrxi+Zl7X1UkiuuAPY+PNfEMR4XAFCb1iwMx
zsY9/VdP62IaapBY8GrGGZJGZ4xWCuIMlPrX0GWWeallfZfQ9u9XRewqEJq7e7fw
EiLn47dHk+mcTS3l1Ibwk9ZYMZbSHAak90gEVyYLOCAw1NzH7bnSYPjbEcQ12cdm
a2F6G2dfd6QUKNVeBcquzQfxs/cwu7XOdyIt5E8z5k143YhNt0b9ZDzrigdu1WPT
B1elrOdeG/zOuzO9cYILWWpZs8fFyRD2fyHDVcuNOAdyNLMyhzRAuT42s0vuntF1
JIlpst1b/S/Y9rNleJuxxYcIjUfTbNZTBRlDz/ogBu6jBf6dHsTDYoOFbKLrimyL
Lz/W5RRQ07wkREUox5lWebT8Y/DhYV5Yxt9bVXf/QtN0DV05ziFW4lKrhg+vCkhe
25jJoGIyCe8+EPufaAq1BsEUJBzg6Po4CuwWw0DUYPLzZkyXq9NQ008u+V8Wrod8
UKGr8oLqBT9HSO/KDMM5T1J5xOqNFPV7F3ZVOWI2EQEk90Gji1dIIPbv/zY4bUlF
naXtJXDfedj+RELCEceEahezqkZFCUbTJtm3Z69U0Z1+YJvspufWVyXiXxk5E2Wt
mLU8/QAyj7fB0bIOqnnK2jzZ7MDgXnFq72pAAukZO8gO/0Tq9JXG2uG9pSirV97L
OnWaJ/B02Y/Gff1C+WjiFV7dXJnrtGfDNQhYd7j7h03fUiJi/GkYqwRKz6gw+7vH
v9xSMvQlqSNmeOKnjQigro6qoJApHc3Mi9ITJ+QWwS/mMxhjjgNu2y2IvSY3Bjie
tQoHyJwszRHSyprbjgDubNuywEEdi5gRWpM+N/oFZWYAG/3uzM3OQxvJFn6xkUJf
dccVecOQ70rh5ApXUbN4XUhzicgTv1xJfuELqJLPlFjA/Nycz0LzTamntP7VcXMA
CTEZnWZ3r1v4sbTPXQIyovHpB7Yd51KysQHaujFvA4ZpdPaXts3TAr7CWiyZMbSs
hLkpCAV1v93Zm01SSZw1TMvIIxbJwMYMFwPY0UtKd5/dLHcNHhrY5t0N0hW4vwDl
z5hH5jmTvbbSPxRMRi2XMo2pthUkY0V+abx3X4jMM3SVKwsDISA8DdLioeGYYSXL
B/lH8U7qOARCn2Q6G/TMd+3XKZ0AXa3Bj2V+UBpT0t4oo/m1Hi/K0SP4gxYqo5TG
Y8uD0QOaYB6CMC/VQKAnQWKwU0g7jQ+hsSxYUTHDIUt7ZlRBcP75+OXFdrW5knWo
O+6Xt5OjIc6VNO1p3yIg1cDuiSWE2PyPduxx29fo7P6EPyS4PXyU8ylBUnVkC8/u
6lbYQtn2xQ6p5ushZwYnV/gekjyPIN9eCVYDZ+tRyiCafZhfoogkTq2cxIGw9ZbP
a2JfpkQWoKZnO2HswoxGAUlqM3YMKMkn968TFyD5GBsrPnpGp1gdH0N/JbCA6i/6
5QfZwqeY+4A4EzUeF1x8QFUzQGwttOLQ4Kk3XQAUMUEfNeGe1GkprbUzvj3dBbOn
10IGPAe8XVrBwF/56OmcHX4qwq1uWvEeWal7zoM1fyolH+wH3Sz8lsduv7ckrxdt
jTt9z6wkf1vAJfFHjfqVHUrTanZOhlDHZxdB4FdB2c+gkUJDdv7VfJEsm5wHl0kj
ScLZEXf/JFH5K4hJOottaDr5nygsUNoN28LDvjVjQ8IegKJxnSundObXVuoU4Xam
yiL+Vngt1SNv7etZM2MbfbKbY8G3OvWG9OxKHsR5qyOLvIoGJ0EYaqDe6vxTm4pc
v+tmbBFZM7YjqmUM7o/H2YurfRVElPL1Rou1BDTbmFpY5uKofMsjLRev7t8EGkmB
9I/QbV7o1j/DNmti31PQAtQfWou32C1TtKHPUKszbeHSa0mi9vYryg+ySwxyCHez
+zpgspniVxehM2gaWf+Aphp/jUDfga7+1WCXaqoGwFnKadGVFUAetx/TUqclLAnc
9J6VpcoXuxG0UVH7p9DabiM2fhmnwAzbdFGBueG65zRYyqNigiKkuim5F/afssjM
KqqVQxA3aUpNHpNqIZtPdnVPG7N3E2wyYh2cqJlTG9BsVwMDaH9O6M+PzKOIDGdg
vv5bS48GLZS9GGEnb2ZHea8AF0+90yxm6AGAsG5sqBPA0BC2cqyWzV8ucRnrdPs+
Qb+6C2tV9wIA3/0XnrbKa8PnlQmzYPKmOXuwhCfWAkn00/JUHvodSOurAfINH6DU
u9ivieeE9qWthrnKcG4UjpFTYQtVifHXfqWfdGxv32YDV5BoVwbxFT8p2YJAoxxE
YkOLMbfmKffmVhOXjbDpW3DcrcljBAecHwDneJ5BT8Rbu7XAngEka1yle+eiiNcz
ZjGlGHVB6DZmiSk0a8T5sGpIRl+1TcqWAd0+zt6t+mhc5gmt13f7gYaB25iDMs6N
KbZWnF0WrJ4LytBEl+24SuiTq7ee/ldgvfQXtcNucsRbRaNAmth34VZFPu3gNynn
xa5OtaWNluyxDPmtzqoU3xcerErdUnBpLqLMT3of/H3KZypMfq+Ke9TCSC0Aa+pZ
9ZmWwAGIT9vw6Q796j0itMb5AL6YT6oGbI2lYpVrc0jAxHGhzL6QF+UKRvOawway
3xFio6QxNQm4UIJCVOsmtoRbBEGcvBDkiCx4CG8to15ydWjkNeQCAVnKrwrIw+ua
yaH4lQxaBcVToBUXzrBAVltFkPwgLw5WjWuM4NgWh2JiauGK5BtteesngXCbW560
r2KliAkBEWKF9pAy2+lipmoe3MwKtwVidwWiz+d1fBQKpqS1UgeTYMg4FtQ78+gC
Fcu0Ds7kw6dBM6iOO0vb1MPTdx48Aro0ZX8itccVPZ0drhZga2VzwA0Z4J38FjGf
XiZUJbRK49E9l42Y4d0scJF+6efmeWBSqlPBbkk6pmnoXF8DL1a/BNnZGF6ecikl
LjusZSaO+5aZ3SMW4dFjmD4hNtg7tMBndS5bnXin0HUwFyv//Hyf9GNjDZxoJ056
Tab8211ZTfJ4nHhjcy0rkZYhcSxG5QRHnh6iTW89O8OHFtPa2lcRihV7Nnq38jgS
88ukWLdBtYxt6yL7r47JwPWGDc863ISb7Omgmujx2WJVMLW8EJ/a46pvN5OOXAM1
s9MwSYZI0xc/WoLT6EDnwFk8qGMM2kWBaMYTHu34CguSIxQTuGKHYpmB0aq8rU+I
lE3Z9SeR7St1xEFh3HDE2qrGMY7QQnVXhQNoFkZfz4UOe+iOnYp3xcTOPBL2MD5C
h4lYb6CsYLCgBA/cqzBgbCov1oLdH02AI6li+aIQvGsh8v+T7FX2HYlx6DzJV6UR
MQzj/0KkEAXF4GAvNg0e5alRc75MnSbdlBDrtBjEnM+Z9rNWex/YznzbDTJ3rejC
q9QZJStFTXAgNuII2t08MnUVD/kNeKDqA12yy7ER07F0xWEj/3wOKHYDn5gQ/kI4
hfzh8G0L2hx5xFEa1LmOp+WY21XtW1/vw8Xbt7dqND0PGq6NWEk2PVLv6fcYYEG7
g69iMZi5htmNfkL+ESNGOTrWA34eiujm+TJGEWBEZR3lstWOtdv3b26IGbjM+B/j
eUwFTnSqs3Nqv3dsGubMdEDkuSs6v8hvTSZeOxjNKyT0GdI+LVvo6AeD0s16FooC
Qv9itgTS0OzGEkwTtuD1f+IVoA9vnohBmjnoXHlXxiks0htISQmg0ObzK494JenX
feyuxXON5hm0jVDaQb7dm2q1tybjPbo/8NLgBqtZ1JJzlsYNRlZxFPeENtUeQfXM
n7T4ixls0SOI6JqWSdrYlj28fvAmnwQ1I1PHnmxpvhBXg1LADhgsZ6S2UzlLbCqY
xSNgLxPGQfCOoh/poHufzsDdX4kaYyAmlhKRedjC7tGEsTjLioFalyWyd1S5rWKl
sy8unJfTaIcs3fwebePbwKJfxq8fBX7YenH46mtsBVj+T0tfZezmHB1gdfd2Ae0L
N8fJwMpWrBmh7MF5OjVudbaKUHbVpWyepJ2b2jvJGtA9HOM7/l8MSG8fX5pmaBBT
cLmHtI2SuU38HZ3GMFmcnXnharw8uSmPqDav7uEvd0ExdQwzqM1nbxAJ+mbz5MR8
Cu3R59bFTxKK1+PtU2nkjB0LCdk0CqwLxep/nbUTCR3sgZmS0Fy1o5liqH8/uUso
X6KUAZjpf9nBJ9/0qctT+MKEzABeslQsgqk7ivc99QbEBCiVF1EdQJe+OdMjK18w
ZSTJgQl/uH5RpXirJAUISBllvbEJJrenJO8Um6iJPVlUFYymm5xxdxDiRlxSNFHH
0LDWyIfr5PLZNRUtW0+VETBp4Ckp2trzYgb9DRXPL2ntFEvycUm/39OxZjm4b/iy
EPCDwTpcu9ay5r0BalDk5x5F6myI4armiGTNIKKpKyaxgvPSFCORTFDMpBSwb9zD
w2Tbafg25ph1EpiikG/JsS5+qY5pCeoNSBI+b6gLhS4mubEK3Pv/iWDDLn66+zVi
ZgNF7Q7xKLDvroGlWG8NUexqd7MGoZKTwQWYkwSJHSuzz27Fp0Xew8QNXwC7dFFm
CaliUjTYi8CmTdMQLvN/S/UaQbRx9u1gPk8IVReThaJZ8p9O/mIM34iejn1Ya+8z
Vi8ibpvIazIU0GKQVR+695rKvLZeb3vi9Q1aI8PS65Dym1LzqhLYCbOQ2KxhB6OW
y22OoHhmxx9AF9bMPU+sdzuSY6zMJ2Vb8Fpq+/zaOWQeTFFLkfNSpOScT6qcQ2/u
5B1cnGHNqelPmJ7OBCf3qrvFeCyVuj9eseOIrviKoOPq/Xfyblv+ugPOKAZ9WACh
/mZTBPB83nAOw/JyyPsI29bG93w5ZjaI08i0YfbNMFSJyAx5vtcLOEomRuw1XuwD
/vpQEVd/L97icJavdf0YFit9+tww8iAQixqwiI0Bbx0Wq8y65M1hwD7BidirMkNd
faPxxbRYROtvUaIFdDGP/vzms1V18LmrbxVTIrjxD0WdKey35iwBtS1f4UhOOIsK
lFPHodcAY6Kt8wTasrA7nIGCRMHT3/3z1o/f33vYdbuS30rGW1KjfiA2aJZqlATR
S81CUFa3wTSq+DjKTeWFub0rKu66zbo/STUmjnD8A+w24VPTXc0btm6PyU+YIu8M
rJehYnq7q8T49tM/CK5FTbMIlyf99Xg4hiBtVuq3XL9jY1DOlW9ONaKBxbduHlAF
RDTFNqKVJHhx5lLMidZzg8i+SqNSMHYoJBYGl9gG+vLHZhMlp8ltt3+yfeAQTmhU
D1Y8Ddb2dzwFlDpp+aW/LxV/tuAw3VpPJZXu34E1f3YUHlKMOLeQrrTPSgQ8iqTN
Q8IcQg8px34O9HEDXHjQE/HuMNYr4YE7cwM/vpL/41ZGBX9mHbbKJjAOylvXzT4R
wrNh211XPS3sEXCXJepl2JPwOhuqJz03zltyRJT/SrGJ4ONpKU54QvWSRa6KIqD9
1GpqS4Evq62Iyp2gOlI+8Zn0x7lxGMTU+qNPvuOdlXRLGP60Cb1RLs0pTrWC9+vL
uioPr8Pvpcz3ZNPPip1q/qjT73d6X1aO2dJqtm1H/RI/B0cK0prgxNX7a2xE9Qqf
8nkag4MTFvtf7UgzHdAAoi8AkWG2U717bSKVtBiwIxs2wvdwhFRjh2KigP4vRu3J
RKJJHnDKX4agrql5oTBsdFfEcyD7TjLAXwBavuvRnyOLVX8GQHDvIAOnctjs6DiK
E/3YDR/i+p7JS8C7hgi6qY7GjIbHrugXLUvHGyMtu9q7rldDWphBaDAkBa8woIiR
tSMclEcoq5EN13vrN24Kl29fYOrwVx30aOe0wE0Z32gD5qiQQeOZSd5H1SwNQ86V
5snL6c6vfO4pQ5T66rDsa0/AWv2jmnfYnTXsFehMOkVYPXPWeSkZ5kO1CdVwhODK
Js4HKWJH6bku9Qe84A8WqcpTB7dwk7zVg4vfPXJCPYNZxcG9hngeRz6SF79KYaWt
TzFTf4jO0YHiB8TqqLsiSTeC2LscEFb/f8a0FKJISqGsOjhtHBhSs+J9I6zaVhfp
+Fi2/6hHbO+LlfFTGUrP3DQ1OYSgYfpR3VvQbzKKCYOn0kU/nnB4i0rH/C6rLlqU
BA8kH8hPpqLu85nR1YHb4k8tBMK5Z5LmY40eGQpBsTa50LsxkQfpAShfV6mBv9ob
vei/7HnxdbdYNX2aghgP4yBfQdCCPzeePtXC6VxNNKlXUoq8R79U5KduLcAkgd0A
V5vdfbL4t4trImz28R+yUKJWogrIRbrmF/oTk9xOOu8uUNisP9zEjq23iiaMCAtz
WVXznpLTAbdpgd5ZikTTDrk6f9fDwNtSFyOenDq/ItV7syAFbZds/jSXl4RAZgTk
YuomjyEqn/KP+hf/V+Japgb4YAcRXlOSy2OuRphwrF390eIj+XBO6p6ukQc0zL5Z
YIdi0VnE61keA5DnQGJtvp7j5v7GdJD2rL0BJHWP0OD6AW1yxuTQnJuNd0ltfDOU
YoLgmKW5KDScM+LLcnGdAk3rv7+5LGlGBM8K0oB7pz2x4Po6IblYe8Ay6RYARlTn
eQIpykK4szEawA+m16kiwnr1hxgLVlf8iil1vB3v3lxsh7CAMDHkza7CC6GqdW3Y
pC2mkzp3MhIxKgt4T/8Z0mXBG/Uc11pdUPXBy+czASv2dXF4jv+wu0xcECCHs4+R
579GMQES7TiZkH41iT76Y/yMZaDy4R0f7iXKVRhKGAIHLeJZ4R2KrA2xAh8kVmvL
brcZtydd1nbRswPSpa9ZhriglbngCkCQa9nqVbC2WGsFzaN4aIQwFKb6+PdG/O5D
PiIJeQHGMYOT7ZttuM3Bx3HJwxbz3UVJSQLv6m8QH7s1bdn7GPW+AwOZ8+vDlDCN
k3ilbwZz8YUGi7lVsYSPjT0K4wtKUo1Dgdb7qJ+Q6ycdgQo3ls9BvpuUhxAGiFdZ
gtMwaoNIKR3RveuvHJJtTp7AEUd+OtvYl8IyjY5btuQcqc9dxDcB6ggz3RTxJF5u
4N42XI9s7uQnrVWVsMNFXcE0w6wCpc9Kcg7u9CIm/8Qy8V9f0P07wKABsK6Fislw
sfCcV8qB5UMgcfrYnzC34GjSNM6cYVcI5zFYbyHPGCNkAqDJYlwQB1we7D7xaKHW
KJCNBut+N/zlQ+PxEaUn/n4A06GS7QmX4sRak5c/aeNB6DjmOz+bfhXqQ3v0OGFD
kl+mkZR0CrFeP3a1ldm79ekV78ybNU3AuO2d/PzkIPSgqET8nod/s9KRNMJuoXQ6
sU0aeN5Pddl8UUnTNFU4iWnoG6fb27vM8HjQtDKurkeD2mWTNb949sazjj1ypBip
ZSEfw8+S6dy1RXziR8C05y2fePiISA0suo3NMYXAeR5FRZMEwzE+kXuNf0gQS+w6
/a+4lrSWamExCkSOWBsavkG8VpkOK/G8WeoaW/amHN2XpqGsAb2UwVQn3BCxL5NO
UUsi2OvPKyQK4ElFx6GpBd35S8jz74W/r6hil7mVTR1xjA6/tvhi7LDwsvnBt39D
K0P38TCnm12eIp433mphuZCfFD80A4wYZyLMT+2sejDv0pBw66M9yK+U9aqvD8PU
96uuw6WpiKRjupnlA2ir8/vWW939utsqlc43zLGNHDwQR9wzt9LUzum5bLCwIdJg
bQIpnxhA2oP2ZLp5ywBpzXSRE0SXwQh0CSxyMAhErmzVS2IrJSMlomTpw9gICVXd
It7Dl77W4egIk9BXsFMtguT4Rz529Qhehncgyjp+2AP7tF3SqyO/MFSTO9ikl1q1
CGpH5dUx1nEMQpOwxQfl+CdQXAZzs/zl/Ylh72KXRueRSVMhJc54ti/3/LD9t+x4
dgZ9rIAVMCbZPoT78eLCbLsmIfy8Y+8NPPZwtJpZS/af1ove2PFLpgPhmm+66ya8
xCg9wQkyBFi3Fqg5TXVENOxmkfUIYnY0M0iJG9S036RG9uSMog5ed5VyZdGB7RL4
FvMHJ/a8L65u+BcVVq0WUtBG20/KRiWPziNu4xZwEhDEPt/MazKUau+umMrcMWzQ
PM6iCS2ZVwgX39lpznt6m8V4GrNP2dowyKnZ/215BMjEkqKgpAxRLqVZuOG1j5Q5
PvIn3tHsfe8kpMiRSjBwBp7fwOzWfi8tmCTq+cqntDF9pW7gVzkZLEwXI0Wt58aq
kjk4MaiaAA946zNQMtXRdpEtLrzPhqaieboyBwhQRnYBsQ95xpa0EisEA8+eNw4h
BLCqRa2Nlwrin94XtqC/CyaJWjYncG4XBi3MihqtHgrnf2nV/rBWP+8u5+zL3jsU
b8+f/scDdqyank+l3THyAmzf5U566GqJhY+iDVOHzvNM0SlYtHcRb9+89XscSAEe
MzaxrOLU8r5byk0wmhtBM55aC//mCZfg8K8jKbH8d0D5+5IhUVkvgxTomekFzwwJ
3qmHCOdorPL9RTnYvsZokFjgYwE3GzWTLfr6s8wqFdG1/1mweaF6ohZ+M1OUjB1X
nPKzQ6nOCKpLq4ZelyLiZk8PTKh26ehBklULpE4SFTVgOT1a5Jtr/PmlIZVkcsJf
L/jLvW7PCegFkLCivfdR33Hmd5St+qTsjYTnP9ZkinDEEZeQMCuJgxTRQuo52E8R
GZE5GcR4nulKXpUXtKJ5YPM3q5nLHdc/Kms4CY+L8iI43GdxiYhdigKM6dC/i9ik
4KmWo9Vf3XKxj79BURwunFS7QesK4yIKPRgz477Rr6n25NumAjy6bPCCbUFyjmf7
MfeI1ZIfZlJR8Ptso1tgg79KnnORmKGBc03YjY8EDb/uYVAkpFeZqRpiLadOl+ZE
+giz5qyuwgZx7zmpsNPVO/FDKc4uiTlu6Nnr3WDgQohMtNi7Se+3bIwDlzoAEpFT
UuW9K51AukHyRsWOtzDtYEFvybTH8OJdzviIkI+BA006heS5PXzvW6DxQqMW98sf
LdmAF5gV3mBSQ2jPZr3NDCl6B2Yyc0J9yzTG165Hz4xdNNtaolKP21vVTMOsl/xx
Bfkbwd414+fJF2C6HnoHLNFziRANLI5+96ngyC3/NbhxpcfDT/HnbjrStusnAuTE
gZgPM5rHz0BnOYnfhv3sFowux6kVJHGzB3OsguShCxSBqTxRg7Ez7IrYCM0KQTkp
KjR7XBIpDPhrYv7EehhNGZSdH/9OnjCMyU0WisoI2L8nIFsKoshEogLN7JbL0LVV
GU0RI9CLf91vhowtVvhtf8iNPlZVA48slCX8I8K9RhsJzYAyOiq+cFHbwf9fmdyN
wPegzC470gzrUj5/xzhOMUuYtd5mDW7xAJKVxYuIc3csJWVV4ZhCq+/yX96vhZ2M
G1QwjcJo5eY4t/ZWGnkKM3+IOHG5i7MElWWv0PN52sczct0r0SsgheSgrfqPl8lR
4Rt89lCGGyACIPcgX7Ka6Tm4xK0WRJR+oCpM6qhGrGYr14UpSriNrMlZVxashtDB
gRDeAF5Q8dKjZf92Yy7akylWhRhct/oA0741jhC25RyESVzg+8Ng1E1RT7J9mUIm
xVzwDQ6Qk8smojHXP8o4ALOQyKZ/tokWH9JSyvESEMxTqvoBIut1rOWUI78xD9bs
EckA/T12s8UoifSZCFiUobdy5cQtFvk8DrvN/nj0Mvn9ldesebLHZLtEt+HCQMxY
MHf+tDlI4cOgVCUWNW+rW915XGQla7UJxgs6ZdVAP7uXcfR8q7SkI/5Yy5ykeKI0
A0Rz5gNo7FsaivMbzl9e6YBo+G05+IRuLiKT+qLJYBOwxoopSt+ZN1qhSr0/1+ER
XedbldjkdJ2RG2q22+Y5c+TyRM6hPSrYsnpNFAmpCIEfvpoekAvlerKyKlkEMTMD
bagaw9qMrqE2KOR6QV+7grZkSTi8bJyBpyZCWXprtjx1fz8GZA0HCNK8yJtUktAP
sf3L1fRgtW9ynuXwk7Z46XFAQM1D9A7ze3ZZ/jJigwx7op2FeM0DpoZDtO5yPBFS
hxSKtAqWys1QSLtUALPPJfRjJS2eHX5f/efjfBbsKS+RshVxZ3oUdL3Es7oWIDIZ
4flUrsl4+eIiL4y2cSiQbhwHRweJ5IH6ZlZpWKGEZ5WpnO/Xa6KGkBpcuWqyR6dj
xCfSjZl/tMRTRhh+0KngjiwRn/b6FuXcocR7jkEN7Vl8+QM5BuHPQexCK5K3z3Vi
rjcGAGZa8lWZ0Hg9O6CeV6idZiOWLeMk5YtPsttSMUSqTTgUTk6QDsUMvt/kmfdI
aw6RQZTkmVw0VvTI46dilBFCvn/iPKjVVxOLoL/hzYZvoDdBAv2rHo0QlqFTdB6I
UrKRncuvslJHkYoJRTvq+pebP5ciME+7YPj6e5bSf5IEeafsatkCebqvcbx65DLP
QDcIzvxtZ3EuBPnKoUqP/F7R8LhvOB4IEAruqNUgJzuwW3gGSXQ6DslxRLhWM6QM
oaRIrMu2g4x8rStl6J7kLHDcyk2Wps2u8VzHV9dqtGdF8iJfjAq8wj4ODLIioVoG
2OrITXrlGig7QCd2oZ9W5tmG9lhAB91qr8chvCfq9RIiLrFPceF+JDC/TLdHHBBL
dbCuVYJiIbsrRv+PZX8CSI7wyNFAy1QLn3MHK7JNZWta+RsbXwOSQNRvdtuxwd/A
lwFfAoP6sxGhchz/En4U0xf/Hee4Ciy6u3GAthO6KiWcmnmd+BdMkWGKoxcMsN2W
2bLJ50Mc07jbDUsOh8yNDm1w4DN6DUtS6O1baa+r9g4CS4Uo0fxeoGBj4sf1uIP7
vQRbw5YwHcGC0Y0yhsbPOhUYuCd89Wnf0wj4OF0pCfV9Rx1JZCFdmJfgIh1u3uK/
YRuZEL3pOB5XVDjqs0tx25bQCoMpX7kAgBjulV7TNAbshKX4XlwIWkGz2uddHdYi
w4AF+aBx5oA5wl8pM0xN20h+3PaSif5l1cnyQhBf16DOHKBHBAYGClbsOK2w8e88
mjtUUuCQkEearC+cK7595ygSv9n6V1IWaRR2l0as8Gw53szd0aCHDQ4tDk5c94DV
SrWjroIH72nhpHEGhfnffgA+oQfW7g7GdBg2XUc2Nn1x6bkQeiu6u/MIWJvd6Uur
RvR5Re28cUm87GeUpqK1Oou+nVKiTDOr6R52lKkjfq3QYLhA9GlQLVDYixIiL82w
Si6abzzNPkzhIRDq2dAf8cw6anlRzb5EyEBCgqpdwGQfhAyz58xh0Q+unkEkfaNX
kE5NU+0Os0QFgdKmfQ9eeHxALfmgWBKM4TyDS4kTdlxtKhJhxSZMGDHThU/Ylvhz
YBxdi0rihVZ7/0M5KGkBH7tQN/ob3CfLcljbOR5TPac1pyTpt4R9NdqpjgTUfgqX
ePbkleUiXk0D5fzTKtU0APYslxzq7ELqqZrSG4yu5WFakGHKFl3HLKaID7qNtOEQ
pw4+ifdR78WwMjRmpjJQPFQX5FVTx7cY/ChFFG+aluaEqWb5Uamv94iouyClwFrU
EUd0zbsJ1zlzaMpNMHaoyR9lbVkTBEhvfxFBhs3eKrpzr/Gi3UI1RoNQMO6CNq/r
UCwaQS63i+Ntu46za6qvmkrkd8Wihrnee8dfppO0L0jh6RyZcMJ57p1tQEhht5FI
nQkS/2iLf5nx32jgm1bVOXCtVekE16Qi8ZneSo42QBJuvYMYvXCkF7CAEI1lWGTb
jZRoNwiheS63pUnmNPwqgtNe65BKN4OOnf6tt/qWFsOruPw6AP6PydJM0cwk0s1c
jlos/WcYcFUcdDWcm8E7BDAl2312nQPlmsdS0TgXfe33lA4f6suEhR7kRQPyhVSt
KzvbXJnMaeAEGQ9VNsiIAzTUHbgXpsa2duMa64T4dFHQgCr48QfC+BE8RW5dacUo
SL9byQD3cSgjrDVeYt7BeD6Dg/M9UXItBaToSPYFblfYtTWiPh5lyHxaLGumftNj
tC73j2qJ0tiVfMNrXRHRYbDUOIxY3pMm0KV/lVPai3qbSb2JHcLakdE2tFOHrCDV
jClFRZYUw1POXYyiBuDYd0rerfRSoI6zfvYbd62txLF+9okON2d4XRQDtTP5Gpok
F2ROB+29Z98vgit8kqjCwFq1llUDTR9V88RJBFNwZwPYcl/bTJHD4x0AnQMYvZ2w
oFqFOBR3/f4qlYUdsotQPKbGeinjJGSYKVv3kOoY1ZjeCdikBZO4tKCgFnPyv8yw
R56xNQ6sDMZOc7xGRtWN0JDqM1KsTcS5MmpNKnP4EGOzMvBiQeH0GQMBQt6V6Be3
o3oRkCrpkKPmaQeCglbVLAzgfBhBqkJxd1sMyrQmj2yszkVqki2KiNyHmnXjX/MB
WgWUUWPzrFlt1KgP60klRjDRSDhU6meZntUL04N5DxezlXbTa9UCGfAvGnvScGro
wF/kPGN/EsS1DfW1ofsskw5spZzWpR1bKTUxoUqZafNu9Ptja1/fQH3z7M05Sr2F
5xB6sifqer/3rlShsJNejbxl9XavLtzOVr9B+kwClykcKRgQhm3F3O2J7F/t2Jyl
WZ80MmC9WaugpTAg2nPQ+ThbW/M5d+qylkJMEKKBdJkc9ZoXMl+dMKSbvdTwkhS5
r3IUrhSk5FZPgJv00jR0KZusa/ZPBzWqK5oJ+AdabfqrFHsKCnRUqyh0wS3kBZ+i
tCNIeaUekdoZo4P8eh6rUR8bJtpkPDREEc46/UX8+4Twm2oikOQ1L39bkJcosLH8
M8ByP+r4Uz+IDMveWHBnKr1smlHLjK6GHuR7xrhX/+RH3TzOP0v6tJOmTCluxYhY
htnW87HUUR/a373JxyGhcupOcH+XSO7F2dlNtegUeWWSg9+WblrCzqyvhekiDkrB
o4PaOslNWMKhJIPYoayKVqVz3mYfLoEZHrkux1cUOXx3SoOkj8KaheGE0OUyrhyL
nczsDlw77Z43i9+WgiH5C+dG0DsoKnKd4GA4h/GBbINihTiBxmL0jqHboj/oGl73
oBm70srihVG7HndIC2Gc1t02XELCytGOa7BtUgxRV3aTGZ7OLXyN+l3aHGBFpMLa
xEbafPkjXDAOSStWN2+DwtdXXgSUPqW1LG69TUtfui6N0U/wS5cmzkNFsysTFrqn
RFYstNiHgxxrLjhLSPUvCIy/UvVJvnvnf/dWPaU7bPIZxq9zY2ibJURqdKojo+Hr
HSMFZSGxI/VR+UvRRhDDnt+CNKGsKwBf5abimYDzFbWLEJL9odmcT2E7vhBat7DZ
t2rygL57h0iKGJ+zs5IvB7r/nqSlNTWZBoqN39QvE96bTFgNyMInQp5k4FsSGQmn
9Fy9G6GyS8A4sb4kYgcz+ehfucZjC9BOqB1K/8cPVFcU2117PUrtFSdJ7zOMquKO
jIOcXsLvbW8/D1QtV5c0BFtMsmvrkK6O3ayxZpbS4DCw9dMJpFLgoMMh2lqOG6AX
5VuQxHg8PVjf1ct1WJ89WVDa/wV1Een+v8DknhoKjgK+xbaEFRV0KPyIeYVfMn7y
2m0n6n6ol3T3ZMJzPYBulgOn6rfGNgdwR2Qd9rlBYDT5zjet3pW6KSVXOblcLlXJ
V8qZca7evUzytJPP+kWReLwkHSN8hoGnHE5X1iir03sLx6g2m6ToNLjX7Tat7JEC
iFuAg/eNZQv/ugaArTZN8Xt0DYtGTcUh05cw3mCVw2ACgfdGKf0eY0TZGOm4J/qd
A1OwaAdhvvGevqgj8mKnV2IsqxE7ErWa+piOjPHH6JKYkYK2ZZoOv0eE+1gKSH2F
I4O1693NVK8kohXa1WYbCRS4V1qT08UwmB+c/qNgSboaaGNvFD5j3Mzu/uT68Avb
wpqfUXrj91ZZhEi4eQX7XNViDDMsEZGhXFaeRWfWDPKuE3bEwpeUB6QPPtbqXjnf
Q2sYSYCOllnmbnzLB3MUmRiTV4rdvWZxSExAysHvBJZfyw18QOjcNF5zUo2DW784
8M/d0ZG15QiRu/ysl27vPvVNMlYGPAepbpW9TXs+HMxO7xOkfIAZNIW6AtmvNPAA
XnF9gc9j/xufgzJHG17/QXByDpUQiLq+K8KPqHZBSZs5uX1wxr+m+1nQS58UYBI6
0PH7pMCsnJi8Q9Ff6lZbmXyYXbjLjaPcjT7keiD3wAysi9oLbJnjy/KbHxCDj4tE
+n9WJbvOqwSJyXcH3v3na2MOUiH0fGExsmp577QgQZdCe+QrSMR7Q4qatbLngbU1
7r5RuZkxPcdd7VO96BGEevQ2MBZiHXh8+xPpjaK2IJcywY81sx/EX/mYz0hbAURx
AgvkuBxEzHV6L6BLRnxlLdFaqNpeaiG93kYBofO9tXutqEeOOJeIunlxDYHAHK8b
rQRBZoAVK73/aCWtO5YCygaiGOz7JAAiLdzkSq+LLTbg0Vu7hibSF6Fu5QM1is9I
+g6itvfunLrTUkcHV0H2aILofdm6c4v7iKPxPZAcFiSD0ajfWVuWTlOEN3AN9BlH
/ijGY6VPv63t7ZcY7/PILhaIhqjO4thLV4kIo2nOTJKDc0MCm1EQ62ylwRLc5eYp
B0XIeN/x0+chSuZMvqgGN3IkYy0U3uuYf8JDUXzOKBITeP2CfNY82f7nxhRo6tRR
yc3EH9RxAJaLaf4e9HQGCdYBendzE2EyiolU/yFSdbxeGbF5EAGXKVDM4+KvUVJ0
yGlJiQxUD7Sr/n+8LVTrNI7rorloDSsJ2eHtqPumvK5v/aqKzYigsZovVw5Y/txv
CfF3Yp3XzzI3x/TkHxncy46pji0lMUlwee4mAFHch0qb9FGZPs36AQfotBzzjO5L
uUc6uxg1EjD9EahOux/M4ezNv+jbgZbAJiOZFCyHW9I8ObH1yA2qYnI/8q9Qm77B
22dZtzQknCfv0yWnx0Ypu350loPmiPA9/oK+Xbb6pt+MPAaqsspwzaHUIi+BVjF9
Jk1RKDScMB7VDvNsrC4lyyUI0G1s0R3FaDf2yydWk3TTcAYZxwAbDqYgcILG0CH7
9R4BE2GBKcDuAkpkdlkVQG98T7ORfIOdsVklgxBCUtz0MvH779m5szO60iVxgHuW
suih/Dts5FNzDrlkS/NGovEfC7mMmvx4KaMuQqcpWK6Ev0+TBvWRWLrmP6ozVkIT
XhVRdrf0I6oKvyKOx5JG5aC8ahcmOSLYnQP3WAAT4jQeXCR2Kda+67WXZPfzmu3z
zvjVIqUHr1o4x/foEGzPp2aAVzedT2qqEqPpDAM4+XKH/JDAreM4oGL4eUG6MalC
DspTozv4ierKofNlzhjgdsL9qumnTWtIVN/NdkFVKQvYUlLPEcjrhHd/lcFlAq3g
di41yN+TpkpcwdmENv8A4BUeyZEGzuvB3T9RZUHUvzzh4WD6FZ5beRnvAhNszddy
RfxtqZg0altzrMjslsPMP/Xm1m6mm6DaQ3f3zAzQkRM1GxPc5Rn+MVXFUZBCwh6N
BM+/y/n+uvEmBM9Ctad9ZaMiXLaEe3Cu0XQkXeGIJ25EnCfmKbDIgva5hsViyJnV
Urz9vpRNPkYpWvaFvao0JISLgX3xhUYU1gyCU+h/9pJ7Z6223MxsNwZOB4rljwse
3PN1aDzv8JwNazCXqzq+sSObV8G20ic6F6tWFowB7eh6B0Xqmeb9gdBKxUnsaP3X
pU2WAaotfJEaW9LNk4FSsc1NL7oH509PSuynCzZ4P6kmueqeNzpImylMEK4gqu5W
BBANvXOvRiubJZlPpgcy0VpPSINNulpO/QiiFZe+Q3L5DurZ2QixGfN74WlF56KH
fkKYV5BRRVzA9Nao2Dpxa8Yw+t0QOc2C9Z3NegyI1azodaVrk1IK3EjE5t3kCr61
jOrIWZc0stEtjVdww67urbmbAfc+PO4zRX2MKq0ImTty0zHTl+c6qoFXr9LiMH1o
l0bIoteQiCfGGwwq+PJ9L5H3lsTlXKj+3vOpzyLVmE/DEgvuN7qFiwFSNeErJNuW
PUhArmNOfwAS48fJCJ/lJz2BuAOjVKDpUsB9gCBBFT/kLj89yMbs55JltEoJ5pAM
ufn31jbCoFIGDjFfjUGLso3Jcgom6J88xqLAe/NjvCZ4rtPhVXFy+avsf6kXweiH
SYp99vwZnnKbBKwa3BCNC7gMjWiu6zcullnuyQUKkZ06XrgaBqWnMB2cLEsIt2tH
WRHXXYZ5psgpkela/CIAF1DqmeDW3CC3i1bqckBjrBEXmqBW4aAMilTEIUo/Es8w
JI4VR+GlNoN2Gz8sMFzLtJ3bwt4xJWgxKXXlC/HDM2lcbMxb8yG6WZ/m0bndJYwS
Jy4rO61tgKTY3U1hUJKiZlK1BmIiNu4SFfWs9C3LzevNd+K+/T5SsVRxty1gzHWh
s9aZjhhZGu+j9g/ydTRsiY7K8gl+vAJTdNp61niFi91EegpDl2vO4EvhoHRTo0ND
ggAb13s+Xx+X0dtCqR0Ygb8RbrCFCmwrqODs8vPrySzQrGlyuiL2sCUiKsatAxhY
1qvCy+KvE/z3Pu+o+vS2kmo1C9KIMQKPRSXJ0I6Z02Z1pDo8DBriPKy3AziUwqWr
wTkmNl/Apyx54aqbzyQVXYBZt4liAY48MJq4Cn+KgpCCbULST5VN/E3aqjTIyEVO
S/NMXRMGkD/XPHbits+bUAStojeXcMEB5UPhzBhEOTlRlfGRA8SIySIAbM4bB8Jo
8Zj6zvU+780H4zn3NWY660Uw+5ql+67yHpT3KiWUNLJNfpnwrVu/vpo/7011mSUm
SBx2PrihFGb6SsgNDu4F+goByPRbCQLGD6s7SmBrdpxGPCapTUKZ65c5wwFtkgLx
jVMFToZGrknynpSs9zqfRwG4rktc+e9ofaOZIfBni5Foto5X1HDgxJ9i05X4YBoY
2p/fr4t54Mxw2kNSsgtUsYxXyKECkM8YtMYO+M5WqCDQbN8kYYLW2nO5XjaXHMrj
NkU6PwVD4XCteqt961FeaQWejwwSaT/r4kpOW3yRGMMa8EpWeL8Nr3ZnEhW5X3ga
LTC8mRa4hNWXOPsyWAiKdZbW60471gsG1o1KJv6XJzrA6hxxWoRqwBWCz3RTsh2z
3Wv7Hf1tJoh+Gzu/biSsjuO846MJBQZG8jRc1znjGfKC3lBIL7bp+wPpLPxjraMP
Z+S6FJnFpF3M9vjNc2X9XyR/wYwMDMpyTt7xA5opgUND2yz6d70nISgCqgqQvCYp
IKuIBxfvUv7pm9FXh/MgAFVAhYw3K2BD3ifCm5PoUvzp+ejHB9lTpfsAFuArhcC8
4kZiu4aiQwzYvO5oN8UBtWl+4k/WPFiKmxPah6NDtvrAI1mAE0secPJ6+UJGX5fu
gvd32w+ut4Cti2hZl9R4G5BUwMsdSOs7MgChYxzCVYq9lIOKbNqHIPdUOBKgiOAY
0r2FyoVdOv80OODISbOkcddNrGr8VQW6ZLubHrVevWR9aNkVp306oWCQfcmC8Glp
y2+allVMhzXzQyvuLamfBbhpSxtHAJEdRcdNYFBuDZy5uRSLP12K1gCYRELEu3GR
yq72qF5GzzEejZhJOprbvblUN9bxkEzUvlkTR0UOJH0uNfuswXT7qdhK5+CzXs2z
bwImZWrgeX7l8uJUH9TJ8PSoTjwlTa09xtLpX51JHn1121S3qAdbr7fH3zcGTmEC
ApgyGb49IW1tSRUrXR4cuR5+fDsHMC/aIF7rkl97GPO8F8NrLirXAIY6OJkgg1H+
JfHYTe5YuSJQi9PeCFdsu7nN1nOd9b+muFaLYDs5DsVVI59619Rli92dtfhWebC/
y4413hRBXlNhX9NL4caCX8stxBk/qPl88Bpfcf67nQI803D5LKyGFvnaxfSf5VyW
9R6lPlLyHH1c2qnCWblzVyVz6u/NpZ8bSU3BS6RKiA1A8cHeGiAzOK0NHMCEH1sv
jRQ7ZN79obPbVIqG507GetSPDVBrhfhb6jpqmiRIn3rzQsxiuxXZos1LkcaSV6A9
gS7kcs+rJUU7so2T8q+0ntj8XTqxBVBMUntKj68hITNGQntbQz3H04OVJOwGsdqg
GhmKFkVOHQS/yHrHXGIG8AGqpyICqJVnNOI79GW1YmqD4FnKAjtUHhFpvMAenwjt
wpyncYuH1rrCc52PBU8ORvA/7P65SfZaLlGAOC6ZM8svEoSk3UcRbs0xDFX2omXg
MTe43Drg9dsg8Ma5ozW0Eh0Gt/IMdJzpAzWYtylWA5CHjBuDW7Qbuz06SINs7KX3
pkygryhiiUSMpQbYdZjMXZzRiRllDca7k/IrMwAEct/3Ncay1NYgI7pkeZDIu/A6
vjiXYj9tMKPSyzd5TUSkZGKX1dIYFfIYpQNiDKZPxG7Tdtd1FyubZdQmLLMobi58
RvqlTolkApPqig/KL3GiyE5LJFfPj5pVauyj0WwMCoaEDxuTv7DdSGWKbCx311yy
hNIBUYmB2OQ7GLcEjtP2pNCZdvOAgmOMBunwrp2H6hrOX08GbOuXZoRP6G3U4hKm
n2jo9lyUcTWOJan1aoSLhRK0+kOm7nYPlP1JSBT2rfTnddNq/P3j2Fgnrsp4/0Eo
j5BoYTjbYG3aa2+tfZwjHKboS+RtKeIldabZAz+LoUZ8B1hb+S/BBLe1402vCVOy
Y68Fp7iCZ7ls45ZrGAzFK4sClh3yJJn/HCqbotyN7ihpRH6cMdrtTZbnZQN2z/Cw
hA3gq9mdHNfmb5K/r2+9NYKJ++vRGuHQuzlQRTZ/NUN+6HJ5maUS19KgD39184Pe
XfUDeLFbz1bBBOjE4K/W7mt24+/1fXSChkedMjml8l8IxdUSb9WKiSfLZYCJJ+ov
hWuRj87/Ni1sDYWK/uEJpLwwjaOIlr1MRvgzZPC7uLmTzAEqmQOA8wC4t3UUyJHz
Xzx8stSFN0XAv9j9Gu75tWiRud9HJ65T4StymQSzV1DmuBAUPbMd2V2Xi7k/jmuC
ri97HKxcYDnmGRn9uDkYHp2ue24Uv3dpJoelHXJzcyBxzB1i2nnF0HkE3oHhObh2
OQBtMET5tQu0jAwfCmAagFiIG9T7nj0M+L1NMCdHwUTi8aZF9OfSjug3SOWrLPr1
8f//YDGoyJb/z/kwz7u+2lKRrtz4mSLRji9ZwCgam/8fn1+hlUh7d1WiP3jxQfS7
hRoK0mXr5mg2RUFzVqObs1p02qExujX4SrYcAasZ+MUNR2xgNMANZh5Bq/G2yRUG
3IvsK/AiQ/VM1FWdstqpGVnir6//urbOHrm/pMmhDDPagxAJCvHKIeHdl1eI35V/
rFQCKINOF0Gvj/XF/wpeRb7cRI1JPfSZKwB5C5IDmuFld9kAiDi/WLZ8aPBzbgJm
0OfV5Iw2uFIet/vg8PXtmYXyqYTa+Sp+i6Dcii+xPXeCq20URsNZLrzvYqmZurlZ
hBUXB5OdNR25FSVdQbHcdln3tAmd9TpT5ZNK+DHcWnA4dRxG/2Cc+OBrT7mHxPu4
Kckh77M88JWlnRWQHuDBI896eN7N5gkRpNVgWXpKF4a7XfYVbpF4D7OZBqkg+3px
iG/BFHPuGDViePiDGfdv+Qh6XGeyMC3psOOl0VU8fTebZEgNjiJZCUqfLx99Gljz
BLi/239KZDQZBgRXYPW2OIFrlAb8MKuRoGtjUh++JbzI3etEuJSZCMncfwX2cBHM
Xb1j7OS4+KR/Rr4wZtM7omssxFMr0TQwAySBAab9rRLRTQLtI73IooYNP4eTTfSM
Yu8X48XEJu+O3RYGhhWxweuw4MkHxvq/Cc4znyaHWB6EMx7LBsEv0DiDU/WfQoyw
4HPQm4tabYHpKIgp6Kmqkx/Ikv+VjIhE0PNQRcF4XvEzukyi4Bwfx1vziM6w8FvP
yBUVrFH3/ILQ/Y1q6pzbE3EtyKxrILz2HZUNXIRk1C/I9WYNjd5F96RGS6UQ9GS6
4YHo49Q89Z1LxCvgEylTtd8jMW8iMU+QNTwbWAkhMGr/6bmMTGNjB01rzFQeX4Jl
LGkKZCgz0/bcbMz3SCyT5q5bzcuErLI/KYdPzrvMn37jQNiwmpcFty/a1ple1N9I
Qmj9cj/sogWim5CtDUJsUVF4ZT6d1J8chuujmMhCM+X4b/kZrtXnAfxfgUkvdv3x
akTRcy32/HcBBFb4kYywe0dg+JLpa0yWShnFxLc7ehoLxjET4fwfADF+yKsWFS1d
th6dU1kvp7Lfr4HM8Z1EXYCWB4zX/iVGZbACbVu2t6twyIUhAu7elnOpi5te9GqK
qdlbgBxZgGhHMrbxz95wpGporfCJ+R78wz2pp2muLCgDOysUTwUP56iBuPPGwz2M
98m27WXpV1AxgVAB8A2LwesXjOu2/QWBRQ6wraaSWNJxZH2GOu5z2S+ryajBaVup
eDM+3Hpt7Ts1olSsN7/Zh39Zsrj3dzcqovKnLkQtf8nz/CmX4+IsY+Zvyn91XaVZ
TZ7Hf/9mWEcrP1wDeo5on5MUtPP8UH80hsaiykArcKmSQ8z45Toc0utXreplXDWF
aLBcsuIYrNGyNO6MfhglbFSQHWDhVc2FgrVAwjKxJoYyx8EgnbjOxhrtiZ/Hg/FT
+G5ubdw973OJX7AB51rcIyGA/jpBoqHh8ecJjIFiSsOPrRvK1xdx6So5EhftLrkz
VeFgWDYdECekKhqUSbsId5BQfoiQns+NjYt2AhhAjaJ0UqVbDYdAHajZQppnZDh8
lES6RqqCk/GtFTsRCGZPHrTkS9mnugh5vuTHK5Z2N0UgnNewjVJG+8la0eBlT9+T
6Gb5iIQyDBJ4Cjx7kVmc58fxQESPwIqXHgCKee9aTAlKLLBJWFSJ/x6JUq30rIp/
Szd4t9ONpW6DLfeyoI9DcvBkz9Hj+bDUBe351gJMW5zHMXwQJ5zLKgL/iTQI1PUo
1QnbktjTwU2NMJ5BvV5wxgScMCZ8iWVWkqJkOItMQJB3dqVoUpdy3s3VOGggE4ke
tCKXSP+uxDXWG3YVv1gAwdIdC6Djo1lJqqyfJYc64cxJ3z9899CyLJlcETGICjEI
T18Wp/RUmmCnM6mFM6BSFto4gUUpWNWHM0yWRft518I947ePo5ZunkY4Gc7BXCR7
8piZ/HxHUVB6cyhPTTo71+lo4jNTDGlXJGbSZYfwJlhTJh2kH3aR6ZJc1NSuajNJ
UfPMXJsZuRVTKLbC3K3vESrOtWq9jNfxxC1rbPvi8npTflZEnu9NfuoR7eCHUXyu
osCFNKQbF3Gw6tvYOnLPsOJsvM/nSASrAUVJFfrZCIWeJTyEc2jDF1zE4mkD4dbf
A7fKyBNkdZ9cJJT/f4izDIj2lPJUTIdTPu6/Okg6cNsbIXNeAsXgtwuozR4kL0I0
xm6WKqbqSJzjATcIkcHDCG5AvG7BbPuC6LdjENM/JCsm5F3YXkYNuiy0Pb9hAPpY
fBqzj96Ja8Vlg+juzfrfSn4yqOcUZsUiGu+eqnfVSvmGouk04tHH4DUVfFu60hXF
jCmpmYRMz5uJoGC7tk2jDmcDmTB7J7SWBuqj/rbokj8fHlcJMR/mMFWXyo6uvzFq
wNPcY3gbpHeV+oTMZnRkjEN6hevM4Q/I5FTq/i/4eL9gdviNGKSX34HqlYSQ+0W0
e8lMy7BzyChQquqU9f4sQ3f7W2TH+GMI96s0FhMDgJrHwgKe//jGEwr3Px+IOYyb
yxMVCfY9jJwqK7r1th1p0Ld0cRujcgaRZDEj2kslUVUvQMpuPuR125v4Wk0Ajefb
AaLZa9xkkJ3HXYlWvwNGyrG5P4tTfMN5jDLO55oSStYc7wPG4tTZcQ34K+niwqbl
Yt/8uTmzR0azm0z6tndk/0ToVQOSM6K63NZqU8PCV7ME/w3THd2C3cMjHkLX0URV
TrIGsxHzQdFtZxCVsM8lmmNuG3CLeWZZKX4R8cpI80iTdnnXWoXD/fIhiRnamThE
Tss9jLtyRg2Zbm03qDaJsFPCTwpIVOl/y0j76xvm0s3xtP6k9nCwZve55sl7inJB
RRneI/nsgbXvRb3AEBBsxdAs64sCO6ohQG51O+/EIW2kIOYHI8rQmXEdOM9wz1DA
cXWggglD8Ynzs6vrEiFlTXSrT1c+p5oNc7S7HqiOOp07ssSWi5mx86QIy6BLHRO+
70haksnwvtfElX2Q7ACvR5cNhgUCmyExLPRbRGXMc4pR2NgIq1Ikl8+PCVtiVVlR
hxQ3ScxiWKcB1l8fJFowjkw+8vUQdr4EEzJU8CdLG/Z7Pfo2JFtVE18Ao16z3qZ/
vxVKClLbbReoLq80m7OYeifKss35f/sVa44mrXOv1czMbzyI0i3w/zkVFbo91Yt1
rvCp+ldNlzXIA3iMkq74h9gWJkqbcHjGM8QM0tZWXQBhg7S3iSdbWkgK5l92npGb
ItshZvGixFyn8PvVOrIzmM3DoSQ+iA0tOUGT/SxwTSQ7sYWOZAvEU1C7+dCP4TVc
FfkqtSI1ho6EP5DDh+QUQIIH+LeTgsyrMdc5ZcDVwmAshxmNGWyvHAjpFacQEuQE
hmMcmSNXgpi2+s03cKzmYUrGkFdSkApoXfJPCTyjl5hTR7Wi3dM4alwZSU2e7C3A
lRIR3JLLr5yLNbPpBCGVK0UZ7dYuvRcM2fKMoS2/M1/wlXwRmeHLBw43AQgMVweR
oLRQDlXL+n0K4cf5MEpAAPJE+f4r/Y24JutFOdEn+z6C/TmRF3OGNkvYBzKWrsU8
0RqVvs0MrESGswNcG8XUqAp6dGqi3vk/BW3uCVq3CgViFtb2+jOJP8eV7YdyEGkW
VOA8czm03bNOmVaaQzXj0QhSjw9i5sUdfRLl6wawq+KwL9O4Atzu31MW7JOiDMBN
swZhm627m+6RHstDgUiE+DIVPB3ANyZ1jwtuu5USesSe6mZLoFxYN8KSXoP5Z3L1
TapLe96Wmu+ru+H1i7334LdBeq68yvhS4yqZi1WyQDGFNsARlHBXQ+W1CHceeJDq
UMgj7cs5Nr+RQt8yNY8ndNQkdrKUF0IZGPh8O6c713yoVnE/dWj2W5+dfXKMwrDR
lQfeWrYGC9HPMXknzYSTS+0kJXsxOd/a5KXGyyfGPEh+gqSdiPLGZp0ZyyKfyJZp
Jc+2+Vbj2Ukc0M0Da7lb0lKY4D1CfZNXAEDuyL4mR9qWh7AAR6BO43tQVpuLZzlx
JmQCyqdNfZ1gl7TFgfeNtKB+UOxijXAriuGNxBng3S8iX9FVFQVQQKHQtItdXhMn
GKZxo/WPB0vaPs4XJ6K+T54po9FxZbxLR2M5S58JF0GnfqHbtgeLN7D9s8QU7Pxn
sUP78ANrL/SMF4k1D4WcIEBCbcIfEuPyRHwO8FI+5PtQiIC7NXPrV2kRUHfDrW6e
Vc76gq9kAmKru+1MR3KnKFNgr/Wv8gjddU9ZvLLV4Au3/xtpiMa5KCC2DmPjEK4T
+cOuajbf/ECfh19RulpfU+cYIc2s7QqNG+gJ1WwgRlW8Ho9BacKwb/tPVxpGnYGD
HMq1mk9BSl3pPVsM/orCpHIgWmOHv+E9L4I33Eu1sTsducicVVrJuL9E0aP6k7eD
FLWyOvjTB56xKJM9KDQ/7Gbf2mr5l0HHSEBS0hJ4iK2CNNgbeKRYYY2L0ulDciMj
JA1axjo3ggevFkOfhllzEgbCCWIR/rdXEHpABVMghV16cYuESZigFQ4WaT9iQ42O
QhwCRl5fRTC7FB/fi2jEqozipHidzLS1FVSG91PnM8h5d87g05au++KlcoPWsvIU
QO3hPNbngIPFCrbAjXyb6CD7zOQCzcOa3I3UOzXMGuAmqpsZVpx5Liaq5A5+zwkU
Hq815EAMaWmOQ91sVvjTHkiKEDCgo7IEbVJ9mJPGXD2Q8TVJWV+opSFhkx/Ktrow
I6jk00+qcRGNRUIajA7HaRJ0BmCq6Y75oJHLqAGIaFHCWn7r0lcgQdj1DFGrYUbD
4HYGSM2Izo7+b2hwSfRi+EjPU3pdVfKCnXhcslGuGYwfYIJo/ZRMsytrym6w0V8r
7b1UtsWRPgkfr+yUwklzCFpnK7cJ+O1d6vrxmkUsdinhEBcDAU2ywuTL6yN3Nis1
ZLYtmPwInqAaPXqSPbWkBiGDTa0nRSztmLRyvu4mDRuOfYEZDUb5B44MNQEaEtFa
ifsT1E8iWfjjr37SAneyU5QhlR2N+cna0imdud2VNnSamq52LXXWyz9Wq6p/F04X
qdl1opgntOOnPr/Iiy8n2y5ntCd8gJ35yRWe9lTIw7vv532dfmTpygR1CTPdU/At
vUFOY8w33DUSVJnmHVAYSVISN2TDSIxEbF6908ZIWk/lfbbOOiMgj/TcyiviDeVj
LClyzq+LqszICBhfz35GyvEb2/dmxG/78H3D6Wwua/U4jFw3IC3iifNItFYn1UrK
SxKG5mFH7k69FF9AO4S7Cl24hLGIqwTu4bGUM0MB2HutQY+cJRiL7luT5sfp8e9N
EUjjh9vy9wwW9bwSG9IRYFLzbdfYeWY07KbxQkig6bvH1U1dT9k4qg6kjEFvvWCb
ctBtBb5QaZJVOm3AOLV/VTgr5uIcayKyL9imOtwJZUxbHjmo0QZ6J+vdSCS+RRXN
Wo4BNm1D3Bk6D1boX9Sq9IhcsEw8sJRgMrKx93zTg4R88NMlCmIQSg5BLTGCVCMz
V2NVlGE62xFoTV5jBt5BpPoTZaAdsDT+xal1IVNAhSxLthKn9H+pnfOa529uBFid
fBIcvmhLK0JX5oQv9/PNleEFPEmV8y9/W/sA0YS1BD+HnrDt6WBgfIMYztXQ1IGC
84tzUaz6mLAZuEduGynuM3+sehmoeU78mmWVCLYaOBROc+d2q2F0StFXyTQKiTR8
tWsXM34kUayraEdJ+07OG53Ik+dimqrWvc6rDUpriQnmAuVNCotMU0CwPVYf8B+R
zvPtBnvaThPmlxSrxd2LX0nSUk7Z1JEp7E7BidkFOZmrZnol08pDppROneoEOIqY
JhWd7GBzoA429/Zy9ACNSCmr5q5rjIFlon1sg763MGdrPE73gWnkMinZMQQ1LvCk
ybZOqs4kpyl6EX5XqfdKabWmATIE2NGzXCBprrNbS1iuRH25z5EzfnJN2A4SSuOo
YnJ9c6rm1UfdSpqBHjH+/80CHhb27ty6dbLi3GJrG+iL+5PBZzQYY1Mg5fd7Z2Y/
0sRqk1fZfbqknuGLxbccWcAfKjj7lwIe6/tp9fwQJCh273SUoOv8lCEVYT0YrNDh
QvJaAobY2ehhN78kGPGuEbyz4UK60AFTgQWtwje4Y7oNzcvN2NOfGuFaK5nYISst
iw169wyNQgmJoqwLqKKiBiRtFrMwuJs7784MeMCiki1zp+fYqCvyTuiOIxl88LWI
5NLlmpp7K99cZdk/vYjfd/sV8vofNF4ukBM2FMSXvdWInpj2sl/vqAqX5buTKJYh
hMdT0qwrrc7iW6NwAiRiEkPYvDUxW5JAy1o6JV77Zb4iBQfpVgnkZP9S4R0+l2IJ
iEUdvrYE3DW7jdl3F5oKsfkFm2j2UBZcQxSF2Cr14nOlJIKJiLBByc8h7MvnBMMY
1ZvR5eTY/FZMZqkxMv+MyhFgfmfiFRxzvNrZF45jQS3vlPN6goiFn3ON4RiGa58u
Z67lshHRlBMwNE0m/G8Z8NkWJVEwxohHl7SbfTfBSTDfHgppqZurHumbBCVUlFqM
OubBLD8bAMebFYZO34DFYWJU99/PHaCNyb9gdKtIBITxBnIZZ+sgArMsYlSEhz9p
tHrS0Nw26EvP+YKNt/jPgtyZZ/tHSBqqw89mEHEREGzP3HmBItYB8gU6lXuWEX2W
FOh+mLLnVWMpKih/F4bOWMQ4I12XU66pxtdGs4W/7sdG3msT1rhpi7spsvs5zIwf
nzyVEU1gobakbIlX79oyHjQ8BhxgVn9aQ/QsKfySKOgmwBZLPnXo8KkCRj0++INv
L+oU53ZUSA3E2WtujRcBLiXIr+qAhTyK0gmJLBF9vmZidH4iL9c8skW2IlNtGIry
UVUgsKsS2OchEaJM+hGr8NrrvnyYwXiFXZJFmmz1NBzIBKAr4YR5MLqfx4fH0wlh
YsMA5vxua/d5nWbHeN8Af75HtSiQMSWRt87M6FgP943/q5AGaENH/h618sXU3Imm
0XOg9dvDw3C6rpuCJ10ZTOkE/XjG0EJ3pMkqHBjqcmQwJQBuHsCzwxdsnkJsvGV/
G36zL7Yb8wdTHqrc91gdxFVHj1ZIu8R8M6z9X8EBqR7BJ9QSSls3i0G6KNcsJa/G
nZ7GRw/zikgzfs/Xz54tyAXZgP8nFdGK20E0t5rUFI4UEk5iPgoGp41go4mEE6jO
Q+jLM1F3rHeqB1dru3W7xjvWcq5xWrEz5YuMTNBK85mwSp60cvkgjXtYjVV5ZULe
3YcCCf4x1SflXTXICpHaFgq6Jj01hnWUNPP8kVBjeDlJn6lz/T8cbiWQcDL4Lvi0
T+aARQv0VyZJKis/ACaWSvFYe/FpMQdsJvcrRpOVQw3DrT1EQHykHg//nt8YG+NL
Dtt0whkb6cmoaBBp2PqbxpUD68fyHITVQ4vmu4E43FtJ9bwann6lEvDGq5iER8kt
+xBmfWcqUH9lF0q2xTvoqleNjOAdzt2WhLPzwx0R3slBfndo96u9MIkcNlpfgAm+
EAUrYtSnRWotZLHOV6rkJAHLXS8CMeuxqcKZwtOrAOlCRhrV2Dxco7Uw6q1gWsKV
OIsddy96gXKOSBFSJ2WYGXxyeFpN9XyElJfmQb08994Adzk8g+LCMluhoG+vqdyk
piZ/D+cFIhaUOtNWNqTlSPJglvKezUPnnSZ6sCZ2vSynj6awkp9sMI6my2A6tsK2
6YXpJD4X/063bWEX0dqWGItHjyiGv32RXAHBooBUxH+gg7ut+AxnBWsthGh/ia2f
VM0u38H2McL3EVWJWeneJ9tUJiOYxd3zhqgzCSFG+xr1wDYgpf6zcSLcVedtgSEx
3Hbk/wtU0UjtlidQRMD9P+xb+7PRkF7QMtF5dpLvPGWFqvcUBmXL5Ob1OET1i7HH
eS0mFwdZQhdGMH5oBZs2BV9D2n9yBTkcdX6WoHoSX9p9KpXR+XT2XMxOvX0iPMxt
0JkfZztjXEdj+2lOmUG9SLvZhaFCzed9mSYRp66OVOgK44x1cn0p54DrAe+I89vH
f2lueo57fFTO3ZmLebhpnsVQNxWqwGwFbTDXP8F7FDPpB/9XUELCyaI0uc9lve7C
QYQ4Tv0pvyCkooHXrRYreeQsbUuz8oQ2nzL/nhNeE3rDgyZpSve5aoUXfRJPq6zr
rQUMLbDGQrZbRwzz5ks287ozq7uxnu2qdLnK0I42Zm5L28d294MpdDuj3tk8reDe
UvZ7guCdkMv2LUgCSq+CjPeABzZYixQkHIJ9xCSY25ORcHpKMrFUjb6Liua+/3b6
1jyuTE2OxWiI6LxrKIAv7eY0kkBOMv9/PcEzYjiDfVwctUQUNL+NdU9d2kgSon5B
2slxAbMDnlW88kgJiUYXbFpa6ScDBIi9O9aHtNYHoKggyDxraaZWujpTKjB+TGC7
OBH9fxe1f2EE9TwFnmr5YJCNEFfbBSdOb7pTZbUC4ERb3FEmqzBtjHvmixhG2YvF
2jyQWXPgzzGTkWfA4PX0OiQJOMJySwtCxr3YLu2tODuixXQhxxb0YqrHcD//YQVl
mzeS5B2dvE/6jocTBif2yTwqV0/mC8B7vq3tMw+WeANCE7UJCycWQIVoJG6R4mcd
iJxWZbf63sU0NBy3Nq2oL93sEyGAOf/g1OY5IMNhO+vcK+5vnlztT/Im7/zq87tj
/Qi+rdc+13NY02PT2ccTJY+TEXNvzoPiAvN1C9mbr42tDLdJsVcpUyVd78+s5KeU
+T2JaDb21p9CivlTJqgWU5PTTABKb1CNuL5oE8YW0teBcNhH/MSRkiT98jrUmbzb
Aj37gAaYmJkhdmn8fdLFSrd8lR5yq0Vkn5kEXfZNfAJhV6XOREGPI/E1JufQUrjw
ibio7eDMLEk4t/YJMzz6IoVM80ybaziGyjcr9tYMHFGXYFhNMC1gM4uJqQfycTs4
iBmQmDMFyp0WC0FJsriiJY5e52UvfvfEBAIhbnTvqt+5JS2gFkfwYGS+IVYjxV1b
D8R6B6hVSrk7T0GTDZiEDyuwHz0bpTKMidE4datT50eLV5X9pa2Cm9x1Ep4jrDyE
tKh1IVLdy/HfFc9FsQ6dRzNVknFDavXCd8zH7E2aCzxrvZkpA7yd3vNkBjNJWaKf
qa6bRuyZ7cpGMF6s7fENI4f4vneDHZml6VGF0lVKKudBl62Fh9tGpzPo0XZwrJIa
UN+vh7ELP8QVUW9vHdcD1RMyEbL9Vb/PeC6/NoXc9doWv8pIb+EZXbHU5c6VAb+x
jsf16TgJ0x1N6AOyO4AZahbaKa4j/qARxgPs1x1j7p3Ky7CzMitinPS3J/OEWm3K
tUsLp6OdC3HkpHcHmffIKsY59uFXR5AxsnylQcXcuSuNi1/SsMi6tonBI0GWe8n7
Cg1DaC7kJGOVtmWHN2XwCi3SHzvaIjPQnZsLKrfi+S41ijBstzDXdO0JED06hg53
LfG9kVEskQdkntIvqvPFM8x5CKGH3RSkEWB25mNQXUEO2U2jb/eNCPOx0TuwlWtp
0HJfE1NPtnlAt7EwXyfLOnJRs07KarbfRZxfNwdQEan1H9Ms21WbGR6seSLdBbq4
KYMn5ipqmSXRU0nL/zqTjP2RLVl9CNVtgyr3cuMNQx1el389mwvdrQISWfvaPr40
9xJhVkgPULQJg/azDQMHTuDl6Tng3lAnYAbZggYJ7jLoXvHl7RlgP/MiFP0+CN4+
iW6W7blk7XjnmPtxFognTW04wpP6W6iSVKWQZ4Y7xY/9HN/5sOSMEluStiyYAtiH
Fche9frbDiWtc/Y1imHLTrZxkQiPej6mD0txN3+7fYzgpPWB6+1F4k0H2bgqshdq
6H8MYmKvRLfnUvi95STrjRnNG4GwGL4Z4d6Qrb4/HW2uTueLmw4XW7bIxBfvt/Z3
3HSriftlUqQNLQC17oVnL1HmSzQBtYBZHZ+wEV6EuUmqqFhkxKfVaJDAt80sDuok
7MMyB3n5F/Ouh7KdamH8GLW0mFj8zmivlVgrPsdZHSE/bEBeYiz6ZHPlP5LXJqOf
1Ul7DsHB26JYGaJlY4CJur1+aJZaiBza1wf4zkD69YVkSeM5AuQNiPQYOI1pQcOP
D4ZULWX9Bb1Ep7hnYtabDQfWLG+DM/powSPM/noXXLbWwlnevtGuQ8FuOcXHAEbo
4khvDjb37nG2Wx0f2uVAlDmzA6I5zMkikvEYc8Mbo0tiRd8Nt1aLW89AmerzkwDP
nWAsjZciinjUO+5SE1BwpIZ8qGaLB1IqSs1EzUVHKFlZBQx640uxQ6lNufThMNHH
1Klwf8l1gtAD9cEfs7GGhLpXmxNAiBfnVdUkAxBpB8O4iCEpupeFV97Tg4bJvN3P
GPebEsXJjcbhLn/vlbpzcvR749RNsRUjUXJaxvGRUKzWsaxu8svK1PcNeOuIaIsK
fMvIpYJRE2tgYITV4fDfRA+DAnorwHe+Iqo4ONpolHPKPkBxdoE6X0HsgzGVdWVV
sY6xGZp2BklOQKTaC3LTN9WR/fqfgeJHO060FLbqreBjWvRSuH+4eiTssO5GE/Nv
noa/zJb3cQQ6WEQesIICA7Ahnh77FM2ZBo66XrD109ddJ3/5eBGPciHfS08mMP2Z
S49zFZmhQo83pI1x+POhZO5ThWXE8tJYWSXggSDIucNMUgh9hN/F+IZVMa7DgBZ+
ZIMoX27+pKoLyrwkBPY+PItFNGqDte+gUjDH5RvyVBOS30u44TimNAIyCc7eMRAG
JxTaUFhEvVvR12eYjfwe8a7W8AJiBvUHqp/FTllfw/t3ipD4qV7sUFtbbfCVSt1g
ErixxJt9RGJxJaXSOOZ8b/ebtWyaPt3SEQGAcgwCWt11Gq9d7nJQ5aDL60RJBZRQ
HYD52mqQdscoGMe4MTIraCWXvA5dFzu6TsN+T2rZONiBDg+Tp4+9Yiku3K+hkETc
bLxjWA6pS6fc1AjvIH9ch4i3rC/qKOxu7TBMo5FjtsZDrfIoVSP+jZZoHyecH2Va
F8vnFSGbGnJbBO5cUnymF1xYznWu8bcvEr6VQ5dWXd7Yx2uEClNuFFWkYVOK2MDe
pY0pPtPutJo//w93byiZljrFW2gpC8cOMHVijLRo1NAPNyNeOYtfFV0aMPXEP7Rz
B92jkPxYeZmpy9fI4QfYFDlaBz13GTAhKKg6HH9OwWbIoM/nJi3LGfobhGXSk70t
7yOSBaGfjHFV+tC4uUS24a8OWg3SlG17o24KInL2clVyPIPJhed+ykOSl0tMMrkk
fyD2cHC28rVtGMLe6PYFvS38ZPWTvnmTp/1jqtTvsveRV3Nx/Ow86nNxCC+EK/tw
AalMo0ViRKgZ3lM0Daa2UD2FFNnKd9GVD162d7WH1fh/0O4gye8cjE1Fq1QMb+iF
S27WCfFK556MZRb3Z2NnyJUtKhPY4l7alz883lXKXXhBnnCCpKDmFLvUA3wNl3gL
vq5XDnE2J+GLldIwvBLMHFvrHRlLtuOAtkAU8zqUepQcxKOr+qVARuOWUeymIvX7
lTvKEBocJrUUWAe7F9lmLRe3/1G+Q72qYDngPcK8W2IorWiqZqhwdMF/uUnFbz7K
lg3uxvAmDJfJYqXtIEC7ZvpZFbpnpF/EOg6SlCc5jKGh1YCCh4qt7E2WP0YA8/OS
4mm1d/Bb1LMGFW5ZJaKpzxx/VGX/wzo+BcIoPCRhMqzb4Au0pVB36V225FUeeg4c
64373VagoQgEv7bGRbzLC4NxeALyTmQynRKc2irPNIsw0aGt2L+pB+54hiTlRpyh
P+tLmlVZOfD8rKC/VyzWc4kuaE6UrhvF99hWPhoRYdV58poqjwg9XS7WrdtHLR7Q
UHcSKYvbksq7d+dyB/CblCAnwn+zjWn99wkHU6DLeqJRNDe1U1gcbKeBWx+rze6M
0H2KUplARCV3c80mJtYjeV9bjdt6oiP0MA69b3epYCMrYZIEZEkNv1EMr33v3lRM
xOdVyRhvZ7WF5bq/B3armzY310SWoSogGvuX3JDQteCdo4+ymgmSNOe8YIdxhccN
S31qPz/sxnl6JqxqElhYvrTuB7S1bBKBExroNBEuBojXd7GkE4TAI2KCYty4oKRd
iDz6KXdXx9GETxWKOAA79yReu0YUSdI8ATGAV81hSEoLtLiGCH6jC3bbPiaOgPrd
FycstG06GRLUdtQ/pxG4RlOFpMWc4sg4HPhzVNo2i6kEiocJysWe9IOz8IGI43Yi
zRvytJdFUOY9taSUsWG94XCu2UCzmczJkHR1xDOmgfA9V1vKy9Vqid7Rg4rhE1by
DlDo68kRTIUu5rvTZ22pXyFsn/LFm1LTinNm3NpE94+2yBcW775/JymiBGxsmcaV
80GrMdZ5cTB4/+zbjzVHAXHjGzLKawEjR0Np8krjz07Mcy4CXLQTQg2rOa4JCQ/C
22DMcICc9x/1S1M96Awde493/r+7sW1gL/yoq9T7YaGsSSq1jxvqXqj/I8Y3qPYx
rmkBbTDxfCEnZOY6Rp0RQgYm38A04W9xaeHPXwKWp5P8KXBg/Q7xhOGM4dQ41ggZ
bztnshlqttRlokuL2Px8oxIx4GMOulkTrMM1h8ErjsCPnBHjPufC261ourfFex2y
f+s934nMqVtu9jVsGpWiMblVg3KtA218LTGjdYpPSw97syx/OW8RZQsTywC1YHu9
jorq+affOw/RruCZb7lPxdf8nZbNVdLGiiaBrJbzFdNcLrQU5I2qRMWjPiLWqGr0
7SPd1kdCf0yd3cV9PAcXUDmW1don03yPHfUlAHPldoK2ctx9QO2QIjl5t2VVBukQ
yW980qRyo7RHQJAr80FZN20QOTsOMUTdEW3eJTTpc+VP3oPFgs9OEmJnWiCL8tQw
VI5O2Fa1GitzoOydlZ7ajF2W+mrzpewr1TOimVC99FqArIl76z3Ya77m60jD4XuF
FfW3gr+X20ilTbQUenhL9+Sv+k5mwSNPE0fkp+YcSPK9wD3BzTnDgUyHmaVX8BT9
DhMNykL0N/HerTQKg9CnDMFV8SvW6S/2U5ZNwwyMrPc8UCcKqSCFf3d3ULfzKPvV
+806G2jufbXTDF+c3TllwnpFxTKetNFULpfAbNV2Z05OOeeKkUi6KqXSYblgkb6l
IJuAU5qwvvrXFdWj3jJs/QX+BsWoMF+MKDWM08tEMBzZoa82DcjxCpSetpDQYZMc
vc6QceGhMHCHlEy29e8ZQ2t32jcIrACIdeFIKDdCXgp5dHl5qcLJaVQ1XV5QKLHR
2bqY6WQni1hfmJjTaWMg+34ufoiEbsEN21od54LVF1kybBdwg1+0xCNqPwbpjFFW
iCOLuER7ZL8bHoBfvBmwNWYY2FvP3lHNPhDpD1L03vyCSjuktgzLJnu0euImoyzi
PJu+5y80Zuiaf01BEebtRcz0wYBno88yEjjFCq4j658SFKInXW95jVdD+G+/VGh2
R1wpYRQxL5OKhQ5ACXjyDtgHMUS82BVGavtijnWxyr/YRTc/WwlT6kE35cCoLJDr
adR1uSPOda8e8bd0Pbgn13vb8sqlSUjTunKJMeptLIEHAfVr4ZtLG4Jlrpor89Fd
4McfrbMLV1pligX+aqHYzUsvuJXxty7H368PrYcFka/qM3uIXCVZpKV1krdRr5Id
tUyyFUL+oJ1+3jJBCI+FUPHW+6T8ykuBWjEI85F5x7QIf3NsfBzC9FiPgk4MndT7
j5qCR/Gn+LjgmeP99mUIf8XUs2qN9JTz2bukgzoCvAOZnltViFkyO+h03TyzWaU5
MFRSHQ61vAh8zKxuKZYhRO5+7CErYOKtdu4lHMBPiWht3BlfCNGLMyA79qOShelQ
Lj0aVgGxlQH9rXMqO4aEY+DXER4JFCkKilgoJV+APrCRqScWNG6b9HpvM1VBZeit
/THTl7RqLTdM3cPVFcjX2//jNhO5EPeEyK3a0WXpbMEef1k5+iW/wMGo3przpd18
8t8RD4vQ9VkOokrl3xKS66SYZCZZ1ejAKjnDRj0ygbP9y/XQoPqqbnU5fN08nJ2W
WaYBxLp0mm3FLFWYLNPEz9kOQ50/MGhkltTi8lDV9EObmv678Nqn+jYCRvd6f99e
iH+orZiq5pEbqbr9KhbxroNYeSNGPQ2ovQGOoC1Ux2BS3NdwLdK3WD2MhO9shYfG
2dJS0PII2xOGP+4dn1DS3k6tzObGAqVeEOzYS7ruyR6Hvv5KHDmoj7xMsLi6fGjM
KCjDzN56R2Hi9CNVTFaLvUdKacoJBbshwJhY+eQZFyyJaL+KjdOSxd7QC99lr0+y
K9O+HtUe33j4HjCAoDErbkMucDA7eThSd/p4Ofz/+atRkFYoPI23XxJasJFh/Td3
/gOJqM9wZilqmnclMPfPEz+eO8WSEsERjKDGtA1oYiKBh77x8VcAhSXngxuhlhV/
Ll/Kzr2dOmM8DZCMdtZOBdVs75w6a+4bxKPFVWiCzvpdSf1reyXFWUl5NjbMfU/K
B/WYHKgnAtN6TZQN0orZ7rT26ju+BEbM+v1XzZUlLxvi68xLZhd4Fp8im83waIya
tUh/uGzjluV1Th6NZm4UFknvLMUQg8p7FkOQIA60oVrepGSgTuIsG+RXRKwURcE5
s9UgohIbaJGyb/Q0+MP1xFh25EKf1nZcR89DX9HjGfHyu0bJxygi7l4QFVwfXSID
VIl7dWOPkKQAZGhFHHzK/O7PSt9bS8FkSpIEX84BiN8XdQgh/LaP1U5VAaEg0Ob7
wdVry2kKSPniJHA/D6tcbqnBKDm37CBuhDBgnJlAs9AIrFsAZAMLNGCbLHp8gANE
vBsK+uMBE7brTkcddjG/3usHW7jH5EBcf1sChJFB+EXAZdAndbcdeujVlGBkXdcT
YKi71WvsOsAnhBQm9iDBGrrk9XdPrz3YC4+jAAMTt3tG0V7xjPjPcLjTCQjzedC5
zxc4tD+9v71cHHphWEnKd9ujJDatxND/PrOe2Jc6Z0SEFq6WOh4yiCx0ETcUjJwc
PmKXfl51dyj8XGack4M2VC8waZNwT1dFh2J/0y77p+BtINW29nIddDaMRoJSAbfV
iACbY9ycSx8tdZ8eM14mGP+Bs64WQeaqzGlfvCMNJq7sWLeWNLKvpuTD6bIUU2Wg
tZldEOmqMszbIrWpn6b0I41CVHH2xdD9CtgEvhX48riwCdyg1cRCt/CMX6ult2gx
ia/cZsPbYQcr/x9p6flHx3L5PbiNnHVCy6P2I5LAnfXn0GfNRW7nzEgaAq4gzbNB
MQhLxsUuU2Dloy93C3W6nnuKwzMemuRGS2/BLhmLI731G8qeGRz5blCBtibOd4f/
xNL2qklkoU3S65Yf3ujotldSwDvuGqrA/jtpp8braOlQeLXBxvjnoekzYLhvS9Rq
EbfgkZR+CwCbjLm32o+SVPcaeaiDscNRjmvcKnxRuzENkXb/mPUPh5eUwIrxIP4r
kmt6kXkEFPKoRr+I/MwWSA3Dm2MLjBsiMOcbfA/QXDudhk0oxcCfdikRSF5SkGyU
ZSd92sv1sP+F9I5UW3zeX8h601KOvSRJb3915Tf+TmDX6KdgPBQuiZKCi7gxZEm9
paEi/8LT02+LviikyDvDs+QUxF9XtrEtsKN2GgpGLgtTGvvLmS8wQYzDd0CHONGu
sonZh4BDP1okoKw2XlY53gmYVLiEUBOqdkhF831z4PCYfZi5XhMsN6rgTOD66l1S
nHGN30cLay+8wGah590jOu7fIMSb4gXACPpBngdB8x0EBGtpAKMWGjQnVS6dgs8A
C5h5+F7ZWYdy+bpJiHiO5VIFQW6w52BCvhIuFWQLse5c8ImQwXgABddJczvpd4ku
g1pyM4Rgneu+v37w6hiorNuU5vVMm1fm+fqaBla6Ebv3lrzDqEafJPsH6/BbiMhA
KvXETZ/Urr5FfjjqL5dl/yvmCOpoecJLQVH8hfXgZC+1v1omCK0I9VbpTybIIqy0
M1jYOYDssU9D7EIH9BBydFtHrgtYx7/GbTjAVmeXy4vm4yfmOf6p6lhEpJs9G4n4
eG9cYbCNFkjZcZpgxk0xoNO/f0U8gUkZ5Y2uD1txNKQzuunoX4RicHwIe5J94tl8
zZuQz7IFxZQrxlAgEnlm33ss1Tu4h669wZsNAYGGmKubY+My2Pl60bCPg42bj72N
j+g17Z81EAgg3bSkAxCQvCqUrDppcHrRCOIb7r9s4JYNPdrwDJxgR+Xcf4gC8v75
RuglJo6a+DtFjcMG+8piz6S3Vy5KaPtA27OjCMU3GUXdSBViEAKRqElc5k39mUTc
ZzPMfX6ODxbNQS1NwOSbssVk37JP0Jcit+SLPx+E58Ybf1B/hh7nEdJ0J8E3GhsQ
kYRg6imbo+tGhXd0BdlBYoi8KtZxEjqSpc7j3bYsRC9ygAae/mp3GriTadn53wg2
tZZSxeEBp6eKJZqNV2Y1G+ujFjycBAoBP0z9yg6iY9OQ07iEV6YkjmaXmQUxSjMQ
but9+/uJCEoWBHzZr5Ftxpd35F9rWKjHY86ZUb4umI+vLtL9dfIjSXke0lBaIyoC
mkbKmB5Hw9RQVatVgo1aHhGczMH5DaLkJIWPmnFizt5yutdQEnbGP1G6+joWARN8
K+ZECUnXn7BurKEIVna4gkH4F4SfdiTUqrvjjGm0VKm+iQQRA1GfG87voEgzhrGO
JcH5E9FrWPmz5uSQ0gIQXTEs7cYoOWNhr5agjQQAvDV71BLOFebXEIqI2zVVhhbV
X1LQLsOXecUQ71WP74XpCy1x0FfODZbfSX+2UyQIFvhVs+tV0xgARd+VlPf0WOIg
bnvcwp7enMkM/465egO116NVz20U4qH3fj+woPv3N5FaAhVdcUouYQj8g9KWZoH+
+N7u2Ukf4Pm4HQzOnKjq3QvQbkqhHYHHzlsW/qFmy2iroyIiONC5joqdajMy87Lq
wblV17wGNLcdEQZt2TAhCmn2DlTn9BqeXL4th/MhcMMkVwZnxCdAyxCwrMsCI/Tj
C/YFMk/VaIBMBTgferXrIK9zL0jWtMaXOq3h/ofO2DxpA7ssmQQCKhdZYA6VVfZx
jHirQLQ8Ls7pe4owk+sCIqx1Zm3HFpmmzIu/jS54PNs31Vi+sr3HHMtlWjsLOS3/
wv/fH/xmmRiEaGKxIVtEiN7Af1N1F/2ppQ5abkJmOr08DfImEL6dzdWNi4LfnuOK
cW52tIrW5WXANqP+tVei5lYwzEaoZSpY2RLVNaMsqatzvSn/Du7KEdEAd6WkQKzA
FMOz94cxMEMFiXEuJ/ctsLYy8gUdtg8QD86gGR643R0KCq9q5csYfYMYz0iTuSzM
8LbAPgIzwvvVvob/GWuY/gVvCmgmItwe9/BedsFyRJ/aiS5IHWkBKA9bt9Mp90j8
NAgshzyysrXNQUry1Mh/KYGwMDqxncZ0Y9qQCB7mMYVQEVHk0JIYMCcAvWURnMii
oidVi+E51s9N4wsd2jtrpjpb80XaDnJeuPqu913bxocnZzXoaLLOJIRXJRLIxt0j
hQLvbNdAVzs73Qvq/aHE9dkksNY5dGusOfPIMaNW1qHUXyT3BfZ/son1gnJ281ZE
K2gat7XA8hkDMmRPkteWxdzsCqS3BVPtrxHwPeueyFyx+pMHwaF9t/px3u+DsHOE
7oSAVX4ws0IWd/XldrQHOZ70uVjVxk0M7kmY0g+fV1KaXpVmnIkPyIG8S1W5MLbs
HXNVuuJg5FX0I/OwerfiTp2uJKzwT9v2r1thYHwM9MZyaBRC0MdoXT4blxmSnsFZ
qoPRqT8MheEmTx+Wube879/Cou1JLwU2MQffZ+Ar5+XetEo8HOpwQXMGBdSTnGX3
HyYITKYK3hmV+uh3GmnD7GdXFpAiS8uwsLxgC2VguRTkNasnngCpeZYQBf35UroZ
KmFqOtp4l791GmvcLd5uU5lX6vvtSuaCPfNzj/dkju60Iivg0Z1/LRRJwssVopIo
FOSYaPUanYtVdEeq2ZxV+nWE5uJfZc7TSznAJjSjTZhxnLHquWVgCbjRkGsnnfmB
SYFy7ufEY/CL2IfvVvlHywQoP51UAW/PjiZqThCslI35mh2sm+QgEQX5TcBX6lds
v1CIcGbzolB841HN5ylwnuS4iBCY1X4EMW5HWssBWhJvGi5Zp3hpD5ULkczLD+fh
NzFaHJfx2qMUGXzqZt+PuP2w4ECG9sZMioYgPuWQn5YkYOIcckzyQDL/cyuWq7vn
I1iadQQVxkVLobuptvdWuiAoZBl0UAZyayVNG+7UHxQckgnvzXHZucivTaLr2uKZ
to7by6NxsIEMyMiIwvKqCEwmiaXx+vEIVl0rvaqBxdyV4x0nnd2nQqycLCwVeL2u
t38al+w66LkvCfGYK7iAWo27ket7hXEtwbLOleJ6yXJ1/pEI5pZWX4W1xdslGjFP
CmfnY84dOQQMbzUm8snUtRhFHFJX2C10bozWrw/QsR/TFZEZjIYpqxmD4e4rYdjb
5rrX4RuFBCvc7iCuzyQUMgqDYhW3I5rWnmaKfnpMpx8GBvaTdAV7BAcwelOSTeXL
Y7NhOjOhrjn6yNqx7jxZRM6SLPax2hg2DOXQBBUHN24PSjML2ZqC7jBP+VKCjjth
taU2qzwvx+PYrsE9tewtP2uAgGzOsVLBTCOh9d+YDIeAtnUehTzjWH7SOHsb8CW1
zaBZ1J/LkKLfrun3Vdrg7SO+GvM5QwhwEeAU6aFDpVgB+7hUTqviYM+yFAlYl/Mc
bct9k1D5KFl+tm3Iso10OnvWvdE6i/+KomJtKViDehoambEDS60h4zLiE8pgfLKl
McyaDss+E2gQ83d+sK+pwjHQ2sF/jbLY/aYycxKqU/L9zmCDV73MwfajUUVXtiwa
h/7Zi1EvtLDlQpL9PEA/kEEe7WHK95U0kgbifei6Wi7unFYsPj+9mN763AQgofmF
I+RfjWvTDWuAtSUqys7FiHp37xADOyyPtNWMyPot99mj5M1elkNLOgwT3Itcg3kb
rLvuWPfMFO8OvDLLnbq5L4xz87tcfsrZp6oMVTgZ32j5R6uhChjps79dUPlQrR8p
KDpK/GgE9S9Hv3MFzIx4ScdMmtS1x97SXitMXbq7wF50dH9We3+b90WxOpJ8YzuW
05xGdrj4z5U9WJjolBdXsH+4DLA1K4XroRLXg5ruLO0Wq1xOuBgQeeKDU/GIde5C
svQ/04ULb1iKZVFje4ZqGHcO6ycJy8+2gxAVVvjQQtul0i3d1DiI/zeXAhbfhwbU
vMmOpIcv7iKBCNxWS+c4iSS8Vx/BkJjDUE7+gPHjqJMh0A9XttKqZIZYSLYK+wBJ
Qo5RN/UKD7PqbwjQskLyxom0YxbEdjprOAVLLc+IN9GJVE7D77+MYEycoCI5rCwB
5O9yb/KwKRIx7M8yCPV/j7W2x5xbenMOOgBdEVdC57Y337rUQUp/YA0YZB+rwMSz
OkckzZmFDPQZxJhTJWzVcOIbpaMVzn0VXGAc0BosO+fMuSLlWz04BCsgE7yFJpiD
oQQWz0Q9drONo8Dk9AB3tqi/HSsaFUwaFBv6mMD2T2rQZdIgYeUbEhiFf/NdfJEj
D8JU5cRMoQ4m30zpiE7vB1yECUigdZ7O+Hc1qqgzX6iKU+thUKlNDhb8CsgOlf8t
cTHH6AammfHi+qutElWBEAtBJ50NkIIk1S+XP6nz2xOijkqaygk+uoHtUQz17R6P
2gUZ5tSmluPL6M1OW2h9Ww9rtn7520n1MMmYyNvsHQ+ZQ5Rs/64bsZb//M2mCWJV
anhn15SKTIziwm3W0rPllo1nH9I2Ppw3o0fVdgPfWZ/0VcZYUcZIWlI7hKedd9/u
y7eBIVhOUWoTbR4Ga4xehk80DrL8xZonse8EiKt0FHH0VxgeGF4C5L0bGQCttDNV
+1cGpiC32j2Sz9qhbJiFhOT49vxU5chQbqfbTKanuUL8agHAGGAR77ONBvNSjBBu
MfmR8Iu557kmXySjxBDUvPqHKGdk3GjDH3F3HQ+gTXNettNrY29zQhNF0Rczaf+G
hRKkNI/XpBFISTIesVK3wv+qdEBC0tNMsNTaf1FK53nm4pw0C85x/lSq0NBD9iet
IzPHWNCzGhGU/XIkXZ1bYBvdIMMgRq3FskX9Eh2vzeGUo05AhGklI426zXZjpZVT
89uD8uIEX4PfPuf46PoaOVMHaGN9Bquw+0//lEcRDSP//gMc9eABkdF3ktfrNtiR
iAgCpE59TmFb52MBHXO5MZ8SIhPP3wuYUywFTORw4opP+4gyd41ZVQkcT9Z2m3mN
BQR92jNEIPLRdseWzhNVo80XLsT8wZHdPQGw+mOgEiv9b4XTMasMGljhWxJycSOp
HGIpeFs7gQYykWhR4dd5DhI/MeC+5gCopNN87neVNvBVbMn+V7vD0nx/CS5E5PVr
VNoQtn7Zmd8WtKpMB+8Iw9wVXDyIatah5O9zkvTXcvMGe0AM6gsLMFPB/p/VahJ3
LTHp7doelKoMe9aWv/p2gG7Pg9Vy02AGiNF6Zu7jVD4AX5eALahGOXDXOzhaLtIT
2XogCvBuhyd92A5J9sAKSYHxbCNPoatRU10Ca4WsG2HRKe3zUinzu6uB5EUceNjQ
GQeujZZclLqyBa+ZWbn6TAuY83n/+hdL66RWcnhG1uWAV0O/2sSBvUAzv1V9P7H4
IL4O9HWmlChjLcLuWJIFrJJz/avUN/YPcAJzE0ayHCnxyuk7rJslgPbEhXZge2Qw
TS43xeiY265i/nvCs1yYt+S43duMx8x1z9cEfYvNUALEAKXKCDTjCTuXaz/Iddwq
eUlx63/SblJayEPfZl2aS+tBif/TdbtS4BpZlSaeA4hFdFq1iOdmCMjILD1C5vAQ
/kgsgXrm0rVq4dxR4Z1/oyTKxuMFzssS4U9OgG9MslrHB3OwnEZVpMERyHdiplPT
ZqpXlQ+q08QKpaTcyEVYBO9eK4778xB+Sauj1Cc8w/VBq9iv3kLwAxpZQ0xJR8iJ
BAFOMR1w/ysAVH5mR7rLrd3ny8nxPRXBzk7giH1IkDayQIq65mvsH7pKfffN2IiR
oJoFZTXnkeayQQU5tMxM3fsjaiyqLr8b8t2gUMsu/Ojo2RjtwpuMGTFRAvtW3FU2
PG5kTfi/vgW+hajs2alqnyzWyXaQg5+AV+2VrxCQ/DFGGDrsnAiWeR6XYObmgUfj
r6QGCS5MYw1fmAThI6+PzlK7hmrtzDHPBeg86uxK2D0jZtGsYTi9lP6fqWeVMeSg
VERuCy02RMHHtzH6v5NlVWU3rU1pXuA6HjjHrJHeT9vqEoHINXN4Al6TXmj3xHe1
jPlVdL+NE8gqadrDIOVIP+hSGIUGX2D9KpjefZ2O2CJdtaz9N/dSvawejJBQKaI0
+Lx5/xxfbbE9Lep3ZYLClRgpTLgn3RlzsFdNSfrzHKvz2OGjGDXyX//ZM2fHpW3A
rT4hyiUc0GqagwTldO4N3m96sIP0K0KZi3PxzjzSgG1Fx4xZLXBLIuT1wkHjFK+1
lUA14/ua/v/EwTvFqmxrYP5GGWWBKTQ60TK4Oe6HDhHEgcMmIwxfjEwoAB5NYiNF
Fvtr0uLorsQ3XyaphenzpyfTaFNFOet0ppsshZXewdPL+oMHDxG8bpGnLyYSeZBM
lS+UGvpkgPTN+mgKo1woKulG7DMkR8bO3dK3J4Px2qHEjh/mkPFWyRtmE5bg3UT3
5M9k9+Xgm5WWf3Y+kPrXdn97+CtzJJPWmrHsMxWrGrBoJocCKbY5Qtz+WKKhVDi6
XyCEKV55XSm6fwv9TcGX7d6o/dKjbPO3Zf9R+/O3R3LkJkSq3mgCJAp16TJb7z/N
76Ju+/oft6beOPRMLX6xhLvQtLIPZPjD4tWMoob0PFOOc0JONAgDy27WEhuMaf8f
kWwGXOPJukjHSldECo3xIwnASynFWWQHdTl/W57nUXD3sqR+zzhzO//aUGPD0+n2
qZ3GT/GD9vs32ksIarHVny2Swaip1u5uAnX0xbi6BmsiImshRHpWAblwdRQHGbVZ
H16GkmMGflfAxK9ExP039jcvvWL/GEkH14NoZ9sJaWuFITkiU6aGUVQTezBU9rxE
1Dn8vVC7YqZTWu7ltSZEiqfp9TnxepzO7+4BIdILfBTN+dJKScFI+XKnTa12w4Dm
WtWZH2zj/te/CDrsaKYXP8fWvo3QUC8EydhzHF3RydtCeouzqEHnKIA/L+MmLpWj
heY1YeqTLNACZlKh6PE3Zyu7wT2BugIXnnhaX1IJEUava1A1y/uzPnrk0QyIFFsd
X2fK5QMCIL5wXlXajGTXIYxlfwf8aLi9yeIqFCpLnKUfuYMJN6f1iE/5mieaHHOo
8qH/kphTNeUd4wnNLbWb34lI2xZqr7VutsIcft8BIujQH4aiLDfLfWzpNHlNgEYB
il9SX1L29ydqRTBOujfzDL+OuheNFuMX+A9UaTeVVNHP8QV8hlMycFiRjIS2oUQ0
9hCoesUNP6If34vlhYmuwxTZHTdRTGzbmghWMHEd1xCcmUm8ca3N7BaIbXHuEzDi
Y/GAmILT5BzguUwjRI4odj+ca/PaUyLKMrhmkh5MJ5KlvOEOI6z1ThDzPztCbPTF
QXaDmKphH+HoW5+W/W/nF59PsfUhSChf1YEdTf8hTpQimMAwBLfU8uns5dZkD859
T4pZJ1or9aYiPusaIflpy85HKGE5lfhsaXY6SOsU06h31Zk0AZMii91e2XFVMffz
WKhh8aC2Hag2i1BntCDde8ouccBidtYmnKGyZkDkrF8C0gYunGYrkxSb3kGTooHS
cS/G8i1C1M223ESnf8p6tFnFPkpExeJK1sAuYJ7IxjB5Hx/VZ8g/EM8nABD6WzxN
GI0hfE8V/JTRO2KgOROxZ3LWyNYHH2tnEBUsJgL5e+gI9ORXO0pRlChIAviK68T2
BLjriVTAg6ujolXUNuLrGpaWceFF/P+sj9GAHArDf758koAviTy9abSDpeoGUzew
CoYo48ggPNUGOXcCHe0V9V5HNNYhkzPsOx80vufhFYLBVA6SOMaDG6wzUY/q7uxj
PVrzGmLPkEAAHTtQkKT5KbEpBH6NYX1lsLZCVOr+Pjy2i6p/7O27rde2x42EOGK2
xDcL8po5DFHpLFIePCvuP+iYuXjKz7ZXHJTMxuMvZlyIzspN97kAK7ZE0EM7pXxR
rL5ccOeHjoTkf80lgqY96xu30yy1oRIJ7MfbZ6yo+eosLS+5aAVOqS9BmP7MPNzL
wg7HDI8dkx5MoqwMqqL/EJCWLhBcV020Gojrr+QkmRTbhnOnOGtz2c4Aez3sW8ho
q3cWv+Klg5BmeRl7bnaedQxB+SrlWPNOBlP22hP8zUvwFTXLbi8CJarYYRTsCuZv
2FRpiAj7+3xO4UJTsNzVA7we5ThxgUOz0fljgL47qDm0pyvNkGe2SbTzSdoQeAxq
FIqgkOQaW55IhgnuGN49NebJ4zUzaNKqhGbckumvFil0uyqWlJm+JszCCGZQgFMs
d7C4WshKYz4/FF5G/ASCqP4OQWFbIZMosU5x8PKLqN0ckKgFuDyIKMVrshabVCCE
rmeTVFaZow7I0KU3ldOT5oZ4ZG/jb8ZGO89ide6T+A7b7JpvTAuHwBTJNa3lXqm9
YZZfPKu9gqvSkSoAUxPYVaCcADolCDzcmAMvTI9keaj971XDGrgmOPV+yfrzZiBw
obpLw8fvtCulIM2rahb3RDZdkznK65e0WbSVV85YKlnMchTQdDAbPzJCflzbVtJp
nawn176vuSYLeAiUyA//675Sa21XEhz3g4A/xnHcrG+GB489k6cF+sdKOAXNHkfI
xFlgTGLd0KiwRBsj+vffFJG+/vCaVoCZGn5icCg+8hjn3pvMwqa25E9ZJhuMolQb
0DpAjBzAqrXid260aqa4qB7AmgFvotgrhxYr1L3F/yk7HwySKWXuS6qglSum//nt
TeLPxkX8Jsr8rAipjapXlOwf/gFMVIMQegXLae+Sm4ysOi/W0AJ1y9WCLW6aolnO
904yM+XLXbPjpaenWFeCrjq7DzqZAB4DE1UO4mZjVj4CwkBCvQTQXYtc+Lyx7auM
mFRkvbCPJ1hyS9xtjjAHZDVlgVK0YSJeJZb05dUxS0ym8bdxfq0D8CNQHd1gFHkA
JTMjdl0SjivKcoSaquojh1Xcp90D+rKVXoNPEeae52K1jCWDs+Y5YXlp39EqgIYh
/JFM6YJ5K1uFAW6k6bPFnN0q3iL6ZblIe8CUN+dvMNTEXlAmVdBsXFTchOHK1Azx
YNfMqwafnT1HsT0fTxUk7D5k2CUhpxQTaVdsnXl3ENl/o+oKqVzRz4Tj1iy6N5rL
OQaweJdoYIeO5u0VCpCDp/BFzuOf7KEnvOgbqKq/QwDst/fdK69/asO+8Pwofj/z
aETzvLnylOusMBeBNDGZF6UkaJzyc6/Ql5PYEp7emDlnYa81lo9m/Bslac7pEsCJ
Ik7syV0KD+78CFgsQd+bumar1n9Ks9XZn6wG+/ali0g86h0n3minr0RmiAIKlvQE
KAe08yvVKB/ya+/9FHGsAAW4IrsKBzp47TevnNdjMPQiydmzvw0S/e1ml3TCkLs1
ZopYGAne788ms/rWzuCcT+zsLFUKcjUGADyo8dLpQ+DlitZpFoQPvxUs1ZnrBxZM
U46LnIvZ9Z9IE3EMPGVPmgE7wsSax0RPcDxJ4+wY9CTLyGRufInLY93e3zjW/8Yi
GNOW6bmofNADRnr/RnfTEYtGkSTQwO8gWvnvmB99w9KUK1pmuIIIQxDySvt0H+kt
JWifZEhYSNvI5Kj0YU4yLV2Y9qQ+YzeET8VqvBwx7mydg85WrcDZyTEXZPVLS2N9
Kq0QjDiVdVklIuU275lCDSivl8LyoXHMvQW0hEaQ8jMSi1htXa6mwh891dUfaebX
bX5dzsPf+6kVxiW9ArwI3xc7+HHwhpzrw/kWGtFjAufM8aS4PypJzluz0Phhrucp
F+Rst0OQsbPRBi1SVcE4xoR5hol+cia4gYiXkMv81Zwa7vIrtNhJlf+xmtsbzwne
TiYgmi+1UYFNxsOo5VaAtPFTegx2QyNnplnI44GA7WjQn+IvQycsADcrH2oUA6gJ
r+os2cmd6GukiLXB3geVaJh3wTVvNVWgx9Yg3zszM0TMXPDsFRtUrpW1OAMEoE4e
vqNsGectICwetEx2/Q9Kpmh6DQAGM4C/hB7p/Czziu4nE2t1UqwCAEZUnp5HWnNh
vh76T+A5ioDMV4irn8M8XNRRunvy/a1ynkl0E1hc1Kxs6Fl0tGZGZK+tfAXGQDtB
Vbe/W7h9nRUk9CioHy8qmTCHp5mq6iFSD3nqcp8oAcikmWr698q+O4T3xYKaKLSn
sNexT8s3GlG05A4PPgOAQ8Bq0ztoFz9b4b7QOTKfutgSKZNPOEg17HcwKliCUldi
oDYTvYQDoJDTNWRc3RqgnSphKDqjONbEARMgDAvaTj0O1ScvYHwaYCcSN3J5fNLc
Xxpi2mHdkTjhEeEneq/ECBaWSurQUENu0E9+FLZ5kw9rWmttw667GFh7rfekBo6j
GLF7ZrvHtl0KqWNUHyhNnpE9Xdb0CmVbo1fqcGLh3uG9KGyJYbPB3gVMufQeLmIU
9vtHnWlpYzT6wBjDsnAJrHbOR1Z61c2htRhE4LEeGVTCxS/Cvvf7KiqjsY9VhnUo
CwuDDXxGg81eIevgDekNv7UGT5UeHpOe/+5T7OkM/fOrQwEhBu4gxY2uXvNpG8N/
zrncTYCLJQFTkWQkNsKdWnG0ndM6mo4Ya5Or/1DlZjf9SNxAKI6QV+aVpfbnSlSk
DwaxQlBHbuEuXUXyQlNpc4iTZh+h7NXUgIiRTD9CnpW7IfAJjY+7nQzriZf4nYVs
ew/HSc195dH7WmaFL7e8tQ4cANH7OHRrWUxsN9MhfccWNDJEE/drETSp0oCwxiBi
1JipXRQMjCT2ytqPFXMaeO1/BBtCm5NiNW3PspUBhGVm3K0Z6CUE6VfiNhS1iRgn
bE3ANuGDJkoFZbIFHKw5u32xytQQby8tvvwKTMtFdhsJCAzlAJWWtHqKj0X+V7Hi
F35eIaocCNVGugLj3jLeX05NckeFOjuzFPVqMkrGTyQALKX8iwB663LRDGvSrcuJ
jR5d7KbCsa5k6orDUkIbY+4hSMofFqs1dR+b76zJEjnjzJCgmxE61ymQvY4HLNvw
L9g56CojMB2qFcIo1Qtdn3a29vCDh362hYydbdYDFNUzcjSM8tzlGawrQsxsVFSA
koCmCVNCejrp+89Zof3bdOoTq24c8kH22KKmkpRtBL3RJ2sk1Y3xcrGLfFkyji76
8t5qGwfmdCi8sdZ9n4dMoghqK3gNiXOHslm6VDN9Rsvxyi1PR3jy08sXgjIFP0EL
8zOt9XL6nllb3xH5FAop8I+6UrVxBNUhzgGt4M2vpi+JQi3Ft4BoKRmeGmh6j7rn
YRWFKAi/7DuAQ5e6r0JgjQ==
--pragma protect end_data_block
--pragma protect digest_block
H5f7D5hxLU8iZOpULbcqhYisEJw=
--pragma protect end_digest_block
--pragma protect end_protected
