-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
PU5ypzM+dN5vvmLe7UMlfiCiAsiU96dfxjksepHHlGoNf85KmxDKbRIPggCxAQvzIj4lsTYNjfbD
ON5P0B/oC4zEv/vO/dK0akjN8Qj2k1oTjgjF/L/Z6ggJgxhTh1n0LjE2mKgqYrTH+Z8VxLpLueO5
DURCqLNwTl9740TBLX7DjrtP5q7xr5s+Vt0XAE6Qb6bNwmICB1V+Iy78HXba+zpuNPbo5Dty81Y3
KClYW69Lw6lSmmw5LEB/kl3XtXsmOwuvfV09513MOx9GkCZ5W3JeL8lVnMUksmewgndIKjTW5uzG
Fvk5nzIQ6qztsLrjn/Bq2ZKc/P+kXf674/fKRA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 1040)
`protect data_block
XqScTNfU29v2bP07gay/dV1vnonJnv5rqzoAJFrRdvXNv8Da4+iYP1KbOumle3BajVi3e+T4WTZ9
+s7sqYzuwwUZGDoiK/LXcVyCiPpX6ZUO707BPEtkrya87wjqZ6VC6MIR8aeLPTjPC9nFNUCD1c8X
ZYmMmtaE7SWIpH6v8HSFpAshnZjuI7BM1wIXmq9XHXlAo3rT0xLCDCEPAbdG337/58P90pI7L1PR
ydRtXbo6pOJIJat35mJ0FFtzrbl428F0UgMZZwjYzF6gE/tVm5RTCrxQQWG0NwsKI4pGpPgh1dE4
PakOCFjg1RxUMfKXguwCIz0lMuHbzcm0aKH2JUYAnnGdDx1He8h0Ky//7HKqN2JtavmwqT+E1H7d
KmDhGC01QknAfS1gXog6f72EQq1kmxYQfLf1/pzl0gfkzkS9xyrJIwHSWtk1tVFsg9pgvrjaDEYx
/6Q90dGKpgTF0e3x9PkvwANe+iwvcSYTPDiYZWr4HsL73+0pAFeLINQKBvvvxxfwo9jJTxZUsKJW
qajgwCtSTnzy5Wdyzr0sgeom9G16qj/niLTrHvbcAvBLMZp+RHk5J+plTAeFFp2xKvhGXCpdn4je
KFxQkZAUG85UO+0+yuB7upx/6wuQ3h8HIH5rPnjDl8QjZ1ZK98lGi16J+FT+Ff6/gr0+VJ+iLKbN
Cp5Z4xP633qbmvIEsI7r8clIXsd6NkjRvaOsdiUqr7oyydfLsfKve/SQjFk5meLCG3Kbg3weiCP+
hZM+XNWekXnYB4Wb9tjiDfxxX4LxIJgOVswxyqS8TKF/DMZgUCStbo4yXMLs3y0YFEDD+/lcHh4a
kJjErxeZ4kjJA129l2oPbEy6glFU3hbp4AOxQKcuFVBl92WswoStJMNvOSZfCegKbTrWPj5uf0FK
/eMepkakuy6LyZBgBXCeQ6nUJKwf9J2UZda6JOWju6EEkeIgWAZyiggzrRNrKXdVzyjMUHD1hK4u
e6Pw+g5rKzLCT7hxOvgUUX5JHxPNmla8cwxT3IR66J+B4lwj1Fz9aawFvOWWdwTZBfF0/PXL3MIy
QDkS83uMv8iJt5bnnUn3y3kKIw4khNYvMLkqV2nJwKDc8W//wEMT0qSVxyzQZAuIVzO1j/ErmETW
usFsSrxFA40DvTXVGNMrST0Jh14Kahp6pDDQqyLlZL2nT2Rp4TaJvvvJcPclytPKZMDKX+96oXUs
3TCrRkgRVLChGgb3203kJguHSKJOWeWnDz8B9lkSbN/lD/gy6YpPtryD2uYiNTI+RqO5nI7Yaw4c
0ozrziZcF/YyCO+27g8vxgiW8LqUq778fboYqnvI75lRdFjc6uUxGMaduAxyZOD0qJkeVauzDoNj
MvW2vCFclhxYx2FhiaY=
`protect end_protected
