-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
a3wUYXK89ElVEZ7XVn/tbh1P2C73J35KDu1tMF5Gbpqj/XS1h4/u7u03Ivb3pcUc
3kF9p17uuxjkEqD5DrIe7cxveX818+HIrX6u4+g9OVzwRQiHfEajnjZcY7FSoNpY
x+r4/UJQl5Mu52mRjmdc+OFu0nVTRf49VclRI99kMag=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 27747)

`protect DATA_BLOCK
OUaAz8DjVU9YjJmkQn1ys3/7jNXlREmargWjRMNEwwf0muu2yoZ++FoeZZouA7GP
GPvNOwt9c9ptLd952Xc/GRYmatlMMwo5VY3mB7Db9W8Z/fr6zF4qVGf9OokAmMDO
5ZodoyQ1ZyFeT/NfoGNDw7Ihxd7/PwFh8mPjn+GQ7H0+5VghAMh+8XWRL2L5n8zJ
U6iVMIevXOsEeFjZwy0GqNJ5/RJRNKqFp0w2KdGjSDz6cbBHdgo5s2aQKteWPu/Y
JmQzY15ykQSjcArmuYBxqz5MQys6kUEFXtcqIrz1/ghQZI+O0RGJoMR8IsVBXOjl
MuhREL9D0TjsyP8aFsEUa4USZFo58/9jCBfaZaXz7gfzHmtDRQ39w6UlLqKmDelp
euGZdHa5ekFMW89F45uRTK8/8kEJNY9UHNufxJRSUSSaxhFF32QcMcbHlTd5a6eA
ALZC7H2wTzh4QbV/0Yk/5dncmSXjhVwpm9hFIQcvwjAqWXWZTDK8zj4+qHc4v0uG
cNF5KEZbW/U/GCGQ1PK80jS5IrDr8N1WVoOjPJzKli1ToTgpA2rtPJXF3HbheoQc
5/N4iaLP/jdTXXppol9SK6mQlqWi8dinAgfat3rZMeXupXxSNcTFBgfkWUoiwRQZ
YXoa1mYDXiqE04Mt3OvPQ/cHGwobirb6mSFRnYHOPF9i2Pkd0wFNoraXmHtVEn5v
RT+QPKHtXCIcgF9EYnyf4NYIyVJiAloCSWgScFxc/ptqaKbicTzf4m8d807qZQGu
1YDoEFQdC64Aku6iiQwkZFpn8Va9HvaLBEorVNWUbeXzeh62Dwq8fX+EF7p9ncNK
khQIAD304A282SXlAoCHNB+fMl3VIxAd/REfUfOeBU0fA661X/t7AHI8b2DU4I7n
DMFDvast6wcIH1gwmtgU6vwN45MGpEMxn15FDjpXfJw0pTxbBpbqVb0RhBiaJmeR
ZAAd08Lt9rDbGZW2+tJtpgJleMbYWCWkHDBQAXRqERveUMq1vjs64XqdpIzLDU3j
y9qiVtoTi6SJamPTUBEaPX9HdttFuYadnlvBsYJnmdtieu9iwbh/k9fZf7yCRPBU
Wnnge5EHjJRBUdMQ0np+Ls4Q3PVg5rByQGRfUyZtsdCnNJV9EYAuBs5QyVqappN9
ZToxd81nsZCSVH/WR666qkMeOEHcjIamv43qa3SVkn6TrzHD94x5HA3hWPTAO+Wc
vawK9GUzTpvhzi/tXw9Bz0No5C9goreZczBrdVU5ANA1Pk6cdb5OCs8OajHAq4tC
sAMj+OWQhzfpwTNL2ZuATIy3eLmcrQr9Fr3Tux2L17heyMSRtUeu+KJ9fmqKj3lC
CUtTEjUF8Jf58aWHC3ECm59+8FjnvyUN1GqtKsnUJITsybbbZ/aboMcztaqBUbQX
aj/x9Xyb8ngiiuk8IitN/vZdcW0IP3tWex0ROh9A2GyO1mZOeSNa8TSYsttoiKEV
VVWIi2Q1pJJCslBJIGMBPKnVuvIuS/WK09hMzJMCGmi4+6Ki/iSlbRRsnBkfTEgw
XNE75O17d28FD62ucaFsHoF9wgdwk3EKtqTbmOSGpUlD0LgDe/n4yYB0hGYWDOZl
DCcuqex5l7kFamqmQPiHkDu6xP5mbOLMItj0mgAEseZFOdv16n2rHsCVOhaKNokm
lbpvhAygOJ9wWyU4ic4rLOA5+0CDZC6XFhjDtSDGPGou7esHya1Mz9mxwXzDGumc
p6wRmRWCXI33daRHCyaWqm1GPfXWSjkyZDJnvxvtarXNgIj8ATRNJVZTng5rE0tl
C6R1Lv1ULv6mP4llGCOfYUApE9Lm8AEp9jd46/pwKfGRqni/R4vh2CrI0Jxfo/Nm
cFJ3ksyLbCryZHPrNh9z1d3y2Zz0R6XLCX0BLoLfYuuDJtWF+673pBi8JyDoVdOt
e8s6JANNJAtwtvrSzTzdfD2HgkuyEktQUxvz4gO7f/xpJa42/K2KZ9UKmLfnLhUk
Jz6Zze8bjIBVKu6wXQfmim2tMoRliqBc3K2blQSXCqCwbtnNRNXGGv9arrJdoGXG
CUUkP8WvSDrCknAWdtqVeoQFQKyyroMY3+hoCKGpg1L9skr7+4A7p7yGEAqBYF0g
2qcBUZJISEDPrkseY5Y6rN1j34wgdZzTFQslY37ZWZpdQDFrSIz20RZXS4I6XGSa
Fze2IEARlfNkM3CSEi4WrRN1JfAWm5gjpTzULR9HYrFdbIVk1ZErE0VzbjfWKWtF
CPDo3/Pd13a+4dMImpDcuHgDA+QXLVCMougy1dH7Qslgo66J+/xKQ061Scb3mC+M
e8svl2Qn+PWh0m9dXt4DAwLfdjL+SLl/VWzmcIZQQvhnAcSQM4NZBSlaaQZ1k+bR
aa5K4j7Qr7MH3NZ6UkYecql9OGlLJ24bnhxXjWYory17835Jr16Sx50U91ZKyWmy
oOJX+5BkFUCACBg98HNeC6BVBJtz+Ao7dhKbg9GQh/vkp6WkjuYCRVpppZ4p09AW
A1CzRDMgNu4hvZnaIXl2RUoujjxvYTpbH8dxQD7WP945hZANuX39gXv/2emG+b3u
a+IgHt7h9wYUtxo3O12JbFxIXXEl6pgcnhAd+t0O6Ua41qFp8znB5kGJ0QgOOxm6
gRy5Kxt7duWYeWHnKy2AyHmjcHlxiAB+U1Chtyv9IdnsfW/68RX9ksnscoIzGX9U
wd/95e3vsl6I7NqNBk92GeGmoNVuaGS9ikruz1Iw95o/uEWtbroCISnlUxWcw3RH
2FkwHl7hqwp0tTeW24Xo5wy0RB279cOvK4ymS1AY6d7sJUBJAMOssCvZY+x7Eyqu
+RX0mPsxYIHwtLElz5+IlAtwHBosaXnz2o1W0hDab/U0JnPdMD3BPKFqttNzqKek
J3S4/eXphqg0QybSZtqU1IW8O5r4q7r8K4FcNcJf7zs9VAE6GEj2+Qzm+lmOzsK2
ud3KTA0tVUdXeMIEdluN+dlgm76wD8zUfQlyU1b9B6/nKUGdUnUqJfsdf35aXkNV
hwNJdWA68Rswc8qVXsSv4I828+YzToFApbRMU36Bn1VbPP8aZJnCt2hElTsrDuN2
WercYit+tVpyRORv+9IaqzyHSHNMZ6arhd3fBPF95uS9UObWrnXGwzZHI+TYK0ah
hwpyDigEui9XP3/O5cwSGBVtU0pszhSLo/x2m7P2d4EFBcioB6FXkRKyE2smoX+S
CtvRpUWYC0HpMjR1GdqFTXp/8gIJYzgfUaL+8qjK2o8MA5NQPo7ubjbt/sfFlnZt
A5ztuH+WWD8r+yyOKU4KM6fRM9cQbDMjY7SkobWOn0L6hiobgdJhxVJvGsxTAHSQ
ftNJkzF2lfgtHa4Rwh6aQKoHJgnT9HnT/JpXtULpshp5mcsUgFrFHZF1ISry2cIc
Sh9bB9UvhLYT1UQZo2J37lszlYLOusbaQpUPt5XEHytsVVsGQWHUwXsQI/wzXoA5
ZVrb5whrlh8q0abXtEFLKlBagLXN3OG9Hj3tSiMrFYZgyn73XzGLwoMsIQGHUkh6
4gtLIpjmVLgWuudM8T+tmj1F2Wu1boDvuX3Dk7OdakWxByCOFpxwWL+Muf1nMwZj
QhsChpxHmShNw1YL8j6JufzPF4Vkcrnu8pyAr587LMc4RyVjZVfbuGxTJ6xEq7Eq
1p9tuVbKX/zP94iziJuzKibLNMtJ6WFbda4xG0kN7nbwVnUK02panKDo8QzZ6eft
OxznD/SCDZ1gqQPoLrwK7hvIIUS3Ni273gxfJKNEn3qTCS13oCaN0gmKBxEYKQZc
sf4Tpnrq/j0EZ9B1SQuPqKBDhWf7AFcqijQ4Di4eMBNOceoSU+YnCNqJMp8rZiM9
pJI+x1ch+gVccqqoac/Ad0vsXy0ruf3Rcutg2jvbZ6AQT1chwlPf2TPegUiIisRt
V03Cy/czHdG1XUCp0TEIs03ES0klZeCjMOx/7QmTt184vA7EtLhnkFBhjJ6a4EBR
IjdYn+pLMAb+i9GD14AWS8GWfdTdrFUgm3ocpNCd9Plc06MHT8hI7HFONsmi/5PO
gX/PUiCGAUIC6R0hdpL/4NMpG9WL/+ugrTee2aEjXIlXXrO3dUnBJkYP3Qt4Cotp
KtK/DiWUTsraYQQQSkwgAV4CJ62h2zud8ub9w7uVnNxbFLlrFdSSNo95GgcoOuvh
7SEJbOE+SatIFohlcGbWR+3Ax1UHEkaS6wB0HAIHFTLiydiclrmXYQ73ajEH5o8v
CDakem055mu6HZx7YNmBujGsiC9XG3i/35JPB2MjxjbuwSvAR4/DS8hcQhkI+x2l
SvdmAF1HxRwe3A70/DnTeYZfIw99QNRwdg6sJJZmEQruwxMYBVBIxgjARvOPeps6
DgkIJxINAOe48dNKsOeAniDdAHtuiTxFOkrYTuqJlpO5tg29J40upwzKXfHdIdUw
DRfEjSHd1RYRo1DNqkw1rlvJE0J2kCYnd4hdjlkOwg2lDOzwY7S11ZqnyMxoAszP
u7GWSksuRocTr9K41yhBsG2UaQ5eILEfbK+0A0jMqvRdKeN1d6ikPdi9cJ+DJVB8
Izp8ZJCqrCW1JS21MhSSAIYtGmp79pGnAlQISsHxgwhaZyWUmLIoqfzPDAiG5UpJ
DjkrNQpRaU1SnRKX8pghBqws33Iv/aRT3L59RbBR/o5Jh9+M9317SsAInSmP9Ilk
0iRGdhoswkN63F19gRAfv+tPN94Lo1ZGqAWx4WDrTK4qP1+Oei6HnVKdc/lHVHWp
y69V6paI11KBZkX6ouUPwcZux33XeyYCNceisV/JdroCGw6CD4mcL40u7AnwTpwI
BshrbuckpyI5uQMIsNFuZVCoThqrN/KwyRlktuv6BXmmqWJx0zLvfNuQGUfCMhxj
xJahB2YthoPQUrWtQiQWoFxulLMChWUj0A6/mFsH3VYvmjFSmWQp4yTVfsTxky6Y
bmTKpfD6/dhHjkICFngaKrSrtqskVVzOvkXFpOA0ryJNo5lfilpaUGtRp9FzKnG9
gIw+Kjkb839Qvsn5L/UCldjRGzRt2bR5LcAg9iqqqm9C79M2eHOPcW8DqD9lIbdy
h/mb2rGfZjG5aJcksVRLWAP1NLCppLkVOWErEKkT3CAidRxuqGbrhY/ENMLYUmT8
ib8Bful3tWb0Mm9R/pbq2w/6cVAj4KQXxCZhcNKW9Lt0AgKPC/R3wRnTh7g61esp
ViCpDLrtjNsdddadXgHt0tMF9byxUAnCHtc4IgnJT/cZGXGqTadJWxNzLT2AuF4G
cJ4a7dSY+xvDQxWgr7VZafnj+Lvz4rA72iM1OtqvTeJt3DcxyhaRzzVrIpAhP/W5
gIkPYN6Mkv2a0V+WMbjimPjGuFfPfHIV5golEsXQEzbptdR9TRPiDJEzIqtPXO1r
j5WjZOkKLprieZQ88+Uc+GjkcSpmnmNDuUUpuu/PGd5DKwr57g5KIu8yrJ6/nRXA
/7j7omDpEYSnH0aoq61eqr4VGoRc5JJnWDlNky2BrSehj4gfSRJZMV4OUg2s2Cyx
KiVwWR5ZSvHwtJcJagSwEbV7NgfiGnnoNsQYvaYawDOxFqhYpxK/SOO37w96y8q3
o7q2RbhQvYwpV5WDIJYF2L9TendI7rqpAmC5E5BM0GEC12U+6saXx0xmDQAKtWed
hPJHLAmFLRpILPNC7ZOjAbq/448MebB5TYaLejBkdeyX8mutT19aKNZs/wwCu9sF
NWvPlIl6oxiAhqR0vzPSCKT6iael1Tr0QS+Xx0LoEwG5AmpIrnDXR8kikEuHGMoS
QpAL6+i80G5tUNc5p8/vXjfFsNdl5kFW7d1nbsKKdfP8OhCnu4H6N/G0f5KdzLvW
X1ItEsHekbzckBDoz7Izw8FejCNo6spPGpMivFilmDQPMS698r/V/FeeYDl5z7Ta
DRIFTJqO4WyldzKigy7fX2cGK1LNVsunGLxeGH0ONeI8l6LMbb6eC81YG2BNvtqN
mXdg+POvHONLTPzcPJFnblAYx12KM6HGBQMzyyoJBWA/X60YcpXsykkdPWSDYGt3
C0NMlUKvBPh8dpE2kBeqh3Sk4sfKgmG6wRbicSXPwTE3OudG2R2hSVAxDx9UaJBN
wwvNoLGAt8co1a2ukf0FSssw9bJ6hDMa/2ubym/AoGxKuRrky4+o+WPxSGynWNMJ
pTmGZliapENasSM8oxraIYooC9ZR++8a7wa8nJEfzHK6YViF5cNUNXDi6+QcjfZW
D1DOVcptlHoVUtvYztYKOT+Pjjzn7hpg5xIEu4Q8V5G8bXJAfBDNWxqSKyyPhY0y
YZEfPDVLqmVFzVtvHzEVHUx+LWYdg4wfx1/G1L9W9KzX2KYwMQ5t0e5YI9V366I9
Wy/6/odSjg3r0t6nupNUZep7O85BD2wq44Z76fVNIW/8oBAv5EW+4VQU6WgrreHO
y0SYSjSYQ6hDvxrK9aP/k9RbzJq4huoG/ZFaBwlyi4Z9tokQRtbTjwQki1zjEeio
Uf0Dd0Nt42MiazVOXuvIHVXbJDpAmYC7Fijl8jUHPZ5sLfkUsYrJjCoEhnBwXIi7
Zo/gQKHBkX09dMaG1MDCg21r6jFA7dnBlaLqqmBagcbFHpK0dzFwLInCl5ffnTb9
eeJ6c30qyIKYstRuS7JoOxDlsvQq+AHtNcmrWMn3MwEgGKMGnyTiItqtgpWf2DVe
O2lXZpvb4gD6fMgAobnIYqZwm8krHmKNhcB2USk4D8k6GZ9mu3qp/ovbLQjlCSJQ
+eaQ94YeOBHUX/J5S2ru0v+6QNFMyorildB48SRkkk+TfkJj1hVMS3YenUsz9nP8
+80YJ0yKsS621zWTNY6KtOqC9wD27tS0mNXjNRZpng4VJYtWhqZ0zu94AUfEwSRW
wXTvtpa+bBkLWlQMoHa0uQCAtqx69/0CaufyqgBy1tMu6NbiQdjoMvyawqPeDt94
Df06Fokw9m5DXMzKxxRibNHeAvRbqYjZ+qSfFX/gHEkxFebFU2LzSbWXS1irW+b+
IeDzg96SoqdNRKbyOSMYmzYT41LHfji6zgQFe7nKqqiFKcICTgqzzvUmBK01UKL3
+IXRaqrJmnwBOL/q27X+uh9SKiw0/u2N5xG49fOiVcWtjcalBKOpQNLcbNQkgN4k
hyfQKVisvk68kSP2QyUCDK72gaLRon0Fazrzs261oGShGimda7CybODbd9luM5az
vcN9d1DW8R8nlHTwTFSdlyu1JlVy3tYcDwL1dhz2FQO3HvlyP0iIyhMEXq8y91VP
JEky/E0e6x+r73kn3qc8qlFHM48h7+6RzCcqK4nlUOZ/X9W8usdy9t8Xdjxpy+lX
b/+PlNcZ0O6ZBBacqvO0rJntJf4cl2eHVfEsWcUpY2ZWGZTKycapE/CHXy0glc0K
ZL+fNOja7unlqsJ/6anK7G8jKZr14n2t7QqAVGYfmk/iom7dmA6RHNw7i4Puk3nL
FrHEj7B6CiSVpQo3xlQXpzOqj3lGobN4nN/pDqyLrQfa6sweJXys5CHdzfOIM5F+
nolKi2VY/UhSUohqsS1GmGKBlxancVy++CAxUWkkSZhPiButfAhU+BcdgHgruZLR
6WnlsGswQIgeukUamnQUyEXNmlOuH1YtU8FNM2RuJeEUk49nNWlyAJFnaoNR5RD4
hc8ebs2yIMkXCPIGFjfw186M1hzJptqfG49nyJit44wCR01wfmu12ujL6cGH6K2c
qLll2nPo24hCOoHVLv4XnwJOEX3HbOEh+rkgAO0DEsceAFM8sv1pTb3GOHiXB5df
EA+eDDCVUS8B33IElh1YV9Qazl19B/+e2gVvGxYrumBccS9ZRAgV0uYsVFYP/ice
ClHvDCoBciPgTTvXDbHr0/sHEvPWy2Tk5vfrkWBbXqbJoJkKCjuJw6/BNrajgMNq
PNlLXhG3rCq2Ils4y7J6BoEpa2QJc/lBTMC7esO2sLsrXOFbCGNM5EI8+iO5lycF
kWpaNOAzZd7W6b+dy4K84LSdw96cxT8QoNnyLSndb4nv3f4cmy6Jg47N5+Sbykji
tc3chlOW0OgoNW82jC3UJ0HLmC4BCEUczd0d3tHRGKQ5JY2FBjvqYu/6kSM5OwvS
E6lj4zH7blCx6OOg1Xwq06CV5+/nymW1sZzNJsDOzob+q9O57JEDOD3d+QscrR9z
inUuqEMCvNYCdQCeUD4ZL30gAmxzoFRvMsAnv5V2vnJ1CmUzyREDw7Qx+k16co16
a8KhZlDW2Ycg5roki3h6obBiirTU8iIBuLbhxzLpWaq1k5B5hMJVyALQ5T7wBli8
3F/91b13l4Cclp/cVX12w/sKnMY7DrC9uBFw8pN/dt44sHj3hbvO4a3N8TU1fbxt
f8+VbZnZWnN71U6By8aA7q5X1/ExXJrE9wmT7iWCvv1LblMbx8FLcoSjpZKb6hN+
FIK5pEPnbB/HvCcGdq3Wm4kpl7iayha+swjwlZaQ49UWkkRwFflBEeQw4/sKKoWg
8OtJnKg8xhVHtwNqr1jma8VKr2WkQHYlbQnM6p08Rxn6S6v11O/BukmEeV93STjk
eE95HaYZ4bxpnnoxKDSwmnn3hGko2ksG2gHNumlDyVfgkwnp9gGIJUoUzrmME9J0
RxuoG9nvm8DyKb6pI227/HGMV2ps2pG1ejPmZDe3GMeCCiWBB3BYZGl931A2Dzk3
1jhQvd021joGHx6DUup7ubx1FZL7NNZZnkOEiPv8hXYuyAHqCEzUDlqI5zM6BOhS
1UtNLnoFkv3Q6UNyx7fCruhL0hanckmJYecPuZA4yCL77i/cNk1f2ICJnqI/3MhL
lvRjLXiC75zsR+FkWC5tdVImY/Ctd2knUyWstTTtRIhGfbGeamqvQ/o8nvcB96mq
rlCGHUO2YSBMtEYm88TvP7q7b64zi+fy6NixGaH/M/RxAN4umDl5zAGxYNJgUSyV
PmKOih8uTvpZ4ee2gI8ceTW33X3yVVII9BR9FmB4G7caojcBkXRPNrOwZrxOJ3Cd
L7xaF6Eq7Uu8On0I8lxKBbXltlicTPB7nD8mpYei6oQa00z+VzLEUonysLpoRJDH
tgDWa0kuK81uaju2cS6jofQxSjgfEwcRxOzacJTmk9SSCK5QfyJCDzwibr42RWoi
bCf4tE0ONvvcdkbiT1f/KGeE0SzhtsJpEYdzYfdgmwSY/tpfG1LQb1eccTdG9mP3
dDAwVL9LHSHmvIcDBiK2jgRagXAaRNOTX2jgFPCwcfdho4GmCmhbJnnlnOUYgJ4H
ExsXEKbZpZMfDYGn1vIfUj4s0XcCzyWiiwH65O/zVcwF4wCOEG//nEY1BEu8I8sX
2uwMwi9Wsv9B93t6Sc/+HQu/w1/5n0eIEiiWPhNUvhho1bvtdFRHmGrt15RLLNb7
483OIzmG38BkiDZOFDWPaqqDIVBL5qgmMt+aKJ+phMRbu5qQxq3lCGwxVU80vC1o
jTJhEXxZ4kh3VVOt+SDqYLNESiqYSvWYtmwf3YLUygssMwDRJ4njlMtjgqF3J0Yd
nqXnXZXIOi++Jj7KOQ2jAtp8lTOxjDKc2mb+k9K7uoxrbMlCY7sSp1beELzTS/Ne
JtC788C7CLnT9iqfkzdHaqGVmJPWLnDatpJBNJwUWfaPRD7FhCpL0KRcxRqhOQBb
of0FFohKcA5CjKhRFIz+U2p/0gPP365Mu73EtIJitvAZfphoN8hvpKp+NUmpfN15
5znHg5ZK3Af1hD/4s6blD38QBBCIiTw2Cc0u6EypRnHcAz0s5MDWylipiRcge247
JKZgqUCbkx+QTXqT/5zYFssGCqEPXsPfwQb665FuduN0DhCMyt+JKdHgeYPsSZM/
GFkS/8DxFKgXi8anDZsXlCD9aGAjZGzoNXUofxkDL6xD7C4Khn7O5C93d1StrOlo
tHCBBpvSn/VLIQXeeJLOO+YYw0PqHn9nL9nJT1hYDDOC9YguclROs29/tKLvdYx8
e5UDj2JxOVgCbpvVa0FzqA48At5jGtevDBX5yfHpgrQ8ms19nVUG1f1EFut5IiBC
MPw86vtOQ2ZCJlziTu07JEU1NV7/FTyyLbrH4zh6260IcESEyV7xVKkNoDAI2EbE
F1Y53f2TPCTrl42++81bmeD+Ncy8FGfVL635VH3aYH8KiOYydYCQwo4EOlBdpoQu
vrUbo83KZN1lJkKS5b3fxpBnKaMVnB4dRiC5eQTMIgsPZrg9KZUQEeec4Cz7HRJq
g+ODGVahUFMNPaEc/r992oAVbeDEoyBpKroohzesEKA89Mzv2fEf1ziBfz7yD3RP
jL8ZZhDZLNFggdLLdc2dRihCTUGGstOnxI2YDfzIEunrq2qu6/6ffhHGmTSzKbzy
YHfqEcrX37pk4NffNkWnctZvzCzGZn5W1Y0lKKNsI5ZAMnGTt1vdlZANN95vEQPp
YXploVyjxUP6RMz96NyD0bSlcKh3bryYfsPtZx2EVTLa8+Js+G+iB8HIcJ5M5EEB
gc/dIR2sJQCICEj6KDZLt4AtGLIF1ZYtg9zSDiMGynfAxalmB3y8rM4l94zG1lvA
H2NV9RnDxHXQfk8kpUnAyKv/ksgcs/LetCKVnOXGL7NalDI2IhrIyunU39yMkAz7
sGLSqfoB0CEr99/TJhXEi1wCRW/h9bqTgIMX8O1/l1sP5606y+Jkdmkbfuu/0Bg3
c2uEGk6FZIEsCpCdQTUZ3KGddp1mkr8vC5FfSmXaM1hbGZhgJUZP3i326iu/dct4
/aEvke7Tk4V003jK7qiDR/QtO9qZC7eU7A1ctmeDMVdEEa6dx7aNNPdqODL5sFeP
BF+ePRHulqDmBSe6a1efsTrDehzpf+tX+oYpLOZSVNzjR2kW6U98TOUj+bitI+jm
VtXDXaHqOCZN8qx+VGxH19F+j6X0mIbL20KDVCKEApEFaZgHdbT7/ciVFKdIq9gX
/lPHZZElpBgjYInXmYwhrg0XpdNZICwCqMUDS4jKVBmbpJNMsNvqp3ONtRUC5LDf
zL8GJUufB8RovHFeLoVIe7/6+6sLZDXuLAiaxTLjIcU57KodAxMdPCfrkoZJB8cP
uy6SzuxGoV7IB0GIPx/faBzkNtRriLVxobJh5npAnkqmd9at/V6UqjuyIM1U+pFP
x4WS1amvyWuy4TpmJ9XmxO/0xxl66NE8q5YvN6FfIGWY6mMSrSFRqI+I/WFHtrw6
kAt0bmmS8hprn1atmudDAdJmYzI0gC0m1tVNeClH4DuRJoXfCpvj8QeI+GOXicBL
2WolgzudJWSm6oQgOjk/Ay+GdfDlLLiiCSP9OXGrvkyAlm4COjhFvgx/fBpXd1iy
B6YI96kD4uA1Kfvf3zuLKmrfijnfkaaIrMlJPRY+HrQsoxk4E7PmfKj50gNib7oD
PcxF+stuxgfdHXC/f4GDUzwNHv+yVEJmzndeTpn+RpYJ3RD14ILegH+kLdF9An6h
htPFGW2YIB57rtVCymPPBzBYX707Tud0s/rZIPZbteIZM5hscAFRMrbPRIoA9zuD
hX/N1aKU1ARSoZVRnevoPaNsKouwyhcS1IqtkjJcCVaX/E7UJUvbVOAJmCoSj+6d
tKLIC5s4AKsO/FzucLSvpzhWA6ibxKRAHQwYhSYJ0bEwXd2wBtvxdl6RF8JGEDig
UB/qz2vs6EA/Nz0tiQvFObR+5XscCjVsrtaPSlccU2bx+qugFmH4b6Aay8LL++iV
RxRSFg5DjdNyVeD57UtylYa6VdVvdAx/LLYzZOS871Ms4imrCVbVIB9J+A4Wgi32
zOc1JlN1vcbjk5RyWLGvQfGnOVRidkNgyDWvjFrN4343KEF0LBODKDTWKo553ows
39lOkKIcHuY1elcAJ4f9dqEAKj8kjx2w1Ohi4+jBWXySUlWa5bBXFEO5wFnU8WsL
raDFhdOPdtPxViQTJvuDzFN6yAx3RTgqP5GG1yi7jFu+D4AFUTdHSTGQkX3owM72
BWPToiHDy0uzYzQR2SM2EsEuY6udfzK73mO3Mkv9SbMCRb6bUr6prpB4VGUYBAQw
q0jD59z1mWXKmI1ev4jSQEYamXHYtwEGKyoMrcMUz7QJmkq15a4/0xCQpaql1obg
p/gz9WBqigXS/6B4AYfQfvYl60ETtSqbSh/XFsPRKkZjWB9jDBIfY9+DB0oBYWin
DFBvTQpwrkkOfDl0OkGqaCj84pV4qnki5guw4k2kjeIy6wfS4ExmqiPyc1Q8k96y
7yWP/W2DGaQTWLYJPx0DNNJ/MbNM579SafECCPDJrdzWnw1YBs85KhyVBNDb3Nc2
2MqqTSjea1I9y5gC3U7b+A4KY6knjaH42SAcj4RVUogR7jjmM3xgVU71rgq0pBOW
UNB5lFnz42WB1VGnQ715j5tyOCEpHHREWFnPhIrEAuPrJxwFy10WCefx7ApZuSgj
NlUvwPSWDFqTaEhWPDyZIrHlvqzEmHWo2sgpTmP2Lz+NAEhTrBxuETX+/EytMkkH
E/iE0DiOFU1IOuXwF8GcqHyNBJfzdiP5CjYf3XyUCcft2t1VbEUiGMgFxdGuOX8r
7Qalam5EbrEBDT6nUWjwUOCcnr8Xdxo6QMM0acCUdWkBOGbdjbRr91uMtw4/baYt
2dZ6aLYAzC3M8P0S64SzPSnxJ+v8/rK7lPo1T29w84peDHYG8u4fnj/UVwgSLi6p
XwVKXoN0gjOdzyJyrh2Rys6G4N8kUxDA6N67EpiY/eaTQyjR+anE8Bj5/ZVdoC+I
42wRphEQwrov4ZRhBbP/G+Rq2xZMWfJobpqq5XWUfOQhrWg9zP3bsSrIi3FtUhki
2zDzYrK3WkryDI13k5ehYN2N531hTQ/5AKAi4S0e7XQy12fV1ClqPWW0uKFR+vxi
VBoPPOKiXesOumEdtAH7JsQTGuG79WES1XAb+S3Imz5vW9ohKG/8ifeI9xQUg+uR
CziDO3F4CDBNQpw/JkVFxjENXxS9B3JDc+nT/cTjN2xcrl5MvAncZrnxy/ZkUDwX
dYa3z1dHWk1bFwL8Nw5fvldYXvGKOGpkAHt/YpXW23erbp9c3rWCtTAZuPm4/j+S
82DmbiLl6dhS6Don1RL4KmwSjxe28oYLlNAnYgPczIQNsOlBn6qb2noj3et85dQg
rXEzCSWgbaiNZbddlayLcfTkQtjxIqdMlkIvhRasUth/lVVqgp7Q+UaZ7rOXnImk
lzukWXToaKd9XFdteHIzrt0W9m1+st6HZLwr/i364w5jyVXl0ky7nvP/rZf/GjL6
+mIrT7Bt4srzVIT6XgXVSVpmAoIu/PsCi5EI+2gdT2ba+my79NgIVIS94x2tYgYA
bcMqAGb4iKrQJHJyD+/gHfzzgep3bBciuZOaTYI+DeIhNBicaYOBb5Yhciigd6OL
9ogkJ95oaYRuJNpEPt/sN/AYULMxr8sRHl6IHn4s5s7LH2/zUdZQLopwuaoL7enY
rsN5HOcXNpUWhnFwN3ruxPQltfBWqzMzy4/iRLS1x7U2PXnObYYQhjD6mVhchV9j
ozQuvjJQ2q7QmjJBRCRtM+fxTt7EIJa+05SjOXFLsAJTlN+Nmo6sawUI52ZJ2XSg
m8I1bdLbuWjeTDBdWwed93FcZzWpe6nEYajV+aAasEIaL+awL/GjNFUEVT3lDIIA
5gftLDDa7vJ6tAdK47Q5iJVqoJOQzrwq5fgpUcMVhppEoI+lLPi/MBl9AXSJTjUD
Uqe+hDn0wspyuJa/dvQe41xONV59zZrS5+PibHLm8ax3qolS3xvPzgLWkqygoUEk
a66Wh7IygkxtdZz2QFhxGP9+tnnVfKMaLcQrmm65jlAv7VGj+qwlRSaWpnV5AExp
RBSjcuRHnXMJ8krJ46qWMDtlGFRNeLVaMQDitKhWRUpi1Ohm1oY780+JzWybLcby
Q1u4AaQVJNm3ZRUrBbh2nFS+etl7B0tARQKIyUm1vO6VqC/SYursXWk3ytjlHfDC
dIO4mdb9KlM6Dva8xOZdze69sfa4lSDxn2JO7pmftAALDRxzksIBfKDx1rRGD9qK
rU8O2qCxtezJ6dSAnLxKPlfTtk0OYXbn7uCJhX1SUeRk60GPawovVuqWxPTOKuBd
U2Dl3orCIaXsrPHbiQoqJBZrQSLpZBseLEW5m7nJXvl45oGlwXbCIx5Pwd3enWft
4g4sbxpOX2Zp+s8BKyYK3SYWIV8gKho9TYHSvqqQ9m6Qs/8zlgMJqFsNK1ghHgit
/G6DFNaUEkh3mhAYB/rcjwJi4NEZeEpsaK/zH9lE4j1IG2+TNKPdpauWEqzHZmce
CMmeKe+RcoYnwI22qECT+/i3XsjvwF5VL2YIZ9oUTLqa/17YlegSNq0aYIZjeZQ0
0RUPnfucc+h5p+3RSYwp1aIKWfkvU0/K8Ei8BXpa5JJJ6RU8K2hk+8GTydPOlGsb
PcHlLhRTbUjK3Ea1Xympi8emBSepX1L2+4nbeLAWiwdLxO7Ot0oSFAYHfdGDCIEn
iXpq9feVvBZoi6sfLTOQAl1VouBYokk+KjAgrlLIcJDv4O/T/6KnOKEOTEXPG5qq
PWjZ1h1/9tsEu7WvMqynB9JjokQXhLf3wGsiojum6gG+XmC3JjQ6yKqxrRd360Vz
UAPX0miaFE9r5c2xe9qd4yeAZR41GUfY9TAAfDkHBH1k4ye/HKAUXe7gkY4TF9uN
B/f0riJaiwXXHBlmImLkMDOS39984p2Y5PlVY1Biv0AywuuwHquAOrptkzJvgXhC
REMJOlJsKgfDVlkQsRSjXuQsIGt8Wd+HFNF1ELkxuVKJSXH23fMn42V2TvA+lTTM
Bb67yqwmhq52u0ORnxIDrCReEy175rcd+bg7Ro/pp3nl3xvzcqSH96AcjbI2NNuQ
COImY6/tgF3FjZpOLzhI+Bb9sr3bsBCfaquVelnMiUsqTsHHGCE+TvaKmjKI+p/c
FFnl3sXS75qs48oMYc68IuKjV7khwWoLCTQAJCrUs4dyh7m89zWvdqN9jpU/gpUn
qCy45dFGU8b218pZCTShTz8jjflvnTFnW5cJxLO1wgs9dNIdwIkbbDRx+dpPqyQP
tkqeOC1yJwNg6jTGQ+aIkFJ7kKRb48zToAlJ0yJQDMYF8humiGy94zvnfZ2oQKV4
zPFssI3T1/IyBcs2ujSvYbL3tvNmGBnJLY+EksWhlNlj9aLeeSr9P7XKb27oJv6l
qtIXa1W0QI4pSsRYovay76BpjnJkfAg3C51FYcu7X7s8Rqoxu36HC0wC1dtox1Oe
vYgxPaXscH3czZapxdbhT+TFR17UJAgcm0tAhuf79HtlW0H2vsrHiwAPfUc/gg6y
zPVxi6h/AsG2U6rXyBsT0AaNCDc/s0l8DeUAxzukcCq1Uwm/t9+WSU7dUmQ/bXpr
gy+Emfok36UWoOfAAtuOkZaLp481fZ7jmtDDay08nHh4Awa1GQ4q2P4BxNh3P1nJ
CdD/KYrJekzPgMo1MeSTs0jrx77OGN+8BXXwKqrVTG/zCVzNSQQU0A/8GTXOIdxc
V6fBAF5DbGk7oAqcBteA1qxNFhjHWVxcIWbG417+pzuIUZjkz4DV938f4Jv9j3/1
SvPy8uhRDO9xK12r1fQeW/Xd45ZJmR8qAZTrZyrTfNJ4i1/82uWpp3nHUVAzomCy
SKVzEjCoi2JesbT3JVvFJyshHymYXgqz0vEwK5aj/hxaO7X2cn4XNEtPNJYNyxvJ
9TaGgaX4Q9uYAXoJTvM1QHwO1WffjrGDnPLXdPPDCS7uSZrNEzkzbYdcMGtsjPgW
WVu1I+50fjZTsy6PU+d8Rfl4Cl+VxkNoXz/iEi0tbdiGnsu24/m2u4ljZtCwS0Oj
8zyKhF7Qd9AglSF7KAiYrjFDmK9zMqZljBlOVYgxdnKIvnnNkKhrkz52Y18l/8X3
RG1RAdUJgiEs+dxJCM5KZUKYUQFlVNAopulhcjL5BW51HG68Nr7dBFMifQV7PVuz
p5iqk/n3FOvkyO5h2bRpXQ1SoOWvCKThNLAyXAK4+ndSTgKZJSc3woz/xCwHOVzW
hWJgM+jULb4/Xo4Nwr0ur1OCsILPf3TIMq2ArBVC0wAouDhBMRbhArjml+0nDwkP
DZjV6BRqrMm/U0FI07yy3dALFOHpfxA1panweWPA3Qp5hPmW5/Yqad4Aen0/pDU0
NSVTO1BAUEdzTMwdBALJcVZmJqO20HeA/VwWhRkW0fZrKousGOVqip9R2bhGWIVN
r4HcxNccyuNZnRjSXhX4EGzP4DLGQ89LgfFybqLoByG00dUHTwn0snUfubP9G0qm
wgVlSFv3AtvKokGDSssnwfaSBoq42zDAmZh8CAptZz8Me8DUm4MGvUwIpU7pqFLx
rl5Htzez6CNqc2sTdoYxoBVEZjJw30rcWRXy5XoUDk61t9jdD4y5lY6rjVBJSe5P
7I+wraAtiV4W3j3JgoJo4QsGBU7rhs/OYlXV220owX60JlO726k6b9yt7npPzGgY
XQXWH5jxvG4aWbHr9NoyXd9XdCbMYSB3tVz4r0eLSUMHpzTm5+O/ZggSmTnEOcUB
r+pBPTzFJSLOt0jF61/ZW5LgfHLsHgJ3dHZdGW288GtBFH0GaSCz/g+ZOrD5ENBm
4KKT97ZhsitwPyAb6uH+y3yogg1rLZtKITY2mpCgxroXD96t+OqmJoVKQDowBnby
n4hS7xzF324bK38vTAXlCqj7nGwoJkVCMXXkCMyvg+kk2sGKyS4Ic2HVirBVrF6V
YRQHWrmAwUYI0J0g2vBpalVbQ60vlce/o6gbgdJ1l6YYYuPZftvweNNvqnSOLYwr
A/q/cCKWDu1iE2ocQZM/dSDiCIeKK52dPi6joLf+YngZr5zgCCdifkMERFW6jfrE
WxlKb3rwEex4GMxS5e63cPriLJx+22Ru4g3OlFlObsYXGXKeWfGO7mWYQ6qGjUCQ
YTFc9CvxmhxnuyxNqDh5Rf/qGvIC661f3QgEHx6D9pZqfn3VwDGeIiBricD1IBxe
oDNL5R8x+cK6/p7X4DG3etFm4RnAzrp3XjYmXukbfT1bCsl/UID9eyKqYAj4MPyZ
KykQddn0/W5VqDT2fy0ueTQLpa/5w3FnY0nj9az/kZgJvt7opNGHbWcyHgE81Ar2
Wy04Od5WNrI75CAuO+4c7VqKXGSjOmYppWblU5rSp1PDBGV5HE9q5DpJnGLv6YJG
Rfd9SZyob/g3tdMelT8gqhAIvdibQ8SH7kTWQgGwyfwNyu1vwwBBmuskakojJTq1
VY53cZJmP4NiapQKGUmKEe/QTjp6RLHYhUDSXlUPIFVxsxObPbe9E6t+hIiWBILt
wVGtK45Bj30hudA27/MUA77J0sh+kVGinYqcjpYmHZpYVMXkNEvSBP3AEZkmExcF
ea+qMVX42vZxPLQMAzwQs4WKkvX11T/9uCSxwH1iSNsQ8pHb2NT6psfYMaIK49am
OUV9lFkbBzX80Ezi0hjUJYRDciVQ24neFlhMpXnlaEkmQqBW9D0FpTdu9E4AA7SO
MWYqjUEg072cEzU9jcp4B9aEuTWFdpUVT5ZPAg6Q9fFsyPYJKaeKOBkD2BotRhX/
MgfLDX1h4Rx5WipFkT+RIBIWlYSnzWZehEIH/L1huRtLXQUFDhmCPwYGdoFovnZf
iS0D74y3c2i7xhtxAJgLqATOPugPIXmC9s8dfu8zuck7cI6uIpE7V8EHwDgM2epw
AsyNbyrtUmlnKzFpyqS0lH0nNGqNDxb54t/8S8I5OI1NZ7IBLgVSk9hkQiE3m4ni
9AELbKzuuZKCxvl+EwVFbAl280RuyPQw7momMKkJowcR7/RTUEogp93B5eNZFIgO
RX/ZyNTWAJ3IYEf3OAHTTrVQsIX9xoeTeLaJrtbhJXImtucFuY1KRAjaCOImaD0X
gfQf7pPCRT6Z3lo9lTqap5gj9XBcMIoow/WiWMHAaqmf6M2J/CtA+FG8Unbp7sex
zRuAPG9X0o7rKgTUZc6R+JyQdaXfSYCFXXG/QgiUpknRVugHO+zlmySZDTEnE7wq
mikn3xVLx8x5OhqEwvw4Z1zSXaYIUdh7lXJyOcC66P+aLdHrsaAyvFAtjfbrGUSw
p8/YRfdKf3W6wd1HJ50sgnaN+TQ4PeyPTRXCZlqKDryZ+wwTA4yOCT8AtYA0H/sM
dO/feHLt5VUo79hFbl86hMUvUS/gq71RcQwE/pE0ttNzLVjvgi/Mpr+2rt8kFBkA
oYCus5MUMxX6pN/ygXOXkq5t82ZZ3Y4gbdvuChWgAKtdFO16Z+p79WNshRUBZISn
mkNNOTyJDUK4lIkBruInmmr2+BjWFQ8qpdM8Et26PyfYcYh2oY3jZqJq259SxxJg
r0VmKGfGsnwDhncL5z3n0r/Cyxf5LaF1eSzNnZWskwf0C9sudXS1yA0mJ1E0dsPz
/syWz8xET85pPD7Y1XoXNQ9Frm6rZfnWG1UAjp7rp+aK7XZNV/BHpwcL/wfXRX6W
LIUhofn37kZWrDOH6OfsacuDDzu7jsF1XlwldECrwItRnQVJj17Lw4U995Dg+QsM
dC3X8n+Kwd6kIAGpZ+ZWqjt1ctWxDVJghpHK7BPTnFnI/yo9qxIrvz7QFLSuxiTH
6UU7mCF/eAor0pKlfw+vYkwpN4QrNKwvaXD+omciO6bnC0Muy0DuSJPNWLeA74Dr
OnQzsM9qLyfalN/CsqDpW+5bw/hoQn+OUGs2nKT7qEFLj2pV51K+fJX/552DYeIY
TdrQVaoYTsD/BsqTrLak7KgklOMRMFopXg1KBTIyRBzEF51IkWxBUvofJDcZ1SRq
2QY4wI0FZg4z+ccha3J0W5D1Uh0VVqYhqNqA67ugMHbb5iDDpmz2w9RFS70VZCmQ
IXEXTKFqVydw3uEwE1fCPaaipGkvMYUuAbfb3BJRlq3Q/k/mv0qRd7NVtvl1mcFL
IG0eLzBLoVL/GLdDqQ4Wk7NJm0wvwr2ALTw/QuUyK5OK7xZgE3aGf/cjtkYxr6Lb
UJUlEdfZrEdIMY5g8B/INcDz9h8H2dKbYMvhZS2PsqKcRbT48OV/texcS0DBicNx
UkMMzdXT4ASSt1cf6/co7U5NvhbUc6wwVtBTC2nK9pn6+17WTfAfm6tWOW/Md7Qe
6J3lwyLPXJCxxQ9Hi15Pg7TTIt07Bq46rmUmMvNb28M8X64eCSLh4O5WdM6jSm8B
3864vWtmWARGyKsPC3P9eylB9pfzep82gsHI1FrHWHFtMldR0poywYuOXDluIlr3
57k2pln07mbrXRAevbyS82FdXL/KOd/VlhNRJAVYCNrpsuhvoOuA3DtOLVHR+Ra5
lE376psUcqXkNksMPmeR/s4HfMHgOeVwS53JiuwWBTl07V4OOyRWKFFA7D/K+Fbz
3wdXcQIUbdJiMQNF3ASW6zk3FFWpftO9Nu/WUOENTwpeYp0+R99x8WZWXjlPun6Y
O88nQ2T7AezfUVn0oozEtW0+Y7jWFLxaK7VU8SJYC5QO650ku2yUwp7XbrqdwzeC
qZuVip2xsX0v/Knco27bqfQg8Z7+upUppk25vExKYul/tZcOl1OmZ+/R7wNQtL2B
XEyx6RT4emMGeG0dwStb1e67Aj4Agus99Sk5G8D4B2BkLVA6EYel+BBFYezpeV52
X+8L5o4Fv/GGar++r/nqJVo6FTzPcIaD21kTcvyTGra56IEHRWlDYlUP0Yi17MiE
De0aaDB9cIgov/G+vkGxusouDVDkDP67m0OftKY3TUGa7UpYXJr4ByaMhJFacgz1
5NVSHc8rYlRVVVbAvhM/v0pbmi4KGOpkBIoXC64m3QS/opycGpB0w/IeoLf9neF1
vTbSwSRUMFuqqFcwktFS6XmJGVaRFMXsAtcvfzAfseTgSQyTfdHMUkUvAzIGxIbW
KoNMAQyOb8NqZ8RKKv1kav0C0V2r4DKlx62F7ZHRPs5crPNlRF6lHM6gq40F0QJN
vrAgzPb/hSaNmw/SkcPSZytjK/jwq/OBjkqpLJIFWEJUyIeFXckB1EcsLBMwRj8z
3CuJXHyowP3p2960HFfakXmdOkot7bLhhk9DBxa2tCrAkghXmM528+U7ynv6NAR7
GdmeBCqwjnSamjEBys7FgPDuzW6drUNf9F3QuZHODUWlMevZUnRrC5Jy/Vc2sdjw
VcKc8ZNXLPkPyyz2dkvE6YfYcmcGimJGGCHm+2qZUvLIai3Wp8Yax8H+o1MII0Kf
tP+a+qU/lVXvtVIYOcqSA/KeIPjnubiAad6MEtVWekyU8f2Ad9Zl5Iw4Nmw3mVsU
nbB86ygmw2CnQQ/a+OMDCwVZvHp5JsIQQqaAyW7UAbgd/W2x8/bzCkoQqj9rHGlj
Tg8NsuX6o7i1VYrMRi7tnJ4jxU2ccaFaIiWawomejwfUFmTqqGNdsiRnbVhmt9ET
GXZCWIME/nKUKmIR/EYMZ8e6/JShRrgx21ule5X/KF49beSqnJaeX4mATlw5ccCA
iPak+sTg2NiltZc7We4sL+3jYFr/wtno2SsosUv5VHc+n2AW/0zHq6jX6OP1TyDy
9EnpajXbFKjWj0RMXYDtFb2mAPWx2JJa/zEfBc3kqKn5Sbczam9xGwZBwQZsiP1t
jTf7unG0zOdnW+LXGYcgn6IqDi47YiTpF2bcroTrnD4hzlP3v/5P4UlIq+vY80YR
4R2v+kUt/yr/OWIISL8nDffjmvYVtPnkvDBaLx1hBtZB2LhA7rZzDOD2NBlGyxb+
+wocCb+Jj4Y5EiZBlepshwQVPSVNWsp7wsdkAR7ZcBvL7IYM+4+xhXqh9iPuWD3p
iAJIyS75XBom5I+Gok4oDYJz6yQWaeTlXawG9/rszhQx+GArCP/YMcrwUPhjCUhy
K6WGepjRcRCcciOVDmbpugf9Bo8fnBxs7Im7wq0TGK06XW+SQ5YGRn5xpn2ENRPV
4awgtxjrJbXcEyb/RGLT/Ag5k3TNzO0qZ+JQj1Y4BwEHqQsvQ99YW7fA8M6pxuc3
LluajslviTSKmB9/nW/nwvu5gzuJPEogp76Zr3X7RC4qNZYSpVQeIJmukyBSpSqj
GlyHxjn5PU1o3I6LK8J3/ZI8ZxqLJrIz5Fd2MwURHDtybnIA71OGrx4KFlbgQKmF
HavSzbqz0DQO5+cEJmtRVPELLNL5PrgyhJJuT7b4UyrWmmM2x/3ipmu8Tvp4+m8w
3NissEJ8jYRe60VWfS4PdEWHW/xdy2nJM6lgMTcjt9zxltHlQkPP8xXM1f6L/Z3R
sbVn/qB4wg7NZK8C9XgALJGDg0fiBhhx7D9/F1mdtk9wFMQkf1AFaKxYcisioKC7
mWB1WpKhw2isxSw2J35sSQcOgdhxFL36sdvSE0q0Dnd2MAJVzagWoEL9jOIpTGqi
PCCtS5N+yv2jU8mrC0s/Cwtf3p/p8M+ILG0Cm74c6cAtMTcEpSA1YsNVAyThTJqj
i+5yNOhzL/JFvhs4xcmwbt/j6Gk8Wg7w6Wkv/fXnKlX0sZgPSPWlIyWvSJkN2cjn
6+aBtda+g+FXHfeVQfJeDnttGEiTt+8BfF7w3C8orgRIyBnesslV1WhA0wCGSNak
hOOKEBxqdMkrdRKTBGIRWRpRMwRBkYM0M50jc1mxZJDBSaFUneffeWFDHWOeTg2+
UYKiwoxamEgEXvu0Fm9Ayejwh6fZ42BU0Lk1n2EBtYGep3ocg4auuZ+xdFgH0udu
eR2nDyXErcp03BCG8jq96qLP8iw1elO62/a0samYhFc+SHMGbmBksQsZG6tShIiq
gQs62L6f3uWwl43s1MvUFvWdoiKWsmsC3/kf8/EQ6XlkX5f8yzb0z8yUGNKR2fn8
OatpJHFsWgF/5i47YSD4gIrsqgbpL35HGBsn/dFVCtSzDIIkqLX7zpyAqhXJ0IPp
CcseykLA4y1QlFSS3Hp6G3Pg8vC4Z25njYQCTUlz8vs9uJyUFumdK56bDWaQzDo7
Kwbozd7G9EfEDUgDXjo+fStbi9SBmzLbdQfacZU3MmDQOHQFysYnxC/50w5tEspd
FGBdp3v63wjjFt72aqRQN2Yi4El9fvBMUbrWelwQ8fLEQFKoQfVtvPbprTpJ+7kM
/eGMRrE3BOhvEBz7ORxGE7lDm1fu3BPrEIPNh+Fzs9e+9jwR5TbtOX1hxWKkOGxz
hkVOWbgcNRakJybTLszQ/hZ8Adi3JwFvy0UUAq+v4h+z23hJvAdtK4Oyas6Vw+GM
amTgv4ebaTOewWjsk+z0zRy0/KuZ1Frvne1P95DH6BaCWBoxhqTr4bdgDBDWiyQm
zJaB53OPDiF1UJ3dZs5lRVs4t6U6/06WIQ5wrje3tfLmji9oh6bcPACLWL+buMZy
WKW6FhS9oBShXkEB7VwCQLliHkw/uAyJANbiPb5Ggm29R4399coaPSgGytF/8/Tl
pSYZrHBK+VIQRxEVIf5BXk2sZkFsWNNJzwhLVe6SZIHavNL4sYRzi35TQY3Luvnr
jofCyXNg+b/LkRLUCdhS3S/kpKBlwsYdnxhCWUlMT/5e+K/z3e8GZaOcEr2SWMmX
urCqR8ieVXJzkM827wI452qUc+mwJx2lD3w+pdC+8T1XoQDRiPe/lc9ur2V+g5zW
QhmTbyQHbhkQbr7UQbBuu2zl7gNqXNedEaw1i4mlH4W+OgoyDrSGTihpyARkdEZs
HsHiMipPZ6Ercj2uGv2bj7xjtBpqwstwsYMPTzL2ywCT0s7MFtrmCrzah3yv57J8
foIgh6AMOJ6rBakATS+ZOZwaSEqc8EcDHZTschZYPA5eic/xr59mEBOT34u/hJrJ
2rOL/h1WS/k151Ov+dDmwChZJvd9h0XndErqEeXfbwOp/GKmdr23MMw+bKYoQUUt
vNFl6oAJBYWUbv6/Zr77oTCeEh9SJUx6PpjCFIPtt1Rwul1i4t6AI/kiwq/qi2HD
Ll9RWQ0bYw8ydEQ5jBZJN0HB9uBJG8FSRtkKXwOLND1vlP2CfhcyVYA9gvtn8jgD
RtH38RgmbzN6aBA/Ok+M+lGk7YyoWltBKZ1K1+GqPwFw3GlJ++k6Xznge8Afv9Gv
jipRHueyMqpq2vizIxCNZFxvTHC6d+WkMKVcmN0YzCPFCII7RXtZzyd7pzZDyYec
EfyIv4Z1KaOPpw7gyZVmWRdfp0b+VhI2lwTxGnQE1Gyzl3/hRqPznT0kyChAVTH+
wtZxWqxyCqaJXoSqFVYDpHM9JjeG7yosf8owKCsvqU+DL9UZdObIY29jh1Tv/7Gk
RuMENlitU9vTHc7I0jogsZPelLZGkhH5IzxImdmKvH983hQGMaBwsyh7K3fVQDFU
HpeDW5AY+sO4WY05YQ3zVqpoXdh3YSddvoD+XPmeByWexMVMa1p1hih2oQUO7yon
vAhJc0LY0yKq8jQuUfJGYXxRN48PzYHaHG7VmFouQaxzN/PMom+EAlKo/8Syn2Pb
Qn3tvjhDy+RBQtKipyYte4iSIBvht4Xnp9VkzJxX2yMemnVDtQBrrkvaR5LP9zM0
lbYP6sR+ZzZFV36dWrfXyMkXeIuJVVWcVWfc4QzT2u7PR0gJvGMRlieWnfzVSPpN
2YRVa/5BaDX/KusOkEGTVM6HBBcXvnhh7cmW3A2iNZb3n5RCEohF7Eta6veZI8lt
Uhn+dIWpYkxU8a1aDHnYdsAQtTwnMojaYHido42rZrzxcsM+ELEec+QUpl6DNRuL
xos0O/RtVKq6sA9MIply+nTBk5fidAu7Mx7j9hg1SRLWnKNvbnZ2oxRTqzuw63Rm
kq2YB1t/N1wOkpn2n7oQu9E5tqP+4JCMutnWUSSXGYJ7xp0MAecmP0lwQQw3ch9z
9dZI5sLFmlfgbgV0G6B3HQyScuSk6cy/RfUjsfg6v+bAkbsKNccuOt0Vr+kXLntz
rJf5qS3kmztbcOhoad7ujMGgkLGxHt2zdh7la5NIaqlEbAYK++yMm1W/EppWkhib
aX1EsIk2xURHyOPYycT4ufN+jjInwfwsHcjsz/f7hB62EP8KozCDDjJ5KGUll3ZJ
xc53mTWeFD/lrkcoZHzxTgFTB02DdE5JqEg+z1cAK7aqNljdajl0f+0dT7xVYOJf
UpUuW/Htnj93FtjVi4FtsTW5YIbzqFUA5tlwupEQdDaD045mOw9bhLj6hgQiW+bX
EOk9ASYt6I/VtbUDwLVGlJXOsSFX33/hXd852Q+RHYlh3xCVNMUT38oUQ5IVhJ/3
j5aGm+SiTVwg8lDhp842+BnSfvpfwk/K2Akn9wH9TarEBv+pcvI67c5SaiceggLR
k4+sNoZP9r+a3o12eFCuy+UWGWPCUrM8vlNYOov5loAWEHRcGnlPKpA7q37bbn6X
FG/pmZZq3DFWei7Wls28nknlVoqG93iYYchnilZBfxJTsp5UplU/9h39eMuaYvUE
84ZSjd38IU1ysM/c1WAUlhi+r9Va68sT1ZidszlEakbRvYhir4eTusooewVfPwyQ
bbFVKA/HvKDrjar1ZNxhUi5eqy+IPOIE57oSCQy2JqUbCo/HlkUmzvZWqFEnI5Ru
do5//X2O+Csea7/Xj6Ut+SBPwiKPQA2C8HbWeL3M8kp8hfkQKfh3eguuBGEEDqmq
cODmcw+8Z9mR4JdIjWi8IkmaVkVfPGY7pSw9mLZnyWeCKMX6++zwPO0xMyZUzMeb
BmsdyBNmQf5M7fj5r8fAsikt7nW2qcHnv+LqJfAjvYv6cBiSnkSDLQUZ4xitZv2j
CudORnXotZgZGIermwSuEWSW3+z56rGzz8bMqfBFnhjqBEGl2nIQwUjLAOosye+4
hZMPfp+3lRQontsgqled5UWiDTD1zGOU7LHfceprmbnr9FhFqfJDgsv0qbzXob4Z
SzP9Lgv9VcsrTgEbnMsqtwyZopSPhdieHpCyziMnnxsiiRdbKN0Dc9MQYA+i4q49
wh23rPaXGTIcTGYJiFm8ssqpGTPGiSDX+qdaIvxZo2oFi+fkx406hjoQ8xZlupxM
t0FQdadC6XmOuYuuxYrOhor6wnrwBJHzlO4VyedqpWUhAobyf7sFZjfGCHvjEmK4
DR+wTZ4sDnOMLKH5heF0bSOmqOiXXErJLGNeR+zx36WZjphiBtqMHCPqKgNumImv
OL2SsjsMzI1YlosKa4VZA6ftxp+AGnj9/eQ/VS7+5sPa2tKHcm0xas+HoALw33n4
B/SvDwHUJNm3Mv/OtWSd91utnc5lEmkhuqrYk64lCi4ry2ypFh1pNVXt3dt2YqmS
Ncp4Y3MsOM74Daiglbs6ETiCCkide/CuY5aZIMSY3//aon+PwBAv0m5qdfZDU0aL
qXVqIXEYDsBHIaY4kTuVtATScEZdI1FncIDfbhfuzoBLoTcRN+grPhmbnqOKWddM
Ev/SK7km+JGwTYnEvKqUGkX5Ju40V6uP1bAXZOiwDXqL5aH58riqUHvXIPhNHu7m
2Yg9xe/EMHweS7ttEWVKE7Ap0Zo1OvRFleP4B+TgLUoT3M9Z5y+c33u4HnUMPIB1
McnBAhAE53W0jmt3MHyM4ILL2MnC3J+yO0iHthDxmpvnFnbBy2VoxNf657fdVQGY
CVhgPxS6VJlqaP36912vcDGuL5XuYS3LgGI9aXDKy0I1rAA3O3CuJ2Z9qf4p688R
JGUqKLMuEDKNLQ7MyslgGN6W3kVL6PFzqlb/IyFviTXAipE5SWYgF/UqNOWl251U
t87iPuJ7Ravy6mOGL8C6HLYqQLR/dcuu/cTc1f50vfzEpSyPx8LkEuaTVM9asmqh
rP8EVitHpHjktr+b0BRj0et0SgQBKhHuZkQmRRS4yJ00QwGWWvBU3wRzQ0Q80ihp
f4DV3I0ae1+TSfcj47frJolXpQgA/238hR23CNmN+6ICfP+Pr+nuwPNydlPbsVVv
vpKFoT0eA6vhhxJiYjeIVwsRPmHDPfXEeUHkw7d000Dczph+/ba4o8kDUhZaT1LB
OoruA0bywmcbaE8WtohsksyFovYY19CmddQyzwvMzGgn7JRaXahegNDNq7/NjxTC
Rg1swxfmvhB6kRlWXnId4rgns/vrUB5pJzaSIUwFJ6jTioZc1gsOiTMDIsXgWxCh
6Hrnzl/BrJvRgyJ6UReuJyxKjo3w6Fp/ij98t7krQebfrFBQ1CFKqWO2y21Enf3w
Z6e007Ii0SaiV40KOxxgSFokOCXfTfEnR9peMSwZAGJGjwhk7epYICxZ0QrphSGu
nVdao9XuTADTocVPLxRP+LR5nrtvImuA+wL77fOhWJdZI8r1PKu7pk7L0+vJH46W
QXlX9kMwv82hwaLVkDRiikos6wp+dTBZlW2Q6BkWUXMxFl+GW0o2C3hnnkMmExEk
BxuaNtVN1iJmVqygTUR5EEHaqEblAyLE784Y08DqWYHd3akauY5/0LuWrdoVK21P
etTlOH43o1ar05VnoPcYo1IBVjge7Gllfcw34VfGNgakWcsDyb+irCwSr5/8gFPt
XgyU/bpCCCm9B9Cfn3Mc+sCaFB7VbIuettRRNRLfXuckubE9Ll8PRmzqrBpXjYGK
mRT/7ULzEud2Zh1nVihqidek6IZsXkg/p89fK2evIOLcsX0pYwBTaGUCjfd0duU3
u/Q9OKQAYrRYmO8EGb3XRw8FycNhvUUWIkWlanHNdS1FR9207Ie3E9inkn7Kigbz
bJZ9pYzVB/Y8cbnSzBrY7ChneFp7c5wnbylCXfeF3RmitRJvVGSOfCSZXe8RUmBh
m558KStpAE+dso45u1mEUoKD1q8uHOtZZIYuFXxMNI6MKqgZh8e58htDzuKzMzsu
mRLewiROA531fxsJUMoMopBxuEkNBCoakFc/uWsJMmqJYWrCBbikk5a1bNJ/olYv
3yvbA6yrcravtmKg/K1UfmzWzuLQ6etjjxYPUwyIuGt2rGCoMmlKJsmsc9399/fA
Wpmd2MLawHyuiHwTqF09XY/+lUGAxHIxb9A/m4cm6juGma9z3wAA3udZtjtp3zFo
AE6BMSTzCGH9yu7HGqROgVVQn0u4UVbn+ZDL0FvIvAs2cPC2LrOceBURs361FtWS
8YkCvUra5NGanhSnVIJc9cR/ii9is6upIsjAaAw5bpMPQp7g/8/uSCSmOeuGGm8W
5yj+CXNz3qypice+/qmGKJ4Hnd7kiFarhfCX/bEaSgxYglz0XL7l6qEmHlEZc1tn
1PpbBjh+iYpO5/2u2mpx3vS1YUoYDh8ZU+x5H9UD75yeiidrKTZv77+tmxfNG/Po
q8NCQFuF7wgkxJPfETBxtLkGbigOyU4fptTaqvwXFobkj1r448pwTpQce19ipNuI
6+xv1fc7CsXahKcDXJoBoO+fTJ7Qoh8PeEzsYclE5xPm1/an+dSKlxYbnFkPHVB8
MCOLzHwj4RhW8WovNDwYHDoKYOkpU0RIv5Ra6kyguPIqEkb4Fk10Q9mMxC6Gc8yZ
JglzdbpDywnb1eqx1TOiLU+/bI0kCzqly8nBszBX1BUQTiShxdhkKKCZ5SU8ZRoE
tqX4l9xNbkOxx6dCDz4Dpd2b8j9Vmv/TlH9pMJqoL+iYSMucUtmE1w3TVNdeNAmT
L4kaCfUeX3onaXDZUXvSUddTFptFrnR7ix5dlMqGLSgLhcIi+AGxg5WyuVHVU8KB
iuRK1HJZX8RZinmSCfLti8/LjjmY+iyfuXkFiaH7wsvZwWyiugzV+RfFaBerXuJX
H2G42KC64JAetGEFEu3ITVRSxx6pLqvJCph8e9GExqLKN8GBITMPvCGT7+Fa6SKe
vVm7kuGWkw0CWsRavJFFSCWvTyzaPy/weX/KU91gP+hSFC5ZnPWbWN4yAMVU5Wo8
PCDNs3GCjKDXb058yaElr4ij+7MStsylCMVSxrEZV15zIKbyXmbGBdnjBmEXCRzE
tP+vHmdda6kr9LHwBWF4BN78/wQVp0CMchZoQ+HCpik7j7WAPE/MmCh0jxDfaKx8
mmvXvNvySX19L7a+hIok3I7/y3edS4SKz04l80tOry4D/vO7+9++LfpuRsNDsAqj
qoTUWITxIZJm6206BuRb8xk0cAoClYUEKMwfVcslfyGuroi24HMDuGWpmYcm9bcS
MKmkou2GSDnePcnAlA6jj9JIYIm/AK5rYEOODmxRP/poiJDU5NhFsvQGOjX81VvQ
ExGiBKCM4xBzuaVRxWyRPCwuAkbq/gT6ISU5KAFLqJSOaP0nGd/gpwmI/XOYRuqM
atg+UvjDmrPN3kg0XkkpBHVtNh6a+nheIjvKE/NEB3uYbkNE31vBSAF0Diu+KTZ8
k5HoIpE1bAXxiF7TVwLoSZfz7QNO4RDY1lCNCn4okarjc5Q+Vzfj/zYmL3ZNWV8+
w18MryX0vFUykJHShhdXVSe3bVb5/WoJMTRDWhNujp/zWcadMiJn+/cJ2kYrucT0
q9eRxZXVJjJ3Tohtb3I+pZ9urzE6/R4u6t4d0+5R08J9dzY/t6MSQqVxOkGDrCbM
42Cl4gG9NY4Ffd9dVimZJviUYmdAq/vnnUqrFrjKpvRHUZ85muA0QJD23soDHkKF
rTKmPVXTIp/eewuFxeOTrd9HP3pC0iNSYkdidILob1EiL2IwHAWO4RbR3Pq9ucHY
QwDQm/ksaoN8g4v3OSYDR5Pa3U7i1nRS55Ghbm02ECAnSLXsdC07YyD937cwiH4m
wh2sqlKxUDaZye1yCGmVs2lszu9G91RxAxqjKzjEqYge/+cRdwt0ZpZMDBCZjkp8
MKsahnwvwxKc6E5xGvstWp+B3t5WiDrCMOYdBJdTqj6IjMf7f6rDZfXRpmJK9Eb7
aQqB08N3Jt0uikdVy3rOzar6FfX2CmbGdlc9X6GJWtiHrPSkfkE7jbLY8OGoktXG
Fv9T9kTxYOBcMcs42H3jygb9yFmXoDuns+VVcoVctH3BMWTwUe1aNejca75aRiYD
K1tKjJ4Ta5n2psf6A6cBAZrlEStA9C97w9zhbXe6lIatHM3Hz4XVEmJ0nPX/7FQ6
tjS5AVZZs9Hr4oC8OBiLuclMbZ2e6SmAmsa+QIQC5SvdyqkNQMZFOxmWKPq3E0sQ
d/83/GQlw+/gQk5FND0ydzus+/ZJSxNoNMReJQTqM7eU2bq5VhfPRCIse16/P6aj
kLqdtVE2CQfwnqUmQD97DB9NzK3nP4Lb17urDhqrD1GKQPvcKztdrB8YpLumjtJT
LEgS+nZmIJm45uFdItmDpWWevXT/2HxPnjaDZdFbBqbD5GpbsD8p4j1963PrWjJ3
d7+UIexkrEcSqLUSWzSwCqrNJQmb70Xi5eKelvVB439OIRNqbPzC7dZ0JJLaaXun
wvTmgzBBrWTmybeuqvGIKswMFzAU1/wj/PgrElsDjcLie8EUX4fSy2+vYDEDcoDi
4iAfhExCrTDMt3SzxFOJI+obVhQJRQdl89H7XBrKSXtXJoX5I+7l8q/WJ/8U1fvF
5vl8w1xwxOu47pFkE2QOfHjfdQSrvBMNAFdfmcuiLdRI/M+NuOn8NvFzo0jY5jvX
MjgdwolciVzEU5OZxMbfvqWWFlP8SUpO3kDu6GQH6HwXfpG7n09LB/IvbyhJOy6d
zrGZIOHgoBdUD2bOGhI/hUuMxE/eXa9931UCS9mch+n07rmiUgSQdh6AvAGJOXuw
syNvWrNAgTxgr7esTCs/Lc6VyCPH6oEkskEX7y8Fak9pXxA8SsiuEQXa4EQWKE12
hjyJrpRgYnGRDoWuwB/aGitbmY9GGLzGGY3RCtX3B3uq39CWYTtA7LzcYPvjeBL6
g4i579c4Jc7e6KC9Pn9SVT2UV0ZO2gEo6jDxpablH37grUN94m5qCOQ/TG9gfoFM
3tE2hdioHN+UHvi38mUyW1CMOd9GZPYI+gecXyLA0t9wH8mVyMq88Jpl5WhmlFVe
x20uXZYsva7Mm7iTKH9rUsh4uCblsajdg/4QlvX7mMQnaV8XfRlzgwvbc2rJKiWs
ySqTwp0TYji2bgd2v/LU4vPNeT/tKBf5xQ5HlORYvifmrw8xQpek8Lk/7s2FNk25
rlHKNLW+gI2hn27cM0NwhGFHAvykg6H3NqXPJz9Jj5brdCqZ4hU/E/gPs/R1tLnp
DThYHxK7AFk+l2Au7+aBpr/xYZEJDcC1biWg/NaNLzgEHIwZuR0DXebxiTQPxpyg
o9/FrDusblWF48Ub8m291/FENFo+Kuqbc/SaIvg6g+8RqsAcLv5jCtsDtj6q5ETH
Y8x1remNgVC8OnarJo4L2tGK4rqpMJvCb4RBcRT9RcQ9+8R5pfcMgEBh+YubJNtR
ZXeKYX78yTsBRMTKUZoYCkEA+yoQS6gb6h7gzcFDuimjIJs8LraHUUZwjxLxgUKn
LLUoSMfRTHu7cNkvBCH8NYrNIW6NdUetSGR+Vr+aDqjPSvsolDvdlsCDnf30yRy4
sPcaNDx9Xm3gaAt25M+KDjRy5gn7sKpz38UX919Qi65KWcHnHZb65pepGIyoApIT
E/2Yt6YAOv9w/2Rd5NTn387Ph/auJA76wyBaPtVGy3VY6gaREsNMtRxwR3pNbKQ9
BNkMWM7xom2c2WXWXyqjhn1LNIFrwpDaKtZ8pD/ODN/rLgMfyuXaVrkq+nKG+lq9
pa1jR6Ypya4r6j2nJ+KXPVak4NNCGcYzRTXv3YxJE+kb1h89ie+dyQDwynJz8My+
njW0e3xgE1Yq1FTFWCrCwWrpXoyJTRhulKaFNjZsIngwNwRU9RhbH+7SOiH5e5bz
j37dNdDxEDCmzBwvVnEGegZpB0oA70NBtaA1Feu20dTC4/66nOql9ePzv2KDbkhg
4Kc7b6Ff18oXtUpSE9O3Js1lqSpQ2dSQCw4KvGXiuIM8fybLuv4b+74Fug5NJZVX
hBxbypAGpJ8cSvNhVHGEcCAnTW+Mz1aZRyK08jLkFETXiiVz65FWzU/BTsdcOzUp
bG/JCdyHOVA2aD0z68xcughZISJpb/DvwH3SP+joUfsxSA8KYI4+j5ta/xAmn+mC
KmkHGqy6X3kHLpDCOj6wAmsj9aCNrbqzaMwWPmtD/jOjOTNCqidvCBltedQjdBc2
VdtoK0gKzQAVQ6st6BzNHvwAtA1LtPLJuX/IU6m5oVYzXvIQVyD+y9j6CEK8hC77
ssZA+zKMOF2RMxMnkASw/l8GkLyxQBBTSpiWvvRS6z+F2DPW9yCey0FbU8vRcO6+
nQnvrjK8n1EqAU+qKAwkF01xiJ9QjM9vbVwbPojFkW0JNke/IxnAG1B2D54XRr1j
EuHfBs4BRYKoWlo/s6oP/LSlzyxZRnd3kdiSV1qURV4eNP/4+K1xRRAnA25GDYDm
8CkrKXIaw3cjuCC0B+IGX1E7Ngzor/PoxSOXPQ26B8Lm6rRbefrwcZj/wptzPgKv
uyCRuTvHtdDNvj3PJDjaCelibqeodpkydnQ/MlnDr1HhrXzFz0/+sxTgyRO9HS9V
Bj1ZPWiN/zTjmajaSrJ9WJ03ROtaQqD9Lxr19O+GGlCOnoP2uUEJ5/spoq4s83si
F4lqZQ+PHSL85cvd+X54/w+XfqRW88lg6LvIEdnWXHUsn4e4zELkNGNP3dUxW0j9
P2y8+2NpkOyEMiDhmOM/uex2yukm+5KHvTPmTDs31aFQN5w4VhpGLsK4NJH/INo0
5klzINY6wA01RKVpc/mKHC6tbvRn9NxYMQFsRaRqWv1qqTY2n5bKqmPQ8lFvtx8q
hxOdUlVFcqnX9eAVUlPZMGZr7Pvyr0Rl78RRABcocj91lYD4Y74EivT1gUC/AF3f
QtF/Xgvx9Hf20twntA480lycXuyLcY5iJuTXy/GrW2EHFLj9H6b8LgqHwNk2ScRa
xlVcLKEUKyikHamf8Y2t/ys2GCxk3mUpq8tig7o1Xp8RK4IDGhISGq82VDlnHb2R
apa7pKHp39RjBuGbHuDAwAnF8vjQpD5WkaeK6rQUPcBuJ42mJP02rjrYEEp4oZL7
Y1EeCw0Y2ka6W8KvDdmlxBD/G4eHjH4cxgrd8F6Yqr9xo1QhHhLqM4qbZu2npbTN
CwGMQODeBU7vG9ggcs4AAXORKaD/IQv/ZmHaqd/RLEv0gYT6nzzoYO6GahUXm5Fz
cd+oVpnrGBGROcV/fskNyRyDhr1J9gTaSQaB+ZfiOPzEbte49hDGx6DIhF6aE7vH
EjD32eYQpI2Rd8tEp7F+jQzQwJ8kRRWA1+OxehWFxNY+RNbSv1xdSzS1k1o7Z/E7
n/BfmC3r/jU1RnhyDKImhvgFcIQm3Jo9Hs5oduDGE/UWTiBDxVTYqCaQZWACgcKe
I04p4c2wvSTYzQf4STzKPo7wGKd4D3rmCR2YfLxohe3/SaSgE+y52oo9Opb3Rw2h
JSx+TFy+f2Omgo9VoRCv/CAaq7xt7mzy/Icsr2JwthNKjO/I4HE0iRihslKex0vE
J4PzrFbCk3Qk58v6/+2WblG2vMB8R4FOHjiot0qeKwseMS7UvAZvLuWR7DpeVziz
kOIg94ldVZwRH4t07btxzKIYtcDJxVsv0im4JXwObphMEuDeINFanrfYeTkcgQC3
8ZjtW2EcTlCXzBr2HQRXg5az0ObnUTX/ZFclSNaYcRzQvRE/Whu39gaTZPaPCsa7
pHtj7QSjWEKLa5cLA1sfHMjOixvx7C1XGHSj8uab39fDVr7WKtyRgurANw23jYLz
eEPt/QTRBaYovfCNlf6G+YfpX02Ym+kuOcf967Nsb0QHvcPXKdQ283W/30JP8R2W
ktwBWeer0z8tcSIwzUt7CcPL+p80Bp1KDtvWJ5q9aYs1VJr/XTJDBFkZA5RRF3IK
DI7ciX4KpBcRmlHMxSA4x7EuC+7J4rwN15r6RgiHeGmEL8U7CZq/W0uudkHRkJ6U
i5/WuttUrSwR6Gk94VNtRwPq+yB9ZQmEsgzPnN35qK2QjKpS42g/soPjjjJkmSr3
SDYtosXJc7xVZBrEzWj2P6Xl/FzpQfhEg7fKaGDy6nL8IVnXAkn320mvVaDhW9VB
t4q7+sp7o64lo3krDyYqoO7NOOyS7vjZ7IbMUp+JBq8obXRpZrd43TSOQGOyrbIc
Gvmt030EBc6EGDHShKAodnygCJsUQ8DtMNCkZnktSrD1dL2ZAvAk7xmCDKMZhntR
5P7BgAJliHf/yfCZgVIE9kaAoZc0rPqc3zl5EEulfLmy/saY75/e4CaSKkyogSzA
APydbF+YInfdJVFe6ZrJxojShAsJoqRyffSUWZBuAduDNoY53natbF1qnM7IhNSJ
kwG4qYp0hmfRoM93665SjIX3gKHMYDf4Z/WnHJT7w377qB12MtjduCC7s0KrLN9b
VvYwArL6xB/PNqDdrr2Ru7ShdscPqmMg30sUcVHUDq84yDvGgFBI8N3BceJjk9KP
discIzn1HjI8Q1yOL9sZe9gJOndSUunNhM5JBEYVe0GvZHE1VEfBAfwz++OIwF2a
JGi/595kOsgB+Oj+nsTTPAFgC4jlCkThDAuKxaw4DMR/sn8mPwr8x7OPK8K0eWfF
yEQHCFAthCNnxaJtrdtWVaZawJVRp+sbAFluQOBbVDedm6E1jQGg5hLMhKpceRZB
Ge+MtpY9iHCVnkJ2BhNPMWq1SWNVVdPdauJYAMg0IMbktPyv1Wq53sg478t+E35Q
dO8HQ7kSWczuwD+yw5RvBPWdQfm143w8p4HWQ3pB4z2r1ICaIZr9BudMVrCYh5sO
OV9Lr9AQoliHQnDEDggZHHlniLkOZD4uop69lnBHYHmstCt6F9co4z1dSBXpaGWM
bAtcO+hbQkxOmbHZ/DuheYToiDfd1BekyCT6C3Z87Ymml4D+wK+fO9f4G3K9KOGF
kSIHS2JqFkvdgf4oVfBcy01la57LS567RdyW8DL/GWlNdNaFObsp6n3hHV69PU6B
pNJ24KK4gMYFsKSWiB4ruvQ7Trr3qHeJ6PTSsuWrToh9/p7eetxE2JXMTaW4eWVc
LW0UjwcrMSsnydrqYBQ20NQsfIUxw0kRXHEn12mQbuZ8pFT69CiZqvwjVZ9gcdTX
CN5oiupA+1lnqU6C2ZaC+yjOfdDkzxnP/8oxCnfIGL3qtRiX9y8m2cqMiWTXrlAY
byOsykQmDMpv46i24bdIGS1El6yArXy6bSUu8AtSMGidzSovMi4DgxKAIbBShMmq
amgadDPetmCS1jE0KYFvuZkyx+N9HJ5dMBpogJ9K96BeI2OwpIE3pw1ogqSslgTH
n92RS/1wRDdo9Ih8bYOn7GOQQsjmQRYbwdt8YSIGRbvMgllCnVZTi50s+vrh7KFA
KFsOH+zlLKPc2zVyaZ2sCigL6gwrr+kiRnCzfCKGcN+jYHdJtOlfM9/Cx7iCvRz/
4AWfyrnpiqtXrl6w0fb+nQvYQIoQxVx8EQ1pNxRvBtlf6JEezsuhK47Q0KaZ1n++
tktBSQJJjvlZsExAPZoFvKwWDxGNGVPJAqD2E8//i7qpvzOhvcMBv+7Ir4YzdP0f
04yc4LBTf5bZjP5SgaK7u3LWGh5Xu02PXSLOWcDE1SUNT71JheAEn/68GyNqj3eb
02oj1BTMhPFJq13loNHpXiO31t5/83fs8RATDvLzOodsYSVf/grAWlLzM2S/vlVP
qMI4gXimL08VWfVyzJEwEQ93vkZBWFnrFHvNIq6HE9Ij1qwT2x5dxIB37+A5p8nF
9g5MUGHaiUAQEFC+mnYB3xUulZUN05tnjhpTWcw4XPp4t8kRgazm6oXCx/rmyyTi
Dr+0e7HepVKgvafT3K8fAt1sKmVphE5bXilwOETFwJunnxBy+VQqLGoKlHkGniFN
47Ced+XyNfZUXUueVbfngKzmWjXkgRk4dibNCMTsAec4sLiCc75oZj8nSpIxI3Li
U6idXM5fE53a61RmdcrfNE1bJiwNgQZU+6c7AfplmbCfY/RaG03hxZDlSK0f3BbD
aRyVonAmrPcidLH1unBpbg0DbHMKimy3nY/ly95r7NfjQt1QXyfUc8QmSG2UCNAD
/63SFcSqoCn3eoWfNK5i3c6Y364NrMof5TBMShLQmagbCsGLy/6cd2EeTxeFGwFQ
5FPgrqUQz5myTQmem6CV+Liw7stKt+le6306f0QSB7vtD5bk2UFFDRcA3gV4yAHa
SZp8UbZx8tKByDiGlhGHTfZJdkune+0Cesc0P8nB9dSxGBhT1vSvx49r4lHNUe6I
RVLDVPbwf6nElbIcPhUXufqMoPRjl17ve/tLyT6pJv1o6pyHsRs7xFDMAKcFMzUB
17uU0fCkqAv0lqH4NyiY7nuRNSzV/KxnztNi/BNNgHuklkfKWwC/3HyNeexZwX8K
etGdDOijH0cr4oUuKV59nYVyirJxAXXZX0UnDE44Uvitxei9fVnPvpvUaUoAmVxQ
GgrFHx2CHul/d0SZxVc11iPrDZzTYJhS7ChLpoAWMaotxkY164bOWj9mTEx5KHLv
YzSXMoWmHYUWsHyIm/B54BrGG4cnr1EKE/Xymhv+jwotSV9gO+ll+hCV45VYk4Zk
axUk2rD4C8yXYso2dUrb2uG5wcbbtuh2rL2kRpvnyuxdnIpXDg52vAbWRDhv74HG
pERapNmCa7KdbvIGXPbZBCOCJJ38BjAseXjVvbPc3rpSjikb5LDsoLo7BfbyzPke
ABuZVvYfiIYeQHg4Z8R5K5a6iEuMfijnEqYQr8jTdYCxT8amj4VaSKyhFrKwSGE7
roJ/txpHlyYMd525e/l65U94Y+t6GvkuGosZzMHoP9uN8eWmm6ix7Y77L1/xAGw3
vbea0r4RzOxDn1x34LSIWUN54kz/LbcWBJZ+ZoOnXxdRy13Y+QDqpWuQl/zGSv2p
eC1Pvrb/VreMcuD5jTGulHYTDcX/sI5906Vh1bE3Cs1CLPaOXRpCkN/ohylprrt9
Nd3lfOEbou8W+IeVW+0aBsQMPNG8+OLGJSre9Tf79f62n/7crFh9skYFUfAJ1oPQ
DM18laIuIaTiQqteBDwehPaH9GFalU3f7bzepNQ65xN7TEbqDK3Vaxr8aP+zAju9
Z+edlw0WN6FHOmX5VOoqs00GUJUmWkfbuIihLSwG8KpaGP5X8hrJMzoGhg8+16GG
c0f1kr1L0jDQ0w+x415Y+BIqS/81oDnn4ugL79GFES7ms0yYFBhkGL58nlnCcL+5
KEquhJMcpM8XJ/Xb8yJpLiPXWs7A7gcJxY68Tx7ovcK89NV6jH93PDILXjiJjGDT
J573cdvrl/l1Ri8mDyISMrEtgvOkf3BQ8oAtAru0v5z1UQc2V0Mz7m6A9kSoBukh
bY8kAevVOmbI0Zwh07OcSFtqQ2PNe4+efxD0y/wvd4zWNQ54Kkn6WQgYipdO9jG3
GWyEGDf4fRv9SBvKU3QucTZ51ZWHvoHeqTg93mDWrD8IUyaJ5ys65UqKlW7ckzdI
tyXv7wHcTgEDXZPFc2OCZ2+Ca1T7tEsBD5oH691dPW/vLYHRBdXbihhDPjsF1og9
sFbBWmYeZN/+7Jgva1xTwdZ1AAQX0ujN9UdajWJueao3crn45t/CxC5/bz/Gf9/j
uHkQ+QmnNmayVsEx9S9o347N7yGTkU/oufPEB6Te3sNhTUesSYfMdx/X8N5WqGaE
0z5kcTf2SYO5Ik+xxq/Gf6V9O2hLXUAK8P1Ugbmr7n9ewd8UPwjcmrhPsUZiW//3
tI8A1/ZTNM5i7cNQa0xKLi9E49Vl9cSi7M3IcrtK2TckbsjSIDr7i2hkW5XXVXrm
oS4A44M00F9MayFWJj9F1lBTu6mFE0NuvmOTHx8cwjHk7LVYzBoxRPLtPJcINRWu
56JGn/jyjmP5A+z/nAME4ficz3LeTV7hRLAoCiXRb/JlRFJdfJx+GOiQmfvYDnSl
xRQ1JlD+7AQQ2McroyB8kkEE1VVPGyc2ndIkREkAvq1yYE52gsz6g0Saem/MyQUD
fYjn3XxvWrTi1mQeWjlxh/TtBVABMMeqykYsjoYd7Ro4Df8GvHTryEehhiOUroaq
uyBjvXNfAbCl+pttARlPwZgAUFDiyguCag/zcY2ew1IscexCMxaD5d2r2t9qX6mp
HsKQNs+7V1YSPK5ZmZTT+4pf5zll4xhxYR29Ws6yIU4GcNj8Y20q56atAZKCAfu6
kNBQlr3uma5afVGpov9ZhX7Nm95ZZdyo4Mo3uT9OF3ADfuGeXB0XwNL97JokKF8W
6yv4PU0MTGulrSRoDFZ/RIpqoUgwppFcTEV5NOgQcmqNsyBbNSeN0K7fV8VYDcnQ
AfEcVQqJqIQ/hx5DRXZbggPNR+Hh1mZtu76o/5Ooo+Q=
`protect END_PROTECTED