-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
mVcz2nu+PSwdk20+5I3Moq6+0nhZlBQMdBB1MS+2wFyfFm80y5q5aTa0t1uw0NLZ
tfed655ZO5sgbNk9Jh+wubIVQ3X8O9rCh21X9TVZUR7bH/n/MbVwBHelZNSgPlyq
rbJjlL2fJYJTHdrH01R5mse6D/2aYCftfDsWY4c02Zo=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 9420)

`protect DATA_BLOCK
105D6XKHfPdoVdwv/w6Lb95mUbItFzz16aQ9xbpmaWTadvvUUXoQjUeMNB/nha+6
m+aTxUtlDNHVFFP5HFXROtdooDCuC+EvwouCxUtb7g5maZfzzl9aZqc6Y2mtwR6S
3vIYV3cSbKSIbYLZjry9cyw3A8RoGHP7ijT3fG66pUbdnKKQyC3OXr2pjANiZcRH
R2ThG1VdEND56ViTHTBmgO9TSCFtYguuv1ugcRnHLngyhEHta5z97fR/awABHXZw
dEav6I04jUcARB+5YT3sXrt7+9uhZ4SFDP4C23knwIlOO7z4b6v73eF9HCuiJzq8
GJoq1PKXG42ABxHhn1cW3/H13ZMfLkh0XWb19MoG9ba14yV0PbdK2y4QALIuT4Qc
CV3LjuMTauA4goNnFhW0/bWV/hZkla9RnAsQ2bkoQVVu4biL97a1/5PZw36UpYsc
/4pz6QRT/zHu5dXj1hD93LK3dgVTDp2VOuZ3v0yNN70BSuVcclYtgvkg6Z31N0lg
2CCJEU4WwUiyGemdpGLMgCG5FNHh3sDGtVNgZS8/Og9of8jal9a0L75tAIgXg9Lx
ePDXm74rAJHFDDfXMHDJMKlX7h8Xm6G7usVa038AkLHpsGCXz/l27SLl9ws4FiCZ
RSbzcD7ixebXRIL4+EdqEp/7sf0LSq8Ge41o+MTAYtM5L8qdlT/YfbXp4h5pTVrD
MOaF1r3BWnz3X8WpoTVnfasDjLc2TZfMzkWHNHt6ScC1SEFv/L/WkZdJlRqJDDqF
2o5e6EhxP/35L0XZzRdC1cLxA5/9K1HJYwd/dD2298EPrzqG4km5dYrcEpotsVcD
xUJfgIgybuy6SrALVHoqC9rWT14ga2yVx9ODewZdJiLyh9+KA+eWDZQKMY3b0Rc3
V/l8SXLiXXwDSiqOG/n6DpkJ83BolBA4KgzrmL71iQoLdCXJ+9Jcwkm+0MqAGy2W
pnNJ/Ab9f14b9XICTmz/cBubazcKP89Nfl5OxQZxiYDh+AeHSE8swzgOcu9H+tME
JRimE3k1UL2rgeewu894WzlHBUKip+BFU6ARLkZ/EG15a1WaJ0+0XDAXv4cpYP4l
ccS2lG/6lncfigU09Y8s9lD96MJ1K45Ex0mrtEYNOpqQOCKH73XgQzy61Z4gfXI+
5kZzvsSYK1UQZ+0xpHF2/yRT4nGKzDOYiQaHsSUMKvSf78bvN84IJBj7jyYeTew8
zTYYyvnEEIQ9yUB1aCFNezzpUKr91NlvYVbdS0XHTqp4AS4tpaYM0tRBAhlmTgiy
hk7FZe0tGoJ8iFRp8X2hoUv7Zlxt3RO3TbGJAFKzDcn9B/eS35Co/wBFfTrwZiIC
UaOHoywW6kjw8vwMxHVKrLb6h8z7Hbqt8NPeQSRyb4LfHVeSU88n01Ts+UZkQvwJ
HXD0HwLAhsZF6nCWMFtZ6Gkhp4WB15bNV0v9D4PkXjRiw9V0VB8lFWWlDG3R45ik
FBCu89NkboPWlfcguYLQ8c4sgv/LcDGSxT9uENQYxzbJMut0eWVLyOOvSiNMAGRM
svvmCTC7avaCOsx7zxIYvU/ajyRIi0IPNnC50mDv56hoHIENEu6jyvsqhEv/NMgh
ejojteNe65Th85skYvxNjGPg+QhmjRSRgf3VOEGD8bGzDJYId1NTfpEY3fQfn8Rg
nXq09r3ZdR9sf4ccD2c98l3eVNf2oEBD0+aN7lOkMULHyITkNm9U9AcY2cZzRnSm
ZEYahlw5z2WcVxVezd9Zo2HIfDlHosOndFwqXzrR7QjUXwb3++jZJAQLbKlRO4kS
ZMfwrHjftR2cwOkFzWDrPxjrq02gzvmDXn0dOt9N1ZidAsc2mUhPPJX92s3hRm1k
3nBFiY5KBUrb9IZoVibC8nFbwgg4KuBSSN8pscF3WJ86VodvsdYpnr8iViiuUz/8
jfGyCSiHGNBRSNFdRsrpUSEqa1N5QOwfggln0x/xEA2A1yxUlPQ+gjWxSoXx4aWc
Fni5hi698rfJ+J5qtnnPro4QajhA2diE4m2hEysxcrVDBjjodiczrrfUSJLhaT/6
OH4J5TEq2bZFhiZECSnn4Lo65yeia8wyOuU7b2rquBTWhZovnV2X6UI9JPWvz4Im
LjgUY8ZSUlto61oVqjDk0+ke3GZ+F8WfaQ3/euRGVNMKHKleQW2CPQIKWqtmuWmJ
IrDXLj5uqUskoPjT3IuKnjAzvyLT36dP4H/GmArVJEeTnXzW+ZHZCvOPeriPNS3p
vMDmv1whMpVwzhVS+SVU2VtCZj0G5loQ/SB5s9uwJmOt9r5UR/HMT/Fftm9wrUFz
s74mudvzKVQg5EnFEfuskNNoyhSmZ3oPXSLrXCmRJZ0pJe3XGum+n6+xE+rkSY8Z
+rGfc9PNyh+cuxeTjbvmmb3p5zQfcsHaTfO/EfIA5tTDuLbP4/Hb0YKS9D6amEjQ
yPcgibUo4kYU3HSvQtOurUiqZcZiobBjXR8rFijFJyTHfRg16BmViAFwZOjzD8Rv
A0YjO/X5cQW5VpmKWiyCrMHeVuXa/6Ym5rzJjCwZXkfVAS/r4HuGREWmVIAp27ma
L2YEw7yY1UkEAIdm/lB72jO0G4ZakzUG+l+KKR7p97gPBVc0jsVgb8kB8ah7eluN
20xzWpSH8ppf2bzgX2vDC+DuDKcJhgJC6B/Pg5CR166HLh6v9u0ggwpmc+eubm1o
Ex6wK2bQH7ANvPuFRkRr3uyVCEYiKsschtM8ZT/Cvs6SwnwQ7HOYgLNan+zsPr4B
8iTHfbV7WCM34Xq0CbBhzesFiHzAJCKB+BgQS8bhXMza9lRNn052Z5l1uZtUhTZ5
kdTIGrlp0aHTMhJ4GirZigyGejyop9HSj27A3WiQmFNsJcZq9+CM/QM7mQfm/Wc9
YqtdMZurrkQK9KhbYbwxnBkI+Ugz9BAmdYLGVnTThRnz/jUfhMDKaoKaRdgJk5IP
QDrVortgX9Ml6G303HpwiZTWPbL9TR7+wzyVdZvI1cxdNL1q5hCwhzkWuPDAFWp5
dap4sDJ7cluDxzydxYUM+729Sh3llL/oguGyOlySWTcQQqHS2ANpDwTnjPplGY9B
+bg4UNGFoQoHzjJIXQvzmIBrQMBkBF7omcPJvjg2EHvqy9PpZD1BH9LSjQlWa5OI
6+4YS+T1O7jVRADTmaNJhEGz9cqW5+Cqxuy1fhCcESqTYm70FG5KgwsNfqJ6OB/V
PQV61VGjhwn07KNltoUr7Go8XNvXohw3Nm+zbVmtziWH3JtkciHIH4NyFf11X91l
OowjWKSAR+MhPFOrelwWF2SDAl8XTpg/oCglZQ0UBQtq+nRG3XUK2P/SIRqjUk/9
EJwv4mnoXHGn57/sWn0i/OuQZ+JQM8O/AuiIGdo8SDSbH/oTnL4jJcW8ifRWB7wV
yAlT0wsh+RkqsDq29nhSFAP0K7jX9KqXgo6HxsvyalNvSDXVtWoja1w3Rm95QopL
rrzlPu+Sri3pI9ksQCGNsqJBk7ONupK+jHq0FWV02VEjYIMonedlsrGD9axPwbLf
M8mPd78IoMmz5tCNItDUOHDrNbIlgznPxVp7VepXxByhIRwtTpIC4aaO0y4kx7JX
SrBJql6eFk9y6iBpkyNodV9jAwXHiO3THregfA6IMxTglIOWnLfzmEsBdAYvxPBt
DV4mGWefqt0LmDNnpFA//ytALJGCHZkkV0tLKMauGw5jnUpif16h7MbwruTbQkAh
hNw+dYy0g4JGZttHgwfRnmBW3p+bcm9iNflsm6K4VKwtJuWwk8Pt5O3+GIdk6LQ4
DSdwshAk5/Z+YMGu1ib8YF/9OlvInpJ+SEcpcMl1Xe+hvEJylKHc+BUSulxvkPIf
+i4zTREgxypsZcFSyqOYmOsKTmpBT/eq+rn2rRv643KmRL3h3S8u0NilvajqOmG7
WkqOB94bGjfbErrNbiPyzXujMxt8R04olHEdPu11ddvqIl10pLMX7e2JU6Zz1eLJ
VY14Y879TGoeqDHrYrSBMvWtd4x7Ov6zbQCChjFemARd3Rdz0QO9gST4hh7Zvpdr
8tL4xrG/QiF0hnGiPyOvbO9H2cwr/1V6lB42Mk2+hNvw1+Fdxzk/gktpLBAseH+f
Ug5e6ZZW5B+VfzTWVPnMNli+FRPWcDLXvviCAz+74MHgptnOn0cPI6zHRhgemmUL
69OjmgT/B/TsnlNqMg/uN2nuVC0CJ30mG/BbpeDI/gLUfbnb4/zOyFcyioHI3xM6
oDwFeBwckyY+skxPGhmYBaRLGOP5VzzQ4JTlkdKNFIoO+9VRC/tP0qr93UcIAJ0c
kmIiBn3c857FNYD30HnGkLpjX13jONqoCZU5mO5jt3rrngk80ScR0oLKwMfgLrbg
edt2erTYrvFeBf5jfg65A8txkRWXzHY0qW3m5aHgQ0v0fsv+Im0MhP4CVeAroS87
btFUdHNCZ/wDtAn/3BvuXnywkYb2rSF1LnwBC5l+4tQLgHhmNOZD8sgzI0vJ7A5z
ipZ8IYJYrj+kBlNTEQOMxne5pWY9UspfBanKVBnJAdAbNj37AAhCDYzIQQO9EeWM
eZpm63pM0DkL5czL2TGGAuCMLGkJuwt1JFCx+MevTSXZfO6VXR7uqhM7I8wm/qm1
pzNYmY0gZoirVmsJE+v8ihK65ZDb7w7Ei4d84/lPd3rloHGe9lGqr8bbBDTTYYfe
5aC2slcW00evh31X2tD5JIg583/0Jp3hadK2Xdo5Tpo9Y1WLo0PdSnU9vuhhoTVg
VElIipq2KKGpUDMcrbg27qawy2Zz1dDYJBzZGTag4+2LQKjEfE/uC4dYyBW4Vg5s
hXHCQ1Ve0UOMC/rcNBiXQr3Ne+xdQfWrnaXDsnMxd+Cqm17g5sRUZXKX/PAhDHsN
I3FvhNWa48RBjmiSIimA/u8MEQ2N/1hRv12HqZsUY2irUZz39Lifs8tmaVlZvh8y
iZWKj1yDSzHPOI4/cyHNjSlEXvN2vcWv82SIL/YUZByxyPR2j5AnO4uGnqKwyMx4
mvCY+/4H7dUiq0uJVhfrKMekGOi9bQUV7CgRo3Wy+jb9mABSth0UTKkQYAoS8Uvn
+lHxvmbIFxlILObyZBEC+x60Ep2dQqRv556rdVOLHZPlJKaDoQb6BQBLGBQfqG6x
LJWiDsJXWK6VXvkDlODdFZIR7tED7/0EX+tOwOuOUeb0/MGcGARWl/MqyPTpP0Qi
GAx0gaJ7RJ29VTsHkM7KGUMDFMjY/JGKlAoXSf4zE0IFLhtJMH1k2+2YcZtWAmxN
s0xsJGAzwfITs8FfYMlv23gVLaOFzMqYai/sPCtr5gp3RtOluhuLuEsHs05f54tr
kVvaFCtX+73ORZchApV5YALaIhyB9f5BRtDGSnJFJg/AioKKTYFmMyzjKMCNUoBW
JSXH/4Oj078aFy/xbYi5w48caIaJgicgaST4Ck6X86gtp+A/MZ8iSEFrOrqfSnuo
aiGX0jR6t7GeSdzMBXQ4i6n5btpjKRpwZqQZd9Lu7v2c4zZMMt1eB9mBTbW2JE6v
2rDP/DiYEcTkJWXPjsg0YdxbEZGtfD6EsARnPlJl/VGXKmL5niIIiqCz/NkM66uV
bTYSUPvE8KKdbzOeAU0t1dtdxUfODYYTsGMALxFiAcY5KXSxB6Vq0U13BhfPC3cd
Am9jRC0D6G81c6IJLiMehsm6uN/S1LIz4jGMM0ipzYE8OWAKkF8hvTT9tMHgppa+
kNQdAduxxI1hkGJ+WE1MAg/GFpRBUU8r1w7+kq3UrDdPXEEoAcNYU5ZQZvPhuWwL
jWfeSRXqOKSi2rvHMSoFIBSX3Oo8P0MbiosRcD4IC+eJ/6ZxM3bszup0Swo+nIc7
eFacg+jGiSyWgcFc/C3MuAb8Xj+4ZgoBhr9TXjqUc0F/lLeu4z7SHVp8uXtnu6G2
yULrcWZAOsMcLg4sWIMYDkq2owFA7TCTxdMRYPUkYiqOqaEkHDMSKZ8KU1fPH9MZ
sqaYVsSqq0H++5mYS33EGFfS+QcOw53vuyu8YegZzYXqEDEzYTdEya4CWX0Od3VJ
/hR9I9lOwUWMi8rvbmQ3IC0/aDEXLCWkj/QPOl/M9/wkjU08MBAUwk0dEvIV9G+q
xkXsQGCsrGLQ6jPHasoTWoomeDNF++XeB2rBdMkDtZo0h/ibg086slsMmBDkB9Ro
dUq1veAZU33RBT/ZplJxJEMbj7CEkdyyS+6LfjE1KyIB64darRKNWIiwT1C/bKoR
LCoq5o+MlATBfcCa2I0bczKig87e8XoYIxPquC+nYgJ+/LP3ck0NoC1vRiN2Rqro
ZlN4iNPicZg1qwkjMq84K4NrWLklwTbarvL/9hI3EFgmiD2uUOl5LHwRKjDgeedW
GqvWJlgc/fKqX8uuN8I48xK2d0YSYtIRQS4MbqgorUPVz3TsuBSOWhYW2u7ZdemP
t/rf8AR5XDh5VqggxIzJjoyAmcb0gNdIjFnmp4CMT9aGq5uey6sJsN+kPp9tjHnI
0HwCDrz1OJTKr4XH1Hc4HxEn3pCBZiSCz9/lFqZIfG+99imrrN2mJV8CoAwjYQbD
ZEo4nehrcjeMqQNju/+hZLlkJ2zvZSKruqdQcUUMIpaBwHQhB5ixVKXblXk9NJu6
sWGhHNq8XaHXamwh2fRCh6BfAhKSiyFOZgUa3zj8oLciIbPaXQZ76l3Dr9ISUyCR
ZNKzfS7zJVUxK6B3CPgqWdJ9xYQyjrVOfgpF4WcsfuX005js7htoIkDNfXAU6orK
bnhG5k9lXeRiWMvkIoLJhmuw07A/UklXZJT2NzaDWqDeqa/ayPjPEwri1wWhsTKn
f8Dz9fxjuO1rEvtN1pMJqn/NtFT/Vnn15V/Mbygb+Tb1ubZqLBNdLlSZiFhYOn4b
m7ZmMMQXa4CqD9LFykh8xbRDK0VgGWXMH8yg2QKuFQ26DpwbXgdES9+RcrWmMxBM
9HHsVRUY2PcF6qKoXBxeVaFSXsB11iOCxvuYZbds1hHp37WjEJm00nu5cLpW7Sjh
N+lBeOeyqznrP1LpAdno2xDS96gf0/SdlcBpH7dBeC1chpTo+JEC+/mqKqBgreyr
VNx76Zzk/N/K4ICxv4E2XsQpEedSPJIyFG6crYnbHqbs8hQEq7MRKCNF9pYn2JKS
L6uEEt0B9VltHB9N6UFA7wJK0Ccre6MCfEEJIH0rAPhZb1nuDwI1tiMw1i0FVjOy
wyScxxeuUd2pPWMuontVFsNSJJso7Uc/9IBJnbHZykJ+CucQhb2w0dn9hBV+DGq2
9Xbt50hVeXnDZgo5E7ZSuSpIYzdIks+JhWGSkcQhl7Dewn9PJLTINcT7GylwWtfJ
i2Iu1mS8Y0i1RaeNVzLmisYMiQjdwuWG39iG24m0AieZD4qFaPz2QAip9/qGL/y9
M4yMpDX3kcsTTZ9rwUMfwSv3V1qCCte0mcuRPQLBbTgreVjbebQ0MaUc6R0uBsHl
NW4wMGOk3VLNbVQfY67Tn7+1JEPNJuK6Uyuh6ugfPInhs8NtAPi4bAX1wfyeI+sn
uIZHc1S5eRHr0EMANB8AfbwveqcAd4kPaSV5Dx3KGZF5lf7nKu3XWb9xUXyj+4+2
UK+YuYB0Tiy/IcfIE2E9niU5lL9ENIURo0GIuYgeAP6DNzztfBqulzh4wOIf1zGo
l6OJttVYhxiyNYMHJq3AED8zhgoVo30ZWqZq4zwkqzH86+H9T2wPb/SvcpOrqIhJ
UloBHLwawFvsuoGNlbQfVYjLU1fTqU83/1Jef+7T5aiAWOtji/Y0ubsTqanMCub+
hhBW63iw35mJ1kXiMaluUWWoxMHRKYVPMsqmqb4LAryi6wSrXf6UvVsSt0Jfjw7Z
8LgAd17TDqLU1OM57Rfcic1kUt1Zh++AuC8It6xFI3ZcxWZeMP62Znh/CxcBjEQa
+Dix5q2SHSoYUWTyl2V7KtxbKt3wZM3OsMjJyBDjsS7bKE2ltNo0zZfoGuNb7UBr
acST4MeKV+ME0c65h4kkxrMPeUrY5D34wLPl1EyWQiDZ0dU9gvUjjhI0TM+7yXy6
UofL+CbPM8AY+gLL6lXzJmzBaU4zeKwyaXE73EnzxOzrRKQfUwWiVlmRDBUhVWFm
sRm/P93YQeES0rB98R8kb1SL8UwUsKi4LA+zjZy5MMSYnsEuwjmqF9FlMYsmMmW9
VXqZvktyAPuTx8SJ8U1z7nifCUxxdholeUE4GDLHho42DyxwCfcZPcz8chwdkWvC
iHHNkIrfmjhNxVZQzYMfkuSZN/KWsIeiAAhd+8wxn4jC2N9JAKtscK5a2G2jUBJE
m9KK04+zKHnCKGPHA+yjz3fuapcM95Aw8sH6JCQ8I7TVG8u788f5HB9eGl92Ek0c
2lt5D80HRzXmTw//TSMYcwG6JkgyAcBQHohWc81Jo7/y6LCeu1Av+5udrVKYg4xh
vYn7kT+PHu3pz0kERWfVeMsldJBgejhDowRm8vW8lXdn31Lt04wz9UqNaYbWmY/A
RA1ZUY3NBXF5s76IcUrbyzYn6OksS4rVsOjp/OB8XIAcSxUfxAPF6s3FNm8jl3Iq
YTFNDFjC+LQTeF+UNkkDeR/UJCwqvCUjUyNYkDEf8tCQWZWOwLhr4lZ5cjSWpoG8
2KbNdbpf/7OkS7Gk5+3AYNSvyziWesqjvndZ+S0dhCqfP92CV79QqG8TYbio1F6H
TCjLFKp2lSIdX9YuMb8HEbhGIg53lEAC0eZ+n7/zX5XhggH2CR0zRxYvhBFGh2MM
tN1Yj/22ZOHNmGgtmhQEvx68Pv2cpjpu6xAAW2yQzlXtR/riRAuxP7wlxwQxswMd
y7K5w32LbgevNkMVjmpLoBSu365EV4sf5uNj0+yK3mEjztMXR0zjzS2jJcXiWbYX
HpfsdWaoCSUnLgfRV9JS/17KJoZVFb4GA3lGgp69jrxLZZK/BV8sIkPyt7Qz3uVv
Ap9uNSEvXFqjM3rZNhWnSqfaYFATsy+yqlk3rK5xMtAfLwlRiK+B9C38j9LZYNBw
AlOnSpcvZNbobBM9T8YuXnD1/ROE5g1WgubCqMnfhXqtrwtP8cBXM+U/qC88wj+Y
Pv962QWwatbbFZgDxTtLbvvCjkusJL9FyLvmw63zNFaI83a3o2iK9rAUAfm5dLTk
RVSfDSNSZppTUpxAxknSrxSwxqNOt/lZsdAjYWfeGY5yICqx85pFwipbrtu2JY6s
TsPP69WsVBOb6o1lyYk8f0oaHvSThU1NrJCI3A6TVNRvBrX4T0ULEq7wTXZiJYzi
R+ocsN13sixBaZpK76t+zv7BEZhzU8S75xx9TBOdhYwXH2eTKXQo2WNMYAIS19TG
AeCdQLdSDCKLY6XtE686fNhXfzYHBEbOcx6PwlOxh7yRlII9MtuidNy2oIZRfj2M
Nbd2Iwtk4bpGTNLsjPx3oxvt0FLbBTNLcYxu1uJha5vjhScGpJnzYDKkVIC5gq97
N3CfOtPTNbHahtXhItCSD5p7t83qmJfp1tZn+YnjlHviP0BS6jVq8H6anRwWLE+D
/dO6XDZpi8ypjZVuM1oyd+M8q/ar4XZn0NtZnHrCnPhlIxelMHoIp+TiWFxmVzQU
POOTlyBSqV3CNxsYSqOLqwflxYMVDyxBXSX6i8GezxOPAaU6s2J7hUwE3c8VHx7z
5ezPdrrR6OrTCwkNwWcB0ABZ5zNGReohwFSEh8yKGUdrBQjYKzAdmJgxKAJisDBS
H/kzKRQLRjS6x5TKCBvc9AFpLNJInw6RS/BKRYaSZYurEZweRc9DHehsJOzAPacC
tWHfa4aPq0WraX6iSQWvHT5atraIcThDGEt12Bx45WsQtyImJNMMmCeNohUEvUZg
+gS6EdF7ePCBD9OgLvsV3iTK3OBlxL2LjixKgLVJY/+ZzIVnzNvCarffh4+xRXf0
4imBxW5WmT4GP+HaZfU9BoqYbv0YI32HKaLUi64I0v9LXFBGhfRIVjG4T3OoPE8Q
ox1od9av2zKJQbqKeN8jC07BoaDzxVW82XPqdjqnqVHiyKT9/uBuRtyzGqLf1Hul
/VXBA2xtbDLmZozKgq3E9/7YKoSWJmYQ+61sR2wRbIcJSu449z+tRFCNl+ADAw44
B/4RWjM2KtYIFdvz7F2f3wzfSEyvxbivO9J4IjZn+LRMZol+boBTNYXqPL8mQcrZ
6AIN2T48S/kr1/KGbUeBx9OIS58geWPouIcq+NJMdlgnwj7MZz8++JdfyCjUjWFl
Ebj2kt6z2MhDXYpWdxfcI8giL+dutD2econoviinbJVVP8q+fmhYYwhHuf9leHQF
v/KGGPiqjFxY0TboS+SWNfbKhkN/3gRIrqoS9GZIRfvrIe4qC+RQ0Mq9mGuCqpu3
4OtHwB4MFIz2sMtPSUxSZXbCjSZ0gTXtpAEp9eiz3bxN5SAJ8bCv+9ytpRJtdKrP
ITYZzMel6LrlTlEYfXEipfE10Tnqws9KPOBACV0bBY4X5LefdyqTUaL0B7DdLZt0
BDoqAUPszen/hYBlgflU5OzOCF4xREGxiHlNiZvAa3UvEML+6GTNRD/JurbEg6Mv
qw9syPgk15EGTVZRyo1mcU0EC6wImKxk0FYykNCGx4ux3Tq+aDW1IIRQTSPrJlWW
iDf1y7N2JmdWs1niSQpGGx9SgsgHTitw2ATnAmvd4Biu37tIoKl2NA/8ghMZ8MNG
1p5gd0Zon1b0RuafxZZ/j1uZ715VyV4Y6qw/t4+JRcqBunSQB4bLhS+l53lXnzdQ
T/t+9VWQWtAE/Fw1sYQvCf0dyXU0hTNIwdGuCfFr3sUg3E9CaYDUGDNSqWpMqgi7
twP+LkwjFUhoxh2U16txlQY4VkEhNsb1vvUbn/0Xjy9+G7FZt6Y+VsmN4ds5UnrM
vUTJskADQ8OZIKnplU7cyOzBw0BLmQloIIWU/QlS1b1N3t/5KjBPk5Umui2Phc15
T5muOdNKkEY0kL/4ihaVDsq+YK5bchrKSzdOmJ7CuVSJCPcy4eon335HGiaqdajC
DKjf7Aw762qNXqAX1Ul2GofayOi/Go1E1XF555C+HxruG1hNl90O9pA8QFKi6cR0
aWv+dqMt6r8o45sacz5IcUPmbrBvCswHt95zqKfdbhRZp4RyqAPIifULarLJjck0
UFlFQxkbOrist1bsYpG//F9ozEKfA/KtYeNU/WWB/7hvNZsmNV5p613aMjufh8zl
K+le7LvbojyTQBrjfkQbbDtH0CBAvEs65QsO/hETwf1j4p3rIlep876vg1Ph7uBO
vi6J0EwNp32LKV3Qt2jgmtRzjTkJGSBsZHazOchBNDeWVo/eCIJiesYrCQjJyAdT
RSeYiOIg+yZj0UX5bD+0YOic7srONpSutbdzbLOH9GUsHxODGZ10S6m1odJsnTZS
fo0wcjR3LfivDP2NkWXjhEzlyr973v3azlTrOAWyTd+RwccZ5edeeVtg3jR14w9G
wylGOsYUeByh+DEpsU/Dv41h66BB9ztk7oQRfMX0dXXGIj1NiWrdy+x+2402ic+S
VZzEGFaHvoKDN4A/c/63Ha9hOWjZG+1mqfyejxcIuKO5blC/USU/03sY4D27RPRn
9s4+jNmWQvWtfQdilEM6gXevhGTtpb6ecyTn+PulFbhnFcQJ9thKIAsRVEDWJNvR
N9tg+yaYFmgOSK1TE3H0tMct5ngfW8+Lo3m6MWTpp53Fo0t/fLPa7GUHQs+thqz/
bdQW6Z+xmfztv5KmkLJsKDGyd3pXB99skw5nZhWTfnG6XognwD0NrTXJXEIUHO6d
BhTRwGkVua+nIJHgpnnQwvHdS0KQK/MQ1M3s9azpTteFraZ0PULBPsnh9WDqJsdm
LygsmYJIzZ/hbwIXtWnHZqIcrjkXwwqwkoYI7xj3gwOYugB5Dco4+eh/V9f4s6jU
xL653RE/iARrn+OhjUONFWlF4EvQXL8Ddb1LZCwTKd5lNF9h9xGtCA3NvJ11AtNJ
i9EKuDitTHqN8CuMNpQ0f8cSxY6D5BjKkK7tteUG0jKzw7yiqm4ODSLqs1DNblEe
OZ5HhjRiVs3ASiIB/GGyVCo+g+FsmG0iewftWtkSGLDKPlIhv1WIZvNVer2D62T1
DoZiCtKF/wkGkPHFu+WFMPgveBHMJ2RvJ9ExDCXbMbt/k/byWDxDIazGBuNuJzcp
ww2On8E/jx6gkKjBhnXF4o4qLZCgABYYUPTPIilirxpqvrUqU5dIseRReeSFdxHe
bsGLH3dP1dgVhaK8s4kXCusRKbI3VYxYzw2MM4Elrveinfk+3nK0TpKmI4sl8tJH
IIvoccIAoNvYyUBDzQ3Kuecet3bYHlPhUHKhdzIVuWpYZfxphtLcpfIbn+fa2X44
bQJ/JqxkS55NrJVeqTIcC0kOTBtfVOQ0Ad/AvoUE4hlnxMWdmTt2MuSjb6DVGLN0
+7d33QnQ3SPF3rdM7+7QWLQzlGOfzx7MYkuocK91pDkrYGunMqMzSfkQI/A1Z9YV
ana3Qd1tos1ZHvWwDB4M7/f5ZnV7ILmJiS/9M4R8O+75XkXvXi4JdHeA4HIg/M6d
DNekr7NMcmAktcq7vWhLv3kG0GUXlselk2XcTQ75i96iKnpAc2dncUduzJ/J4Z8q
5sVLs3I4I9StmvUIyb6d3TGya1QWPxgxvs68Ya079Sc=
`protect END_PROTECTED