-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
--pragma protect begin_protected
--pragma protect encrypt_agent="NCPROTECT"
--pragma protect encrypt_agent_info="Encrypted using API"
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
--pragma protect key_method=RSA
--pragma protect key_block
hMEJBsh5WKB9Aczt3men9KgAjqp9BUsmM5PKuT85O6uY2q+iLqgfmG7XwwnIL+jt
ve0C1NphAVxQyuUTxZbICulezLVCAv6/vcpc3dZDZ/vphCu6oxq1PZn2DMHOtH27
zcBh7EOF7obKfkYhJ+hZoVEvAplbjdpIMarh2Srcc2+8G4LIy3DS6k49z0Blw706
ykEob96lofYMNxbFAbrfn+ipZS7rUntxJ98WuQW/Kw3B2XViKTvVAuakr1Xvw40s
JYilmtsZ4SDHn/3axAJC3FsDkSy7WQTO9P1Eec3GzAb+3kEZIQ7orB99OXbuCkZ/
lHOFxAWMhso2a5Po0o/mTQ==
--pragma protect end_key_block
--pragma protect digest_block
5Rx0c+7SABkE42ROQuQygQuek3Y=
--pragma protect end_digest_block
--pragma protect data_block
vpNorD12Zv8w+XQ18LbCFzSZ03eBPumSjEV6C1JWUMJ90bMWPxpFSixiRz80det5
kZAMfCI5A289CWjcIfMS/4/KZ+9v+kuuRUjdGHkj3ZFEEpZNgUsddFnQNufdKXpk
/l24A3sfH4bCnRN9fjqxO6iS0JAPkJnFChBN/otnZk+9tPQs4Coea4StmRD4ynQp
YPc0YYOmINyRibturymikzRHhXu0MuFBeV6eD+pMDSInNJHgCyifcqTpyIp2P2fW
LCYy+HfXz2CGwD0Lm3Gbux4YlIctOPoBXNC5PGFRrR0Du9mS6iTvnBbAyOW9z+oW
vjtgFnzGvXvzIaHecH+NGchNisX6z+4IT6N+sc+VT0zERsuMLBcHZkB+Qr5aqrxd
gB1+rG86NN35zBnmmpS/7fKpWEYX5m3TBlflENmcOSZ0fJtRJAj543D4Lak63Idu
IU1BZ6n7ATKdln8ZHToX70+xIBRrqWTzXlBgmg29siBzyuU8asRH5L5zjlxnPosq
ahCYoc11VLK1S5/dgWCFxJpSQzU0pEfaR0raMfwgpSx8j/gQvXJ15sUhPhU0LyYe
ctX7TFuUZlFbLj26RMnUDDgkgIAVAeuc+8+NigxW10EZquo2Jfh+wQsEfUZTeO5P
lZcYcxa7p89SO2FQR5/hD3xdK27jaihfcuyCAb9rdhHf7Andq4NHFsiWc3DX2em8
JTcSq5OI8rOx2kExL52LSbcxskNMw559eUptxPSc2BEexCYcLgNULAVgaS9PJYyx
Z2EYihbqC+vs6RdRaXGzbADYGx5kM6YeviBKPRARJd6SVV5G1E97TX3SiO9sVlYm
XdRSi/s2v3l4t7gCjERIHqBgT+tsrH+uXERYK8GBPZznY7ydNgf0gdmxmk0zuw9f
dQVBzXpQN/aT5W3digO75R0viqq9+JvFwT9u3JD3yg75epj5/Itc2xZpq5kS0BmQ
wEksHo+LT3V3FYEeULAjtEifiS/BRbJOQw2+aU+MZXFQT+oObVIc8XHRPyaTOI4W
bnD04BkkMhySOz/w9FPmZduOtnuRVTjLn6AzQYsqkXTYqBi3Q0uc+ziNtsVrmAqO
2lhmUjFOu0aPODAET346S1h5uzB4JJgGlxECaXDe+7Lo8BslmqT4aD6reLbNROWL
QgSvEGkwJ3sSVqz3vTdAlFXjsS7Ov0qZ9qgz+hS7qVZs9iNgexROH1QMQFlJfbLj
aDbus1ciYi207Vp5TisfuK5igfB8L4gPFJSDFbmJqfN/gnJ4yO9PySHJ6P2CF8Ps
qZRc8SBvA87i0toTSgLs9Z1K4m212L8vy+accYbByuAOGmH7fW75ZOUYGujbKWD4
ddonu6qI5h+vzDXW6VeWMdci32Obxgzu3sRsovrcg6klthGCThEvQkksV5l8MTda
wjXtzlenYdWI49SJ8JyQoqIauTHmeuSE+kSCHok2UIykzQCwcfC1DlCMAU4mn+Ym
AG8zOMUw62OgP6EvRMwvM9MvMmKYQd17DNa162whS9w/8UP4QqWbNoHWTd3HMQw7
YEOYyHHZh2cmz44FoC2sVgbjX9U4/NXb/fNwbgXRml4whQWovIHlxwnVI/xXRP+T
R9s0GBsyzMas9zuc/RYAOjl9YGqz7LGJWniE0vhquhKGJG7GGfM52YA4asvixbB6
CVruIO/LYvrtu9I3K83IXv3ND22H+H3vVU/h5LWvCXQQGzzIHQ99XFbpJ+sACe6Q
9dk1WSwA/AMqtStk2iw5IhHjBPKnu1Z10ii8xeEpvO7WJQTjISfURtpSiJFNi3fB
z/q9lJtuFb75dlf3X3nZrihwow8Av8NP0oCFuJ73KLZmRb9SgGGgzbuDHqggJc/x
1VzZ+Id74zvcgedjqeQhHUh+I7srErneEm0b33q0YMzEQlB+BpMxrDSdSdrWt/nl
eUPVSb+aHVSQoWoDdU5uWCg42XUYHfcM7ipy1zvtnCp5k3hNA/By49W61q+0LIH8
UaeYn4f1glQN+wWbKaJuKocErA6f//JwEMmi7StmZKfWeo1NAGvJJh7aoJ5ak//o
VHlOky0aI9kj3o5YYkEqGkd6xbfBZlevGA+MSGnCjW/86lLZArsHECLCctq/lq8Z
RtGhb7rCNutzrFeI8NZlWkwARCbKKWZD45HMcj6F4kPlMSVUi3tJ33cpTN6cnTN2
BlBNsZ3Pw8nMH7dfuBWjcmqJ+vUHfRuv/vITB9imNu9ohI6svvW10uaKZGZJ8C0x
c1qgY3MoUFdDsu9V6Ipv19FXke/f9gABh7LA0vKggONNMHFNQBIKhc1UR4lqUXet
+kZN3LP67dh/XijthSVjEWt3Wt5eseIvZc+AChSbuj9TX8f3z3o4XL8DqT3904EH
8a9HNtitdFbBufg4LjJYHjPHkAL5h4lsiUmE51+EARjODzvNn14DZjhp0HtQuG/m
2gstgUjqdYXjqNaxNYtwixJPCr3J6EGhxRHbePh7HZEsK0PsPBOgxGKMLXOgpxYJ
UloYJJ3UZzMHhJ2L8L/BDY19+clxpM8VN6T+ndyYV6W9CMYu/s7gWfpN34s71Z3P
DJAnJQrXvuq0AEpKTLSf2EdyNkvi1zbu0Xz5m4GpPGHHDcivggfDZJDLaXemqnSz
n0f720UdP0Dwcc5a4qlGf5d7dwNNstIjBiu54VXJH1f0NN/iN0sdW/0XIocH1n17
3JNb4I0TngCvte61fLftQRGnPlk9MJaQIE4Wu50iq8052oQjdyVdsqpf3Pl1hsqs
XBzOzh9UbDi+IFt3/aZCe4hkogWxBrEbnFMwRYC//C3mDmEFR+CQChMrkiOFH1Gm
wijpmhOoiaA4FfsAHs7ezE/LiQs+TxmRpny4bPaSvB4HVlDRAs2bZJLTiC9et0D/
8jK+9m/Vn5k/IEdwU4ED8idiPV5bzMS/Oovjx/IB+YRhY4bmiBcl7Et/qHHwXNFk
L47gASu1eMVW1Jf+ia9PgUpwYwAWkV+NaLRhD7m9qoromVs3xEWzmEKcCkzkMNmE
MMQQ6hb+IUZ7GR41SB403jgaygLTkdliBb9ChS1PJMW/AsDcL406ldP4OnoNBRdZ
lHQrfOEiKOSoOxakzwlmnLlYhhP/EGiAaKS3u3U28kOC1m2M6drxxbi2pqtqyEeh
ZHRp8FdfAhFt0qqznq86wKClAb97HiBPVFD4F/vOwXl7Jk6IcB2VE1QaWvhQQW0i
cuKZp/KGf3jxJeXBMN6k1C9Bz1mUvG7Y7rYdGcfrsHJnoWLZULRe9zJL7gHpk6YQ
g2xVNqbH+Wxq1ajZsT653JGGaaXRHubjJojGXOY3mScNXJBo3u7LAwVcBsMBM60V
buH+6vNp8xb1xf8RA0q/UJZbc+e51qXrIG0tnkQHEcskLW47EVaDjGF3NfraDxlO
dKTPFF0ad4XVu+KA1FAmyuVh5bmUh88L/MXHcFRyPrJ+Ypz6kyND6d1JWoL2SNDx
pMug37kszjdLp/SZ5KsciBqgZKBNrPLumSTa0r6NCFlemTJCWz5hNxdyamfNyL7O
1i/rc+fQZOxg3bJYkF4HvadgHwuNBCZMVAZCQsvt8SRoVFH2OQguZLpMpCkFupFx
Cwv0D5E101nhOIbPdafvFADpCR+GDzK3q/JE483yIN31rdfPuBkbiP/VRRJPTZq4
3fJinzuNtX2SlaaoAdebknstla2u8JlNRXuhSnAyJcnlk27VyqUr5aILAwpZ+aSx
uRZ5c77vnUBI7y59FT0mHj7AvKwR+WhXwu5i0sfzWfUPQ03m2oiFIqbhwgGKFUl7
ryt7tBQGYDs3yTCQXGH1NNKEC/pJFMvJBTrj38tkIQphk2b7vlIP7D3Z7ITxNumv
ykjURfGRY7D21Od/juz/+ewjbZ+B+FVJG0QTQlZzWB8VS7BQ+YiNmIW3jssxNgZk
GRdYRGnLc0gQPBDSksyf/1ggwfLSEbIBSVqIMcoAhmuQ1e/5O+GbMzfzwPboGibF
fNaL3RBs2jAy24bea5A3qdU7N6hBNZ/+g/wgSpMz0Zr2grZtEJIor4ykpi2fVaKE
psbfkeHykxJzrTz81K7+PQ8wJv83CZ0xA9dehk983ahFJ4FK0HjWY2lk2Fj5LR/N
klEtX8cH3YGd1quIUyFcgSG99vGzbMQVAiT3wIT+oTuzQDAgnAdg1V+0rphBEHcY
L1Mw3A9FwiaNykfHZQ7GNJxLl8ezYoCYOuXWUiThVt3qwcTgkkTevlG3kqQKTJ0j
0bghjN4B3DKOug9hCHY8Chmwhs9vyu33EKnWmL1dDybq448ZyzVPvfpn+WqSF21Z
UYZIS4uLdiO3YTa54JLMX4O4d7/pSBFFXPBSolWXb2kId/8oEoJ6s3/pxX81ivH2
O0+6rJbXiBxpRhKbPO7HBwoU6rsGwhvgQy71NXlyAZijEn3ZAaVgB9yD2m0GMv12
/Zuc2p9vtubqIUY+0cSlIlRAzR0W40MmTzPOw+sYAF7rHq/lBxnMEh3JrB4pYs9y
u9Y5kZRwbWDb4/TdQnKdcake3N0hro6T4IC3HAlBq9JjoCOKThgKL76IqYuA4Vtg
7ieojYK7g6Ap2BN9zfCcYXc164wrpeaR3m+HTp7xJuLmLTe7kJXUx5h4npc6itBj
tye1sDehgHT9m7950WM9IiLWkWkZ3P3h2+ZekqrfDEEtUHbEKotfGDNnMytEMhH8
4uyzgvJ1UuDuYEUA1wLcgJZCW5W+57FgYhTVAQolTWrJfqHhLYZZlzecvAiM/fZT
WUkNXfW1ghatGOdqxXuRNc2wCnxWcSmL+geAHm1T9YjeNCTXrgOWXwbf6T9UprfZ
G8+iXEeNLhlqya6s+hhmflYWNFwTZAk+MGKz7eiPxbntHvQ3VExztuy3nQmIcqY7
pxn7Fdan1N5iHRh/VWqugEffoD19XV0C6IM/tJWwpyQu/4i/Be1zJ60Yyo6tOrmc
nWn+eKNn6ZKJC58e373HW58ZKeWAP2XV+lDNlhZKgeCqZ77yTL6CWiNtRoAcx6um
YeY98yrExu2TDiH01GH4RE6xkOzlEtxK09BifD6lrEZLLJtvbaZ5QeDKMfRcbvpJ
Nc0OIeaa59I4MzNlCpLgUTq5FY1Ay9t46vQqw7Rkz9Feas2K4vVtDC+TtavINBat
4eI0JQ42u1KqwD/WxFog5t+3cSB8vHZWttZrQP0rL87UJeFPYHPFnqpX5Z6Inc4r
KQkeMUQreiEJnm4i9pBIYeqyGKxK5SDJEAgczznInMzZNXuXp/KSFyxYy5AItHT5
Ml5Mbz/ICIKAgDyaauXqZ1z2SZznRUj7lMoOdlDMISDkCTKx0ff2R2PE675amUc6
fF9CltQ3mnpAUd8X/ZOjLaHHlHK/g2tYQ0/bdsyoOXwauYWjfwqog+x0BL+fCpCb
Hm5qi+wURXuaR5FmgJrsivUPPl68nyXszTlwjeDPIw20HaN1UjXxwZA8/QO5zqd6
nMn7vmRcZqRuwp0D2ZGz8djia6hAfCcTkuHAKAL8gJiNXycKaGTMC9/QveEMx8n1
hLu1zsuTU7I1h3fzYRMkSn7YBT0jGAIwBsAJ0bjnIJorfkLLe3rMMfwsMwzuCRJ6
WxIc0jU07H1S7/vHPVCXWFk9mnUDc6aOpBwvyeou7hGDXlpT5EbSHmsN6iJOTxk/
Vm9QAabZuAtSrT9+mkxU51lZWObKuu3jOhqBtXfY2InKKYAhuKnlPm9rQcQJHDeJ
j8LKukqDCIbeceA0heZxES6SpsjxxgD+FG1+fs+Hj4K2+3vHFPDLR9uH+MNxfzxM
rdIa2P1sw8XIGAZOmlgDuMhQ2GHVvEFeoBYAtoTUuJGcaKfDw6lGozrq5u/iANFi
hn454hnt63r0ymFR8qQq2DTLepya4QsiktEF+OrqbyfFe6XWQK8EhYZ7S8m61TDQ
SKwE9VsfKVtsKqFjaWpSiAQ/9kkDCiCLz/+kWXbjPpwPRCtmhY94t8+Q5CgKIC88
Mwx7iUl/IlQayUtK2ypIIH0Ge8Dc1w/lBUDBcL6s/nNuj21XidtBvT9bhfiRXzyf
bCjekx8UEFSkUqCxZssYrKpDd65M2dyhxUDpAjKQ80o41SnGB7RbkAaQxWbuf+I1
FadrepleQ42qkIz9wKKMNyw2rvTUu/tZVeFUUxjplG6tA/A/UO0+fe+vZBM8cc+C
6qKa0ha1V53zyZ8Y5zQM1bW7QTy3xZPlBdPdHNV1tAbiypXeetUaCVVNh3vtBm3I
5ogqUXCCFhLj09AM0qG6cNR7QBuSdOC5FPiNSUD9I41QdjcDhcMpcpg9ZBxyWNnX
nyNQqcFxvXjowx41+UGsjqJGRaY6AxS2UmUraWWokD33wR+XNLOjZYp13Gf6LE6L
jv/FD1XOAXGJGm8Jc543gpVEkegSARrHP/f9zwYVDVL1IF++OutmpPS7w7hRbrr8
GfSqPOOeuei4sX6hH1X0HId/pFyt95H0Fe9LssePJtcEglfBkP8M3migQ+Gx6bQ3
SdGC66JxXEiSwbHBwZlKmn4dq1eTZ7dIvHtYOA3H/99ThxIvRjsPuHr5h61TUSOv
u8WeLFkMancfQfu4uKTr+D1BTVkZrIMkIb8kmdF/ndUZPzvZkNMWM9pai8ESQDc/
LcMtBO8D+flbHM6xWCIB2+7PUO23d5wk5zxO8txkD3g2BmCN5vSjob/cDcaEvIPg
28r4iRIuRcwwY9V2ntugIwQkrkrWK2TOeHGWECozThNRrpxYXQnmXiuDBBmTSntY
ZY6OPoQNMCMUH9PpFxLmUBOcM8L6KaQRLuaXcePqyxyBTdVjmWeB7jTY3Qkqvpor
F7QKPnISJ0fKCJUwZwESxt5ENoFt3jgVQ/ZF6pwjRLwF1Xi2ARWtlZlSioLUlKIr
+6kMqL4qZRvBhFuPhWt0XyDLEyKGh2U0TcHJLnZeU/eBpzPjvnLbCpnnKb3WCOuH
f0+B/j9bprwWw86LPxFJ1OupeZPlLNPtMSKUqsyu6fwevU3L4qMkohqUntF/KhTC
bSDhsMTtjaBMhjTgYo8m850gIa9BY4l6UhGdTt5F1QJmjTlaOJgPbDOHQz2N+uE/
mTP4ke7tOjC0yVAAjpoPVoUrYOdyVTOAXsfDybKo1Yeh6pb4FTo/HUjhbTx0n0gU
DqG74lhuEHMHZbXvUXncqBOHS6OrUmf0MfV0lyvCK8Dg/nfj5TVYFEPjHFmfIvaK
EXQqNMlBKAwB1uD4FMcz30OdpeIztuKiRyq9diztq7q19Wrt/2OpkgSC2nyX7QbY
XscEiDUoa/Dh3/kUOYKtRv+X7j6aDJl8+U4zvm8RmqmFeS0qJh9YKdJpDDOQC4af
HXg0rCcPpiH/xxchE68wUHlVzFVgcL4b9ZmDHlaI43KG7BrIWYa9+aBt0S2JfnEi
TOYfM2nXXoC04KyRe+WDKCO7ZkfEixU+KCHpA0B8rP9K/4bGIpLF94hGeaWyetWk
pybokKcM6iou5nOryiMV5ff9HXyHDRDNeLh9WVW3p0DZ5Kb1Ds56wlR/flSwds2Z
EQZN7XrkwfqxGX66prhGrSW1UaNc3oSdpRgETsLntgWKUiNuYgrcTpr/CJpdFedF
sfFLMaxtRoDFLhc9EPgoTl3ATXRRh/N226J8bWUSdcmuVNQfraW8EO4tBM4gaZej
s52mccVuprMj9YsaZHk1jsgtla7T1jIAr8OuJjj4fPc/rDBSIDugR8Geilvut23j
UvbqhLoMgu6ku7qMFBNIs/BVBTVNR8FSZwt5HG0jK0emAmdxb/o4ZoPmNbc7mdJr
IZN52t0wMaBkgWdWRX8m9jjbSC2Wn01hAFXjyfHpSwD8sl4aV3YTZYOsbsTvGKYr
faz26kt5t34jFOYA/4HUC7ul0NKKIm043Li5enCiSeaH8+SbVZ3BE9RFvedzLCQ6
ioIpUbcMFZ92KW5OATYzy4gz30KrjGNOXdJ4fzAQwjiI2ryWinU1DXuujJhJTpUO
gSV1bqKAI77kKJRQAMlEKeFuzqnDLcYJlHdCa4MeVbyomaEiCMcD1H691VJ2HCLB
Z5+1N9fyIpaufahol99UVRawPPsKSTtlwwqzEtq/UkbO0MBO/aa1BC165YhutT7v
35Ul2Ja0dVOuA15RzmPBJePtw1NJ54kr4LbxU205Ya2uTYgQEP95epnT0iTc0Xog
Z6NPku6o32Um5Phl6Fo+huKbQOEJGGpXdP61AkC2/djMR8Yut8NJ2i8ej25i/ZFd
dZUUO1p3vq5sKsKXWWNX9Re4vEjyShSE574YfGWkQQrWNvkAG0ePqDlA0r1WOFPV
LMBzYV2MK5X26EHquHDF36/iuYako8V128q63NYM5rLT7F4+d2DqM6Jcb8Vs7o0Z
z+Q87dJfXzd6ul1hoiWzdjZQCTmiVk1TuDN4EPDULUm5E+6sIPvfharq+EgmY4xh
wrb4+lY45DdZ2LlrB8QttDkdlFmO5o3JWlTEw21y9YOER3IuKqV0Df3LyG2d4yC6
dzFVBv94SqB3tRFeDwcPzAIuNDIE0uaY9ileTLvoUNOwfExQvr7b8eQDDwXgu3MD
H4sIy5xXJj91dtZKPS7wrO+3coUNu0FmG6yHYNgcJYRTpDcq0BAE3EqO/+THzFhh
f/ZXAXq+Ci/ycy3ejozvLEUi2ltRT57FoM5O9axCbGjbwno3P+me96bkK5UszeaE
A36QwM1qmbB04OgVcpwhSmReOPCQcDStbHhQYB1Rqkhzbq59NALb9AyvnM6JWFhl
VHh5ctyfEkUUvHpOfX8fesxofFdGRazRrwwEH0NMrifI2ErokGrXzsGCe8H6Bjef
kBv2iumyyVGsQnc2csFG6HBxsMzIHgIEWKv/eKczXWYM6nNtY495DgPONI6o9BW4
Eido7BYXJP8lwAzMnZMkFpiG8ZyOPp3wluXYE4cPi0tG2S9MhZsGvnu7qKqtGt0J
UTy8qK5u6jVkfx+g7+JghZKIeFbrBgLsaB5r00CZHziOUnFZACKYFhj8nUZYGvsN
mqtrgFfQ/jLyAZIGr3r2fcyK8++gsd7uU0rQvhhkD2TMbH47yqx/ClxgfflPv8XT
wIYghIaHQSrG2JsB7AzrWAyjJ6U6/g0FMhME1Avtk3L/WWJHuCLJoXR1IwD7cg7Z
l0ZyFZRZmO4AZMstfk+Qd3W0SwK0p5DEWOm432sCWCK3z58Nmz8+9ey8Ug3qpiOx
49/ccls4rUvp0L7lxs1391dlwpkR9iG/ALFz9levNPre/bLlIlm979DxwGdveJhr
7IQ91Ly0HZV4G5TtVqoNpzv8ZMsaWB0E6nAGWUGtRLxbBmM99rkvprM2cRaISR+m
vDAc5wUNBiHjBVmEi0VgDT+ox4jeWw9FA2o4kMTmp0fFO0pRjrAjlYJkk+8i+Vbg
6oZrjapHQnjznDjnYeObH463cXC7aEsUgkF3I15ewB08mMx3rtPhcpLQLmIOWbjX
Q8+O9L5AIYThUc6RUMvGcYRKEtjW3niHFe+5AduCZjr6y33EsDYtwj2OR1pKtelh
xDf1tzdt+vQayv5+rzt16G6/iDCZ7RvhiC4cxYsiM09z8sdjb3HDtfuwSKCEE1xQ
iB98hZOLqckHu5CErtj+Na5sQ6qE00xrbYaU9hijhOFznzQ+G2XgcvHrgT4a8vHG
h16MTgXem7w47uPVFWiXyCaeKexq2uErsghBOpiGTf0oOZeZQTMGm8m4Qgg2aDqp
xKHd8Msay/uYaJWploQOzYaN6tI7h/GY64JfbiRqtmY/DqdJ8Ag/RwrjBsldVd0W
VSr2u4uQhqjUs6rcHaCwTd4mxm2LoU8sgrl79Y8TyCIzyxaXgmkotX51IUdu+6qJ
a6iDl3aXpqLiP07DJXWzFdNF8Dshm3oqmRAHLocdtf6a17st2Qtf+5xEzVwKpNo1
3fKueZi6WOQ7ukchTU6eZdK4uBWXOzWxrQq0wfAtw1yT98mc3f5tCVdVR+DCJ6LX
emvrU9cLeO/IjE9ESt4/Gk5JVmFZWkB+0UUJj9N2fI3a2/nRYYdZq5ZC8wetDos2
JFHcKPe3CZf9s6raHEr4uCPeeaafx8mzmBHh8K//h5jP0GbhtF41D9rhvg+ZHiYY
Rke5o9SAkvkoetuDS402Y9W6fEmr7Kvl8KrygwVEJVZPq2DUkQNXmXqQLyJixF+R
hwKTvkGdwEw4Jwg0JxUmIcxk0h2c+LNp9aOg24RIrYfemHbYcopdIiGfyMAlfzBo
RoL4byhLnC4vjVGP7XGDaw9kXpCWqhlnRMJKJbmzVko+gR5ifZ3sZYfChtxCnUdK
lCuFO7UtI8AQhTmATgC+eS8/PZuIPMLYooZDoM1kbxdNUPcmQyP0NUurPW0hvPYu
gQITKsledv+THVksmgLBPk6jLc/cSmC6NhkW4qzG9J5gDni6ThmAAXt91Gjy157W
nuwmqbsAMnNKwfElStZ1ymsMj0Smi+lOdDQH1//SqPEedxYEktoX1X4BvbnPNBM4
bJKoXcMhrid5CH5XtGyGi0wD14jfFeMCmBPMk2nL9W/pUNSFUYGTq2eTE1TN36cY
SnXi/3ee5lxbCj6UFr8uRKdBy/1zqLqgU+CS4g627W6heYcu4fU5CfNtoYS5W1KZ
mG8CJ/vGXnmSDOhI5E61d0P9kfxBi56VFZT3lYMl/7IxZmMdNhrK/y7Uuulnh/gx
ali4QlOBt4gXySo9Aet/atJ0jN/nhaMtGBODISSEtL8KaTaK0neDfJL5AjtFNCER
pVSGw+txJt2Ly+XHJzaLNrH5uD4lNL3W0wLT1HxuF5pznRTXSTCukQbQEdJ6uzPL
7LSFP6jj/SFcp87DLwhxSoosmEQEqsZI1Z7yA/8XbLsQgGpI+LfeahYANNZigPTt
m9oK/MDdQ8aqjkaexD/CVA8m7KSdvhyquuiKQx6yOj9aIQygWlh+k8t6Q9N1OAJG
i8vp1VnhVuUWo/MH9sFboNNFK4AxkiMaT7qEBQKRlEdKo8t/YCzFFAX42k0PCnT+
DuocgzLIhm0bU0QO1PKP15ZcN/ALK6WYiGf547LGERoF8Em7LcAZm9i63ieY7+y+
qqLneD631DU64Sg81QsJwgzZ/IWoW7/XNNqSAilXxWmLrF2YVbOq/sWJISpwvHoz
bXSYl3bey2lqZ2YmaK2QiiAXjCVw1ieCDc9Id3YcOcFweV4JZc7RZYIerwyHQQmk
gcVNAKvZWBsJZSUV9dMml8M2BRac9M4tDzA7olKf+pT+dNZgeZdip5nUNXjYLqBD
800lfIBLUFp6vOAS1CpGXVzEYikyyymJTMqP8vftxeWYOJdsg31sbtIjkvW6fODq
9RMXAfDeW22Ouy7sAMXSYOEqIYEi9vqT9+SBBws0/l54KvdgsXyMgCpjnfK8KoiW
HUjmb0l8U8hVJ3qM4ig4rqsUZXseWvsjbL1hys5xxeOLc3K3vgToLXccGb6qIrA8
Ue4u9NWUe7HNX7czfe4HfTLEbrKC7hncYMPE63GrhP3CtggKW3S7W2TqzgJijr63
eN1fFB9HPofpI2b1EJK2RFT2AAiK1nhpAdUFGKCNIisaIJmlfBqCc0KO+Esb263B
aTc/clmGZswSdIFTsh+HSa5PPgvKQflHFe521Ajxo3D/v6JLvRtAFSe+91REAbrE
2q0VE/93fJMYAkcclz78SNhFpV8oOfHwxY0THPNk+I4U4G60B+wk4hYhHthwUKK0
aMSE8CajXSlwkgZ0UAxoSLMHLHuGxjjdoW//p47yABPbd773gZAjNO3ztvV8XsUh
3CQXhZvLSE0Q7JrVWUc5HaxyPzs31trjRhvTuuprB7ypdnhgGIHGbKAaDTYHXa4K
RAsWSIqcXBMdtb3RWC5OtIyhtgR010Ox++VtFkKc13BpLyv96KMv+JuA+3ptytVN
CmHg1EaNslPN/h0KXYtiN4h5CmQPmMqE2f2hLKVK0qMqVbfxze92r62ADJspALy2
KsMdHcM1VoEN+CFyqlMbeRPn9q89pXyS3st3fKZYJvmGDwJvXY648f2qmoAwvZ+3
iZKDMTsuv3LCB5eAcwz8MF0dNkophUdx16dtGkHKLuEEhV1SpQ2lVOuUmlF2EjCs
trAhiUDq1pIsVB8kCzLwsZeG6TZiINzuP51e2hl0W52XphWKpfptlhoMmwgm9S5K
2tW7dtr5yGLedwoJKHKAWaHZ2MvxB9n4pd/3cv7znqejE1x4nKzdPWtNfvo+0dL0
IvLXs+Ph4s4Oxnz4ukALXhaJzMrzFi/IYsvY0pBpGhKNExoMVvdW7FTIL02ixh50
tFAA6iH0yj+stIE7cpjBsdLm86tGwVy7cXQWcsh8IAFgwnyd1LnT8mfRJZey6svD
ggLVjvuY+E89n4fkzClrRXwhfkJrS4l/M5tnHHMSHRZ88GXbVkaVfonyJ4dYj15g
rj6uCsXfiqMr7dtJ2RCYYqqYRn0a93HzNUxVYZll1rkZL2xUqDpv8fpzxHoV1RU9
hDh7ea94yHN8U4q9p3tG8/F7qbfH1EUsq/hYcTWPz3bOD7pTiSJZ9ercOkZDt+RD
f2r5ixKhvkXEu2cccp3DzMQXc8oRKZnPGRn5Gl0IelBpxzL5Asq8WOrJSj03+vHf
mtybEeFO0BF3GFKt0zkMhaOnXvsn15S7mr21x0VvliYCR3P3pElYUm4g3givQL0l
pEEMwG9DY8Xp/xshuXbe3/U8OAEbvYLJUV8yXoQzF+RImLvyT85afgdNKjemohwt
R748Lso0hp8vSxLqdxD6X8Jjfi4mJEot3pLrjsIfFaFv2/Yz7k37PoDmUJSjsMIs
mjt8Yvt7rcaULnKbNBbwzbnvfHOyudlJfGTY9l+UYQlfhdauJqUzSFdX43QjOfDk
eUkq7htoVKCiFdna/1/WUuBPuWXX2E6JRjwGRbaSt0oMOS6UwbBd/9ozdWLCxBXb
B/D6J+HrAKCeiX6xsiwVhxLr7EmJWexN7vv3S0ZCAY6QwpyqLuklOXgsBcXADNBp
KA+eCXpEzRlRiu9dLmItvIJsMbp+ZIT0djgtppBkAGXjyURr7mBACjssRto8DfX/
dU6WlDDJOKUkyDkT+MxOJtjM7zWDVki/XqL9jNbdUmHbaXQPZlFjM+cmMFgRRrWQ
Qq1kaj5GAOZRF+CVEpleCKRqxlc1mRZT3R8UZBsilNTrVYrHivnQiCEFcfXMuXUW
THx2NEme4TQGUKAW6h2uDwh6c8BRncDJqPEoLxwwa3cyqsV9/jaY2lMc6af7H4nN
ATQO/8gHctHgUTZur406kRF5nb1YJvqBUrEXnglzYmxa10Rm21JtzZpMWQZJ8m6V
hZs4MnxQGFjEe9SernlpEJFKkYIaFOSdxXM230IP7e34scDUYv2MMN/twPzkgyNK
0SrZyenOmfsG5v9BMrMfs6mhX+2ZAHoBCvLVcEihJiocmdjnRMmWAXsSjY5JzeY5
nblH5tCDTqNj0iiYFel9/oRDGcOVbZN8VqhkWLC37aHZRJNaAIFktcf+QyOlzNfN
Rf4SRWrr1krK+PWcm3kN4OLvZ2v3H/gzKnzG4gzaTPY3hhsvMIj258VnrVdfVnpU
WhUYWcLKIzPysIGYQLPG7A/K0VSuBq7j9nFNz4jQn0kBEnQkgGLF3guq1AYawLE5
2ILZ6c3DN39MU5nmZmnbenx/lDOT+fwELMbMIQeFxNg+qtBGZlqpk+IPZf+sT5e2
iZAzDVduW7Di1y33f6khulE3mYMCCqs1Uf8ca9KMCRdRTBEphJrubvFo0gOzn8IC
nM/xmcJJP9bS+cPphHwNLvk006pBEHWcXtSC1IX3E61UUe6nFMkxvDRMRfnk+Vtq
Zxafk6VvXNfevMM8bjB1kMl9g9W5tN3VACmmqOv77BPNq8BIMCOxH5bBdk8nJ8BG
qwGObQ3zIlzbM4N79SAkIcSjRh48G5wSiwfkbu8sy4I77+ULkXh2uXqUjXyRnVtc
Mx5zYu+xxBWm4HKuDCJFAIDsOqKDXm/PSQP8hHyDSl9tKiYEqwuNpCv+/Wgp83Ww
lsJ6a2R83d4+43c1/8M7YNv5xUuf2GufjGWSh3FUBYb+BhQxZN5PO5IJubbUCUBG
OGhBNYjzCNbHIahL5WgqmD1jR06QULG3JNpW14rlh2vmhggGoaS4FXDXDmM/ooxN
Hns6S8BkICrcADFs5uhJyZuZaAMvlIcvHPcVpC8du3AyFqiJHH/rQfWIVymgaLsT
64pdFHM8zx9KIiy5BbKAlhTwTXr6/RNUOpEhfWWONk86Ehty5Xq26iFFGm02IqcF
T5xGJ1tH/o1Xfv9fAUKPYCZ/qAxsZyXg+KnP4CMDrdFlISNLr9mk88XcQkoYx7Io
HpDATWUXGY79pIFKZlMC56c1AS3qdMwNWk2/LUuXp/1zZ8x9xUBXdqBcAV440din
ZE9Td4D9nieFyS7ue/giLesYNb5MQrd5Na1JkyZiEeF9BIPprq7b78wtW1yTcthQ
VPuCI2kS7OOfMrOpE/sH6+5zq2WqqwSyJzCDDth5n0FNWb27vJgUH9YIJPhjyPwa
afe9vFG7v3FF56lU2XIEzrOgN5BhbBmsUA7bz9Jk228lbO33F9WmhdqGytgWw74N
pMt+3nku2JczJFIxMQg1+pnG/y9bPH66xQpRgjBBWmJ4qGq+VZoJ2//JaF1w/j88
QZLhGUvSSYXGp5psqcOPQIqoA2a3QI0vqkXWxPRnnz7LO6uvTT+zZSIqU20Z5CeP
7UJMQrR70CMKqsHCd+fvYGOKRiHhgGkrswU2xvwYT5qYTZvICi6lM6vlCVfVGmWs
2LULjfors6QV2f8FtFkgDm4UGUCCRwx4ISlEDrOvfduouJE1cOLHga0X1MtUwIaF
e75bZBVuw+TDQdt4xH/U6FPhVoTJE6OZHjlVYaAEgk9M3lVvBeG7h8fCnayYWabe
T6Tbl+1qlmrpedpAdeEoSJLaVxDOEbnNYaJ5pBC5GibfBkEu2vFQpIaekKrNRFaS
QEoVD6xpBBm0OEoyXgLvTUkCHcV97DbYaD8G2bZPtBRc1aUoKA9XYO20RfLREWUh
cfXO3u21mpsnnZxrhVydmV4ypiOItZdgLaCow7lyLwyaXIVLQYzkdp6mPVwWjNbg
nH8zaMjRJheVjp/LlRGXbAJ0S7UACvwuQV7a43hUOw5UJjWMXfu2MmY0DC6dbSrT
ZAsw6csX2s0infahl68Q7+U5qBVq1VgJJKyNDhFovqSsDf8IeZDp+0XC0WP4T0KL
GbaEObFaJjcv4vbPUNNjlF+RbCxWSXnr07uSZQMgCFTji9EA3hy044FcLj6dPEhy
Th/y3q2zIqw/nvx4T+0hm3GxI8J5JRdiazEgbk9It1g7PMUf2O0aHUY6MQ6m12Iu
N31mQ9SYlJ25UqPZdOsuWtEEo93J97SmBBbGuDE5Z6qqfgE0TMKoW2vP3DDIgdN/
ucSF8yo1+csqLAJpAkhC3KXn4UjahZHcOPJZre5LrQv6MIGWyGlZDoir685OtYRB
yXhiBn4c8jwZHlzyhLQPCOYPr8rzTTnOC/wNFGGUMFrbAe+jg8Z1a1EsW0G46ZDg
cEFIEs4YCTAtksavEIcMaOMy73W4TT9NJkodDESrNEQUZ7osaVUDkN5xdDhtLxjP
mSfCukjPgtpABHsxYoYw8hOkpPSGZzOWliFu9BptCIInGfPtQ5fh8JBczbFbfQt3
aHLR9nTF0ZHlEj+8y/gHseqEN9BwzuXuL453qrZvSCGNlTAiLJySemzmVisl0+zu
qLLboHBY5agl6VyV2Z+yJsHeYSFTt5g8oEema0bF/V0=
--pragma protect end_data_block
--pragma protect digest_block
vYJbXNstgLzdvjYFD1l8OFLr6iM=
--pragma protect end_digest_block
--pragma protect end_protected
