-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
jtnxAL+J6/0SfxM3f/YzfDgQEe6e+MaVCIWBDjHlGb4uOwmjLjH9PtjH+jI5YnVf
6xNqDIhn/7qfOzPfR5PQ9Tp8y0gHEEIv3WzY1NYNukLdfWxA12YcPWRJNrOtyqZ2
qeuTCWPcPoMUL5aRIPfpPVYDhq5GW6Gp9BG7FReC41o=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 4148)

`protect DATA_BLOCK
+IAYJ3FGFIyG0JT46yhqdPMH/R8sNk24RXnmEHcQlm2ZnU3cNvuWoc0Vw5xJrulV
ItuI9fOwf2rA4BbdwdUku9qczzUCGhJC+NBorBafO6GJksBGqI4lfu3neBRygbPZ
QQRTUzvIT0SQ8ITf2Vw22JoxoLrW+0XVSjoOzh6bfpSkusuY8DgdmeIm25yjsK3b
t3e2hS65b9ZHRSuf6YPhcr/3rQO5D7xfx3wK1u0Z5IJWpX/nIC0mdqji7A0sKFxU
1TCtmtsF0QRaEtHB99uEM+hDfIJrERz+TNvY5WJ6/dyO224I7E8H0PqJUUw6tKDb
fnyo6DbgDGw+pkJ+yICLzUMY0drujYinz/NqFpPDOUxy37NKnQ2tSZwvfqeJAqd2
jF76ygIVWZ1G4cdW82FxjVUN2yMUzjWsq3MI3od6uo+IMzDwOASfE8h5pcW+s41i
pi4uhLez14H9TuG31op7h8CCL/0TcGIQQb1ivwAKOtgaUe4qYLBI/BldC/wf7320
p62FjGbf3YByHvjLtHucjrT8VD4ubb1g8njzw27zhSU8izlP1aHglLHcX3ba913l
kOZGdQXdQPgRYnOoKNBE2GRAlpNrRD3nYzk/P04FwAjppKhNEG8tM4vknNm6CgOO
TrBP0X3rrQH+CmqOhM1FItvVOWOIE26pD8SYvflCnWJ9+oX+lLsTwvHJXpUvGQIM
a8dXXU1uHUN0whCXVpqug6U+XPdDPumv1NUd8ISJfSF8Mgpvgwua0y8hTGX5jS2n
S2SOmxb6uwa7MRdnrtZGmki2SCTEWl2m+EWjQigRLBZR/O/ECodS47rsQmsTDd0Q
2mebLAq6uSTff1Mb3xzyrYh8N/e5+N55saBzQ5L+vLubUDL9gnYzlNs4a5hnq0Xu
gbGjaRSLn+OZRBPteZBV4IPgmgWj3u6uw6mwC0wiMcLpI9Ywv+VWvz7D/mxWUJzu
wQ0BZCDjHXXLo36whbVMuOdXr4TGV2EXuJjsDZUuzRryHJJWCc8etG/e7qjpw+WN
727MOiZKkA9kdHxIravchAZbuCaWKnpmUBtZby8g2yUdZ5UHZ3ThyIacBU2SQDiP
EN9zSZRrzLKGqpM/SpJSVEAovvJy6pOVZ/YpAQW4i9zDZUEayze/tfto8abtU++x
I2KSYaYvHS0h+VnlccoT5YvuBLCSW8HWwU7TmclQ6UC+6z/HgGFZZGX0BLOWpejy
Vz5c9ViBN65Qvy/J6+bueO0YB9vyWvEc9V73oUD4gHOD5TCyiw7i+PoMoPVBNJFo
07pIE4owbOF9+yrPjGilR4RCHcrrBJ83hMTyZa36//NQ5nx08QGkSTwS5i7Fm8QI
06LPw+B9n09dcgrw/TdFmL1sDhJYZTr5r0z7hICdzEh8Z23+Jz9sZEadiQiU9H27
DufTDB+SFK3Q1YPh01LEYehKkbsFGB+GdJKFKyYtekqfevAETE9xUyzPyb0okUlr
NT+omWbvWLsgQ+fB5SFTT0Q2TKhix0+Kn5hMuj0SWJvvMUZtO+PlhyJiWrNuzjeg
YkrY9iGND3F4Ex60XhdLd9ktMKW6pC4SDrHSsAP/zlXGaCydf+GUJtvlpjgjDzp8
6gw5AqLrFtrVt4ow/UUwHimM/9nN/l+rgPjioipREWgSGe33az51p+ixydNFFO73
qQYr2iWkkH8etM+4XTPRQOQWni+1Df8xCpWghdN0W8YknOeGQ2yQDAjiUo4iyfLo
Sd/Y9OwKnrqxX3qwroP0dl+TvXB4ROhkG5HGjOGMI+cqg6anyiMDZX1E2JRUmXOD
qq6Ty2rF7kKuSZjbI16pHw1abBko37qIRzwDfXoM3Pp4F70HCSBEnQgkIy+3pNVG
3YAFKD9HrpoQ36H5jOwQQOBRZgBRQIFptYX2DMIGHsjcOuQ/phc5FvKAMVZWuE39
GuIJs4/P3q+oFV+73/9VLCnd3NfzXMFvb5jn/Vs24CHuNrRrKpOup3E0Q5IjCTWs
egXzpcJ0LxkxXADPwP+Z80JR7X+lTAS2pmJQ/bCXS49sxou5KR7yLGAJVEwquIGs
bv+RPRFDk7my5GkzzfN9mWyaOZB5DkyQnA7Dqmp6m2eXoWDgbR3K93XGr6xrSXL7
dZdRbGbS7UXI50Hka4MmPgi6E+4PwpAjrTr03yU53VCrF7mWOTgY3iHPwJr/8A7G
a9hsGsPUbZYbJv1EF0c1fvhy+qpoNrGpx+SllkQxCmKpuyxXsHtRJTRYprJvax41
HLA9P66XijuO/+uBglFDVCsof7DrsuKCmNvGtK1Ib9f/nJNY2syXtq39EeXBmyoE
Lopf0kqKAe3ePWz+IU+1jDkJVMvhSUo7Jv/ezxDriKhC7MIgkTrOFYmro9ConZyx
FoagMu3YEDr6c+IhY7n0x37TS2Lt4yyRh+p6D8YypEPfkr2W6+BSd8l4ejTJFtc7
o/SFatjwvFxsporELemKD8aEQu+tFFTg9U3pK5OJLIEx2MVjVnPOP6bbVshf1/go
BvAkLVCTGbioO98atYFajda9To71dHPGpXDrAyVqW0M4iLNt3kVMoI51I7qCccZS
IKkFQ0SV1VbOLM4OVDYyPP7fNgQ6ACd82mCBf66XPxY4U4Tiaxg5TixwriHPwQpz
llGeK0dID5QU6SLPHkKd6f/MagXSIDo8gkttr/KVwfbdc2KW5X4Ni/rBRy1S4C3D
W4nhXnX4dOkNCRtyE3nk1okgVC7VpwxngJTayMluI7TTRyoPA3BbTd9KdLepQCve
gcfxqYg0XJIVinEAVjSgY+EPoSJzJiSbQwnEAKEj5hJKk3+VG777lDWrq4NDHyFB
XeKEbaYVl6EHWbiAw5MDDrExP2oTA9tqCBFAwUGMN0WV/aFNXRX6QK3zUUTeQCjs
VvY9Kc1Hnen3pq03rJjiQUBUx0jU6yRXQZiiMEHSTT42LZmnrkA07zIi6ILCdjY9
TIIKdlR/rjF2Xquxcn0EenuS3ZLAn6jVKC0jAwWciMkLMCOa3wjJwsFeghTr808x
6mKcwksAiRskEMu+RrL6AKgLUjHhbGZ+enj6o8Y0yrwKQnHwcQX8uQ800p+idnI9
ZYYRyuox51jxXGsBis05kzmUOzHEsir1axckNDXpE22Rxtl3/HRFNk9kv/yRBcZr
287sqRSQYdeM+R8sK8/Gz3ftWzz5Oxz6UY/EnW5m7/YuQrVV1Ad/TVdSYNE4bIAz
s3GaeSj2TUvVbXf7eBG7xS4lhFZYzc3TB0/oyq2lukAN3lIMJSkJ8iuTcrkAX2SN
KR2ne+WlT1vgWKHLmebiXVEq/V5WFxRK6HQKLET+lQb6L1Fj4RR6nKUg5eiYrknB
UHeoVjLAPqy8tBWuGdCpUh7eHZSTofapUaZImMNAHONUT6FHvev8QhqmBKUyCIv4
UohecXVtSTNNfcqFV4CWg5WRgk7cCiWfg4BtRydNDitLoU4PT26NxldvICfiziuA
DIfz9Iq9t8LMbznujNCZC1npCJ0HcgHs91xAQq5zM4CGn4xNLpsChBSWezL1VXOf
DyPAeJ9duTElBVS1TbvX01cJDuwUMHzfT/WAagfI2Cy2HAu1ajKcJYT1q7oEXYQf
LfAFYS4Yui1V+KPuicONV/JTUxBbdQwd1T64Y1QWJJ1b+55DENLqTv6owdiwSOzv
KsVNaqmk4sGHj5h3frgGRc+/3Bv1CXawOemBGukA2rCAsb9fOGSFBjmoPF7f9KhL
ApwNf1/Y/Aozf2hFAQ/ITzdAJ4ltkRE7HIWW0P/V9osEp0MSyKIlit7Vd5Id0Amq
HArkWIe3kTleSkwtZk9GnispwWLDDmHeYPBfb5YxEK1wLPpaTvXeqh8kIwrNZ2P+
hO7qz1Mrz71pMDtPjayUalJx3IKdqOLPPpUvS6I4ctUe6XVOoE4ansh6+qwX0//v
YQDnFYRsgbV+5G6mBjlr/rRGeEsz8Z+QvaCMKZu5mL2jeGU2/94gji6hdgGRtg6q
1Bz5ezQTZ6E8IqUdnqteve6oRQaVG5EXHUNyQC9XrQE6aAS16vLf7mIu5P+25Xm6
GKNPrgJa1+Q7GZSq9AlqZ7FRjPC9C+k3lmbVB9cNN0wspYGB4AI818VZA6ZfCu7k
V66iyjmp413E+g+jeKo/468VOJVQkKQU8OTCGw4ck2A1B7Bkj3azdmq82V74n045
hjLsXC6fmaskteA/RwOxnulyB6NA/tRgDl7EJlFQHrqkoqz+mdZMz7JNZ9p4hMwC
PPwZvDPtfsXF7b1WV/EeqX6rSwE1abrZLsD4Re6muPv6jerSV4xKfmWATScT2Uh4
SMq+E7Qv9W46FBpdP6HqjgbwFXRgILiBekT8RyEqcDCciIj2wm5E2lTiJupf780C
nUXoDtiGq3ThcZibfvxXdrs2qhfo/iK1++D2ct1YA+sRygeoORooMu1LcKEywvVc
0V6rcqeSOYASNOyIz4RiKk+mgMQt6ke6HbuLqRzAXuvSHYiUYIVDSClr6h2ybOwH
yROaiU49ckDvVqP5Z3tL0CYvyLQkgzyOMkwRE8+PK5sXMxIyxOdhpwxDdoz9OHyL
fNaejI5TPLPCwZV+eV9gY/3Zi2zXvZx+5Yp7MESm7mZHAAHGO+ScVTgunUhGf4HZ
KXGRp5l1hUls+LeCnv/l2jtHmK7utZwQVm5FP7aPARC9Lg7d84AykPRn0hOfVDR3
d6bD7ZKCAILl0bo0o6I4Th8W3yunRYDeZUxGDBD0JywhNnBTI8gMiTqTO0AvGKjP
rKVeNwfAQxfRYS2DgWNO7zYCmZUwBEaQ64HkyALTfOQbZStCN3v57JtN/H+Rr2fZ
e3EVKjDAgam2x423dDUEHeUvDHs+IT5bX126kDTZK4qvMh+Zh4p5pbVPP88FLBqh
YD/UT1jo1n+Ecjy2jLFHWHsGzRFzTAz17SWEPyI61T5X9DCUHRWwsyvqssXRA5Gx
4Ccb74wDIDqDFEwa/tOCoFNGwVizazkCKz2QOi+6opPIx97m+7ZYZt5zDO6BbH+5
ip5fN4xip3HE0HoyHbz6jrSJxzU3zHp8WleYgXw5bln/uRHzH+aF0i0MNbZy7fc3
MWGIy4UkmIe9F38+seUIeVtXABmgruGLbtBBkdqcX5Xyui9Bru4I9WkD43jiMo0G
v+VRizQOZllm1xsIx3PEBADk3Gxe1JZPlNd8AGdlyGtQC6nLjtV3yL4gNTPx/QYn
zD35m8AXWF6HXKzAh4/zTZwDq7G88ozzSQJrMJGk6IXRuR++hJgbwKfsjjqSyA55
sPfbpjoBK0xfu/f7Fd3hoFyMyMhc4ai4gWtXDFP53dFsg3KLYSbENdlI2yskc3Gd
exULE08qfhwhUXJ7xR0IJTy9cMQRHCNerwDwYEVxoodQJ/091ScO0MV/JVfBPD2p
ifOALYVWFNQ7tEGrxZQLgOt5Tq8N/0sBNzoB4j9CVPTS9/A5TbjiP4NVElrWefn0
AGLBFhUPQQ52rGdnzP4w8byzEuP3JodpFJqJVPOb0P9FlOxWItH5I8PqQeqDv/Ao
wDLZoWsINDZkvqp74rp7bS1oc6Qxl3z6Js7cHP2+9bm/i5h40ytvpcZqFJq19S3x
`protect END_PROTECTED