-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
--pragma protect begin_protected
--pragma protect encrypt_agent="NCPROTECT"
--pragma protect encrypt_agent_info="Encrypted using API"
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
--pragma protect key_method=RSA
--pragma protect key_block
Maxc6I+0wR9u75ZN0dCJp5SpBOiWW1FZUM9KaOK8IyBcB4S3kNLePrsGKeIHhI+y
NZ2mFC2rTJLr0O97PShqf77Ezj852VoztVAX2iZyYipkRbadCWZX4CBVM7PC7HOG
3bKQPVHq0b8QWV4Dv77stDSNJel1iHUy3qCqgpUDcgXHD9puJo9RA362BpRhSRGY
Uu6Co3hTse2/hwVBdm7rHZC1KF4TZZg2ptgC6LCrBI6ESsL3IUNbynyx/Umgjqy5
fsWx4E8Mh27Xt460ugsUt3fC5a8NKXRAvemBL8C2oKnlHS0URqpTOaQhRkbDaJFB
NuctvsqlvJUyCH1oqSKb8A==
--pragma protect end_key_block
--pragma protect digest_block
X9i/gHTHYZMKo7SXBABTxEIi0PY=
--pragma protect end_digest_block
--pragma protect data_block
FJvFsj5Txjjhw2/zyWZyTUQz4HrDGUqDYAa2HwsfBMDH2qfyPVAvFapDOT/CzEg2
QP9xjAXyeeAj5wGbec1bAO7qoGPByQtXgOLl+/8ZZwBPHYLGKTbbOnNe8SnSpFDz
pFxoy30ylfPv2mrfBZE1YJEeqbZxBgsYSo4E5OE99nK7aFrRnRBqPUt8R/OBB6v+
9xaeTFgjFj6PzLOMo28T1TafWeh/byXvIaYIkgRLVUKFUapup6jaaJcvycCS8EL4
B6ZDZ1779Szw2dUtCzDkDw+zbxl8qGcD6IANWuUa05lgZ3wxnhsQuQT6lATbJUdn
tt7pjcJdPGYx5fD689aGo3rQvxX1HwGzXyUowFZ6owz5FWPa4A5sTrLOhdbeEkpk
3lsixgZYwj9PrtE1xXcn4upUTgmvFboLe9bEKpD0dODtEhUjCTKMyhXczYlrjxgP
MTkrXSECDMr7Ukho8ENWNFJYZG5CGIA5bRQmCB0b4u2uZHu7ike1w0RTIemUkcQ6
dzXpbmUmmONJTdyRJbmJU1Q+CFX5uB3wDsS5I6LieFt7T0nitYztOEBUYIm6kN+G
q89EODhw4fuP3NdjFyZ5qO7QqwxL0etn+7OEvfATXYw8YGiJ+QSDtzpMgx+oIO8I
3pL7BRJPA3ZboAT1xGQVoWkGWBJLO2XwIcGhRzyr7lQVHE2sW1QKXO69VI0/JtSv
o+zH+gXzqYx+nyoPr6XZ6nfY2/mynQn3XR7TuCotZ79JCr24pbPKUI7YXkaFaVjT
CHYDtz6LEuMi9vfwflQF7Q9hdCVcC2eEfxETtqOgewlyt4rK9AP/IetsSxtB1P1e
daAYHwYybyzCMe44AByGe0WJL9tY3931UI6dFkBVnTr2q1rcjEDs4RnIVWeiBk6C
CWX0O7K3+t80BD04AVUDgAsOs56bW4399qqxm2+3+dkwCRJiz9BF0XOn4Q/BI9Q3
EaBZfu2W4TDsh3uf+/DwJBIKA8weGZGXLMpDTRPMvz0rd4RlMbdb7FrMPm0UxjdJ
6A0DvSsas+Xzw4gtMvVgV9dqTN4h0vHrhQ0nSYTqym1+e1mEm+4UvVlRyUP2HHkP
TGqxiF0a5oJWjBOvqfkzbiVi/G8YhBjpx0ON/KRvCysigi9fN3ZrSwe6k3CJDiav
bw0cuktqCtyLZpsAtw3KUGs85WaT6jnwOgPnesWd7z1GaYNMFEcOMhQ8N34aDJnC
SMN5KjvqhJ4eKkirxGS8ertkjHHzyyGNfHplQySEdC71MR8n6XjRAEq/fOG4t3pW
IyjN249ezhLUTcTojx8xjVss7NRz4m39wwquVUZ/wfApVDDnqeH6uj7b+PtoplIw
xqH1ETrYnGd5kvqrJInoT3ac9Kx6j15KwV848tDKAK2+4oNFG9PgN33mqC8KfVgy
/kmUYqqdMtHwaftE05O8SfmPhCvkGmmg4oF5G9FdUSVJSZzLJPIB5NRFP7CzLbto
idMGaJOweIu/gBksjeLVmsfR8f31LqPxB8+qHSyuJsMRlxSWQcDRovFA5+5Qh8lB
4tDAjHi1sDBZHJj5Rgg+yaTfXGcfV7PTCuKMIO/fXWVmanQzcgi/XX3TuFGnKPyF
B4KK+haUiDbNZbC7aQUT8sYVPBPceQ229yScaDJ8fekI7ayaVj66+dKARXYe9Cke
2tesyNYGQDiKxGMhJwz/7g==
--pragma protect end_data_block
--pragma protect digest_block
4JcgI9HqOhtLzhisoyrj5DZxZEs=
--pragma protect end_digest_block
--pragma protect end_protected
