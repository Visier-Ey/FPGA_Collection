��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���d�v����0�i�=\��A��?��� (��1_B�f�	�Ѻ+|n��y��Q4�]�aY�����*2�y%����>��������K������ �
�D��z�z��C�y�B�� L���,F��+*2 ���n��E�L�n��R���DG���:L��$۶7�V[��n��=�e�ʨ����P�����*�&��VAHi��	�P�[�mY��fv�������}X��q��?:�偟n@��]�ޑ�7��S�l�ENm	����o0�����.�V���6p P����j��1�k�X]����	��WO_�����	_Os*��Ks����^%y�M,�x���@��ծ��1��W�"��l�/��O�!_0�2�X�|�ETL�>Ew�&�W=K{�F�#�t_��Ȣ-���K.��6T���x��Z*��!�&D٭����,cg�[�;7�+�=�Тc��>�N\Z480M�N��A����w����cunf����}���V�q	�F%���+⿖'؋:��!V��<IIQq`yW�Ul���ƨ����]��f��NQ�G�ͬ�5�ȷ{���'"��pHA�H8D01����H1 �r<�6���Y���>�����4��6r��{(���b�t$q��O��6E��Ꮻ2Y��Gr�,ge��AK�:���bG�oJi�	�}��p�^��+Z��|��[�uJ� *����r$^�֙�p��W	��\G���O�Yt~�A>�C����6�jl��}ʃ�qa{:8g����L�§3���y�N�b^��>�T�f�K��c����Z�kB��6�J�p�*������l� �V���%��!�`�E�b�����]+�~h��g��,br����e�:�� �	VR`%b3����^Z��=ӄ�r��Z��'���|�[_ӥpK�J��0��[�����E�zh��x��BaH:
�m4���Ǯ����&����V����X͖��#�ɱI}�|��X���Z��YH��� �W�L�A��2�\�/5TMd���H����$M����3���"�vo����C����v���?`C*V�q��!G�t��*�W�]�n�/�ź.
�v��g¹��S��k"�*cXY�����R�ˣ�������|�H��rw�I����[��d�л�������@�Y���U2�,$�{!��(��@��_Q�p!n|���*��*"�v[�� ����f�l5����|G�Z"�QVfT������D[���^�yА�jy�ft|ah�{�0��ׯH���!�%o� �sG$0{�Ů���zW�g�������� ���/t�)�s�S��H�/�!44�b���2�62F�U/_EvW�t�a��m9^�9'l��FP�4^E�g��G�O���ʔ�����R$\9���;&9�L"��z\��������2�Ӳd�aCv3�Ӿ1I��y�E��Nma��wp��{|�>����R�I��t�!�<±�%�y�e2��6-���νO��*����o�Ҩ�e��όAa��X�Zy��;�Wo��3 �x��C0��ߨ�ˋFnu���)�F�j�a0~kqG�o������e폪��G�F���%W���P�S����N� �D]�O�|�'l��д�m�r�M��ڔ7��ݸ�
��B�Z�~���\d� 2���)J��N��Dz�;��-lҤ̺%����c����G�.�` �A��"A"I�����M�a�g�����k8�?���J�~)�i;P+i�wi���~�gx��-���Z���F�7̦�������HR&@�a��oe�oy���w�K�Zv�
����󻋞�,sl�����5>~��+�*#
�����n�ĺa������|b.��4�u~+P���i���ugB>�jo��UJ�#��޺k2����A6;�x�	���}cJh�J�n(���1ś8=~�GoMv���O�������u/�
9:�F�6�����9��'{(@ͫ�ۑ��k�r��B�Q����\3�P��e1xjF��jH���V�C�d!�\]P�r�w?a������C�Ƨ[ؼ�s�_��윞]�0) VbZ�QW�L���ޛ} ��*2����a؀*^�_:��/�)DD�
����BdI+q̼)�8&7JA#���Y�g%�:�'���5Z|���!��}p�����yŬ~�5�^�D���TmI�3��4S���
�z��|"�(�9glV�Z�=⅕���
w��3�o��@�w�J��^x��Y4��o��lr-AUo]=e�e�DS`Z=