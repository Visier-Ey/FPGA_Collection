-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
cGRWXvjC0PCxzZf+k+rqmkgV+PCJcgIf0aMXSD26fLTD8Kyzk0tBBNWLkAr51uGzPonMsPVIr3ZB
8pbRNaUZML37myH12dnOx4OKRl+ZyRq1WJpZQGBjHVRVdW5geONp3wrU6haI8eaXVH0ecUHbGIhF
BDSDVtRdL60fpnWyTA9UQGaw0MkV+fvcDvze2h9pXpzxJm8B5K8a1929H/LremUq/lsqfWzA6lbu
Ak70DUmm0HxWr3aJppRCB32bwTCrqCMaZuU8dgDUs5C61VWpk3rVc1zQAC2brhmwUEKeylqelWMg
3CI1w5oUgeqQQwXub0jh5VFRDI/z1OUsTMLbCA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 24112)
`protect data_block
7Xk40mUuC1RzK0KIdHNXcVxdigxI0fVE6dAZqalZS8++GKDj0vNesC21HWaLFUkrEpBKBtU0DhXE
BD7Pp/UYITOyMVaF3+ZQGgWh+L5uWqy80JLsQ4/tT5pz8DSJlU/gg7+H0GVZVtJ+ZQrtYA2f1w7J
fqvk5JJmUvgOkF117CLY6jjMLoFickzTTtKrieizRCHzLJLohsj6/Pr3sHnI6qEZfLZMDyUsWGQa
2CpYxeyoOdVKYxWnz7YJ5FLoyMyGQXtr4HeEL/lhQVi8jAMDkzf9c1aKRCaE/2Ww0hgzik/04rPC
kRz4EDMgcACsQYItOYTfsu62HvyLcG9eNMzCFyqx7ZrCXfAfUxKgbZzSsY1wSylTKe6V1NwHQBK1
2POnFD1dSPLC4wVBgxQ2aV7hdCLjIsZh4Z6lkRfpo1eLIfFXmfVt9KHH+4fUA90lFQdeanJ5Vh3N
O4ZznVqy6VGFtveEOIWD39VkyO0EG+PJSzbBftRTx0En9qi6v75/ezmLY8qfmaRhRKerhw016ksa
n2+UyI9uVnBU7YWl+Wpt4cwPIqRDYgcIUyk1eqfzovSSLQOEheSOVU1obntGNvXk/i6QhfFFQ/+G
8IJTdZmX7lABl4oQ65TxMjdCuDbZiIXiusp3bhOSDqmGHDFAxE22FECUcp7K14uy/H5RHrRj+0hb
FSc45g2sUQnv3pElKnbt9H6mRns71USrOOZvBMZ//13HZewQtVd3F4s8Fj3/fPp8W4zhcxK7eT8g
WSJdN3oAtHe3jo0Lwdhri4IH5Fhw/bPN7Q+0uZy1VIw3bx7NuzewtM8Dxmwg2kSUBDQ3ZWG2/hqv
zF/+cu59rpSWvlRkZlSzVD//Mye00mt5Utakh4mgZa8YZnHpLbaeCzsFVBoekUS+8eGLjrYMEGNd
XQs8LsxkiwV6Ph0kGxwkrvLTzdtnDjQreUT+vthLWo4efoz378vrEEKMCHc18c9oE+tfNmK5BYYy
vbi6SfEYPKtrwtImjp4jYt92DFtdhojl9GLTh+aBYsn+EqCFqToPZEFuaXNdFAvHqdzqhNJPzgt8
MGB5JdfmkLtktLLeB9uIZX+pDL9oW8GpPp3ff3f2cJxWNZJ7XLgixWr9uWnk1wvcQh2h9oC3p1G0
joBTWFB607gM5HgrEypu+1C6Rb7Z9+NcdRPBSAnaKIduKNM8y3dYV9EODnRyikNKwZvaLElOziP+
IfiKcYGaSRc3BFIj5x9IEkBOkckoyB9IRi+ZVO1s+agO6JdGDbjx5uMZ3/QzvdO8V87vKAIEa2IM
Nft6JrzmSI8GierGNqBH6ju5svWnZkUkuY+fZrtKOgU/m1lZxRVt2XFjt75DqgAP/NaJz5o7dCb6
emTpj+TTmc5Zr/57n1fBU0DI7xEo4kB3QOzklu31oLOi1SsWBjLWVrYMmybVUJoWzeobR8n+Pe3y
mNAYKNNSWeSdY+AJI9oDAIVKcKA7R/Pc3827WWjJpD2Dnz0jmDsiueAaEI7hCs756rhoSg1cX/Vh
VfnqUr1jU9ygpIE5liGUA/Nm+S9bErZlw7kLLjtizXg4ZBHUOiqAImVn8rUBXJ4G3F0KB4Uhvhx9
wE2rrpDPOpGt5OPP5EieVoI8YX1BLd6n/KPsmri6JL2/xozoQJy7p1KS96C2T7xJYljeBKgvctW7
/X5X0Ab5yaBkkl/WtUmQZKpf/WAHPS9lTGRCvtOIwATLJEqS0iEaACX+QqUlhoUhjpKF9BIkHkdf
Octkm/rFC6MfzBelxa1/q8EyNNIdEGVG3Yyabd9lwasCkuEkq1yRa+vSRXQyWu7zFtIMUzpFL/u8
0KyQey+WdhEaeFV0diyu8cC5isM+jWCuvkJ4yMIHhgSXzz+PjNf07FynLbeRKlJ7ewDipU/FGkMb
/iEXQQ0Dcg+kSyLBU2zXlqlYQI5LnNJO4OnaE8Rn8i5bzry5xAl7Ss2blOVksuLEUFV+pHyhVv+1
Y586em5cBv+WB8ijdoMZX3R3wC5bP2AIMEGuG4ggE8qpN6zs2OkMTZ+RpyT3mcia8GQbWqULgO+m
oyP47hJibpFFXPC3U2dnA7PQKRPOo3Q8oOvM2p/f1NpwTbvjsN6pVkv+2X1bResqAEjSQM9SyCr1
mvKsmSGyR1PRkM1rYwDccGjGoXoY+8ZKsF2Y/D/CJw/Vm0/qCpN/pUHX5LeiMSTwYPQA3kj4eQD3
plPyBodBxPMpelC13XNcGFDDhd1Dd3a0fjTCEiE49jX78IxsoJZiwy+6xOdDwIqTrzgOKn44Oe31
ftQM88IR9P2eWOFb0NOgNKF8Av9wwy0HWjR8DG4BTwjj7ycVuO0/jg/2uO4ZFw9Jdcul7jiMji85
XlivbCIdqWX6lomcY2qmB+RGWr0zOG4u6YvQLfY81hpCs3DYuteJERTgxohxjTTUR+7s7AAFjsMl
tv2LTJXISYatC6gkANL1oOpXxuIYVpI1gaHhDk2qI8mauQRkqc2jNjQWhiTGxHVATfIkWPmU67Mr
rx09taV+OshQT8i9G8ILXN0C8yseu7aEQcYdf/BHAWHFljw1FcU/rip21Qt/oC7NUXDzVTbnDekF
E6NL7zEIUYNdJ2/QWx/TF/QBxv5+i2v3fs83dBw8WjawWlUUZTvWkBnzuAFCBuB1xceCy3lLC3cu
JeqcYsAcWJSEBIxPnZYZOWa+274YADVvFOkYdjbJrUYMtLeSXZRkQZXkTvC57tdiXuCaF1k5tfzp
134ZL/PdzxQg2BhPc8rgdIOQJ+LmIs5IArj3PkEBhBu4XBzF2i8vzUXt95o1BFfjJtyKgS6VH+we
S5DOk1PEeZrCqcKJAkWuIxnPlmJW6Ofy+V8ZBIeS7fKXbL709+BhFCILbQwADsLr90yyi8V601rA
do+GF/woMCxeCX49ZgW8CqwshRh3bLB88ur2ChRMQAPgF3b2TrUqHU2V9WRM1gfS0RFVLxIcQRr9
6C2j8TUI1tsp0/9RBq154ppnAMrtLbcz0nKp7KA3y0ZlflKenqp2bZ822LGqOfbyYOhW3Rg6nkJw
lf3rCk1Hx7GD88bDhw6CiH5UvTXk9jxyo40oJszf6fzqHwRsdcWuX1W3vAjW0GHw2Ly5lh/Afcqf
SUXomC97Hahrs6bcP09DjVBvunYNdV81g8SrlC4Kznh9LtVjz0NGmZI1jO8ikum5AH18XSsF9idU
iZ1cMHGwrbReKda7VPIJ106kq5RXzz3soyG9tIAAsVcKZQn+mj93BJ0+cg9EsOIPAJiF7NoDf7dG
orRiwFwnjL9CXphFsQPD6ISWA69zBJWdQEF4DBsMFogvoM1Rlchg1i2awlJ8+uNiPQBmO5kuaBkO
BU/7VzVmyPyU7RHN6jf2QlELNcq7PIAnfxQAVKoDfs+viyio/M+OItCwKakPm1eY4gZGZH/LFQ/V
izEweeBcjS764ZvwfS9NUSF9lk2YNXMzYP7oXCB6MOJd0xdG9iMK3qDTZqMuM9622YBNR6qkxwqq
n/VlnUNe8/VTHfbg7Ie6L1AtMAUCFtQLwPjSFpoV6yXeniAd816FYMMSGqMEfQ0q1cHBtg8xwIGb
cEZnIdV/oucx5PEIC5mH3DKtKu3KxYVnJYu8mf9SOm9f6M7vP91nh0+1uAeJlNJ4VD+3XS6uUvns
vCLp0Wcl/Qf5R441z6T1CLCBPpVjCXAvxv+ijc4lYLXejf0I4COYmx4WlTGaGP21EblULPHpqV5G
wWyo0sBs5HGZEQ4fxwqaEMrk8U+lmrp6NnMZmRPPVWPsIbYeRoVmot4IdaLSTIhKp9B1notKB5/w
Or9oU4nD8RTamIbc0in/bMNjyLmwfS2SUYm2jqA8TgZdlaHKY7EsrAxl+0xSPVjf9m/mpvKj9BF9
a7nmHV63f1h76A4KQv445g4XUOI3/4Qj4MZ73GMwatirL/iHFI3yvZGBnmOwj8YqCyX1MSnxKUzn
CU1EYHmu6WqKHl9VbXDD/dhYQXpQDQdnBoS5s9gpsCP1IZAKNgJ6nMwJs2MEQ0XKIGD/Y2qKiRbF
JX7xLhiZquGfvFmi4nSTWj6Av4vfJY1SDsy+cduyA1yhF6uPGhP3mXj0MbYucpRwtzSzT9powMYF
Xdmk3T/vhKc4WxxlMdHFITpWwlY3PZultpMQdefnszMutCBTdEjDIUGVQabnmgdjcvvb+c83JN27
QTOnDUu/Mnb6JLPk1/iabOu0p/Lw5U+dhkmYKm2DOcpG9OgDntAWdVXcVgJkvbQu14AreWnEy0ms
gcWK8jt+Qb45VGOZvfO6yAIin18TAC/ICeUgWmd7Goza3JB8tVkiHdReoik2g3W/cJ/vaVR6p69r
XCHeaqBcbsQJye81Gu0ELqVcTTZHFrv6Vlzsl5QoouSfrwY7VLzYaHTpe97bLGMj0RVM5ASP1/r8
hzDmmAB0ZPTihLsCFd9cNuOvibD5nEaHiW2PoAFoL4+98FP6MX2Gq5lWdi6yeIya/+KNgTh04R01
M/Pv/l0bIehVHp/NBfNho65vHRIk+0pnGIE2notIpvgLGtn/jvWelIv+yB8Js0OZeBufmbOror3w
xK+Fh6DYdv/Tc9ZKDWDuTg6uxYdTQDKC/mKl5P41vB/UKfhXeRrbuFQdB/J5Zn2VkOIi9LH96oRc
S7Z+4CiVeLUxX9fXA4X09FPnJxLIqNKv51ZUNF1BY01dC97rHqGSZlsd2DzjIKddw0PP4nV5H0t1
DKXEJRXNInly75Ej6NnD0fNB8NeXxJw6OUpPhMnzxUCLQM8Xsg9BUBy24mGet1ENcr3ud6cmg+F9
V9b64in2YytXPveQ7ErdbMRH9xFSd/SLIqfZc2xL+4XKjIRuil/BnL3zdHQqHVLb/eg/z8L98eqE
lFHSEX9A/IJdtYSH6hWmV3op1uWoMFBaFx+IXpguxoRvBvMUf3RcNMqPyLObNIwbnIDr9K9kSg/z
P389QhOzOPaNSarlvZNUjHEF3G80c509jEVfJ/Tv9QsUDot31DNh+9BfOlmnQk9P+hydv8+zSR3t
gtdR5TggdxWb756skscRpDrkL3INmPZNp5sB06yOMYnVttb7w0bBfVq6mcPqOps1USabmKwyWeJl
6tq+JbH6l73mTjE4Oa2EUx+h5xeytp9RoC7TkVxm3slXeqHo8d/GQ99iXSOYkTwzKOZM8CkhOBuH
saHG4pYqptFUjN0aQZ98WZuy3FvuL/uzlpGFlT3mpQ81kBfc313Vf7q6j+RVGd+f7fQKb46sVvCR
GYwto94fb40d2o8HckpLpBtdHFGTtImI7L7Wmx4nroaJJdyOg5QYexzx0a4bM/OSCyJiA1L54p2+
kHVHdLId5g8CPqkoWJ6RCshyPhfb7vjlV6dKQ9PY24v0MLuZuCBF3yDbJ+zHebI+Q05febNu0YNz
oo0lY1fVQCdLQcVTsZPqvqWNq7+LxHVuHiM1J2w5FZx7lb+GdGcu+NJ/9bkZIF+soan3IJYMbACH
1MZfKVjfidVKm59C15r0dFHHvxJmAcz8CU96y89CogLIzj/siETsHiFUhbfGeKN0CG68e8Miy8lL
4qCsWfnxC8UFlZo4PlWSjlQfWe8i5/yYL3DCAFpQb6h2JEqk6IPjGJ2kQjFTGbHRgMmh3zrdqAIu
ylLnv5MLW4fsYzMKX3ZPfckNaIGReeYnW7xyTgv/XvVG5Mqu3CElbuAsLX6SHezKVvJwdXzfWh/N
3KSbPhoL8z2Fx+J91hUHhWPueFbotz/nKC+M6DxHwx/4awYvjJza8TCfsJCJkEDAj5347cGnYfl6
Iw6HMk2pa/NLSguU7YLWTweVcH/DKdtlF2s7nx2Vr9XTPGjZYN4wNi0djPiE6cE9ZmFpYFSTt/j/
u72TNvfOVhrArgKFRBiSOz1mblMitLfpb+9oduV3gYoOhY71lB6qfS+INJj70o5Jb/Qs6ndYgFXc
F5YeQwfJ/xuuFcwsWz0YKoLHdP2Yw1IM6F+tP1WcU1G6CSc04z8+zkqDc2YLwWVfX9PMffOjhyMp
7EzxL2O+bFnxJu9ec7XfIz+74n04KaBqiOq7kvmrBXIIk2pdyvwKSEwCWew7BUrtNGnNZOHgnpOs
VxvAzl3K/wJijnJdI5vHrHgKuuK4dFVLdgc0TvPHXUJ2c5Vx9LyiEtVq8FvIDXM10UWKcGWcKDfg
lSkzA3r6W83cg8cM/a0E79WW1fTCEv0+VxFBx2Ix22yarx22Nx+6sEljLlnt7XgFlIoWvsHFuCbz
mV22UeEESOYjEbc+jU1HdlqkcscfGebqwd0/ZgXXj6sxBOQF6jBPrivGXJDQDezxY81z5JsfxJBp
/DDpzReqlFd0VVyOxX6mJvz5lCTWR1+J9BZeijPKyLW2rgfiSz3JMn4WokPQ1A+MFi5sGlizttSX
QztCTQlnLQ8OMX2JBtk2dt0UJyteVPdCxoq5F//2+wikPfj6u9Phab0R1ZRcRxDMfkvJopt146eL
2tgKMqez+1hLvlrUg7iOGOWLoEUS+ho4cBLMjAg+LKnJwI3h2jmBROauAihldU73y8j0tE7tzuY0
E43rMkefOUbXgKRvC/tAxHiD1pnBMB8e6nGlnhbQRepGVhgHFXrgHPRW0LCVcFcxgkqp2aHQcD6N
gGj/FKEW286qLw7p4ZvlbH3/dvYLKoHXa4QLZDg1eMN99/elt9w72MDxExDKBR9UT6xWb0AoaDbX
G+w3vTZjTUpFBrnODIKSmUSN266bbgq5G7MXoM3RFNK1nAg8iRE1bKp5FCoLOGbZ3gfww4Yl/+Mk
KoMgi4NtFlaDPsPKC11M0nglq9ygT/Y62R0NulOzOI77ZbY8HPSO3MRLqlP7vqERJweUvEyX7aEW
Oy2QYE63tUjSZBnTAuv2eai737jighUEiEwf9X8xs/RAEHNLOeCZppwr2H64FNREeeXgb3/M+VBN
94RmYHUHnfySXWqSaibjs6MJlZIuLS7TbYz8M9meM1OBYkIZ97zs+m+N7ZYdOaKAiP6F8P73YAFf
gqCZRnsDBZHAv+P7cWyzaUGItgvpfK0osYgkpB6gpspfKXfGOKSSECr91fzsExVlJrCn6Mf/Asn8
BpGaEHMrw/LvjGhlrINnuVfkYZLp2bCvVHsKSrCD8xilOZxttZ+1e/X82xErv+l0cO6qYtFHo34d
8VP+GCRplR/nAHNLuDWh2UUlcwsjf34SFqG6i0AmPKYw00IP/1MPAwnqEyWtLRYjGa4BxG4Qy+Yu
NcLtUoZyrmwFrJ4zauYL/34+XpyxznEmtLMR4Q0FzC69aBQh1Z0ct9CmLFxPLaZojywrcwG6brEJ
lKpaML/hw+OEBI3KVffeUnCn6Awhs0PGnsMxRo3I8nMn9zfEREQSaM99rLn0ssWaAI1y8Buwud4N
QtknASmnbYVPJC6Es4IRLCu/hi3WAVhnvz0WRDbKoes71wIMJ8TCnhh0SHuLHsDaPgOxa1DIs9Si
AGICMf00ylwJ8Y2PoGdHvJ+5zqtCUswxn2zf4DvTb8wxYUY0KBue7wVEWK5icSQXva+PAO860qE1
ej4LQpuMNGU6qY7YocvagQ6zwMh33eaorNydOVMj3e4joJo/HiNRvUsc7C7shTUa5xDY8nKAiNVH
jz3Xe75k6s5AsmQPp7twH0CODcA19/8h4X1FNenYbELTxTx9jmZQTHUuaAIM7H7/cjrs6ZuTFISs
++oH6INKx4PRrr1SJYS8og7nsSnAOczsSBS4n+VvXREclkO855JwBmg4NfjioXoW17XdLuomFFpx
EkIvjXJKZll7woPT9WxPL/r+rgHGRqh/8vXHmE5AscLT0fpTPN5ZTvTXP7kIPqnaZRreRInjJ+7w
deup0MqUIXAVXR0Za6WmZF5wtVLzZ4B91affKT5z2C0+wo8P6T2+VHu6W/vP99kbEK5PWk9GqGkn
rZpl5ljjzRKTfj/ij887v6hfQHWUedGimxVELUDcTlqK11kiqgrorVWWF8XLHyG8o6ZwvS/+0PHl
ihlpKpSCgg9pgSzQdY3ThuexD+tUdyiPG1fVoZOUBAaQyKtRV7aKCO91XiUU175Yl4ZqB3zNZFVA
AzaXW6Zd5B0WbMfRGgkdm3F5QH3uyvkXZStaa/NeQsjAeOM8eKsZy7bKY8FsU9fFO0Rf3FF4DUq5
W2ttsdME8Z2AJ1+zBtUd0vIr9ONDXD+vS4AYbD6iPHK2KYNwHKFd82so9bzzLqq0mGeuL35mD1mD
4SdKuRPqboJMsv83/3G4FiR8ah0Wl07ZF5cpytkz7aoOjIKGkDuP3m4VK6ikq9EFy093U4YQFykq
OR5z/nj2ah+Dho6Vy5uqyQdczZW/wb7mWSB+r9VNIdyN332Ol7cDE9XG49tU1ZY+tMLlzWQ5Ojgl
I6RkbaI2aXjn1OI/WajB9oJDqBhozxGYZXhUO+wKxjOGrDPpXEoKlNGET1JQNbL/b3ZZ6omkwpOk
L6672bZEwgMX4C0bUe2vFNAIEPO+kmyWh2iydPBgbBrQpodKsC8XErF0EhZg9Luocfj0ECFnIwL4
5/9cmpiTnpp8Tq2t+h++DlgZDZ9Sbxfp7eGB7BywiNCJF2/d9rZEIuSkrpc4dGXJxvxfINqtkQ4+
GvcHlNgKeKdlHCUWQbAt+ku8JpPWIDSqqFNmLjMumagiMzBJVknZb7LbG3r77Bn627k/1zXwZwc1
eJOmf6RCtDZQ116Ue3z05ghe3b+wRIG841Zk9EpyFVgmMStIZ2ygeyfN0ohUR+Dsncp3n/Lj4jF7
tucRJUaIwG5A3Emv6PtCtpMDt2v5BLvET8DXeQISDb8jeLD2SQCSjNNwqHKMR9atFR0g1N/c3Gsn
0n80tLDZW+WcwtacdLhHSMEh85CPppH0TVkLxtx0rFPLYkicTbDXzMGV+5/DhnOirv+r45Kmwlt5
2+9C6tF41XMz2YeRRaAsfdvFYZz3mtZFiXOYw6m9iOTHwYrvcKICoH5Is9lo6iXaIbR3HaHlBcVr
UqQBAXDmkOEHRadbWnAFfaoYW72PLnGNvGQ5tuADRAT53qSilPCFYYJpxWYjM8gq3/tIY9jGrds+
9wSVoMEGjP+AmwbihDbjctyy2SbvlOJsnlcV2EPSVaDWGMGlqIrMaodj5j787TpXZ+si8nWtpoZx
q8c+/xWdNMwNzUTUWfaplKLIL4XNvX/jqAtSAAi20ypg4d6dJ+I5qTFdFdASYRJn3QEUdw032MBv
0rxAhgz9exO1FpVoUxpHVP+jkjQ3LLD82UM5/NT5VYhBGCiBOWXEWulo+GoECcXPJ9wnzwYdq+3I
2OdUldIz/UoYChsZ1DxjpZxD8oqHx1f6BMG0iShSHfwJceM3S8xvqbVrWXAK88YnWRbYgheuqigk
xnZTrI6a0FbeNkoKK2eODApFnKt9An9Yl+LqTCcNSRVYcpr0i+QU2JWns2EwNjZxEp9cThDjWGpf
bS61xUL95anwGy7ZFKYzLf/nFHM983t1pwsaIk8dYI1+ZmV5oaxS5J4t3zjtL+BfC5Z8Drkx0Mo2
l788CyJmTgOA34/zUIF3zpk29FdX/ihikvImKU7i90NuVr4m+GWlFx5xezMTHqJVzgSHz0muiG+T
Tt/U0TprhXjmgy4BuyHwUV/G02S/RVL3O1DBuNPT03F5ff3AqDpVThHNc8g9PGo8u1KttwTP4UMT
QPHi4st7SOPkPrfE+p0ZcFNHv80KbWdru7PAeTS5gAZV24jjDEFRaAldmSDWP/KOm4lQZwOE94yr
lD31cnYerERybfxFEed8HMzmvo4pCweY6/JnS0IInwaAtXs80qmEkV/X67za5pjGPz1cDFMr8eO2
6jlScGEYZGJJAtVI6Jtzpnb+fw3xSrcV/E93xOSzadmW/XJC+VuI+kU//SjeOLC1Wv2ajGIeoSBF
0kIRRKgwhSuPFLznrf2AgLU+fAa2Y3qV3PLenvX5GjgAMLRzbYElx9lfDiBZCFSqw7K/k/IkkrJ/
Gozq4lBEJCelYlN8xg0vzt8HmUVyVS7WA+QlVzczxYVXnOy+hLsSkYeJH6NDQRTYq6Meck+QvG+q
55q8YtMoBYdSV4RKsj1K3TWhhKQa8K76x8hqwa+e442WsC9YAle0NkvG7vaCwu7J0tLgNWZG6ECv
97+wPh+4MZsyvHEa3i5sWQ5flJuhADseyLJ5kJbVeCSzXGGun3Wp9deTl1jiWPkhhJr6K1DOayd3
qARiK18qDTWZOFPq69sSOaGUmY9BM+hsUXI+/AX0wUUmkQdSKYcWY3GRVQ1DU49Og2iaSyGifk44
Ex1kfLnibz3Iemcyq9zWJxcLqW5NCPMMxiN57ylC/+kUSfdGcYHwk+SJauIrSvIOcOKb5GGQFxr6
EiXDHiAXaGd6m4w0E/3X4FgINg6VQ/pbpvotTyPTL8Rxzl1wfzSajrs5XC96JP+ES+qA6TViePXH
/MOKqLgS8mUnYQ81EgG2eLjiVpt0qvW/7hKg/2MRW28FDozXroYgxCMt3OeSSGjkI6ZFtWRHVC+P
5ROeFAoELlixi6p6FawxKRA0Ajj5q1ub4M1V9p9ONEGF7ymYJj2MfEDetGcDDFb8m+VK1kdf0Ix/
LsNCGuEzXy8CA7IYdbotdG6K/6WjwEO2xhqCzw+VaIZ5utcZZdb64tWch357Wzz0mNGDf1k81agw
vgeWnfWbIsUh/jJ7FxJTxf2Vi35Mw3QC77KZQEpZ53radPM3Q8lNbJ5UGKuxf8hIFBcotkpVQCPq
22zlnt7tjtsDBamKYP6GpCKFBgMpaqHBtlqO/CWmoN4XBjQYHriUgZOIf7gn8bh51g5nBdlVX0So
8efEnbvJVitoj7Q7Txj8ArRhJ9ZvvmjWB2rDIKc23aN3Bhe08EMB0rQOUqKa8YEgJO0d8vr3zfWm
3RJc27dVcgndh+rfYl73VDsPEBom1q+x+h7s69aDbbakgBRK5udKrs1Jqz/A7Nwpecl+uY8DQKhU
FOqJJ1X74NLZFXBSiFnn8YOuD+aMbJrQ5/95O7vzLhALPbi+kwzbZQloked7nhhErLwD1Lw3sQGm
jF8eDD+1nboUV3PjFE8cjG7gcpJR8QF2GSH3St7XPPP7HiKy+OEgKmyvlqVj4Ng92G7C2fp4+9Iw
SvTOIPqia2vADnsg26HUP+7ZoyEffae6+mMAVhNHe7/uC6QMV7VTe36UX0eFTwc1hP1WqPu0DOa1
wpiGPPqnkockot2QmI0bcVyXr4d4evSZ/Wk/qQojUCqyWvEqcjAItpIaOikQd3EtRrkRuQRTd/ct
L8uLYiFC1stCA8K56bfCvAWiLEPfVp3p5FfqX2ENlaouo+HqOPNaUcKslsv5DN140t9bOzIxcxHs
2ObmHJhUKwJRBeRp7CUbmiB6q+9ed805nsWK1E5tpLe4LJ3+RtLbZrrq1Qhq4ykzTV3iylKM3z+r
eo9/l7w9jPm6C5yVLK5XrKRQ62hMgnle3IZJqbQT0vShYlumzAkLSB038W7EbqJ/4uvGfQOJsKH4
zjsGUUiwhi/FzJCYTrovYINHzOEItQzTE6pt5IwNaxUcD66jDiUc9KMEv9/8+SuT9z9/5fG6wd6r
InZSwUgwD84+Vw/ZzMduZA5dBY2a32Y76LNRyo54TN1iQ1z4eRwmSkVQ+Bv8owVNV3w/O9td8o4z
fs7Ifon6fUzpByEFeP5uXv9Og86Qs51hrTbIAoIru6LcC6CYqyXekEFblgkxbNC53nb2gETBJlkS
7FFmWRCJJUxU/J7nZ3zbdVAFdCfF6YMntQkyUrAH7t67IIePNez33DktwQZDN08Tn2sp68Ap2Na7
fVqrI4j2qVez42LNgy+S16L7CV4u2yJcih9+Zew05jVe3YZd41KVhkYpkmml/Dbd7sEm4b44f5xs
YR/N9DwGY3FgXobaR2j5MubSto2fqA0/m008u94G5eQjjG7cZXGbJyRhjYyS594fVsdrOU0d/YCi
0Mm7uvkBraTtM7qGAU2nmWJ2QkvApKAfBwfQlDDqWZ+eGx7UhUsMzxLOnKIWOTeDtPl4RrG2UwpI
UDKC7ITjBTU5fn95Po93LU6NwAjsNAHbmJo7sdm6z9dtS+PEvrghefD409sZXFF2hov3kVYmdDvj
NTIy9DXiMIVyWERsUKfjFsbhPuOtEkMXB8wtN4qjQu6Kf9V8zQCCSoaSHEX7Blhg1UuIZ0ry9gO0
uRISaGwOyLduzLc1U28mVijRfCkBsLRRrJAJPyaSSywfViH3soncAMTgXb4teaprQ2+7i8mVpvXU
n9/K1mEcawsT2Qzs2z15iHTjSlThZaKSA9j6KGlCnImEfmZH230Put3R0U22HkpUr5lEWmUPfEeS
skpdtvh58kdWtNfpYgh2VECxS4q6AqBZJstHQt0UYK3eAAClqT/R4/w4kco1pnpmEuwRtZn4nUi6
FCsVzy+7Jyt5GEfc1QF3sKeglLdKLE+ROpPQKxdFj41dLCmcelGgrvRfj0tYbpqmzLWxOGcEJlUo
7U7fDPtOwtJbJjXIqxn+S5P7WQ9UypxgBJCivsgTLthkuiqAT8lwVGB1i8ZKLCFzznWeaaIGyWSX
WDH8RhDzsmQPU9PFY/UTT9FOgCsntW5X1uyr44TrRPj51bX/h5XV4aTkvSHEZiGpcgiqDLCcQog1
7f6hIravnHSJzYs79F8o4SGZsXPSjJA0buOWa43u/382000VTt3TFBNRcfBK1QGNGGz921LGKDRP
98aXJ9AnQP3kXWI9Ey0ETlwWIcOrb2/I/ZgIYp3vrsCHlKl7kqatZVPMLKqbthE8miHg4tMcTw8a
crZfpUo60+792925Oj/qQLevLwOz2u/LPOsUUmbpd57QScQEVpJikkaU9CbElkvv8WypiVlUmd+1
2SICH2/iDCpnJ7PihG7j2Tx9XoRaxRoZU6sASsH0UMdJIp5SwIxsVFn1xG7+lWLgHdvNxO2FGUAU
5p//KrXs2Le8DEeQ1mUQBg1FJjaKvsiP6cT6K65mr1ZYImmzqhUsG1KIhlS5gFWwK11skioqXNEb
ddSELNvdqggjDh4mVryAMp7RsX0CwlJONUKVYowzEQ5/mcOwm5yIF5iIpAnxrpfWbediMfbmJKd5
79fOmW0Lm7soOfh4fHIsY/Yle7LPcs2lHq7vvVsq5gTmqOPSDiiZ3bYJZChVZtDrFf9umzT5inWt
TiginTN/iVQV4qpbPOEyMAkZSG8W31MfPzZDXU2jK2WmErAhp1c+nwBjRmiXc/JiB2meRh30QkHE
UcXm2zz8IKphpjXCCADAHLr7uW/nr73VFVXFIKrPGJdxhJkyA1ldlf0PQoyHjHrcidGzL0ChoQ94
f9mGLI8xbDy06NZNIfkjBB4k2fYwhok2N8UMrl71EwzSbXlSjfFA5E2UrbJ9V8LETu6aebwgN3XT
pT1t0/BeZWoCENdp8wC61xrhh8OfUBn0rcoSJSPrCqFfLIwPPXY1dqyYPq8r1Vnd44bRof4JBOFG
QvSbD+VcfgRKX7GFSb9D+AWQo65hdcG7DwP9kBTnN+AJOXtpkpo2HyulcfJRohlXd6iLvo4Svk5e
57v+7RAW7eMQzb+RUEH8dFZ6nbVrP0sJ11kDI5HL+Uuwq9Cy2KeCQ8u5vr45Ufbm+ln/W5xI2nCI
eCFuLlIX5/9mrTKmTOhd/Q7hFYvU1SfJTC28LMMt5Rpjmgg7AtMDyj3gZ/4+e8lLSC4H7s3yPfwi
7W/ekSVovd9bmjeDfWxRSuqU/HnBiAUFR15wsEaCfL0ZrdlPebCIjRLDNJmw2J9teNLOfhK3fuo3
wDfA5rRLLzpA4RC/UnZEJJmLAIOUyr3lYa/Wod5x4l3ywdhj1YkZFpJyUmPyOCWd/CyGUa1kWyTY
SPE9f9g8PtDR207AA5Dw4wUJcgLl6e5pimBGuPzlsIAUJGNk9gNGtQCMURVbd4QDxnZg3fQQoHZ/
k59hxKNWi9VFVxygOdA6atTMrrcM5ucpjsaq4uLq/jNgrrAmSDkhISRGOnAuP4G/rQdBiz1EnvrH
ijRCFVjodJjGu7U4C/ujnKg+nR7a0S2o+zWq76/n7nXn0XjEiL4eLiYDI0gRHLn4nkM1WGOzaMXA
WZCHep/Yf3rn7aLSpxmmBGXqupJO8EgHiyVsQIwSwG4vce6z+c324vTyOUlley3RAhlfvyr7+WPJ
on2suuQTNUS5J7CVcShJYSwBZ1VxMU9FVmhmFipLJwhy3OywQ+vcZOy474X1s2Hv3//pYyaUrRWu
BYLd27mqNfVG1ZBCFwBhznZbyVJ9rmmPVCoTkuvfRQzeV4MdOgCIxb0/1EO4qext+cC6a6rx1ZYk
XEE02Aibe5TW8FKLGv3LBKDeZvT7uYODBC1HYPSejAzemgHMM3dGvxw/mEsCY49wypbEwbG1Mgy0
it/gdlajDfHhrTzsc9sSQi56xNUPe784xOrl5PUNC7mTc17Pvy63UG9FnmbLRzpMoMV/ZAKdONnA
Y2a8KVxcOu1dwnM1BwGsciK5LvIYUAJ04CKEn0X0ji1vOa0ED2A7R1NMLBQzM7Gev7DD8L3pUNsQ
bH6FzSYNVrg1LHyM06u567VPDLt1uzgAGELnhmGrHR6rmoIpYNMYH84cepOuCkXnCvbw/ZdtmpkZ
mm6gnU4Amt+olRNyrNuoX5HMA8Yk+gBgq9lM/kAhehIMCGFLM0glhjohvAyPskeKCAS7rXQgpYhZ
sYyU+L1s8hTUXfsymzdqHoiKD6+GRW8SZ8eh6/P7pyqP038EQbuGJD5EigxeLE9UYWilzZ8Zx7uC
4oiNXPTKGyx4mt8BcpIO1ifSFmU5aUnTD7YKi7ECbjcIbOW9TdFNF9OJsiVd2dXZQUDwRWjKS5Ng
q6waTOuKEE4aUgIjagPlypcX4+PoJaaIyQvKnASJFeO/px9TSa49DyYYAwARbAmVbVsV5BhX6A9E
NkY11tS3ojwNIrcKQxAEKc/CQFy+Ug/bReUe9nemm2DWMhS/t+sh5mWQPfD2XaiC27oCIGlNRk9w
k/7FTabvrVaNiP1vl9PeQENnYzd+pjPhFvC0rRB2YQzCpsBej1tWcOlAI8qjo/QGmpkLUPh50Zbw
lQUHEZmN6keCdMym1HDj5o9i7zTUiR29q3PH2EBEpbX+BNMefRwtW0pzLLuwG+MmbkHerFrNDBTY
YpOoQq1eg3Kjxfp1zNzb8vsODeXjsb/axkfPE08DPlMLddJ1V1tbvCLM0X5KuVQFF3y3J7psl924
o8Y5NVKe2nHuhbOJCIb7zc4R3TMbEI/D2FksJ5CEY2OZ40IRgxnLRDgpOYlMjtv/DV2vX7gvCYNJ
cGpgWzigBibcqYcmtxTQnER8kEBmi/GvYRxLxRdIhc85+NXlJ8MY0aNFHzTqdmxZDT2oXoHi9FmU
1KnHhdp4NrR4ZVhe0EwTCkMr6tHXBND2PqGAftGXbLU+CVu/9+rqnjoiYcRzZjRpTsjrMXl9uXsz
yDtk0eM3YSVPALGUUQeKOFbciyaoChUOxGUXfEICOvT/lT4UjkMXgTz8sZv3f0b0PE8MPSY1/QX0
ATYcVyfIPEjOZk0ii4Ql/cPXIEF1Ma7CQnC/1SUqsXhnO9V4UN+U1eGRPaqwutyaeOoNrLJAWJoT
Hz/jJyoDeJ1wNZmUIU4t/7cIgCllP9bROWqOQUQNUAZXUTi5wy9vsAbprZg2O2Au6mNTI+7dCGfP
tii9v+VdmF/OKEMMeZyJXLX79Sl4oZFW2WlPVz6t4yh3K26M+rNoGmWcvXBdJSVyqHYnYU6VhFQb
9Zi4uqqf33Hq1Ct0QUtUd4ut2yCx+p0cwD/gkA34IIe9XRpybOzsMBQ1bWqt2DsjpOyio900wEv8
UALxcYM3zfxXBQneVWIaDW588OLoaIkj5ytco01lc4a3ED6jqpZGGWNIYNAWAu9W7DInO2daWB7c
6S74cohXA3mTeWTo/o0L1jHR8mAd5MbG1feN069Prd3UmkWH6PLdEM3jruQQPgolp2jYeQ2HgrAn
9J28GhhgYzXWF5Jp49LFfiVg4nLzTt+fK54dxPtOp5muKCzdDExNQBzwmsrt0eKtljffo7eqmL3+
HY+JzXpOjUTF6QA1HvEGcjjDBRaiEZZx8EqYeBFXLmMBom0Pq1HBifq7PDQLFEFQPgK+m8jGRRMa
dmdV8zNsymQAEeAmx2FSK4u6AADZHeqYve19Vj4mKS2WqLoj+IMd9dq+U+/ftAYdKdC1jqUpDgfy
4XCHyIBuOI3HpY379OjHx1QlJ4SNrK6qe5pOzlmNGhYE3U4gtnBhT21xFI5wQ3f4cEw2wWjp2C15
zt//nBCUFLJD1IsrtQw7yPw2XbmcVJNZ2nVAY6V237kiRzCLsWmAmQUGfFHdQoSvcnJspokvuPR5
kVUXCsexpAqWik6qotl3JSTPqieIYv/zmI06Igf0y+TSsfcQmTK/7vwGUudh7U8kqLNKY+K/nYCt
UWINFgyzNK60ygMReVgCq6/zkxfXaCsCzHebgV87nTOEjzTljUgKNNuoSM5vDyaCbCUQkROZxVIK
BrCYiYUoC2RC9vcGdlNNxcTt/ZKkj979JVHT2Djuyux+9aNWMeLeG3DdTs8j4AakUQQKildo2+HA
B2y7iaDOQgut82wAaVcosb7sK5e0iKlmu8xnhVLRbJ3f08sxdGScyiW5chnYYwI3nkfhktPoHEAT
FGZgocD96JdyAWPcVqd6bre61EuIEshnAS36rGw/UtX/PprihVb4xVzoK9Es5/1WBtDP8RyTlrZw
hkCmste3IWoNNxc95jD3l9sWLP1Xyb3B52htA1rbBuhI1r0m+Bd9aJeiu82GbiKvDE9lnKrB2bbp
xTfwzDILupn8a3WhaAVaCuUUveIsOGq6k/SZt1xH0yRfwywmTmLY3bTXRgY0+2WvlU6KDNhvMJQ7
Em+AkU/o6f9xNxBU/cD5U13yxdDON0eXDkJK15hY0OmenjbbTTt4kGJm8Q8a6f20p/33AOt0Kv6M
U9WnapVbdsuLN0y30iMYqaFvjkd/P8mxPTUSek4xyWJ7x9wEPoIlnApc/LPCXYZ3n36fZWOxq/bK
XGl0siT8PMVEoS6bgYyOudFKhD+THNXuwABQeValblcsFhGznJ+ECM3xno+QxdKP3E/cZYdQUyHN
t7Vc3P99emXUsqKM9WwRqOS1ruCd0KChbfl2QwXdn3UNVUnIBc6P3leqeAwYz7GkG3pjhjnbQ/9j
q453jfkXuPkLa21QdNZVuY05ZzWEKubGYdWYkFki1N1clph7v/Yppu7KR0/6go4ndxq2JWYRPeoA
EUqtniaWZzBXSp+tLruIYDre1GSTAlAELSCdq6d5mHJiDBwXMA5Y5yPmbCbW4lxx6CfuPWBCFNta
fUygHAR4DrW3zXohTw1/iT4mIz58MvzY5hJK5+oKf6HFdzMdQ9WOPJhw8CD5fjFfGaloZaAYlVVf
7dOulgcNbeVwGzKdif6HQT7n4mjusgABZjdVAAZuL/H+VBAe3B7k7SHnUvFMkaL6LyvBCOqPzFZJ
29U1/ILF/1cB7TAVvvcE9k9oRAMFhpiKRSyqVcZmzKDy0m7J4JJ98sM6ASvvN5FjKs475TdjD9Bg
A6Cxh8aMe5FMmLqqpBYRZjTzE7RxksS/Gy1qXAegRkWw/EVyKwyqY83PvfUeI6iffD+jMhvHETQ7
S0bRdv0svUYjj/8TkzorhOWj+c83x/d+f95TC8RvTHrZ552mdKVPMYTAzrQ6wh0b2j9uzpZFGLAh
3W0htYqSIeNrPdTGv3+7LTumsO0TCR5Zc8BbGqErqT7LM0I6JM/r+FkBeAhKSg5m3hBH7RJAC11s
f6K9d31uzAweAN/bv0VGlcb/1P4hEHsg/MQDCuJoFuSJX08CoMhjQCMmiu2uTRK1aBWX8VxQ/SeJ
OSPGB1Obm3pK7OO/+VKtXf3jyRN+at3fkyM03jYKR1QTbceasds4Iw1Bo7H2xz2IgBvgvzBJ7KQy
nliDjxe9p/dRJBtLHnJYB18XqUXR+u6IH/G1zFS9tIRY++qd/37dYTLQmyzCyQqStUC/clfBkmHR
yi5bJGS2DmeLxBX56dFo8oqSTUj/AdVsNYMndT2PjW5H6sS9042a81iE9gqTs3TU9S2pcKij5Fv2
IBCiU+MOe8ga4I3XTqM27eu4QB6o+x08vsaq1iZAMBOTmI70TxIKemoONOORWNkXPbkI/1/HP8tc
iFnjHVClZkFX46TnTke1JgbFabA9UcA2P/XsJbXtYnNTr2LZBUOgVVthk50tofmOd1RuH3nN91vi
o09N3W9/cir+eGrpQPxDKSOsGVbgbtx5+XEAAW21+ejfwetHF1J4B/urP2a9Q/1rXfJgM8z13msK
kUI40wdLP/o72JxrSLKn2xJBim1J619OIPphontIv48pDebhO3bCEedMgpfdMvOIok35Ho7Z153u
XxWvs4LVxLLJLXcGliPtBJojl7wEMt56QMhjUV/rvAj2huyxJmmKB79FYcYXO8ID6KGuGniXEdRy
AnucCDSkO7ynyPspPhiazSFN0sMzBEt9DEyEYRKDGZm74mnUJzZCRSQ6BLcLvuJhpja2ijBblyHt
Pc0WbKtHXwtasJjCC/4HdKhE4uoUWNCnl8/HT8LSkXqiSXSh64vVHTzGiqC18lqThff65SQ2eaDT
eIlU92MRwfH+ua5UaT171nG2yEneCpf0GfdnsFRhtai1RtzB7Osyoe408W5ecWW/CvYmRYwPK0rF
5M0aidaVHVQGEJoUChddz4OML658VlqsPHCmKHWb/Olao5AkhsVFt1SY+lW10x63r3trnI92jKLa
NMsBy7RQM9BVd/bDVJ1tYr+wIGQNtGVghPgjXMcoX5zi1CpAWx9j1VZwrYqH8lZLqQ6gKqqNbh60
HcHsCD+SEHEk4GcLqVmZFTQUqfkSTtnm5+TwAadJ1umk779ucHSR9P+Khqfml4voSZjo3QqDG+3f
Ehsgv9EHFLQ4pWJU9QC9e93Xz2qrQEZ+qCJ2F8QqueFrJesVOVEpHKC7Tc07eclbBSxpJ7QGT/La
DHml+kc0YuEM/yMzTuH9k/ovfahs8w8qe0l/DBnY4uhTg8usvW3JQ1sfeD24Vj9yolzG5ldDfnKv
67QFtS6e4SeV8vMwQhPZNOAXYr49XbfSkuqKh0IfOgtUZr7o2cprCjmEyEwAgE4Q/QCNitoWnGZX
YDQkoW4hfK52sv6I8G5M51uPgrn84OB1fYjQK4mUhivKgUMgGWTWcRra94TvUJnCzrs3bllm7Zxu
rfWD/EsBhj03vKt2Cqyu+G+V/+pceUbs7XFpPzBJDIH7vgaZxQdFxLNOp5ZpqI5pYu83sIrTx/rt
5FaHh7ZbInHUIrhSuDRzcWOVLBCgjqjgyCCSLCJ9VLilUmTFXqt+tR7P3SONpOT5jL01OS4rATcP
cXlTHSjfdTnFNctLkuzEmZlK3RbgGQgFDAPQrGctGPBltlTtHWXa44nVVrO0oaGhRLtapsC7h4Sq
HTAgRL/PboseaJWJVS7oNeZUjwY/dWeD8P2qDHVLu0RB8O5FlFEeuCLjwcjzWLvzvCoex4JjnS7Z
sfr4V8FfnRz/s4n3z1v2gd0uXnXZMeiHL+nvq4x5Fv8WkISoil9lg+T5o/88vmumXpgYdeOlJ9xM
wihQHhHwqBLtQfxPdaQIzzuSBoCm37/SPDWZJt/e1H/OyCzk0ygADnXzxWfOSPCqVMflBP232TCl
WyaJow6kW4vNLrqWtYeqocZhbZmd5TuVzE6oaKktbeTJClMs5fi/ulPZbDcqk9fSWRugdNAYwINQ
7Hc7DbvlEWGfbezJx6Op4V/OtuGX1DJzeqirlycpGwApa8tcMiSYs3xJkQc5ZFXmlzHrQICERuuf
p/dpOu/WozGj8P7y2YN2ZupqKFYJaKupF4EI3EMxlsmwWvF0c4LpNiK8Z43rw0s97NjaefjkIk/2
ZfGwOe0lLoqW09L9XNdJ/RqLD49tWRo+SkAXYT2gT6aovWK++w6doYxiGgOcUvjr7ei3yklPoUPI
ASVQD8ZE3yS6jkfNPI+DdLCk347OZFRlvZH4n0r4BwacaMpPP5zbDtzrQDN8WD3DDNSUxnOB/xPo
D9EQ4oyEk2HinyDl+a/vrhq+fCx+VyLpD/SlBL+P5XGNXa4ntntOvhyux6ZHTSDAAqeib4KZprhr
QbmgqAT6h0ElvQyln1tH4/gOsc2JwhyU2xQICiAFcBy8zLcKfWM0aL5CkPE9X3Rwnsij5t5TQYKe
azU+rniPA7A/3nRwxj/m0oG0UkXGjuWfjjejrZp7L/0WPC7k8ec2j67FthNAuc7ermei1TT9l5k/
AtzTA10BzcPQYSkW1jBjzUwg5oZeGXEejcMJkvQbH0NHg9pKgBcQ32jE1FeN9qEM9cyoKIIQJxec
FczNZVH4LvIVsCxNd4sq5MBsSgZ6JYihSwkQ4Jcm+GeUpnpTtANG341glOIzBf/mNAo7d6MfXbs1
bi6JvA5jY+GwWyzHe9io/n/Mg/tS8pQdb3HWyj4H87DKTU8qXLidGyOL2jhp26Smmqlt0aRGTl69
YJan54W62phZFXmYVR8c2PoJRseydARLRmtGUHQJsw1jDFEIrkYGdLEEEAi4l5AbUCFu2Y2LBOt2
e/HIPvU5PQWkanm0EdZ+RkEhHF3dPFafhXhTsJcNyqeQdEnHiBze2KCMe9RSu7OlfiI1OKMW2pjN
YTg9YxMMutb8sedNWGUVwvbLI84m7vOmTofhON1pZksoBe1BZfP0gHdyMvL534NMqR3vyY2aLaqV
jFc4fWMXvJB/j8XuZTfcpepuFsEcDuqgrDRaMQjFhudF0abb9yVv9kCP5Hl3zRELxeLYOxoQZJ7g
4U55gUJNJB5R0Tj8Nrrr9Z9NKqH3vo+iizEV8GjZmYGw17/8AtzsUKc7tfnWxUcSgCwruGLSOB7n
QvBX3w9l7akAWwJrOHCw7h6HW/2lMjtPrcFdZfr6qwsCVQPsQeL8f20OYFSZW8rx5hwnAQ1Ung5o
KOVMrV+AhEFPSu5VHB/edg9UDOEhhpxCh/rLVN3m15pvZoLkXTd4EgKXBaJBz9BYRv1vVJuspLPp
U2FYr22vIXpcFI861fAH7odYCtjz0LEtP1yWavya9UvtrVZkc3y3RZQCXfbMZ1F5l3WyLMk2Fer0
93DbOzmyUxBNObf8ZAXnEoJ5chwTm74o7B4qQEf39D4b0AO5v5DtJaR/Kd9Ff1e/8Hs1p8tt4Ohc
pTAVFjpqIh+YaEuFZ/sPJTuCmPMiCtHXoI6WO8TJZuHdgwgfPSKM8ICnjnhFzAmOBkMvZmZF5oQP
qWrrXn6aKbXAf2v8HXf0EKoRfZuLpP9Rfd8lEopElzmLdzEJoCwW3Y6S28GNg809wUPQ3vsT3nx4
Fr0txxiN6pRFkmmvGiuki6RCf9iuycZYCO4w186Le5nzybIE/9LJ8H53TjMNbdPsR+wEZXeEDQUV
UBJ+y3XeaaaLsTE36UqsBF9AywV2gvxemMdtM2IZjhaxwHxXFrehcLu/j6Jq5qeZfajxzuvfJSYt
mP3vKJKz8JlpZMCVO4DuY2XRVM3nTvePLNxAMO39K0czcSqZodQgd/P1jNdxIiI24rSEB2N/1xyu
/Dvh/Nti1jJPNit6iv0/NzCCTpiRJpYKf7RX834clZyu9aKq4N4ci/eGS+JrSD7h6Q0bfLzlQGdr
P70yhtrAB86Gqq7lL5fdBFIwxWRODHMvescFI7REJvxlYB0egffSoysMbuBfta/NB4BEAVGd0cft
FhptHibp+l5k1GbS0pO4Y7fM3TCqkql53w2gMYwACSOCKDHv+y4SAuHzu9BNACL7rpfL0LnxJydb
ujf5Ih83uBzVAcEo1UhCLv7PRPNtbgI2+i4CkgAZttWAJAvJHHpcSTFLbt72tuWegEKUdqQKaJLN
edOwA+4cC7OFa/eGBDOrIIvDoDcjjo1x+pzRGo/vbbc0utF3n0b7RR1ugITRb1D1lid5Q8qO6Epf
EZZoIIhqmlJAbeoS6aiwaQeamHmkQNf1ae1bx+lvaqD8l+XY6nrJSMF5kvbqbYagkMQkLuliEQwP
KD64Fj1OJzXKgehDDr1l9c6NVt2OLae4aIKmuyJt5uNck0KTRNyNlds8vqtX5VeX72fcWldCAKod
X98C0F8dF/kC4OjgIv8QADBeMzH6bDQapnMm/qqJuMgicKPMvTyT2bJo7RCEtKvSLkwtCvJR7p3a
J118ttDNFr9xa+Lm0KkjVaTcI/xwI2tI5LmJA4lZjboM71eS/oeljDE68mB9fYUPAhknXi/9d14t
i0SQkTg66pE/UJanEa8G8pYLnDOlhB3Inc5ZmJ8GAMPUpjcgcEsAOwLAf1Tcg1jArYqM9asdjiA1
OzxfMDqPbwZ2m9nl0uzKoedaWGtLv97iSNYqtd+z2fC1+VAROJkWHQ9rNrYnbRzyqKRG+n8/tYEr
BLZKQuzfnJgnUyg5JWF4wfin08rtdkpdOC4B71NzJItYFZBKkPPL7bowMcRtrG2s7mtkwptjbZHv
ZRzjdCf79v4FerTtnqYAY88W+5OGvfCbbZ8Dp/z3xDk+nSQ77Ajn7nJMNwegOIsb3H7mhkkngS60
00HtgdISorr2OyHkwFhuL+w388Ii6wCpV4ceejb+vyeCMau5nExG1KOa+wPgy2W32Fvf7qU/x70A
2nfp0C0wtZIOsyLWht+XVIRE8JFrcqTHqQqamW0cP18nWzy6PeY23DLkQ2LAeEPc08ucN5LxU7lo
RZwUMEv09CsRzfB298Og3u1BUdxkOI3YEtAZ9MDDrr2KTVHk/TVc1N1YSoh226GdT8Lb6eUzr+/r
zsQNlYIV5ulZgyhmsKbn5QtyGHNBmqZ7l3gHAgFjmez1a25+qONitwTvXb/SdFHaARF3vLAhFmqG
oV6nDnj47q1pvyxpPyKjeUxxYkLZdPyL2umCFELohvFkvEWLzRPF280STYDF7n2spkG5ikLjdl7E
MpYmj4Uz2UhoVbX71NhreyTMdhlmakQtXLnYS5EhKlatJcbn2uweRpOSby1sCGo3nakr8XVj+Jcq
rsi3cYc1AYH5YyDN4wrTNc0bB9zM+xC5pakqEgIaAO5xrqje57D0wqHoA4ZKxl08CCaRYEKwJDP/
CKV8CAa7qwXQMo7YxveCKErPoD6U1A00QnR44VTWqsmVthAJs1mqkDmNu22MPYUwMhkA1nREQVu2
0bGn7HbAAxGd8tJTxIzoBQqaeKyRxL5x5PaCB0aEz2mowDJhzZFgZQbhwhmOroJDusgmn99qCgLI
wYk45Xhzg4Xs2DxC00Omm1l1xZmNqIr6w03DpKtfxQ9rSMYtZ4piTz4s8okl5ClGVfay3wn05b72
WoF1qSnu9xcJjmKsa8oAYXK4GvMvZy+NcS7lvCg+/hFaW3Bgkg4aygYf0yeecSTyD5pxF2DlKRI1
WCoExOlc2X6ngfJOuxRZIlLJTw6+GXqps0tB/5EgArt++VI0ZqF3T+pQmuAha55HkUkhmQIH8Re7
zrPQXfG+QY66riAUv3ddsqCE7vZWa7F7AscbHJUGkgsAHVOQ+6fB9wvg9gskRf1gn3OqJ6yd6jmv
89vgtyn3dcaOuiC87QXPF2wAMc2/P+pxUJC9Ltbq0Vl3AENULia0INDHQz8ptEtXxHIhr9Uezfev
iwe7CCg50gWklElARUn7gyv0AtwT2WXxWFd5a3uOtoFO3IjdfwXwnFoaZoj6pr9fhecJ6fz2/cRz
00dznhiIb8D4XxwFcp2I3uUwDqXKfBnJtdFwoGHKDP7bUl/jS2wl/Lr2PZE2PQqjj8msPxhrF2BC
fjmR+MTDAaXpbpceDQyIcfPRfQNWPHmfAt7lGoEU5nAXG9+hhoGlgYGuV+5UJa1byXkPLibrhDZ7
VaNCz5HsE3xXj4pjMXyq+prCJsaE1nC/66LVKpffsgyxz9NqnNLsGHy2MmO0yzQ14FfGJK69A4I5
cFKu5aWoEmiIuq3PeOW3W3v+1tE1uOyVMxam3jQdUntXC3DKEq4xM2vAvDuaaCwJVcfEUzMUKsnE
C+QAY+KoIU/Gs7hACTAKHM3aB5TnL7fHPT2pazbVokSLFjMq8X++wYJs3Sd1VZ62dAKEMLcvHybJ
+Abh8474yisv/IeZkkAwW1Z1w/J9OJLrl3gPdhVd8EI/u4Rdp9m0IQfMoeoMZrLd8G6p/a/WfxTO
2kvFHdI8cdGJv+hokR4w4g/KZGZLg06fGHqaJfMxEWmPHF/+HibBcQaKDypWgzrIoCmeIyfqf7gt
/tDi1WzuBRQSuWD1zz8v5GIORKh/U7Yy1Mo0Q7zuZuT0DReED9JKMApeKw+5DLDR2bGadNpSFtjs
812VAbHGKyNa8G2iL5/5uPyJQaAFNMpZS58kP5vhhDEgTxOKafdAQwmebdlVtKpZOWEHLSQ6roMR
q/wedkPbecMkUix/aPPowLzNVm+V/l91UzMJikiunHoMt1WOsZnaiHYPZcKP651KmLrXXqqI9daj
EkkUoH9hYfOg5Gn73P2WzjXTLtiMSJIE98D4jJ5XE1SiqODxJgHkAMM+HGmF2UqZkYCrzm6av1R7
DYiolVaw3khHyIJMu9BThfEw/tIpU40naKBDrVO6DXTbuRUB/vxPtTxZnAjLl2V64VYUkGLa5TlJ
RfILfdoub/Y/QcAU6tuDKo6BejhJ/GXhRKe7bM6g7nzZz1zw+YAKhRKzw3YV+8TaH93KEKyWEUqF
rfSqSY8i0phtmnyxHbbEtENlvmVbah8RHVYPd9C49A6m0VgLqbuLuFwEPTU4xIf9LIJ7+OmwbVQ/
OqJVjDmTycuYATAH6z8VRsVVWIOX0Lxi9xSFrpe90HjEwjHGXDEsPm/eEdQzjgadWIxCswZ6EkaD
9s6cB/X6E2RIQ6gPaChGE/htA1vq++HLwK35CV7h2ZfBCu9pyfuSCk1ilUP3tTj0dMxNVWoMtxxu
2CLZuOk4gmTttQY8iSnxjPUL0z+eErbjizipMo6/+eC26QLEq0XCbtEKvXSKiTqg0GjaKxKfgUHk
EzXruRrhXotXZCa2xfr5xGM/AUHeZoBNckX88uSQqIv7BQcsxTIHEMPrlH0YJqIBAITkhOWY2PKo
5tRwSv1wIQoPu4bqzDGMkHqohxC9ri7UzcyNZlhYNQOgyvk3dgy4eFOKi1Od9eSSOfPzUpHCdjv0
PFyF3jucvkt/fPd5J2ki/759cZiG06oXZbSQrm7o5S/Gb0fvjgkIBqp5FwpMpSzadu4CppPn9Fy3
8rVc/9Jb5kmmhz/aI/RQTTlK70ZBSME405pzS8hF/cNHbDGXOP2A27Z33E8FKIHbN0wz6aNICXeY
HNmKYEy0HooSbUKEi7rY4Ns1v6GY/rZBp29d7/InkqmK5F71wQrUcMifCV+7DApJtT9l4RwKV6YC
JW0J6jMH+JAmnz484fI8FR1iENNmUIdWAOD1B8hal/KPggxXflYOX0pWI5Lak52WrWhNeZ7Ycp3g
7dX/mujtDPodjrCt/gCGCSbjpsi397URnOBZP1KwHfy8ftTg0m6f2S/LjAdQgmlDHj2yf585n1d7
xqsHH6xnA5u0Qv1a8RE4woZYbnNY3ilTf7XAU6jyx5oON0tyWwsMfnf1Gn6TsUvjEW5/K0f3S0PV
DVVwgMAcB1fSXYaobUavcGW3tyEUI5GfT7yO1eTDRioa0VC5aXCg/8iM7cyM6UjLPWaiM2LGm0xn
/jCC3TYD4r9MMnmYtup1xgfE2TG2Dj2lUCGX6gdP+w2Fv5GU6P6fP6aY2Gk36U3uWN3ogR9VhWRx
u2ykxU7ubJE/AR5B79SkZyI8Fy4y4eeA5XQI/SGYngdzqzUq5EpjJ0LH19m6ObtqKSpLsxIHM83Z
YCUMS1z0d1VYzNouaWbYQbY6+onrljplDPvw2n7KNmNf/fPPpBXgWRBSW4yvv1BXMAiOt4qqHaE0
biyO+05AT/TXj+ki/44C+5RUYlJREUvKlqorp9+HtqApt9UxNc++URgxf7IvxQZranQIj+D4CX5Z
/VLnmolvI2L3n1qlexK01jJ3u9EO0S6RxJY9Zs7FIKTG57gdPqyS7CsFEfPosco+EiOM1Lgw4/aV
NqzM0tILqIH2wB+LNrfJ8VY+HeIoS7/iUJUwFBliVnhvR9gbdxPVmrZvK/vMERpn4Q7DOMuYbDXY
2ZCfC02PnPvX6bsatPAIE/dGD8iiKo1fBNch21jTUnu+6XLikOvOJJhwbWJWtrXiQuk1vsaZLF/L
cbXf7fj3Fh1uuJ9BkRgwvBTbJmLtji48REAp/cz6t4UY7u7SwStiY1bkkIgXOS8yzYQZWAF0Tj0t
iPsbvYGxQ8IVZQOWVZOYXLpjHRoMp+IhBx1ZdZEgakhyiE92+BWtTXogwHz3rcG2TXTtZozCKbmY
PlGy+H6Hg0R4QBX6y02V2Z1LEwh1fvDzXy/gVSDE1c+GvDouMWIgXZQh1/+S3pAKlic18ONb/1v1
lOvTaPdZ6e+Q/Ys26axFsF7l5RhKkr1vMNUf4Qvzk4IF4eSFezKlxOPSa0UEUL7WNYi3L7OTyIW3
IVI+36b1YNuXpjQLLIhLD/vUcG5Oee3QYjOsZb0vepqsQ/uLTpe7E9bZfnnZyd3cd6ro8Hphy4sc
uCc/CRMQZQVrf4oqQX9ofa751zJYuiOG8FuLMFkzNhKCzBOcuXUkE9XUosd4cYx4sJAiuQyXezhU
mPPAo2rIIH1ehDu2GO+djQ97Iw5qOfkmBjYbaof9fpO0NsUdjG7vjZ+4FzZ3mAHjRzrLAWmNqVpy
TKgkIyphpj71RW9434uS07WPRA3k2d6nibcQaTap5VxtsogDczdVwo3Y9PO7agSe7tJ2jJSgxbRx
RVvDYD8O0pm1BXG9KtneSeTE6XqhCcYwaT3vHqYCccjl5RyMrkDfUkq2Yyi6teQ0EBjH4sTXTPCO
EwZP4pCwXMXbClJeQWSScIHom7jhJ3ebHYBkm3slCRkf6T5lriG/CzDavoQK9HAGkXFqDq90FRLJ
kC77D3yRlicmSUTPcSwT9Hk1Vq09V4taRqeWI1OjlXXJaLgVmDZtUJdQwJyG50b97I6bpr3oUmFo
xLzT1Jp+Ke0yLbkZBt0hJX0r7ytkG5cJs1UT50txr9SQrsUDoK+e241iGo5lLZxrtG1wbYLVOdYC
ygPUzLnj07seraw7pZ79RvAaGO9dOVlau9njRnNbaC4Id+MiV0+bTGRHc7DthZofnzDREnjPQ+Jf
Bjj0FuXTAkt7y1/LVFHzYwyy3ahtWwIWdlDo8GfBWSMaY65ycKdE9pEbzCD76RRxpl0Z+x24NgBb
QpsP0ApFyJ+TwqLcWUqtuAEt+MZAL+GJop2IMaXvwRueS64yj+m6dBqf/nkiPM+ocWSQ+JB38ynC
obnqiqYXJhu/9knPS/3X6HYLElyfgQqUDBUqwE3tJwcTUwFX9CYHLCrsIPx8SCvspVhzbNtBzgjb
pAPT3pz44bi5Er/dZlY1FZh86wEd9a2rk8L1AHKWDutFF/lzFr+sRp0oQ2Oa3A5ipUE7/wWxAONa
lN7kFoB03ATTN317KYCElIsYDq87pYnqbJyD1Np/0sFVPHG1+aCCNkF5ze12lnzp7OGh2k8OEoYu
9Sy4L3cFgEaK38ypqSxbkoolZ0rEw20dYMxDQ2GveehKrmSUQalwjoeyuPQBNeJ0cax9FXNREFXo
rVyN12h76nMz0SFN6X2P+c99ggYRSSss8Z9Pelf1vQ0OG6hvwXpPWTns6rZW3FIxrfnkRdEFsige
A2Wxwz4PPfa5CgoNDmOKi0ev8TXvi4k+vcYbYFvkB2JUg14mKEZnFkvkEmIBDYDdRVlgUgADuMYf
sxlDnatXwlZXwi0t1e4WQb4YxeoMdhNq12qzY2AMM50Co/ydXwiBX/j+oFnkttpZlLIJgWBeB3qa
TTs5/ASX28rl8P6FVMjmuRHY+Fdyi1kAn1bub7ylV5jcxR/nNAhnt5Z7cGhD428h2+u56iO/Epbk
Yz8LAYYuYYdihGZTdCA6F8JTD3lg9rDE97Kpw18mlBd124nXsyHItEkzGEkvYTH3ca4nculswkEx
ux4+3ILR4CZmh2kxbS0EkSZPxnvkIRebnm8L7rqaMh/Uy1V+YUTnedW3ht93ZSD8+bJubFXMJg0P
+uGZ/2Hk/TUhxe2g82mxBqUK5cLAJYc/YOgDH+n1xAvfs9TGQJuo31TmKpAHLRpufDIWt3OMQ1bt
0UqNW0rFVqCZZ4U/hP9MeQJ1nunFmQ5HBuFzOo+QrNGdWD1gwYQiP7cscbGRzOgKY5Nrn9lm6PlP
6DPhU1rdvcdct21FRnRTylCXJSo9bG5UMvo3MN/+GzC6nmyhVhHuDHjwCmVaI/llmqfDkSk1r5jX
p0kFrIPM2XjLv3YL05CnuWw6WsHvX410BFKbJbifmT3+WC6ANDt5lfNZWADqPjCkc0cPh2+lGpo4
Ri3v96NjyfdqkPjSWTi+cUNMYLnOaKRAApECSqbGZJeR4owZPaifSHkKVcqDAqJPp6JomqqYH61a
EtFKlKBUkIbJ6K+IzRpGYy11jhFfI6ndqQ+/EXEhbKG1l36akWzwA6oawfMSoFdE/4FUohFKUXuX
W+fZc/8YE+QuyE7iOaPzG3WtXwywYzG53AvxY9enU5YVj+PI5t3mE4T35x+KPvMt4H3G57dS+kr8
GOUEPthErX4Ss6mKndLMuJl3DHdO3OPt6sEU2O8zydBqBKm35PC9MjkhxHWY5fTpKGOC/SqL1SCp
JYbGSBN1RjuEb88r/3CDime/g5Cd3Dju1KQ+YQn8sip0N6YfOSR38EN/u3qps/ohzix28fG+Ode0
uycxlW+QTzWfXJKpMJ9FYSoo0qcqz5r4IassW9LQaSK3MeQqXguBHriuxwJKZSvLmHRBVoQnhQB/
6sdZmMIxDU7zmJos1KepdR52bhO3h9DT6vZpre5EyVktMVJaPCsh90HGVWLxuz0c7XBgKbZCutde
gptc1ZLn4rmu3CMx30NPBTf1e5UQ7meDdM4LwgMvz+l8cwkOp6C0q7ZSGaGNqntw83FIWjvrE0H6
38g5cEOJbefwXbkYMz4afSJY8f1z8/JQQw1M9otNybZAc/pHv/8HB3GjS6jMi7FeVwVO3+uobJyg
KUUzEW0UMsmFnsFWlyvYg/z6lfrMqtgAOGdZ5FMpn93mTcZ9SlcCvIZwNXyBsoxuYXhGPsYj52ej
GR+go6ViXANiBjAQDoGqgVviXxhuQgWxThsGH6XdAs1BPJZbaGFanb9oki98i/Vwc8G80lLmUsLR
d9xM/QFYFKf0EtDlW5XWciswWO3+jNkNhrQ9/aTcwl3Oe5/8jeUAVx1NSXlKJuHsUL61MiRk4av9
09D6eL2GE4B8mchG87XA8SPbGQ4fWGcZg+UQUaNHXHGNiOhPJOVGmP+4Zd6aQQU3aXEJwlN9+htG
pEq6r2Zhi8hncj3zosRxyPOc5RQlMJFoYTOA+I9B2pxgRaD2SLastjFnMBuGGqxjEaehEFjFxdGo
JLZgQgrgbb3fVA4MiVoEleo989gG+7OayxHZrVe/+xsRJcwWlgJzbNASMcr7EuvhYgOxZEEzhgjI
P/oYquNuyt5TE5K2SPMshNYSDJYMqvMSKl5RpLUmAOE1opQbZF86ATFVhEqTw11W+n5n32q2XxmL
JYl1tupo9jqKH+uFlE5oQjmH16ev1AZbX/G0JuvxVymy7Oz8boIyEFMEpf3vdq1yF6dNcPRdKcvG
c9HiGksABS+/4+gPzPd/RMSfipS3V+V+iH4M4cqImOCOlxlkwZhdSZaz/pr0fvhZrCd55j6MkC2j
1zYexzEpJn3Q0c5NlbnQHUEDtYYltdWHC5cu6bIQdgmKAniG8mQqWlUjs+16UmsytrLiXsufgsw2
mhfofd4z4iJTzSlFfyoFbBoUvooSv9mWsGcWjCdXNeBQTQN/fS1xkIWBE6Rz16P7DmivsVd/4FTJ
WAJHG6N0tiu7WQiBEfiV/tCZ2Ww5q4AZT5QggaJapUjaY1Mp/XgVi6YdO2tXsmJ+FzxovR/LM0zj
+KbybIHFX1o6TN3hzdrQOyPS7XF5cPTgtgfGSZqnsAWP16XuJ69QggLz4O7GHUGmWcaBbXZc4oDY
lEt4PC1jV11ztW2IYa4Fr9io/qENDWxg7n8Ch3RR/drPq709oFuBI/GcKay9M2nKLWN1G0KMDVQO
HZv8uEeonET3VelpFdg/+TCJZ7R3mTQlMlnIFDRq55lkLKmj39jy12rfNPHAXRlyxhtUQiSQ7ZWE
nZzXaKj+DHDWLKd1w2JOwqMbS2DlfmZOpBUFh9e9dpcCXtQ8Lce8/Axkg3uh5yZCs0kO99oNLJjg
HB954rWHAnY42Iq6Q93raGudOOIVdrQTsj0/0sThfvolOTksxagAlH0HNCgnyPPTvpqwGVEkHLI8
JaneP77hSdLujtd8CjA//MYz2JCa1fltLM98O0wSInlVm81HAJhyQR9JfgsKjyGPXNdl5iLz45Uv
8rZjOKqg+1d0ypDIUSqE9nWesyWFs76QCd8LIrMFMxh/U5rklf9Rf/WdTy1tR7+ji/RMidVF1RYd
ipL6J5zA+Y87XAvCEqKHkteWBCLNPzXkNrMKPjADRYY/gZw2Pz9xjEs7vO2dydJk29N0H1R1J6l3
TOOVBvSPFYpyxA+weswuigp1Gk3JU4jHQ1rc9uEiBL/9Z885OzqhUUG/+zdyyjzJeoY77XS4k7nw
UR1W3WB6ZO3mryJxQR+YoQnFUrqB2mHXT/ztxz+4g4Dspa34diP83o2l8vu7WJR3Eb2neh5b84ni
kQMiwTOz5j/W1RQKuCDC0VCAGS1b5vgqdJVKaGtFMvVMZzXUXh2AzveyZd6t3yTCA69v96eDzRiy
cUR68+ugkXpI0uZjmAyM0WC2Gt16hGpahkmj53oL6oFYs62LtPbGOoIP6sRyp7T2ue6dI2XMc9lW
IvwpuA2Ut5GlOIy8T3jFMoFojm2NIXGTXqJsXy4I1yyjGeykfF0NaZnQWBFWR7QEtn9AawJ/5yoP
P19cNDdHP6vwgErWnMZuc8iKOhWwOpM4p9H9iZFGgMS1oLTqrIEm4pYY7GE74MMWjA/lqg/YMmWT
+uv8mFH5A535PhBGSgy9lpPELn0o80dm6Xsv2qm1DNSKy9MrHfI5sdlZkXRjQ6Ye3YL5653ZGzDe
YAuaAN6qr2tNnJ2qJu3E+AZQtyVzwAAxRsWvDc98GDQzoxXnyA9jpXScZ8Tkrx7uhoGCrIvX81Qg
iyAVFqyP/Zmva7UbQR+LuSFMQVSPcm9tawm5nyHUhWBe9L7w4PmRL7LPsrDK0x1wLRCHGJbtnIUm
ZuVG9fdwZ3tk11UZw5UqccGsMUHoEfBmqfWtKMqhHhjqvzYz6jDtf1hjaduIlfy+zPy0KpidSK39
+9C+rOrFywEvZ+96isVwvAp84hkezcjyx9cdsTFD8oX4UawspKxL3vafCi2V6iGH0KHddrdkPEX1
F2lTKT/CHQ06/uhvgp6Mj1wBgJPcj+VyQvJz3K9n+jQIWtHilcJDR7CuTZiqBV7KOyKs4T6QN8rK
3/CfpGY4Cu5TAICvm+M7RQHJWTKr8GdT9v7nbWqIK1kQS1vY36Qnz6A0DHkfxriNfYhoYxAaHMC3
aomLz76BySgILTbCWirx+DmczahCbBX4M1TXAgqnNvn4quDr/OK5wNa8y7IWNDFDAGEKa9gMtKrp
ftgz02B3oAg5jDduZg0rA4vaPFc9AMrXCS7VUsMNISswjkGohIs/yNDJGdQsu+jY+pYSFaBxMs77
H1W3GPCRIa9+ryh2mEjre+FhmgEsiRu26/UZ0YtS5t96SFuffCFNnH+43OXoeeImLScQdc8rqYUc
XdDj3i225Wv3hxII4js7r7xYhZP6dV6axWuiCpn2Yx4HOh4lfvY0yQZjfs0lZtDdlriOL1uxKT+w
eDyCpsDkKiC7lryf125gdcKJRFM7J8RwAehaZ8lqDNzWPFk9b+u3cWZGhMBzUOqux6+SUeK4/LWH
z7wXsrdR1NRAXjUDnQIOvignrXY0ZnHWKTef0i+H6sC/ME4dMKiO4n9AynhrGlVo5bGoW0xyIs6z
iOJoXh4Kg7FaqiXcZ31y58IDMXORLDjGBdeBA+b00v3R4TSulVFe1SmJzXFNgLthd1yfyb73SbAs
tw==
`protect end_protected
