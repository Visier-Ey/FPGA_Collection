��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@��D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F���Dx�hH#�9���߇"�q��^�ኤ��Ί蕈�D5��7u[�j�����t�
�T���L�4��������P���F���6�D���2
�q>8�\���{3JZ]���P��`��P�y�7�SZe�U�)D���H"��W�)F��Ó!�2$��mcmtD���Etg�)I�Q��j�Y��p��Ԭ�D(pG���(ԁ�֝�2������g"�����dV�@E��U�70�J�ss�+'>��g�ʀ��������8S2u��}��U�f�w�����֎+I��e�q���k�÷�c_�}ȴ�;���_�s��k'�5)M���چ6^����tR��	���v��]�D��i`V��R5ޘЀXt�� hu�^�F@.��}ǩ�X8�~������-z%�{J�4r�'�eX�a�4A+�k1j�g�?IKpdwc�hK�E��A��ԧ7 $b�!�"��z���M(��&yR}a�@���Is�ݓѩ��Ps� �~혹�����0�4�mj��6�[	��4�`n}�ЄAh'�����ۦ�6�cOX�z'\/�U-���g)�	klB	���c��4��W�u �� ��$jG$Ew���i��e��ޠP�ƀ�B����VNh���v#�#������.�%r�z��r�"�6�n��h:��6ki/'-|�U����P�ݜx.�������\��˟���V�x�Z%�6*�H@�p7�B�4���f	�5v��d#�G��a�Y��˄B��_P��j�v����Δ�h`> �WjL�T^��d�l�F�&܍��G��C^�xOv����й�S���9x���Jq��Ί~3�J_&���W������m};G�c���u�m�6����Zi�>C���w���C���)�h!�rE��jkx���X�a������D``��%ʂ�?ϷϿR��])Q�.���Hw��qlۭJx���b��8����#/W!/��:��yb��?sGn�BE&X.>�9��x�{�Pw��;-�n�`��W�2��"������ĺ|Ϫzf�x���b��k��q�H�����E��?�������c��!������m�$�&tr��1��ulFU�\	6�;��?Lh>�>0`���Xk^���C	�J��0Ux�WA��IX5]�Ο����D�"˕�j�;�lC���D��^�ꞯ��;ڲ[����bj����TE%X��xR$W���z���ȟ��Ѕe�b����b�,���+'�^ޕ����/ݯ�!�p}0uKo�Pd��n�b�z]�}3��f�H,�p3��,R�<��``�f�d�u�8�V]����2��@a����X��ٯ������&L��V('���t����g�w��(��u�v�}�a.�`<��� 7	\#�:Ȩ���R�l^�,�����?�M_�61'�v��i9&^��nG�Kn��T渊
5&��H�m�x`ć��46��0e�����(�cѺ��HP����W����ԁ��N��m^X%o�})�Ϧ��^{F���](T�>p�^km�8��j�K�|+���Q�0э��v������df+!��3��4}�Q`V�z�H�5����-^�(f$|Bhn�7RuVv��+G�9�l?��oɤ���T;�jR%���TDJW	J�aA�'�D���J	��̋�-i׆r�䣐Xa�95�9;��]P*��R$�l�tf����Cz2O�H���kѵ\֧�L�"i��kO�*��4�V���E��^�b���S]M�VYJ������O!���W\�t�`G�a@�}��Ԉ�����3�z������T��5I�M�6ڦ�Ƕ��#�K�?�����td:�y�!B�|��;�X��a2hpt$D�5�r�1�(�X�B����Qe��rV����Q��x�J��q��A��9�Vi���t�>UXh���q���o��$�p���SFL)j��wA�҃�$���&U�}�'}|�_���נ�6'�dt�F6/�տ3� �f"n�	�oKd�d�OWͼ�/1m[1���1�NRΧ��s����wd�&h���	��["��Z���g�~���{��B�&�P��U ������b��m`�~j!!��0[�S*��:C����1��'�����s��w� �~t�vpR�Fp?�U넴�}<�#L˹�p/���@v�r����D���D;u���[@��·�hpѹ��(�&�˿=@��e)��6W_w�~ܼq�e7���v���jDº�:�_FƷ �����9���
��������p���&���9��kl�c�$���Ԕ���Z��=�n��x�0W�g��/�e���n2���G'�
3_���H;��N�"B��5@P;���8R� nc�%��X�Ho���a�wq�Cu�%�^������H�%��;�4�yoO�H6~2u=��q��"6�T6Ғd5�	l�H�k��V��ŏ7�l�L�����A���{M읳�~]-$-[А����ס�����ө��]���^*w��h���D��i����d��:��'V��� iB�Y��v}��X�,)>TC2��%�7�U�aXec� �qo��Y��3��Q7T���G�[�:L�1z������H��ƫ��88���[�v�K�C��������aarJs�C��3>���� �gS	zR7]�f�RFč��h�8�`A8=-����~��n��N�|c�����ǪTF�Õ����!̇�X
i4D,M�ī��?�+\ʣ�z��O!��P�$p�p���#�\vŇ?�����=�0׏9	���q��w_�F�e�����7JZ��9@Б-���RBqjxd.A���R�Ux�yt���g�Ӓ���)!,n�x��֩ZY"Є�1�}�	����)��������*+\�Y�0#�4��L���.dʆ���VD���N�Ҧ,u�xX�Ly��7�U�L�1���M����Q&q٭S�9W,�������]���C����|�[s�fv����ݐ,rQ�I=��IXKdY� �U!|zwt"��=�dӝgr@��:������غ�q��ޮz�РX<1熇*v�]��۵
P-I����G��6�f�yYm��O�\���Gs�i�r�djF���,}���"�,�V�����",���K�#fF�]��smh
��Zs�HדF�֝�Ia?_�G�1��O;2p ��}z\߄� �W2NZ�1d�X@�MWӛ\�|,�)�$�I8u_KqML+��U�b1�%�:�@��&�����hߏ�ª�0?DCYV{'{�x�N���㌁�XP��~'��a�S�.����g`�� �t6.l��q���hJ�d�A�7����
[\��b���*��/�Z�NI�����6Ȣ+$(��`��Y�D��=��MـVqRUѷ�g��Ņ	���)���yw3v�5O��ӽW5=���. �T=�icq��j��77�htW�z͢��d��ף׋�ׇ
���z'gc]�W�e��x��~t�+��3�ϻ���̫���q��93
����?(��"p�֞wc����$_S��:�����a�>�g���������lk�R���I���݆U��#O �,3�#��3��UD�*av��b�AW��x�Z��?>=!b�ZP���p�3����`Y�2F���.w|�Nwqϳx���wВVa1��+_��x%��fZ���ߒa	K���۷�qw�-�K�����A��`�2t��7���g�C^��4�Q�<����L%-���|��Ch+�8����dY�pRrh��]���o�RJ7��ZH]b���O�%U�ӣ��wa��B�Eߪ� }�ҷ�T��-��d�����1�������c��&��Z�h��oX�擿��i��xT�Z9��U[�Ȭ8��f%a�`o;:K�C���Xy��z�Qc:�0"S�J�Q�����ݴe�,�Ŀ�<_�Y�<��ay[%b1��wg������E�Y�9X�1�g���
�ED�k������Ea���Ju78_j�Y�O�����3��N�dT7IW'W�[�Q`8� ����9��F�'h����aw�[,&�N�5�t$6��%m�jL�������H��M�&g�C�nI�
����:ߤ+���VcE�� �V��\��;��U.`�1w;ӈ��dqلxmS4u�{$ �QG%�%5ϢGWV-@��e�܉�@�����4�W1��!����za
�{4���At~�P����Ȓ�%
��1t��(W�OH+g6�����֦��a<��$.�P֬6�Tyr�z�(�b�� �E3�8�#�B�Z|T�Q�̬l�ͽ�g|	�a]�
��5@�����#�0#1&6��O�yX��TR8�*��ޔ���)~S��Be���rD�y�H�m�'���L��0�ke*7�7.��է`��F��Uaw����K���7�?2���;,+�0[8��y����8u��N�`�W}!�WK*����'�5�!|̊��'�5�"`��y�X��faЖ�=i�O��ٱ�`��DU�@���s�ֻCW����Q����C��Q+�0v���^�h�RD�BN�����L��'A�.��nd;��'f��9�>��X�R�3�y�����ɮ�>?F�T�����_d:b�j��´B�l�6v-t �G��\�Sbg�ӛG�P���_�	w0f�G��Z��>ݕ��� ֵ��#�T�����8o֔�d��!�oP�n'�'�F�6b?W4S�F����ŚQN��(C`�_Q����m����gܖgp��=�(�Q�͜�e
�3�+ǂЙ}sΊ~ �e2o������ё��!/�2-���i���8^g��]ߌ�`\{�:#�_:qg�/�����cɏ��n��r�n	�6K��T+�@�,�3f�T�!�A;�N*վ��|�C�'yhT�3��y�"��ʨ7R2Go��>�2jڮ���q��� �Kw�F+I��'�����Ld�����7���xdX8Ǧ,	gR��/\/�B��>!��;d�}z�7���t�G�ê6l�1
���Kk�O~�-��;@���$M¼�9�Hb�t^���}@o7��л��`#0�FB�`J:�n,KJ�j��qsR���_�'��1s���Y�5�'{}��u	2��{�x���I�� ��J�R�c��X����3�z�'=�Rw��I����*4׹�ˀ�mo��s� ����v#���ۮA�u0J,
]u0�R}�4y�gjH�dz�%�H_���z���7'���1E�����9JPCTFf�ѪQ������@`��y��ؔ�Q�&�ds4Ld���CF;�To}BX��6�#���B����-&t�n$�e�\3 �X�������+�:G��Ro�=�_y)�9@����*eC�w5�x��0V�qhA����\0��0T�/ǬܗJ�	0fo*&���%�M���n'��� zR?� f|�jCq�E	cA�e��j1��Z]�;�8pFx���)�G��^��D�b���	Ua��us�.n��*�\�K�o#��4��{�k�Q�DSA�����@Qv$�J��P�-B�Y���3�blR�}���j�pS�ɒ��zK�>�>O�sb�ݾpw��s���|��a"h��!3bK>cvݻj�)�H�7UC���5�G��>
�����y;{C&!�scΒsU*z���!]���M�Xh���c�Ǻ��7IP�s'Mw��o4[V�\Χ�� �]c�}|n�Y�: �Q�>>�8���5�^&?{�ߙ
*$���ۺA-��LV����������A�>*�䏠�8���eC��Mg�]��r����8���l7B'l����k�æ��?�J� x���MhǶF�:u��τ�H����G���Sn.��V�0b�e�zC����ƥ}H�F���bW��PȔC:77�����R!�~U����0�{VBSh#Ͼi͓ٓ�z���[9$B)Mw�8&��T�I��v53ѥ&���w>(/�fk ��׬���no�|>Խ�@G�����L�-o�.�e��=��Ҡo�b�+z��?��Mqows�F$��:'���o:?��ƟO�޴�̂�ۂ���I���o>s�0LY��p�dIb?)e�Xn�F_ъ�C'ZB�1�~�1�_@>Oi�/�\��g���?/�I]� �n�@�� �Ƶ��BG?������2���3+��A�p��G���CR�5��f���ۋ���αY����/C�C�U�[r _l�X�=�L���ɾ>T*� @���û�Ґ�=��/����2vu��'�����9J�oW��JA2�Jskt�u����4b���	�ඝ�{�a�{�iC(_�9�ʬp�S(0�}ʌ�-���]�RLQº�/��K�=ש�ɡq�t� ��M�r�+E��z����4� �y��q��`+��Ĕp��%(N<��͹0�c���˟�Zᩃc)4�l��xw��&�w�<�i�x�H{_�i��'g/�R�p).j�r�~��u�h���Pg�?u}/N�.�p
Y�s1�J�S*� =`�re`���3[�D��X`O-�'g����5�G3uj�(0�
�#���aآ�b*��0x���d@Ds��	���7%ǡxU1!5DQ������E��+���K�_@���]�p1�Ⱥ��*+���~��:ZpY�Q�?�֑����ŝZ�F�:���Rb$4~�!Wl�Z?����?��d��	���_�gBE�Ix�9�.��0qƌGl��L��D4�X$j��?�08Ln���xy�:��=ȡè�*�w#�鷶viYɕ�d�g�l��4X�yi�3;������E� l~+k���oY*;мSh ��]dD�a2�Gm3��5��|C����=Wf�0Z=������{l�(��3E�H����.�iK�S#��/�#H���O�x���F����$��/�Pj"=�@ַ�Y�s��߮�� \۳�g�h�r#�9�T!.�5_Y;3^�����A���ҧE�~#�#�s��wP�W�L[�3��(�>�.��tŏ�[������� �HWmJ"��[9��ӗ@��'���+eɃVX��W��a1O�ܹ/�dm��$'v�����y�sl]�����~�*����V�W�{�����GN|0��a��X~3�>������}���YY�[%>u�o���;&�j�|\�U+Y�"�z�ދkeJX�#��S�u���7���_OdRU��bX���X�4u(���4�t���g��du�usmP�߰�������&��mK�W'�6@�S�('DJ���m7�>�6z�oŧ�#���.�D�9r|W�U��>A˙3�.��K� ��JM�'b�ْ��IΫO����Y҂$Nq I���d��h?u��Ʒ�̑J��,�x����h*g�g$�Z����G���Q֩{T��T��R���6>�Ѩ�j�1�K'S�?��(6��};ۃ���5�9��X|G��aۛ�v	�V�Dh"|�.����傘�@[�Pw��S��/��W\H�%ȧ��.ځ�VD��81iԳ֊M;된�gK�;�#��z�r���B��9*V�i'1��	�X(<�<���d��H����D��&�@ɫz�,�=^J���+>Q�4��p�(.P����[�����1�h�|h�!�o^�UW���4ƛX�/f�^K�x����ZC�b�%����m��<����r�c@ĮżM�6v���($�EK8�W���t͔��`���9u�҅ =��}_k-���;���B��6G�K,;�TK�V�e�?����\T�NqR��Ӕ�6���#�fO~�lhÒ�Ug^���UC�b����i������L�Z�E&��'�~
�ڼ�����&�����'�M��3i�з:Sm\P� �N��&P?A���QU`*�T��5e�͡F��Y�B$45�)��m�����-�}i����Їq�p�M�ϑ��mvd��J��p��v4�B�5��Q���<�b$�.�ny�K\շHu�au6��zXP�5U�>� ݰh�s�ʡ�I)%��b 1C�E�2s�٩�~�X_����΃�k��R��g_U���P�]��\�Ρ�(���M�����'p�ة�j4Ω��[Q(��'2f�70��k�6�<I�.O���>e��)�6���Y�6����X�u4-�uo�`�d�,�s�ϴ��ySx����T�mVX��c��!E���Ī��2H �t�ZX�JOu!� e�3w�b�TԈF5�^��U�;��u�G�i��B�7QL�!yW�~�Z�i�o��c4�.�m�g9[��;��v�������
����rxͧG/ԢK�K�ZxDt:���`�C{�33z�z�%A�$�@�6�%ց�1B%�/AG�50$^(\��%Sx�A���XW�PߕpN b�rͻ]Mk���X�ʇ����x�*Y^A���S|�8��p�����
�R��_�}E����pЅ�k�I�8�H��*�a�p�;��=��᫰O���;P0F��&N�>M+�VO��&�[]����q,����Hd��B:k�E��ẇ*�������/����rq��o�
��+�O){"k��b�vX���(�J9*�c�������	A&�[�!A��"�fL��sbaX
�%U	k� &Q���B����L�=Sk�@��΋����7��J��3q�?��4�,�=�2��7~K�~�͝��=Cp�MS<�/��@qem.����w�гH�~J�X|:(D	��x陀�I�;vr/��.��H�)bK�!�+Y�C����O���=�,i	E+"��;s�$�i���^�\纨�X]O5Geqb��iP���0�����1΀�L�Ul<N���uZ��![t������Ѵ��y��m�x�������i<��d���̂�E�0���
�'|`����k��䗵��ʺN�@Z��V;g�wW:������A����)���������̫ȉ�fh���|{���|g�Ծ��޲��� ����!� _�2_����̸��X|�D����뤫 �F{�`��paΆ�y��mQߵ�#{F�O�Ђ
��� �QP��FuA�.G�5	镽e׃��D���	k�9�i!ԴH�>����J���~��2VfȺ?J!��t�f2�Xg|�!6�<uw4��Aي�v��z����Ż�7�_tv���	<�8r�,c�Ι�$������#�=���6o8݀U�
�@sD���6�kޛVm���ݒ����j����{�*t���� �E2e.��yd��/���M�9����s>~`���΃z#�g�Yb]�B���$u���Z��@��|���9�h����>!4��n�ƓҮj��D�D���Q��}��x
�]���n�����&=w&ff�||�#x{O��0w��M��rg�_T�1{�:$�V��t� �ڬb&��z�QG^X0��DK=�],*���j8��ښX�k�6�泧0Q�{J����`�؜�OgX%&�-M�,ZaD-]-��m��R:�GJwsfɽ��b�/�ĳ��(������3*���,���7)�4�!���<Ԕ�ҽ�oQ"�՘մ�n$p�z�;��E*{�S�j��dm{0V����.�Q�:8��m��H��H��K@@�x7�2�	x�[\\y���-rv���(8������"�k�W�o�*����0b�*ʢ
�tx��yi�v��=6�;9�%�ǧc�|���>���Qk�<�������X�����|vY��R*UNw�'�v���n��;k�����}���.�"L��1�2�.��Sm	ȅ>]z�&��