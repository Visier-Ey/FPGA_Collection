-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
vuRLlb/q1ckvzlWuMaTLZpXWZkpfn51GvdbZzQ9z63UJvE2nmX6JGhLU5Yczj2bYkzHwNx1sERlF
j0dce0I9l5hdeDAjGgUA784iHehOlpmOjrsgyYFcK5Fik24EjascqbCRU/zjLFjkVlN29iUCsAOm
KkNC5AGDqrP88wPtmefCwY2OyDby11oOT+iLfIR+OFqrrthdf3s10S1RL7ec6tkrZ15+RSJl/tzj
nL3zrjZhnpDQspIgnfFjmYqAVd7yWsVGFmrmzVxC8Hcz5VUYZ2YnQRQGW6WaKctUKe9inenF7jHj
cUqPuPEQ1p6JcdM0VC3ZxfXsQ0iUrroQpGn6QA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5584)
`protect data_block
BMCGGBZhOQetdJzGxgnAedpJ5WfVFee8wQRgkJF24QVaYkXDYlHXv7MLxnvW4SBbVeYBSTMRczi1
MedGF9YXwonBgNZVei8zW3dK0i9sYtTkF/WZ5x5uHoA9UGmFg67sI0PIp4bRMPyqGAQEgyaEvJKi
WZ2CcIAscikT7cc6RSKTUB/8GGCeYKuya6sifiUiZaNxpVF/vVvQDazXklyp2krZOBfpRvuS7Fc1
PrF8P6tFIU+xn2m1PDJBi6S7NCKoPQkdVFAKeNJKp5rePG67jFAMmY12BptZ37HgAewySNHYAUTW
s62SAAHy3cXAe386KT845CKgMGcsm5sZTTqaayyaCB03ywg+a8RaCgW5O1z2jwM+13w8j5w4Q8RO
mMFJMsUnwKJO5+nKniXNVbRIfBtXsKoXBJ2z6tPIlUQ+oSMUknbbfwdziKL4tyQcDeIbOIO2OA2M
wKCad5DS6F2ECvGYe4BqWRyXNse4sMxkIfD9xMbSUTfAtKf4tJQo4SD/GRimTk4t3ZODTuxZNysS
Y+Ac7USU928JOxbQ98E5gd+e42mX1e3GA6ADKhKibtUATGiBh4e7j7w6ZKZhpq9W3ycQLooBX8OY
veyHMN/LxRu00QzKVHXm8crSqDRvKAE4U/PNArKVRa8oVdZ5LsCaZ4gFGnrgT4exTFz08Aavnrp9
gD/zTSK5c3mKuxXcZbMVjTszhN7Q4fEG7Q3rmo9BAc3XELJiPFC5qvilqzrkO2sQi9pqK/xzdajY
qypV1poWRGxT/47OWCRFkmv1bgifis6WUdIdanqlr6bIK3QG1XzQz1D47E5npBYdopg8lYNGxv57
alXdndP0bffu3r3CgmLKCWwQnkHDpl1wSc7L7OqsA5UkpN1EhkszNd908uhHGJ5oX6m1Xc8VBS9G
fMbhoQmrzTH0/BLrnUJVaNZgt961yjGa/0IR67kEYN/xqYyKICN/lU9wnHWUEDbDkjbGJW7rkteR
5VPTsj3iCv1xecIbAfyD8svGcTuX8zSmC/QbXRHLVd9di/Cn7ar3VD7bcjSV9dYpNrskoODngJN1
3h5Gh48wdG8GNdmtf/EPonQTlKSF53kFIzcR+1rPMuwILWKVy/K+0q5+zw1FEo7GkSciQtyaDrK7
ja1AqgBN30Y5v5UMJBiF1wP0DxDgVwLsOpTC2B46PNMKynyKgVT7UPoKAHW4zG0Ajv7KkACrcXxt
gVz6mRYyzbYogI8cHQd+PdFlx4oJDipnGY6AhoM5sGPoe9PEou6k74A7sEEkJax1Qb9aeyk6TIsj
lRQuTnFnFRcjif5eoK9P9ONhcaK2s4gI7339Ny1JskhEqTQVSF+/wNbPSmdHUDicnIlC7Sc+y+wS
lUME9jkXgxzi00BrLag0ca5w1kuqsSOmo0zy3NRNlF8mJJo7DiIew5AYfda27SOVVL0tIEs0O9b2
T97B47kM0YaQoKOQUWQfHxcr2MRG5BQv+84dUKJEP5DiKKuBxDi7MbhiSnG5f2UeNW13ZNnfvJ6m
Buhty3J+O72Fd9/3DO3t7jm8AUbHwAGAF2+P6G7ozvMxU4dKaCx+xIg9qTu1w0xALHfwHBRLUhwS
aEPNf3CJGpbZxqSkVt3Pq2IZUsreANa61z0fO0IPbATY1MyPd0Cmm4Ak9Cwli+kXV9CJaGO6Bu1i
dKSO1qpUwUXeCwcRXGWmdZbVWEsB3JYoQ0UALWJ0Oc2g4WI/kDi3Y8Tm1/p+22XHBpsd9mEDHv3m
8OJIjId8mSZwy1bVpDTIBrk5edjkca2mOzbG90gCIJfqcPxm4UscDPKkobNLe5k8oP6pUETRrYMF
fnyBOSMQTdnnaXsq9JtAncfbZjE4wgUN/Aj0b3jDY4UA+7V/EFLpLq85fDeNdKUnw/i3K8X0IomR
2ANSZOqAPZOUQzvJqZbVrJuRGYR0/1guVL7ZKlMsNuUnAQSdKbEkD6ezDJqEwS0UkyhB2r1qq4So
xF1/QC+/3+mX90nHNh1Dq1/3/Km/r7WvLg1XVfn05y5CycCxzmfMxNyDnURW+leNjQRTDI+b9juF
8ONJyL2d5op2pkx+VstqBdKqgzuJl1LBi5I/F5JoR4vrEaHlzBLGMMEpPuRwE0/HI3h3F1m/cd3M
5G7UWWd3fzDlm2lAMbEsDZlbCCdQXCCOfnEm7wLg0XREM3i9dOVhIkwicsS3Qp68Zry6oMkY1IAP
3cDyldYr+L4dhw/7avnbClyrQX6wNtDQPaU5TQnw7OZLGLVbhTW7xM1m8A8KMQ7NhdV/c12TcuQ1
77PrAis8v0Oc+Od4vYETjpt/8BgoLt4qg3AauwttoxWXDV1eEkrYo/cIX+PvNzkj2Qb6CdijXVWO
oRnvmE2aTo6GTyyMGXKSm001QvAWMi0ok0Chd+WP4gWJQTwXtkyqstDXJXlyBApVXgLWEW2t4y8Y
oACKy+yxxqlC9atFGlEw0JfUDObnn6AXLclxz9R3e3I6H2Um3Lefv/76kweb04ujanUrDQlo172G
o4byOgrbgjW7Kqb9EE8tG0Qpn0DMpiqQS4AEaDd4rtXiSiz++QIl6I/hjzmRvIpXmhNJ8oVnnWbK
x007Wl4p3kHIcsbsmYXPvGIyYJPNUu6ny96MFN9JXy5V8PjhqT21sDmCFCAa9qO4Bh1ZKKcB91hM
uxeH7/J1NSb/vyo8D0HriLV2JsI1BZH8fXlkQn402NT0GFGZ8KbnO1jokCkxBfz/ShRXGCEDZB8W
DYlO9pxcBvR33CBUjj0d89FEAwiwXZc0TQ4Vh4yrSTlonUQpTgKO70HQP1ftw7r7SRcvVy8h0CAb
47nTTvBoAUI4Ge/zx5l6kHZMOegiZpRt3Qi1wXrR4izwmagRe9KdVuqRq6NVD3oxiQ+0wvqEZa1k
8LGyfpIEPRcY1mNjPcjb9N/PoQjOU+h3My+1wZjH+ly9qUCAYQT3p5BYJqTFpZBduS9nmMnbYzw4
sPmx+kwW0hVMGbl1DmBZRq+qVnGT/wPgkYQ3AA8hzOognCOsGjna6h1Me6lzkoow+jcmcndfzGsm
nV58zgew9r3O49mqmqDm636PkUqXa9w3uKZNsgn7EFTC1ywFzKtk/Kej3AVfztItLkGa4k9Z0oA8
aLl1MCmy1a5hPbH65zOpfVkn4NQ/jBQmywtYsqj+25xcCvdJ5uhhqI7E9VyuUuCWXvoenfYYHkF7
Ovfwd6/ltxwyCZmLzCll+qYhe7SNh9NvNs6PBuGSKiJrvKGsMfkUc6ovcZP0L7HyBAYZxb0V5HGA
n9CHU5ErtNznXzuezV/Pdo4d3jbsRtywQV052R6s/mlSvIP7UrzNVGfT+pHAYoJQaVwAM1f/ovuq
ZuewzChBtToCj+bZOe0TGu3Zq66BF3K8v0cZTsp5yym7j63xklZ5xKePItpVN5Hy5XdpafW56+bs
WO6BpuSus7qOUz/ZHTIiehjjMaMKy+aeuj+2p1g6BTnvkrwSYRmbjNLHe1sCsRKCpTVOOMwrABvL
zlyhKS8hv/xnGg6JewEb59zyfeRpQJHfk+RprAy7vw5UQQU5M++LqeN+gFHRtI3NMU9GTLINpQs5
8jDhewIV/lJTF9T+YxxVeRqfDfKE+9NAgpQoI4sPMz8HiXwTA3wZWfJaUfwkQQftIuCA6NMs3Rlz
IWNgsM6XluTV0Ld41ACGlmaSioHRzIf3pLNIht5zmt3NwsaHRtoKRX+n0xnN7cc7L7nT1LZ6f+qR
S7VoMZHCDneAlk4+9xn+dtmH+aiEtR1RIWZPD/r/SoclEge3XmGeQ7j5MPBrKR1lVwhFZlzdWsUH
drOXHrM3oVU8roAu/lLfn4laC4zxKscSeZjjKfht1Fk+1cDRKuZpVU181DlBzFPsZ8ZeBrf7cDNU
/hyVs49oHOtdAT6oQu9FQhNWfllZ/gQaz5fyJ8OyihZ+058ZixLlmkbPnPeRo7Coy7wCoPQx3ppu
4ima7atQbMRtx8ZJCGEoEuqRD0LwcqiqzDObjkW28lQTYNLr2a6pfn1zSacaT/BDqGlOKjodosoO
QAPiyBHcRXeKpNKvvWWjhqLjd92KN+J17zBuwiiOl3ig7lnhNI1Yz6c1BnIdlh/NT5U3ibR44t3g
FyFVX5qdxcrWsDCsqnvMf1jNaGrlvmjbF+B3fpuYk+Kl3yZu1aVu3tQJPVJRfPYBdg1xNz/kf5GU
8nGywPr9Qsm02IBPaTZSMPvLQeuTDNMzP1Y1/uTnmTiv1M94iScAEfYnxhjm48AAkluV0O3Wybwk
e9SGAnub9oF3/lcMPcDc3Bf9Y1ir3a9cpj0RESBySNGRwcOQzEZd2GGeLW/wKIjBARQSMI2Huye9
NgVgyWzcP6EuLnMUcO3AumeDB8uHOtSPJXaFXEMqtoyq9VnEQo6wXTgm9triHSCLgJBLXRYGefoU
3yrUrq1ojegQAPptpqQGkvHI3sHmplrQmH3Z2f9im55+O2LX7UZI7O9rxeyIGIBuASQTj8vZclYQ
+qSv2jh0Ggm9ssJOY4FZfHHlm2qgBUDwhSU5SiCSdqrmbR2YMJUC7QKZFPGgGfliqfQpsrCXpzGN
zC1BdjOekjJwNmGM0/MocimImcFIjmMGzeCeBJ+519+o78NWVzlcBuSa/XkwSS0sxDufN7ymQNVq
Ol/1KSIY3qI8JZ3bvSecBlKH4y+OBHvhXoBcIMWswtLK0wiE6Qrkl/bumGyUbVIKQkA3UlGmtTSs
iwG73xj6e7x92vzsp5c2AjpdW6F3bHA/q6C5rnvLDeXW5CE4OJvwSkgdcOV0OHPJzNI9dygpYBUK
9mSrURsJjptyl6QYshIyBz5jpiMGVyHGgavDED/KWstJ04auCXeqIJGdcvJskHlE16A1UbbmuBvh
uBzYdsRTdDgMgnP3233z5uBUV3SuRIzr/jsk3USmQum4CQp8rQfx91Cf9VvPqRrhU6DUnsuxA7pq
7j7TxYfnZe6u3Rs7F6RglrDdCL5Z/56JqN6M3tiuUR/DJDDvBNvagRswVIzR3zDHn+5E3JEUHBcf
PT7Z5TmgPTl4KpqiVot4edGtfuxwRaNXtKAFMobi7w8HULOdVrwK4RIokXImhmm0q/ZH0oM8fr8l
58D05Ddbl+/+cIlinfiouhXHeJSGfeGZtGl7Vq+UHeg2TxqKvbNt+Hg+d8V4K1Lyd3tas28UEUMi
x0EIWp58w/a+0jEotiFAlym9DnKzjCHvQmIfZIkNj4AYvK+CqrlnC8amz/wcsYbQG416KnNeBklt
4tIMlvzLc4QAcXhieQY8po3hkMPhinKe+tlz6HKTysI+uowZs7LoMO/4g7oP3o8ZiD8JVTvM8HIz
HFEomCXT16MG+6tZdZwKiShyqu6pX+7fHosCBLN+McjmS8V7X92J/SmBJ/DU1hY88bEa5i5am74y
anTaOV2DOxJBIKFOkbJyv84lYQF+lJqlNR2Ng1N3qss7VR/XZJPYuGpmycQ3n/d/ZpQ2OfQVbbzA
n9DAqjSdCfOp7TdH4UjpIS86xUA4bMvimpEOMKAtiDouYz29SvnKVfSGnoa++OD3Njgr3m6kS50J
S9+33DJ1i0T/Pp9yJ4F5uwzGqhyxSm+HA7iqZUN72wERjmZ/bLkIsreh0eTiLbJqyJhyE3Amz50B
jm01zcpKqQ80rmYZtDOLN1FJNmp3hlj673l+0yT4Lw1PfKh3yE6R2uncf8qpk0liyNS/tIX1yj5r
aN30d7DSB3QNkg6yANgBhulP8smdMC8tPeZz4Xv0QpgzD5+yNMBHrauYCWunHq1ywf5/JSeQbarf
sF9Bd7U4W9CMsfRf/vlfnnSAhhihTAzoobuASs4a2pYogmqotXfj7qsmTJwivLGnY95PawESvlxt
3Y5MHiC8uKzWvdcSDZiCHlFJRW5XIw4ZKh3hKUjeZPI8gz1qIaznS8BClHqUJkP5LfqFRdEPM4XN
PK4b5WegOBksT4JN/cax1onkjbSLZPloev3JNkljU2WSmVKoyLEx73DmLzJZ7grCQqQTbRZq9U7e
8XCoXH1F8ocpBUBST2l9pA6EAkSRtC/tWBJY5Vp69VBeWG2Vt/5VpRNggqXhROPq7ng0ddSN5oo+
xyafw9NoD6l6/dR2sm23Y9DmTOgMykNWWOn1NkLmLQtdUgnzO3J67AoVw5nLPN+7Dgnl13gvzKq9
npi96BHYbMn6EVlzLa9Vci/urzTuyELRY5WmaFpXo/fKRCqY4OvPGciIi9Pps6wPDgUv91ANns6O
TIHlTLxJoVxbIG9MZKYJ788TWuwPmlxzjbLLedpUvnh5CFXko4/3lNntdACSkdh7eAyrxE862sm5
czbojz/L4nfkvc5ta4I03f+ro2uVg8yDpWKT6a86BlVqNO7oUg5ydGelLKNksJxQMSMJLyIr9r6l
ddyAzARedy1loOB895eLH8uNJ3O4qQq3tFrwInePCifgrsh0LI+Y9R56jG5R6ncvwrjKzo+BncpA
Raohdx/mGYAhX7IDfIFbzkYVqFcaMXpt6LDyXWmMXyvXXMFgDWf39uqOz8Zj/ydYFo2mXwxMi7yf
T4p7cCIR+Gu8vDJp4Zco+qa1DF1V6mGx3UPYAsvb40rqVvdA693IE/BbxumQlaE3B0G0I/af3EtT
wd/xUVIjIIhg2jCAwWvAWR41fF/lAQgVG/xmykkC1FbZIWa43k3wruh0xGO/iYiHTYRr3DGG9cji
LcGnjQvf1XVhOF4oIVKS5GM8VhjiNsOLpremqW1Mfgox/KjOX5cVbuLtYl1AF9FWHA5/NcVxWwdc
aw0JrnHXRTFfxpUFl5LlVDNxOD5RD1PtzCZK6FAo9hYTKhBQfY3oxRzlqKtoPK62Z2Ect2mnzDhi
GhDo3Hl5e2jizi2rOf6EBhrzTTAtNyhKh0XHBULVK3b5n6F2e4c6qCPnkEQ2jwoRxWZ4JOGFo9qs
uQeF0Vji/1MRhsg4LpBQRZjx7b/h+AC5+LDT81VB+e4Q69CD11AgTG1hVzCXUfQmrOY5ze1dZC6Y
CPRYlgx20pnUoCKyeEZeCDRx6VkLh4bjFRnZDxeqdPYsA7oKg+tRg1hAghn/GaSoggD4rqFmB25p
mIcqB0ajkPI1ITFkWwTsPGto+dNTikTwageTlNQVcbdmpezcs4oU/QoG7lJqJkpm+CDT/7zQlBfp
D/WwAzDoi+EN0PdjMHIo2smWB48vUG1pCQ0YuxGbWU2n2tRSKQ5xYTcq8biZ2Xo+e6+mHk4Ec4+Q
avD3rolJC96r8eZCH6MdqIBiQ3Im0KVfoegxRrxxmE8Nra+7SJz/wcV+FBWdRb92yg7OIUA/NEtc
yvWopnW4G1D8ohv+SAgkUkxpY68sqZEoTaiPDyFZ8lDgTawqOko0QCAKbykmrIbkwpwpxVs2jDYd
rIvWqaWFVthHLx/X6sn/eBd85avY4njilUYe+dIE5DF+x3qPt3Kghg6EQI+yDphTms/q9U+MGw==
`protect end_protected
