��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���d�v����0�i�=\��A��?��� (��1_B�f�	�Ѻ+|n��y��Q4�]�aY�����*2�y%����>��������K������ �
�D��z�z��C�y�B����
_�U��hkF<�~x�ܕ�c�ij��(�������̫�s���֊v�@���PRĎ�cj���3�Ŗ����i@�y�Yמ^���(:~�]�%]��u{����jA�
x��[�}�1W���)�e���`OI6��bDs��x��`؜c�Ǘ�Sø�8pY�m(��PqsQ8�(��x��+�|;a�N���Bn,���N	`�u���@�
�r��qJ��=���U���dH�TC�g�/]o5^��������:���L%ڐ�?}:�c���C ����CM0��?"1{5�wh>�M����.4>jZ.�l[?��sJ��㓥C��z�}�.m��!�p�� iU]���N���[x��W��ɣeӁL3Q�����l�##?
N��gӖh_{�oa�ž&��
���m���h���,��p�Of�Q����a�Y-�	�C�U#,�X�)�=�w��@�fN�&H�qF����%���s�$���(�g6Y)a T�gN��1g�
A��'1{��f�XW06F$��KQ���=��~�7ft�U��V�ǟ�x۾C�	��/�~vt�._��3��'��TI�!�s�u�����j�6&P�)mp��0�?��U�u�ߨB�.o���Y6N����AW��bֱ5X���k_�+����������/2��d2�̎{]G���x/��U�z�9���;��\{�W5̆�mq�x��>n������S ���9�T��,�:;iI��%zቾ2���l�����CA��ِ��'�o)��5�c� R���xmv��9�a�3O6U�l�&�0p�hy�j�
a�7"�[΁�䁟S�a�@5-�Q�0��I��9�'19�aNQ��G5�
\φIOB"aUa>����Ԕ�k��]���.i��
YP��F�h6���19Y��r� ��?������A��g7�����,������_��d= ��jf:�#�`�Q��g���;���2��H\�x�6�5��RKvৎp�k�@(��Hx����I"��d�9��0P�֍7s� �$m���O1^��1���Aɡ@���T���D'Y��K��;��3�?xA���*�f��l����|F�	OHhLan �ϜJ��h��zAQ���f=�6�Fh$rq��BdS!�ΜD8vV�L��;�qsjewS~g�t<X%u��+��ey�H}J$хuRĀL�|J�F�·ct�6Gه�/Vc�D'�J��s�>�|�ٕ���J����8�P�W~:�í���C���3L�9`��Q 6�h��Rϟ��W�QAl���j9�{@\�������T� �%u��L:R�����O��!�������%Ԍ�5
9Nz[������ڿD��h7܁Is3�ݺsǚ��]����'�X�%�$ �K���%*�Ϧ�B##}����E�=�ꁂ��eǩs=`����3{��'(�2R��%E|UT����:�����V�cӘ&�cEFe�?l�ֵ)�D~��H���� 2�����5���,�ܙ�����6_`���i�? ��:�W���ޒp� �wJ�mV �f��&d���'��յ@�_�R�$��zG�h�B�_�41�w���ȩ�>C�Q�71�Eӻ	E Xٻ�p�����U��ޓ�-�Q�}��0/B�H8�"�f�
�L��_s�Ͳ �QN�	I���JT��L�\���d�gyY̺Pd[�{������Agw:�CEa�m�e♐_�de�
�ѩ��!������ pѧ���=s�~U���5�?�D\�x�mɡD����j������kB���A�"b9�U���9�ΐ:p�������V�q-���_uC���sj46;%n�ٸ��8P��{�]**����;�)�׭����u���:���f���f#��{t^PI��>Q'��p�u��d�)���0!(DE�=GwWa4/�z���]��[�q�a���N3P���-��c�Ң������b
a5��^;J���[n�YC�����b <*A���O�'��@�.�&31�-�.�ҖG�oB�v����h����������1��n���SN�'$Y��$�\���E�E�pW@���'f���[�h�}�2m��I�{�C����]}*�;��W_u��L�zT5ac����2�I�"����5�Њ�n��F�ؽ��A	sj��9��W9/�Ҙ%ft��Ç���)�c���]��T��!iW���ks�k�Ɏ5��Ij����O�96��q��~^�C��V���f�r�l=��H��������=��Z��&�6�I��Q��K�C��G�u���ti���4���]����� Gs�X�o�uT� ���K�i0=��U�@h�_F>Je�,v�c+J�텀O���d�QUM~��(�h�S|G�N'+,Y8H�h+x+������C�r��5%����4���7�R����k��.�bQ��PG��S��QVT:���N�2��N�BM��H����lΖ6�����<�h�
�W�AG�Wm��z��_4�B���)��X;� K�"��Yrݘ����Uʿ�6��"&��Ѿb�ݎG1ՏE�e� ���{}m��|K<�Gqy�M�>!Sg�����c�X(��f�讑�g�~����a�0mPC�eO7�[��6����k���t\�a��5]*i`�wj���P����[ϡ8}|�W>b�+]hO���]�����V[
7*N�}�9��-$=��B������w�s�Np�t�S�[UV2��>hK�U�O�xg��N�⧕���z�1�v��OWY,>�`�ە��NI�uK��Թp��ԣ5�ϔcQB��vH�tY�W~}������g9���������V��W��LC��6U������y	y�~�Lt5�x�ɣ���zϏ7��y!�7�s�!٠���+$t�J���&�*�WI���g�؅�h_�1�,���߈ﲣ#�X1�����&�Q"�l]��� L��&Y� �g�Z�'@�<���c����ʆ��mح,!],��������-��ED�-~�]:h�[<���k�W���ژ�"�I�TawvA��8i�ؽ�*L����ʷ�%^f����R�����,T�J���f���`�ͪAc9�6��;���^�GǑ�{�,��O��)[  �?�o��N�v�RcS���p�0�������L��sT�����b�һ���DR��yb��xr�5NNjR
>��ȼ׼�B��o�vj	���&�x���vVP��5�S}�]h��w,k����� �?���C7���q߫!%�*_�_`0��"�iY_̮�|�����ξ;z�ѽ!�	C��e�����9"3��}������/%�;��#�u�!V	���'8�췚��Z�Q��[M� �Om6*��"Ꭻ�_.l	B-�􎍐��A���J��z�cW�46�+<fts̢3��������,���3֟,�Yr\|!��=/�y)��H�F��{�w�dlS#-ǽ���p�;��ʡW�V%�{+4�Y��@}�i�Ѡ�>����\wN�SDɮ�������&�"�JJ�{#r�)/�v��"�8I,&3(�$�ve��=���G]�E,+�P\D#��*�]�p��2LПȧe�[6���v����g�"#Y�Y�T�;�J��H���gv�f�ܗ�~E�L�RI�_m�u�"D*�yv���˟�(�ʠ��/z!����s��(�����.�f�l�5O�#N�o���ۘڪ�C�<J_�F����m�GZp	��9	P܅��,��<J��i/_�B�Z�Tq��&nPO)B�oI!t�5�����8Q'�4����W�#��K	_�u0�Pnl�8t	2���-�;�bֿVx7�ڷo����4B�ɔ*Y �Y�m5�Cc����O��;�p���za�3����pB)�wd2��)Q�,w��2�9���/"o��t&"�c��������eA�R-.\o�F��J���0�k<�Q���I����F���`������ $�(����8��4�TQ,a�*�cQzj�} 4|�>�ύ��0�WK&��C��|�zj�NϾ=�Z������呾
����2�_�����#a���/��l���-��X���(9aW�F�}"���]��S�2es2-�br��������,�l� m4R�Z���8� �D��p�
��d�j��*\��O�n��N@5��p4���
�Q��?6���%<��n]ꀕ�������->�Eހ&�-`TÈ���6����-t����QGz'K͂�9DM���3�=�{�B�p��(\�{#�c�,��(߼��
���D&���m߀v`-%v]�Z�Fk'KW��!�q����izQ�er�"}���5����7��aE�F>@��(Y<{DF�tҭ\ZIh?4$g��o��e r��8P�/�^����"*LВ��R��%�vӏ1�&��F���~�B�\2Q3},<���dh��ܲD&�en���&tW�o������\�$<Hf���1��S e09P߉�O�� ����"+�aO�*�.
�w�o8�/�O�Ro� �"��g$h+?�����U����7S��-��Ӽc#�Q���h<f�]_`�qc�Z�)duzߣ1-�����k:Y �RwU*��˃;���7
�d:}�ک	��HP��T�-ʍ�v��co��I������X�f�V����K��!%Q�X�t�W�/Y��Zb�6�ü��ȯ&��/:Uo+E4�cƣO�Y���۹���eͭ���τ�3n/h�k�=�
�r=%{�@���\�Z̎f�]�KiP��C^~�!4Gd����ӝ��2wk��ś�MiA���Z}N\"q\�g�gTn,�~e�`77 �3��2J�)�7̽�s�?��QKir!�q��
՚�Y�������9Q�d��KG��V���X��c�bI����9�ЖU\e�����F�n��G�r'LA���gL���碬;>���Y�Рh%F�%���й�4N�INs|�+��)��cf@��f�����@�q�)�S�0�|p6�w��ʄ�
o��gJ˿)��ccwNZ#���N/7���Mow��)j,p̸\��b�D���aJD�	f��e��:/M �9V0��q=���=?���Ǔ�-�q����9�`�űBeI�;�.W��-������5qwވ��Q��n�����ke�7B�^�X�:�q[fV�e�Z{��+ $��`7�!'H6���	O|���X�>h�Q��9 rr�M�o�^�,5��_B��!��mQ	�����+�&�X�+�R*�t�ϴ<T�(���vsr'dQgWϸ�8�a��['�t��D��İg�V�t\�.d-k�����]�P�����t�y06��sr�B��pL��f,�����T3�yƣM|����wY�=������{q��l���0~���>��H�G�Q��)�O��H���Y�&���g�Uq|�\]���
�o�%Eݾ��{����� ��Tv/)����dA�B�㒹�S8��p{)�V�-�����gSք[@�����J�T�r�����Ul����'��x9��}j�Ʀj:�r�T��	�c�b5���#A��cZ}0�Q09)S��һÊ�7�T��F�(+�>I���b�c�����5�����_��("�^�n��U7�����7�*/�[�˧�rL���?�EV�����)�@�"z�=z�B9e���<�A�������r7UPW�&{X4� ����Uj�����{�M��#�I�Ԏ6�8׫9��RA{@�{�`W�Ҍ �G`yҚ�-��['H��b<T�T	��r<}#m���ǰ%��C��B�E�GTa��Ʃ����q��Z%��l�3�2�F�h[m�I��{������p8۔��<_}�{P(M�QW�����s>��K2��f�s�w���1�n�0�����l������B=�=Z�k��hL!��]�YB����u�A��Si_q�R����4��jΚ�p�i=���6�T�EC�+�H֑t��@gW���"-�6��bV�;��"�ZЮ���s�@�VXm�Fb�Qy�����s�����ȧXL�H0or�-�����bq_;�ñ�kزv�#3�v�Ӟ��V�ҫX3i��fB*��M\댣��uj��k�c�a�����_ӌa�-�v����R�Y73O>$�
��,S�|����2�1o�>։Sq����|LO��vK�*�/a:ۙ�uߵ���c���ugV����Zz��y�׮���3���[�	B9	�K��^{<��8�7����L���1-HW�k�2��]ŋ���AB�p6���0$�y���UVM.�3���i��<�?�{��2��g�^�Z�����U��9��r�����~��A�c�Ò�u<�J����4�޼�M��t0-� �}���h���,|5i���OhNǓ�گi��P�	d���j�̧���G�&���^$@`@�-G�����`��Mq_zr4�\�ܹ�NL|��c���f	�0z`Ol==f�+M
���}�=D$O�Q.�Y.�xC�	8���&=���9���	� `/0�z��W�H������E	v���nq8�W@����w	͑�J�����y����7�HTa^���GͶ�[���ǽyfY��]�]��a�Kȅ��p���?	?Ħ�r��._6���ֹ�}p���s�~�^��t2���T��YC�������T4�Y��&/OW��s��36��$@���Q�p�д���]�_�KZ�(�ATm��:V�s��ġIL��A�p�u�)5�!џ˹j1��[#� z�z��gv��a��4�a�2�%��H}4A����8f�g�1b�_ϧ�ɔ�!_�%T<v�֧�_?pdoo�M���C���#3#��Y;sv�e,�2��ج�
m�=�5'�S�����$;
�'�Ӯ��<m�+�!�I>��9pj�0�|�F܋ �0��`T; ���L1�c1�Gsh�$��UX��H�������eU�n�L���g���P�^��9]�4������[};gay"xW�r-L��>�����I(.���'/����SO�� B�_�x<�:C�gEvS�@�Z9֔�N�@���C[�z��%
��8����@�|�PP��!3�YΗ�a��R�Y�Hy�w�_���	$mY�q�bi"~[�f:��Gt3�lz
�����SaM�ʨ&?U�:���G�[K��K�sXQ�1����Z~ R+��m>
m�,6����� ��p��+T̿3F�2*B�U}u�;�S�XE���m��/ɖ5��MK��6b%�K�[x�_�&,�������N��Jd"}�E�X�V݋�y������H���	�J5V���{	���+�8;c�b�h� L�Kk��F9è.��Ve��ߔ���
�w�6/��ЋQ��L�T�"�B4`&"���mÊ:g�O�����=7Po�e��h�.�u�u+[i�F�W))�ug���~o�[��������p$�k��g
O��F�`M)i1��2����W�>��!�Hȫ�p�V�Hc����	ك�Ӟșe�x���-�u��d5�kI��ae樬��6�]oĳ��@FFΖZ/_�_M�N�{S� ����f��zR�f�"ek�w�VRi>��A���������-@6���4^��16�`�*�5�M;��\v�}�	@\�`��3$_�HmS��L�&�%s�Ĥ��?:��c��Ў����?@���Ƅ��U��?��>'��-�E�f��W��tt��_�
��8���$ �����e<%�Y0 7`�D��@�N��.y��kzP�w	����5L$AE������I�9�,��df@-��'�W�%>�3���v4w�S��{��d�{Z�1��L�T���DJ��0��&�5��h���T!%ڻ	�=�W&��������3d��߶~�g�+�ܣ澞kbg�!'��|/	<T�!����[-�pB��x�3�|1�z�YY��6���)�"�b���b׬��L�0<p����e\�|�%J����0���������p'b�-�`�P��m�aj�+~��#<� L�G�3	�Wu'@��a[S|��ր�Rcv�W�ak焘�7��/�ȩ\����N��˖��`�aa�ٿ�˟�p� �_X�ສn�3��|5L��'��� �`�!���?͓�ce�UB�}��M&�:�뇚��O����o p��P6� �ۢ�����?��b�ˆLr���
j�fS%F��7�����o�I�?Gvѕu�P���p7�u gF"�)w7S�{�^,�d�N� �<����}�\S���e#�~��>+���;�R&�,g,���#��dq�|j�uQ�VzG��Km驠{�f�E��:(\�r�ip}����=���eo��!6����K�������_Y�5<��7����'2��]����E� �~9T��p��%!����U+�9l�#P�ڹ�%l�MJ�HpG���;�{�23F�h:�1��y	�󸧁���m�b}>ZJ�����g/��y]�k��tk�'�B9��}uA���2��U�S�.� d7F�o��� ��Ļ	/մ�n�8��0N�B�6��Os�gpNс�(��$��sg�s����oƿr7�km>�B����ܯ�Y<L�\�?pg�sQqː�NW3��J�c�DB�y'�V�E�m���"��-��Tȃ��?���;*Y�ٺ4�ד�ֶ���0U��޲8��G*m��ka�|�U-"o�e	uHPE�\��%'A����F1�W�1O���n���ʩo���7[>�7d�0��ח��T������h��U���
�,�����7��p4*R>�Ce�/�I!ǰ��lAy���KDTH6y���
'��i���%�>�
E[��0�5�=�$�w����zQ�0�2H�-{�a�Ʀ��0Q�2��I@0�C��@`�§���>��p�6���������� :�C�S����|�7���Բ8S]�_���[��Ƈ�qO�*��u��l�P��U�
nƣ�N��ɸ�?�'��v{�r����ᓊE*x8f���:	�Xq�>eaI��#;��T"!�d������S��95c5)d�v5����%���!��)$�}T�Z�;:�n�þ.�<:'��չ���>��So�bCV�`�'�7\����1��
�d^v�rG�����C��!�-/|�Üi�y4�ƅır{��G�7���;�ՆVO��P��PL��ʻ/��ʁ�u��m�l������i���E{}�3�O�B��mP��,w#�]I_·���.ֽL؁;X3%��e@B�2���&���S�3�2)�$M��vў|b�b%R���������\=�����t���-�xc��^j��Z!D�bӌ!��*��$��
a^^�Ik/(\o�"V��cĞu�#㺢ƍ�T[D	4K�I�J�}	=^�A�o�~�2`�M8B�k�^����7� ����'DƮ�`hNԜ��}+�D�W�'Y��[�	��O�#�lm�u=Ͷ��r\�Gǰ�3����� ]o���ϟ����Z�����ǧ�t����4�#��<G��'�E[�Y���~Z�aX^�*�y�zA$d8`*y���"�+.��!�SW��%fU��?HqT��t��'7��}{1�bU������K�$�6Uek�����2��z ��lnZĐ����M�R�5�A��#���K%0Ƥѭ��2�s'��J'�}|����y��@u� ָ��i�^-���F"��� ��i6.H��#L�g�-[i�"F]�YuZ��W������%��3�6�w?�rW�!�S�I�_���p�v	а45��p�*>z��ϻlcQp��2K���˰N�@$]�%�$�������h5�&T2�}�5I����&�� ��{~sl+��۟ш	�Jhu!�������0��2,���a<.z�8<`��{=1N}���{g����Y^B��520�$ȓK2~ީ�n} V���#_&�G�N�3p}����#H��A�G]�Id���DB'�Or��9;IQ-C�}�T�dnOжU$u7�o��:��ڦ�h�a�1,\8�69ݝ6�2��_����}�{�]E-d�K�*���o��\ĉh3�Gq9='���r�I�O�{]z�5�[� ���f�,6}��6���`�B{�)e��?���7���������L91/�?u�0�.n��;C��ßZ=kG �H΢�~����Y�ɳG�z�bm�"�8��mƎ�0^����sG�Bd<�#��R���5:ED����s|�u�.�l!���-뱍о�� e�j��iy�]g7�w�����f{K9rcw��qaw�a��S|V�!ݔ�� ��0G<�C8�}��M���˛���؛AE�C����8�!t��`� sh� :�ȴ_Z�(�Ϡ|Tg|�� �����Bٹ���5��9�_Vƌ�[�,Ô�䯴�C&��eﮧq�O�$��ML?q6�r��Y� �7�'g�_#��@�f�i�����Ft� �R��os�id���ʝ48�X�k�W������F�a�C�f�a>�x�U2��߀Éq@���������b&�����N ��,f�q����G߿0[}nO����2���p�;��xk}r>>t��R��%a+�m���\U�37C�J#T����5�\1M���Px�n�* ��nV���n�j�p:�fY%���������nu�6A�������{ �wLn~Z,]5)h�PdA��U?-�8������T���73���f���#&�����ĚE�Co��c~=K���C���NQ�[������.������F�XH�VC?Z�o���;_��
�њ����1Ծ�;˹\jxY-!�F������4��,ʀw2&#�^:�u�V�{�+��҅UQ좥�{H��Q�Cp�v��v���G���/���S��J�c�����IjҲQ�=o�%���d������"��Y~���c�0��!5X�p�	CoFۨ~uIz*%��� �e�<��B�Qv���k[��d��Ax�+ � ҡ䊭�*`�>��|lDR�bYv��@!>���h���2ݼp��p���aVА���Cݪ��`���8	�p�_Wn���w�ъ��������b2�,7۩��$�+P����S��!��5�#H�0Nz��w���8�bͫ�E���]�5�&: �"��/�O1B2)`��{ű_N�S� ��1��b*�\?����D��X_z���J��e|ᘔ���l��_#�]�r��:�I^Z@�4P3kFH�Y��T��(-Ro �������i��y/}ȵݙ�>�G���m��)�x�vb�{�y���4�ݷ$//J'�oE�CE������
�۟���#�9 �0��+��+W��!Cj�� %�Jy������ŏ��`�f|祫|��Nլ1����M�'��T�MG�o��Z������|�ib-��?G���Bo�ǠC����E������*�r�n(��r�	/��X�$�T��ʀ��X�X4`�q��쩬m��X(|,^�(���	�xp%xV��}1�OR�q��2��%y��W[�^u�.~�Lx}/�U%M9_�a��ME���ON9�J�]2Џ�)�F�8��t��Ý)��4��V�T�1AB$g�@gz��	���
���ts�PL��6��C���cLݙ1��B?_G;l��=<<B�f�+�T�~����Mgg[���$�9_w���m�=I�,�����d�򬋳^�f�م�_������-��I6a�y�I:��t��۽�ʷ���Hm��H�~��5����	A�?�j*�B*Gݑ}��*<\���)4�`e��Q��^��{,�$q�?��CFx��ـ�m2:����0:mG��lY�'c�"��g�OP�����S�����[Ҝ?�#��㳒�L�H��x��s��wd��:���(����Z��L�:z����Z�:��VT�r*�V��t�#�=�����M.�\��לA�ҡX=jc:�hnq�f�ݾ��l��'`w��VBv���kWٝ�nk���ܾ̐�Yv��zy��L�˪���n�됍�9��ׄ�N�tC!�)�s��o��0��X=�c����:!V[�w�>�q��0\&%��xۯt��}�<��~4���%�G��������}Z�w6_�������eH��K�u��w#6�֖�쫅� V�Q�h��K��.��|�+0(5��)�(���<��֍���&e��ɱ	��<D/�kE���·I��+3�Y,���I�N��"�H5��K=��h��MY�T����((��=�d#��4����o���R� s�����I�P���F�){NP{��0`��g�]j����tg����|?&�[�f��<����Ag]�wt���Q�lxQ��FȬ=��I�FB=�{s�;��YV||xm�uԫ2:�97����`c�)H+'���V�f�qd�Q�T��
r��¦ev�u�w��X��Z[\T�p���PFGn_�NF�=����Y�Q ���.U7YFM���#��J$�X�oi�.�DVpl�����3�&�vf��0B'�w?��\e	�{��FT�����xD赽[$��^��;�y&�UC\��<{2��&��X`��]���]�<��
������M�o�����.���3=�G3��[�:�֔|�}���bC�0�/�"w�S�eT�?�;H��iě�W6Pt�㧬��n��a	�C������lVv�R.�
���.ᚓMj�	�2]�6_.�@_G N����"��(n�Q�?�]��`EQ���B�A�OI��Bȅ�D�;o��M��į'o��[=�G��'�tD�87����Z���|��l0�yVQO�jE��G&Y��2Jg&�h���O� ����8O^�)�!z+_�9!c:�o�jFd�Ts�!�X�Cp�hp]I����Rr����d|~˹�%#R���ĔWbę�V��@���'G��4�RT�¨�%q�,{�Cg�}���$̕3^ � �X�Q��ޢ���}o��.+��+�{_���܊���\������P����RY��tx�Ab�Gv1tGOl��:�eb��@2麲��!v.�ZU��Ͻbm6��]{Â}�]/`��݁U2�Ids��v~���p��b�y5������[�kC���e��O9�{ً�A�@En�ӊ�z�9��0A8eF��8�z����o����!��F�N|��1bzd\��}ݐ�8��	d�T~I9.��:�w0�r>7g^8ة�S� �����$`��6z�n�@M�v� ��<T���b����/�f�6-�dV|u��Ezc�-ݬ�b�P��GΓ�@������r���/,I&�5z���{�Qъr3�7�[��{Z��F���-Л�Ξy��S~��Z��U�24r$o�|l��rK!��Xl"ȱ����b۵���e�� �~�tU>��HK�r�T�wX�|D�� =���z�Fe��j�ܐ���|tanZ`�o�*\h�� U�/�p-�{l�ɠ��>J�f:%��tJ�;�W���ٴC���cr�Oh%e���{\��KW�u{��e�i��1:}8����C+U�<e~E�+Y��p�1�q���N����)3�*����i" "�Shy���Z��8�ˎ��'��Dȩ{AZފr�1#~e�r��w����g���'�fQ���U$��7��<`.�.����֙�7���"ñ<�ie����g��-.2~Lf�&V��؈�����h�@���M�{�)D��X��9PwX�#T#�Wa3��ݿ�"hќ�K��M����Y��:Q*��Ϻ;	)�j
n�66A�5���-���5<�8Z�r��윋��x#�N�������a�b
Xq�q�����_L�i�R�����ή>�dg�5�!r��3O�&��O�Q������!��֗Xn��J{tj�e�쟓K@H(,	 �&e;K'6/�_���
b<��x�W�F#*�-	u�X
c{��¾8�4�v*A7}0k��t_�M7x��r9bl����M�����s;#�@=�3=p*l�;X����X�L�i�tf�J_�k�r[��\Oi��`�&��@3�Gx����k�-�y��{[��<]�V?�>S���{��*q{��V��Nʡ���T �_	G8�[�̄%�_��t&z#�,BX~!���.mS?5yP�?��̻�Qqy�X>.4d�R��}P�br��!�����hG�ue�j�R��fERD�dL�@���;r�DZ/K�E���j���^Q��6���v´��).!��Ϫ�8ݿw��G����]w�@����V���x҈Ԗ	�1Iо�+h/*2��FڳF��k#�𦧡WDb�ۍ΅�",F0]/�d1���$�&:k�Kn�A��9��K��cCO�m�e~G��E��ȹr���b��!��M�˶ޝ�
�]g���m^�R�$�Tw�~��Y��(�xʫV�Q�j��&B
?yqQSQê�+�f{��WZg��Y��SOFt�*�h� ���K���U�H�ʜ& &{Π�-��e�)�kTO �a ��L)��`dI~�Oa&%J�������h!�eR�2ye��}Y�r
�>NEVY��\[@��-�Zp� �e����tn�j�Y*��� �ڼk{^ʐ��BI�Ĉ@��{<͗�����u�� �M�vI���C�!����]�N��~D[���y���Z�	mgK�P�u@�0�(6\3�`��6(�������oC�>�_�.c��E��ɾ?Y����m)h�����:c��*���
����qDr�PD��E�}������Љ�
�ce�xƱ�:6G��ʸNc���l"�����;���^pS�UC��i���ͲK�/p�&�}3j*% iy`����
�"j��:�	��zʨ/����R�&��/x�*|s0'�vF�
�df��K@!�[w�2m�!N��ﶺ:;���60�uD�����ܰ�x*��b�Y�2W�$�&�.�,'D<Ć7�^&��1�|9�ٕ��h0#�����{��{ju�Ԏ���t^*�����>b2����|؃��H�#�z�+��Z���;��N��3�����Z��ҴI�6��ϯ!T��LO+��=�&�4;���H%K�bA]������K�J��51��W:��T��aH�~�ͦ��\�j1�`��s={��a\�A��EĖ@��*�l������Mu,�i�:��3u����e�+'��y��
�0���^,��X�~�Ve����Nn�������k���i��Q��`��P� �G��M��$���#�Bi�Oʯ9I���/�ε/-
� %�L��`'j��pl�N@�Y�{�P�a����U<t�17�Mș
|*mY�]���+nD!�ܡ'n(���/��%1:��F&���V*h"Űp���yw8s�L(s>3V_���
�Yj'����BGD��c�(�$�~J��1zΩg�� �5�W{fFt�WG���u2Mה$�l?�ЫW ٱ�4s�b'�H�+����W��i'w]<�T�1[�[�O "3�T�$�rwa��-JT��<�J���/w����V�rW��BTyc�K���)E�#�ſ��'%@�&��Xi��{�i'�s�ݡ��k���[wq�e*'ǽ�؜M
���E[3�sٝ��[onf��Q8�v=��m�xQ�\v��H�K��$*���yrK���$�'F�ǁ�M<��{֑N�Dd�}�{~��kg�ܭ�1�c�n+�ߖtj���y��Cxe�ôFݦ��)��m�������IӅ��iV���W �ߦW��s��R����/0 ?O�L����dҷ�}~h1�̪���ě�R����}���O\	���nFb��B)���G�:�3x����TY�%�za�)1�o^�@���@�U�a�Z]+�1��*0���|c�F/�bq�\m�#�E��ޱ�9+
W��#o�Ҁ�b�E��27N�F"8��2�f�6��v���!U֟0@1 6�Џ��/����XD��7�N��ܓ�N (\-��Q�c��`��uܛ�et�fG�*g/Mw�'����z���4�Q�����P��4�b��|� ���a%{��1Q��ePn�ͣ7|�m]6�Mr�l$t�ו"�!���+�]���.�n�m��\)�%�aX`j�Z\i�_��Y����n���Xv`r�]�:��fJxF��p8M�k��;���߻��Z�[��R���{�f:ǃz}��P�O��8�wDZș��}�?���*���0��E&��3W����X�P��V��]�X� =S��e%HvQ�dˣ�2��%�';�q?��&�d�Ԑ��(����%`�_9�fr�ב���+�H �$N��e�V�ڛ����6���R>s����!H�C*��	ٌ�Y�b��~1��C�8�A�Z����҉�k}W��\�����%�v&�[~ǡw[�wĿ�^L��^���}�� l̜���S�fč!��	!�W�b���LΜ?\��ļ �_��A�B�N!H� 2_�@��u�7����l��A��B����Z,_,8��`��!hhA�jD���<�#�z0_A/�����61�>��>n]�硎2А�wHa��<�}ь�~�!Oԙ��<�����52�٬�ܝS!o��9���M|����^v�s�d��6��R��(��u�X��bv@!@�f�s�7Β���[f������x�+K��� @VN G?s �ArW(__��Ȕ+�-r.3�a>�>�
�����T��B�X��X=��5qL"5 ��K�&�@{�Ԅd�_�ҽ��W �y�����]�C�D�emOq�p�&l��7;�·!���q���8�;�]H)�J�/|pm^d��r7���=֏���b`ݰ�����^e�e���fЄ?�fBԤ*g� \��Yk�O�>v5Z���H��+�`�L�����׆<!s!.$�=���q\az�����ņ�ۈKIŌ����m�C����d�R?V�a� ��KW�4T�>�V��8Ä�˸��J��~<t�"��E�,��s����t�0�~hd�xc�\Ж�Q�(w�7�~�g��3x��y<�y�>���w��yѨ��P����)��QtD0z�a��8����Z:Z�)�c�a<�\(�c�����ߨn�m��g]��gV@�k��΂�[K羗#7�.����`��A�s��0��iƶm�hd��^��eܳ�Os��c�x*�x��p����s}���D��t����?�������Ŵb�v� ��-M�+9�L�#�q&6������V�\���M�q5��;FV]7��@SB�ƴ@1b�S��0��3),	0�	����m�;�k�D!�DJ6T/��NJȦ�}��GWG���÷����'[@�{~�t`�[I:A�Yƛ�j���	V�֝�dB��X
��{�F��2�
̅)jP4찿�۲%��[��g��,W�Sa$}^л9�I���.�t����b�|�s�F5Kd	/r�0��5 �!�Si'��Ǖ6)��u��]EO�P9>o�Ƶ(�I�s`�6�8��5IK�m�������zݪ����t~�.?��,��K�gU�ʭv�{�Z�E�B�@+ҙ
 �(m�5Ό靥�6�
�J�<��}�;F��?ä��"^�8�|9��D�$��u��<^�h��p,��Uq���Mذ=�BN9|�s*�˰��C�iK�ɓ"Mj�H��/���B�ʷ�	nq: ��:L�$�`��}����3@ػD̤�Vq1��r������4��f��R"�r+5>ݵ�(O��(�KҎӱ�;�e��m`��y.��Bdl�1Jnr�ط%�@R�Wr��y1C��E�k�~!����tRΩwI�N�"��G!>��Z�4K*����id��g4�wS���K����|qdi7H���2l�A��@'4ex;<�f���l�|�Y'-��X�ck;#edk.��7Y �;ELz�v�	�����ev#%3sQ���-?`YƢIt<:�S�ǘ��G���cw'hzд�-�L�w�<zr!�b�����o�i��`8�s]�S慘p�I��-�p�A��T_��U�dR+Bi�&�p7���j��c��� �)<�G�f<TƦ��������1L�C�Q���bՒZ7�VV���̵`�C�v����x�B�.�l˼�rc
�G��S��z �
$��o�"�yTϋp�Sc�����-��3E�S��6Dʰu#�Uh��u.��[�iU��V�j�x�>yl��Ld����wp_w�~"���N�x@�I��	��o�M\�m ����f�n�Ε�u�!�lr�&���ޜ)c���g����7��R�:��oz��I�i/�@��k�e�x+�L7��j�h�޺��F�������A�&�'�Ƈ�B\���4�	Cd#L�|�y��E^�RҚS�"o�
쁊_ʱ� ҷ����
�����y���/�%�^��f��ہn��Fᗪ�����.�I����=�~�v�z�|��Kk4�E��)fvڮ;�e�9������E� �D<��)������J֯3��^ej� ��(r���7m�Z��{��4y�������f����� *��
���6�),*w�G��"aC�YN��ZHGI�et+�+����I; NY�w22��=
�"��ƘsO��B&�T���{�fh5!�Qh�f���3	��6�k@ 6��r�[���9ӌ�T��-Ig�]�D6�G�^��IU���o[U`�ȼ�y��C˧AX_*-��ǌCZBv��5�@=>!�4a�>Vk��y,��;z�HL��<�Y����0�O�e��}��y���2�Y�m����k��3�1��9"�ws����J��k�NٲY?���T�2��8��M�����+�%}�<��$@�Zw�?�7�Ě�,W�:�����|�!0����<��	�L����٩ݍ-^��(X�W�^>4��#��hy��(y^��F��Sʍ|@X���֭�5J��+��OW)_���)�afa��J��;�'z>Ŭ>��\�d���o��?��ȫ5O��C��ywx1��6���Z��K�s`��8��9�ֽ+��)Y*'ӑXf3��p����ax��|�[�L`緾���?�P2�����_����B�i�Y*L9�������9a�6-4z�A�)̜F�M�m��tPI���3�s��o'G⎚#���X�u,�6��f�����|�J*�&l-�ꀽ(6�^)�j�Fd���6�����PnLrªS낀�u+�}��[��A`��� �2��	�Ԋ`�i��jXI-áK�9�\��NX&�q�ur��Y*U�?����_&C�2���5��<�(���s|�q`�����%g<�e
&�e���+q��Ol��v)Q�g
ǚ�17�1�.�0� ����|�р,N���烴��N䐀�ܩ_/�'�cX����p%�ٍ/f��,@�x2i�h�Ԃ��1��s�T���h��^p{�f��8�aulBh�D���q�
��-ь����$��c�'k��5!_�a�`�,��7�g��W�$��)ǻ0�Dsg�{W/��ct��{\ak��i��mn�=%���%f��,������1��=����yOa�b~��!O� -f�Sz[K�){R�p�O����Z(c�U�W�OJ�s��.�:%t����l�xk|��o�����{�{���0v����{��1d����gO`-�%4�FEw��S,*�a �S��{�}��ʄ�!a��|UuOWP�m�Y�� �҅.-�Y,��A&2S9����y�7q��5F0%��;]��p������xH8`2���sΨ�It���k
��!��	�����T���ݖ�XjQ���q"mt�6o�c(IX�A�/�=�}GՈ|ۭ��م�g�>�!�f���:�v��Y�p��n]�� PV_N�B�O�}A0�B���X�x`�s��H</��׫�[�(u�d��?���&a>y*��D|��>�2a�ƃ�+��I�z3����h�s�5F(t�j��3,�$���v�@�@�aN�zQ����{c�W���mm����;U���JnW�?���������w6e��W���t��r�.Y�A����?����Nn�ؚ��׆[X����\��_��^Ď% ��"*����;@�Y��1vݵ�@�GQ�ܗM�v��s?�a��-�`���b��s����(=���O`7����xR-Sv{�wye��������Ɵ*$���S�@G-W��kq�{.��?ZiZu4�y�k?��{��1�4,��*�o��\�V !�~�*��V1�p@�C�_d������#�S��5�(!�>q���A����ҁ�RB�v2�m�^I��ʐl� ���<����k~���r�Ds�~�T���BM��f57K��;�̤��t=7Ke��I����6�kw������W���7�%!f����4���-b�p
�+5�uS��qlB��9i��V��j�B S	s��
��������y��Lf=y��ߐ�Ҧ�����8�gN�^���t2�D���`����Z�7�*�o���w���M�;�"����S�:Au]B �;������Lc������6�>�ެ����:.>b⸿αǰ@�[�9���q����6g�
4�������	�WPi��,ɃZ[(&�f���rL������A.��6r�k�h둬�$!׆�9��J���w�;�ϕ�/yY��/ۦ&��FzT��o,<��X} �Y1����h}���E�"�-��D����L�r�$(9^�"������9`>G]���p�aI�O�%�~x#�q�#b����-c,\aM}ꠂ���X�)�g)U�Bh�]�/��{�c���b�i̛8���I`_�l+i02iH��b!���T� �F������Ŭ�!ju@Ge�7��>�>����m�܁�T�k�E�}��ŉ�M�C���}ݮ[�7t��;�b+�Ѩ��Mc���8�����޷q��WD'�A�i9��I��Q-�]�/7��zuO8�8��3܇Ї�e��K�l���
.�[�v˧�ۗ�n+/�H�S=����W�Fd:���r<��-LZ��%f�h��t��.91��� L�<VO�;�f����,e��7�D��kF*���?ini7q6��)�n��FWx��3��`=��F��O2{����N���g���,�MF���fj�Ӏ;\� ��$yQ��q͵W��5��]U���+�i��Uk+_���� �,��bG���©��^9R��ܰ���*a2l�}j��eH��@�p����Sײ厶<]Q�3B^|6��U��'- {�p���X��q�'�5�r�/���y� ��$~Y����o����Z;y���sM}BSȗv�\Q�Ş�2�Ѭ�t�ɪ)�?\��
��֙���6�ڍE #��N9�>b��>�E"��ܥ�x�~N�+���d\��DjA�6@$�0���"ʚ��eUi}��r��I� ��'ے&8i�}��,dJ����f#�JK6BR�5���!��3�.c��^��Q�C�����/����&�?�F�h�YQ��{�^>5|��_���tm!����A�ˆ똣�gK��K<&�!�VZ�����C�t�+E�M���A�S	�45]�쩥�Ӗ�U���<R��q9y���6b 5���T�1��=�°�8hҖ��=��R�H/^�7Cυ�W�	Hk��qv��}�	��X������7�[��<��v�5�'�n�jx�k�-�f��
eR�.��Q�rY8��f��{!�Ҋ�ܷ�-?��Fh3��% �v��,_ܑ�y}��Id�ت��B���b���a���4R�Gr�5�!7<����1ct0LF�]�|Ya)�?���Ys��faO\հǯ��^��q�o�c~ΖJ� c�K���U��4���:��U�-�	VL3�1��#��}L{���2��E�Q�{�����״���`�ާ��(t�!�U'���_�T�V;��g7�!}�VΔ��6Ү}67R$H9��CSQ����V]#w���z&��%�;�Ę�A0<�x2�!��?���S֍��A� 3�]>D/C:Y�~�?�HBX<�Nj�x���(ѓ_�f���b���cyT�ͅ�Շ��qE ���x畍j����E#Y>ѲHW ���������zV{sl������K��W�.n&2����:s�TI�[�_�4|LGJ�ǋ��+�Y���k��*�/Ë��v�@�Y��[�*��7K��@�=��Ҹ+�.��=yJM����x�K�>W)�}t�s�c.c��7�U�+AP��~jM�a��=}�� ���@>���eh�A^��k�8����� ���}#�Yc�1p�nK���C�H��-��u���l&������H�iV�&��3d�
�Ő4���b�솷�Uh�O, S�E���Y?���YJ�<�Z�L��ɟ�����묱l�a�O���2�5K6U�(��K�L�b�j:#�Ŏ?5��V��S�����#_�6u�ГoP�W�d;��S�9U?��8���`�9U�������<k����kT�j`W:q w!E���ڄჲ��֪���c ��
�]���T��+� ���Zy���`1�{á"nO{Ӗ�J��\����U6��2��뮸QrgT�X�5P^���aˢw�*U-P���s�l�?��X�'���Uc�'�)De��(��3��ؘ!03�UNf;����BT[��`G����KH�>�J�`��Y��F�ϰc���qF?j>�Ϲn�W�����l��+έ,w~r:-�&5{1�����wI8}6@ԧj���-�_�������r*�E
d��aA����ȿ��'z:��%}�h���{� m�
���F�C8uJ�fB��v� �[U5�~�k�����	��̽�)�D�m�@)iѸ)��c�v��2���#|�{�^�BAb�\�~���J�E�jMs�b��ơ^������i�z�ʴ��n�Ý�?FTM��G-V���i&���P�v�Y4+��$%xu�>D�р���|֛�v���g�)�{}a�uI_*Ä]l\\�,c�e�F�d ~Q�U�=z�����X.,��-�_7T)�̎��C��i�9���z&zu���|tT��E���%H��oF!�~r�P���j���^qI��R8</[�ֿsuT*ӅR�,�w�ց��G:i��F��^K�GB�c�)�,(푷���3�\�c5���'h^�$4�9��<]�{���?�u�hZb�!���y���S6wN^�ft-��NKݢ�X���2ͮ�AS��D2Zq~ꕘ�*���xW�|\����,�]�h_bR��~fk�=��T|��o�*��(�
-��v�Q�:_	��v\l[ag��X��/�632�����QI�+AF��1�������i�,O:0����?����"!Y,�/�x=4$/��U=9�@�OZ��|6��4[��h���\��f@���ߝ�	ߴ|�J�9��wgT����l�V��|4z8�כޛ�t[x}��p�)T�$f
��r���+�Sa1 �i]���!��0�M��5�cQ��t$qc e0�ȥ�X�d��i,�9��K����!MTfqa�P���׷]Q��C�v�ׁ�j���(,�yGA!�GD�.(��a��W�m2'w:��ߴ輢�^�����&����<1?l��^^k	�����
��#�;0zݬ
�.�|���G�������/�P�`F�A��W
�7'�C*ٷ��-��$|���<U���+��d=^W�&`/s�dl���3�(�9Wb@�3����b\`�!�ҽ��4�m%�0�KF�)'{"�����C!e
4nT�{1�]��h���*�]GP($�);G,C��[�aŁ�Po��ih�h���Oة��]�
�L�[�O��( ��V�L�F�l�(�g��Nb 5��\� ɀ���#P����OyT('�Ej�R<E�K�,0�Z#(5�$0F�����m�����V�!��QRM)����o�[Η�(��˛�q��*?*`_B����|9P1�w��r��U��`Q (���_QTz_)�b%)�NgV����g�u���e�d�9>�P�k�bؙB�N"�'�G��t�f_�`"��(���g�\'ꞌn^ex�9�]�7��t���"dD"�E��C��C�43���|��y�9���R �賎�8��͕ͭ�A8��f��v�[eh�j��O�oԸ��KW5r�#�"�AE[�:A�'}0�b�(x�j�Pa=!���Pl�k�S��o[H�M@��|�t+��Su��I�8�&�'���ٕ��3���W���nW��!�x:�C!8=�p@��`���>��a��,~:�{v�z��$Κ�>�@BbRw���?e\^%�n�S}/a����K~�dL����h�PF@�mg�ϣ;��$���F�k����j�����f��b�L0�Ci%�����Y�Q0�+3ڑ��}���҉�죖6�TߤE}\�S��f�����5�8�j��R����v˙��P��2�␆C�|�~:�#�$��K�X�`M\v�0�c��,��~y���b؟Z��'
�|<�*-t���AX�H�(@�Q�%�S|�����U����;����]���aTt�Q70�� ��������}��k> 9��'�ƞ�:y����f��_���������tF�2�y6y����2����0���x�ﳺ����M/5T�[ښ\㛙��TӖ��I�!]f���k[�uVʌe�c�''45ӭ�d�>��^*�R����ت[n�mw�9�iS�o�k;PL+�+�eE�����Hc���{�4�/[�� ��!�Dg��I5���v�@���c���Hp���ח�xd����H$,��JE��V�U�i��4O҄,�VL[��S-9��|�h��de�-u�w�BA�9z�,b���,����GJ�pQ�#eks�� �iєcghJ����҄�AXV" D?%$��d��'�u_���&��_K��Z��B�$�<��Θ����]=�b�>xEbA���'�{�J����H�W�K�� �ǟ�Gq�F%�F�2�t䚲�F?��n%���"��H�ɩ����O05�R�	^x�/����j2f{m�`p^O[�g���uL��/��*Ͼ>8��M��z��^@���#���G�|��`ld�̺���B���f���v2��(�� �$����cGuG�
Y��?+";���0�K�i�*�L�2���Dn���l��pRA)��2�֦J�SZ �}��{�USk���x�\���uɩܢ6��2��L�G�(�t�NT9���]�iG�cp�&Vn�q�x�ȸ(�Xޏy���Ͳx|���q#�]�=]����ȿ'�����I��^͏��������Z�@�>t�#w�Pm~��c�{{p�w�����)�����3!�j�{��V����l��f��M;�
�<N��5޹��*�-FЀ�*��ֶ�~�)�p#] ��AD���̒rj4�<����rI��]�I>BA���BӨ*�G:�"�D�$������(���#��o�2��X��k��HS��.��{Āܜʠ[�/Պ�2J�y
�nE��G�~���\:2�O���u\`���B.["�ID�.�'<>W.0�Tk�V{��[,=������ۂ�0]���-!<����
�Bt������Tm
�2�"�k�&]Ea�iL8�O��p�{4�`�63��?����j� �g�oLZU 0�M�4�l�Q}׶g����-�=��Dx��=ڳi�^`X	z`	9% ~l�G���VS�����W׾��O�Yz{Ji�\Ν>wG=�_8�3�9�S�`��� ��@32\�Z٬H�'�}s�f�RA�ʃ_�K��|:���k`���+�L.o#=<G��À1/'!��V���^d~#8;�0&0�[�o���ہ\J7<���e�2!&o���]���?������2҄8���7�.��1<�e�3����ǎk����MsJ@\�Qs���Ҏc�(d-4����
o��2���R{1���u��崪��MWp@&�A��"H$DVx�q�qz]AW����5�<`�5Qhr]i4�s�%<w��ܩ�����
�6%g�;�'g@���hڄo��/���:����3Ù�˶@��&���EO��	��@��Y���p>gc��5օ���l�}.%�&7�c}~�x/�}�-,u���1Ev?d�:9� ([gX���e�F!��r"��9�l|1q�� �m��� �!��g��f>��UyQz_��9�h鳧�e��ÿ��U�|ߐyy�Kµ�kåF����x�j�0	7�~l����6���iA;6��t����|��Ø!J]*����%�"p�dWSN-�:�?7ㆣ�޶�K��s��d���n�XDg휝