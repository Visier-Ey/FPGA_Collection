-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "N-2017.12-SP2-4 -- Oct 23, 2018"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
inArqV2ildHTOejhBLvPYNAWP9ZqTUCkCcI0n2QNYtysE3q/u/H1ZZItWx/8Dgdu
VU5dlFZdu/yG/1sG+bgH1xGyQ6NsQMvftlXog51HjNv3AWtC8vpMDlEwY2reuy0Z
IsAdSlvr9G5w10g320i0V4Xp8yhfIgF2tT+hpPhaP2Q=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 24080)
`protect data_block
p40dHYaA+X9OWW8lHfvkDNJrbXiemOr+/9eA8k9IT6Ar3WFgx15BS+JsWIhfx5x4
Q//S8dAQ09A3IQwmEYEs5Lmro4UBeMXOmXoTuWRW3tpaOiSN53I6ilHvYpF/ci2h
OrNmvLG666K28CWBaUwqkUOIl2MuvwV+/X9o/n+MBZKxN4JeiAUmng5M8GsszJu9
lUwZkwYokcAnOTEqxT43ktbLl20d3kjN+1tsdVpkrSGoPtLHV4hINfaJ2Kg22wqY
UnFsNI2atSgzituWaa+RzDaFD9cWhLI11lGtJlSVS3/on5o+IS+DeuzwbGJaE2F6
hEnXfP/bNyl+NrTpAZZIMt/AhLi2IjCOcmjffmuaOH781vvaPz04buD7iqmdY39k
pVjqgLJjqS2RX0MDJjDSNOTrTjwT30W3bLVRMbD/J6bQil/MW9lxPBp3YPuCNhTs
Cy0yoCDebYGsPrgm1gvEBQDqC9ZEYLmqU2dqzT3/8NaC5ipKbUCHcM3eLnDAXOb5
JUl3kNAkVHJJISG+aPfO0QX3N0RwhaybuLVrdnmXPoo9jH3Y9crBoJCS9ZPfFGdT
hwElQSegRZJQrE3bCDINttjVgxQbpD8ganh0v/HQQKMgo90yne7MluG7Lf5i1Z8f
DoPxXiAYoErSIELq+Wg6Ue7WBqtMtNNaWMYjNwbRHdt/H3fdcRAspAqm0uWxYCJ8
HMYHM/sGnjpvAaz3L/LXSKn9npuF4uyW89wHkIHDC7IEtWngH7CxP+BSzV+XaFVK
PQ2WaH9+9Bme6cr272SkKRhgqrgy6XSENoKPpLD48EuF6oWwDaBfdBo+GiV3ekkS
fB69HiKmtYStrdr5Ar04WK6gJinmc9GDWpIeVAvAMJ6Uhv7UFyJ8t6dzwVW34vDo
zt+yS73i1EWlp5IWb6vhiqEpHngWYBYOMScJU+MQ3Tiwfbj86ClUeqfQBtCNsdNL
k+jtGXlVXHrQaN4N9gNP+BzxqafYojQNIoMDxUb8KzHJu6JDTj3FG5dvSXwAwpKj
9UsxS+UcJgsMHaisibFN0GKTOjfqsIIMFKrYm3WqLioK6M4Y1cMBn1py7FZQtUy7
klB9kzLS1ISkZXpNu1+sdmvlbP8cbFfdY/R8oc958CJ2KLXLJIR/h+yohcoaPNq7
K7ZIG3711nfQpmqH/1x5UalxHFFDaedVOcGub4xdg8ifrPMYfmprvYOe85foOMEW
4TP0EYyKvhPhsMHe7PWR+i7dbkzlGSL7+iS1rt0PVADbhqbE0Y7vhTGclSEhGF2/
OoX3oOl+2CHXIgaiPTGakc5T2ZmCIQ/K6ZhErR6Siypnex1cmSeC2Fndqh7h3HOB
tS6sAVxU//KQRlNKAfvKRIOzm7VnpEptBr1+G29SGorql/4c2IyyDaHWXYh784Yq
rBjYvpvI795I0smAfz54c+F+sJMnPKtvLPoaFmCBdaBbvXUYihriz85OsUSon3IE
CnYrSnGXrVvMURO//B9t+EDfCRD0gCl8v0ZFKlzRTrTC+SGWJ58Whbcmj5/1RYkY
fQNvfCbNk6vwdbvzIi8TFCJdw16n3l8gdmYu0Dg18uYWAF3+hSCiXmxBm2yT94eP
uDkL6I3Eu9QLXSfwquJq+TINvPbxrpYlWLF7RSSB/1XeOpEFsO/CPzqlveJ1cuSb
Wd3tLK9FV8azWIhoYWIVNLBgpxk43MgSVwdv86vYjl4AfMVtJYWj1WZ6DyMUaVFg
GCSiyd1/mc4dQSYjg2tYkMjS/AGsNPO1iLLCRsjMsvau7fbBKH2Xm9rEaj7T7gJM
iByFw2eC2Kvx1ubun9VpJU62BM47GsJe6iFDgdG2SoCP2KVAcLMupJl8Ni3wG1Xo
hPf6AUjf5GKtHmX2H+CcgQhmFfy+0VLZTv9GJVyTZNrhSoIF8RssL5Du/5VfdgiC
VSnGJLc6yVEikhITv4ADNE9dzpQryK/K7WKCW2O3ggWUoMV0U55MFf3Jmjgpwm85
1gqzn97unXFGTksfNSPU2clLPqOIs8J5+e0RxYUFpQYWWhAFvB7G0X/fP2cqnpdf
RtW2kRfC+erACDlQgeioCwZ3P8lXiqBqr/K7mMFpapzwTXGlLZT4vxBBaeCucugg
hp/yabuQJTJkMIg2AtdmWYfIfHoBG298t6slLxVjVFIRuN6QuVb2lHttI6K2ZED3
BypldpVZpOIndGfuKlAyfhtWZb8IZQNUv0GlTP6DHS+ZMovGs0yxyMQUuicHIymb
/fUiBbhz5FIx4QdaD3dME+2DLb8ioRIGbyyiDubP9tG/z7Af3jSWEn1+Osf8U82V
qnU4yKpc3LsBHV6vp9T7/smBZGeV/I7ypmKKFZVqmdAUhJcqB4i/VXuQG/JEvFCL
EPHQk93tnXMRbeJP3+/p55AfLYDmDH9eHb0HJPDFEby+W4SOsbiu8G7+kDYqSlog
VSGj6uoGAersiieyVURcJ96n+0UesFPctIXQ+/gCLigk71om0HWKnNr5B9exaqwZ
xargpUT+khTl4Jed0AZGyHRM3yQm1uYRnj52LL9HWWQIsXQBdCmXav7LIMepT78X
4v36ROOZpe6eEgBVhQ8tbvsxFlnMhnRaR7zSQ2azGxvN8VAlBoT+SRzVqv7HA0mK
6kqbs1qivpl1DrHSB+X3RhDXXh6mcACQND/mQ+xRMNhiZZARiNXo7HgKFmvHc/oT
IuLHZSETkZafMuI39juVkwcCD76dKNWgU3Hot3rnhFgGeX6yI/SJ8NyCs/A+wd6l
3Hb2bVceCjaxVT2oA3ML2uP8YZ4rYsagJD6ZoykKrYrEZxWWiqEQpkPDg8s7khVS
zg3B6UeLdRfE3aa2ULsQqvB0nWZiFIyf18eerFuucHUXfQj4oRIHIzkhPSw9xQ8B
LqR1G+LVU6EtdugwJX7DvBs9uYE/C0nCwZm0i1e2kd4SOM2dH+uE/uHQAwPPm/hC
Qb1q9OlvvzGY+yYSa002NHIu0z91G4GLrJ4hDnp3+fQOPpQcIiyDxIJadFdG4drY
Nm/WeUpu9haIHNS9uT9jvqcznr7Njs0LHdItE6vAfpO8OzjLpmU9MeojBVf7HGAu
u03k2x/rFupzxPNLEise8Gr3Cax+BE3yDgETWDbWXSTkRxbZvh69Gj3PCHP0mLrV
oGAPtJtJa/VF+V5CtwAs3CRYMeBckQBPNdrU11VnotSMt9AvxUibAb0XQ7uxb6uq
az2/OqXpGu/Zhhkkdx146nHkoF46sCSXZZh8eKX862ixB59Sqw542C2mPt7WTOrP
74KAb9IvMh1dJhwgVc/nU3YSxb7HVZAj0T/dnoKMkDDOERFpiSxuKeyOajirKpub
wp9cBd+UoAs6zjrvUWds2/lixigGnbv2JkyYbM8vh8wfnuw2KtUzWO9HX5gbE6hl
MszQu1LAfTs9E/Lg2ta2BiQkUKu2+aVtlDDKqcY3UxrcWa2yp7SV8gKVKlmmpACC
V8gt48oYKx9i5633R+Q19e4A4yP9Jj4k7cVxqZgqpkODwZ5aQoXlD4XzKLju+H2A
oU5ekyg7WRZeB6MF/beXqyKnYXJUw78YmZjpn0ff6ZMNhfLIFV585hh5QpN+P9lj
JWvJaj6RWh6er68QxsUjVld28XCtrX39cSdvsqpiwYyhdfrrP4P2aTt3bMkarsTa
X/TqfFjAZ6Z9U1Qwi3sK9m+Vj8g2M1+atGBmQQ9WrxRud/7KPFrTaVlJiplfDzMZ
uHzQYryzLDWZrJMQ5W+9TmYNst7VUzlO12Ox8MTwPO53JZSPPPrnv4meUX+4YDlv
eLo+LwBwEHB+EoNCbZkeRngUWsl391b0X2glQfmEaQE7TXSIC+VzclkxPIaScsnD
XznLr5Y2YQPjUWYn20mnRLLZ8CVL0Fl5+VtF0mwpM4qNU1CIQT66uSARYB3EO26Q
YaVinH4VLSyNpS57sFUHxKL+fZV8ZJRiWFgLgarXjumi+x3SnsDpjavCne8yDGMD
x5yS2SZkikVgneUz0YMgu1ooBfyAVINUmQci40dT2y8AT3ALJUWb8GGBNRUaoSWN
edkVqwzRHRSdM25B1oy/D3/8s7fNRxBGXORluciVgABvLLt9hYRZBRrRJ1EUc2ww
Cse9ROcxPrB78AxZIST8Qtwc7g6LnBwXykieKIYiShFbRjzevTLqHU444BgI1TsZ
6A+wfhM/JqwhaFTPMAvT8MvTiOfWSoT9jZDNk0So3zJCjVtUVSay8mu1bFhYLhAp
1pkSSndwqSufZvUmSpRQ2xWJh53zO7rN5FlBTHTpFfEpjATJ4+HfWnulwS9SMUlF
hURE0Xdv88/mcarFotHwmJZeEhHqZEpb0lzNgPx0WzyusSaSDONQviYxxt/Dvnez
BvWjY1scHygXWMGJ0WPiLhZXftstxPo4PpV68OwMDxT/Z8LNr8t8Yu7Ta2qjBLQR
ZBKt12aKRkOwFGV9pfWy/Hya08R2XB4ZOV+/cYEZXbrJjaXv+bF+FohcYxNWa9+r
agsSvpPScqJX5lFJa7dHX1mIILptbriLUpXBVTXnk501hLuZPlfGnYwD6fiFf79T
6JJElH8jxWD4X3KxAsXL5opVXr83rIpK7V7igqZOQ6np5ONfkIbUm9V27Yxr63KZ
gbJrknlrptr9mn6UZUI382ptTUyji6cl11wsnyqtM+3/84GRTNbbqXMbR5Vf3/xk
pTqGHn8CuvGG69QnOwB2+aKYMrGs0ig0QTs6M/84qvgbN8beER4PBqcLES/YUmen
VQ2qh/DeCCN5UY5KvrE5RtD063/AJDoGbcFDlzPzNn+gJo+wWXaiTzJxhAhAOyHy
NNVW4xC8H2pjEpzKwYqUTZko/tUGt+w+bgJYw3vSJE+GX75Ov8LJAcWRdYJBGsRk
0fuACwQ+sh2KDYW9zX0YZEkkex+i0ykXiZSmXeS1TdD4+2paFK0beiXwdDQ7umZA
tEeuBznBwpTK/Z2If17nvHLTL+PaSyDUon3B+NiSJuBKb7h9lBx94x+LeEhf3YBy
QXSRYa8yQ6rFa7qF65U0qg4F0YvSYBvvybLCv/Kr6uE606uZrUi9b+6koBSGJ7L0
SI5xbdK7881T1HPMSo5tcGViL0fxx68IZGFfG3LpaCqebX+2IApJrKjmwcTl8Jj/
A9L4C0hykv0pRsplN2TVO6m3ZLIPjtfKti/2RcYQOV0yP/v/63VrHPMJDt/TAEaj
ATF+uFfVShWg26IOSIudrnHEDT1lnewV2RnmDvhxWT7329GOQh4N+x4f0M/PvvuN
W/o4VAAdKhn7qwJtnFLBR4S3DsGmacTLWlp/mWjn3GGNFrAVYBX6+YyZAaqIkWbY
R5zFl4p63FUZnhiMzh63Ci5PbXrYFd3XzReafIKibXNnuA+ls5lBJLfKr9JqrGRx
6Iv6zqg5JPaFgd0k/rMRMeoSGn+lGtqI2u7IqnWqeqfp/YHfp/4gVsfl7woHjKCK
MOvlQBrVIflWI9Tww1h28Ozx/jh7Xyg8YTqvN4WW7pGjEuWKsYYnuEbGiDyYVOUS
Ts1del05MvP87fEkRsF5k6HlRFinu4xeu8fugaJJ/OwfolDzD7yEv5gdKaoD2f/X
qrAG+c7ASYGfYlescErBub4DtRRlUO7z7fT8cGReFrW2L1y0fM5tU+FpTFuqP8ho
EXg97pyPy8DTp+cT6RzmvJEbBIwBMKbEjj8S3KJK3Ry7e8o8OKyn8LZ4D1+9oNsQ
u6hS1ZXhYijhBdtuP7qBI+TXKJ9R7lh0yMH4WFHJAm7XyxW28c0Wu8TbT60GjC+Z
8QpblFzfEs/aYCnAldv9EPas26ulFXbG0liBndrll/SEqCvvH28gOachNg2nc6Gh
j4Hl114ipQSxoYzCdBrjd1kqFBMv8p5QC8CcZvS71MzL06nFCPY58pBVzxSgePN3
tWYKBJBK9XaBdBTB6D9MdTtZ/8KGpk/lSMtCmC4yjPTqGPU9xMVbfycCWSbopQKE
AB8vPaRAoQuSnnIiI0N8uAypFifRfaGgmZUdqbPAmpLUYTiXMsrY2qPFMbxNXDiI
2ZOxvQG9K5d21mkCA1p1SnUPEg+nbmWoEHItHQ0UM0O0pY17Knf6j95VSIPvtkrv
NpD8H3BwMqsXpAb94spNxkQt26YvK8viCAo81AIuKQyPCy+a59/W8qkXq8aTYC5c
6lWp9yzIRI3JkGJRetKpEiufRryxkUVvKqnE3x1XbsTAsJk4SWaJ+sbFRlIyOKDP
NDQMOy/g6Kwc69EgtwVXcBHnNIL9DCVbRHU0IVGyY03FdeTYBmKCvOrZl0O5RKCr
uOnAotFzc1XAmbjGN+I+uOtAvzIyZQyQLsetwYs4jWtVhL++IhaI7dhWDZs8Jew/
2bpVCzOApw+eZ3ik/z8PMFFVKMTgMJ2CM9X1qbok4dYZM9gU4Q2RxcUGuHEIj+R8
XSUJZc5/pfNk0Mq1Z4bFBVK9ADgT6qWbc1vF4j7Paj1EEv+7R6B7r27OucAehySB
/irScGiejxET5H9cTan+fdTljpgfVsmRf9lXWMTZnjyGiywVQWFGreqm1Ec8O70H
tXSBmDWcyjkZiDdWENwTIbxh1AxhnfWCPphG9dfONIiaWRR5/GQCBR9T8esIojBt
rRlXdUhiA4zjo75zN5eAdG9I531Bq/r/nEoROVHt48WPJnV0zCQQwN5jFWd2MUxN
zFNh/5KIbGMXcjwtEMHKOeq7hMsa3ZRSDr09nNxHLddCCY9ShIFwrD+KM5qDNfDL
X4uanBU5nnd/RneZ8d/45exM0Pr9YS9ImsuPPq+nFzp4SJiTcGaVJzLUfw+LF21p
QIgXP91V8PCSIx/pmbWvdGxOPY6TDtN0Z0QMhqfOywzyo2I3UO+Mb1CWQiH2blr/
plGVZp6KYCvILY80Bec1tMd1BD7cqu3OWuqiV/BKjahoo8+tcYKW/4IRymYqoLkD
v3wavHCt73t+m1XNsyLCcBaR4eMY9+qsLI+lXUnX4wOGhA8MByed1H8hbVGpdkjX
GviN91zmJaFYsNpP9oh/wGqNpdc5oDwxd2JbOEHppkCJ6rlkA+D+UMA7sI+hN/hY
MIo/+IWPK4R0Fi2Bg60Z2P4kolgdjcvi/uWdBmj3NN5xVU28LG3Z7PCTQ2V6xhhD
cykSVigGNFzHgby1u8DzaXFXP1SwA35maEhQ82uV5aJD3T5MKZc9dBZ9fLMGD622
+uIIiNlk2gZ6g6+PuypDHMzVlDDUXCnyIgKSg4AcSbdYvn5a1K21raOLDsz9i0kh
I02ZVIVcQ7zixUhJLvGOXRJrOQ2I/wDlPyyoIJQAUM7RmjBSzjef5vFJObtFzUxd
tXeU4jB0T0lWPNqI8HFjYTDKv23kVrjzzaS43gA94EhxvjdIodoeiBRGf1F+HwqA
nHRr4jlIBNpyDFacCPTa2BGMZSJCOyZzCUP0g3Kv+RoXwa4hFvkEH/oklXJbLBCZ
Ao9Tc438IB5q5xh/6Fa+sDDobd9ng19qS0aljKFEJYqfaR69OqWdX0RmUOnbr/G1
DP3VHXTD5aAjmYnMU9ba6o0sNTSBsUAO2xiVrB9vE7eMBIyO5lG+uW2jC7BgoCYQ
JT9V/pw0OV1QASJalvIVBlptdSEKkom0NpLsfr5IzqELXiKPDEHmBQOOyFcywEfx
cUyzuQBA/6mGXOtFwdy0aTSXm1jXEUEaVFoZRAtbJF5JcPjrAIi4yk4bQgPgB2Nx
wF3Fo2kpeuEJlok041LwfTPPcmxl3guLQOfJY/5NY/yGeleuerpiSaHmXUkxMU/W
J0k34xy7EFQK4hTINizjY0/U+VRqrVep4OUibpMKSyO+uflR8ChfWdkUJLE9leex
zAeuCBPW7sCkRXSEdxFj2zrk34BH/CG7j6Hfj0iscLVpPNJ3hqBSYTI4Y0q+JxoR
XFrwxlEyNDldvKO8KSjiyDiBuK/XDu/Fa6WDRsX5O5aknjdR4y4+znbUk/Y3N6Qt
vaTOFhekqQ+8JvC9H4stsLfOgfLrLHnVY6D6JOR01HgLtWgEwKAUA+x6ubZ1weyc
ax81DnREws2vowMBi5lA4JA4Uf0CUi2bFTId+vjpvB/MMKZrEv1s1xiHdtUQGm0q
X0HVW4FvYgPrYHVXg5HtrW1uv3PaemDQCEZMGGOzca+L/MBhhHD0yuLSWGLGRv1b
0NnXDYWq8UdxGBmkzP/GD2S1fv/v9kec9j+ezvF9Q4rBJZYPVHjYwXBdbNdFEFVE
DevUCF7D7P8g6kSsRaEACbcVVzzRPN0Y0w1EHYM2so+5QsPK+4uY/fuPDNLnFAWr
B1cQ3fpAmNfdcWa5p8Wn61i9kbkw2AHyC/mWiFaKudlMvrv6l2iAsIF2EAjpWMtJ
mjuUTTV9rrmAyVnE4YZmG7Tw3xL+IL9ZAetKuTG/Qx8OXjqr4BqdKEPNncjlp/hu
ZGtgFI3tRh6IjtwehtgYMbnaVWblBAW6L/ERSH8PjKzF59TerTeb43f9g1EGe8Mn
bnHNvk4aPWKX5KSXU5IJh4F6jyD83X9SiRv8iDHYKcI1qqp5+KTmIayOyCM/R/ec
1QBWGO5Y+CkYf092afzJx+aYgGga5NvV5U9ElalxazwLN7olANUHyPRvmkMe6BE0
OVymg/5FDsw0KrQCHqUZ43sRCfL8HHMj8kZ7X+a9d9PM7HMlR8ivIgL9JFEBH7m6
uDVkjUjpPkaivw7g5Ho9WD1fX4O13AhbT2mFVXbik/Tz3mLqz1GyIC2OXzJVSJ0z
CrHZ7Htdvbar6lQwUaG3u7b0nk1Pm9GGRo4Sc3gM/gyzn0Vjj47Gcy7SdcQgTzKY
+ZfQz6cC7v12wbKhdUvS1Ium7HJ47iaBI7dmMxCWWBHnLSaPNVuk1ODRIUfFdifo
Tblv9BqYLpPFxWaXD6uwUGvdYkEIZc1ANGDNvyPqm8blEol8z7ysfBf49g0kGqD9
88rv9ZPj8ZsspzcmrZFAFG7Bxs9EjTxqJf+9pTUzYf8t7k6LCgny07iRS+idTn/h
dndw7yWdstqNXU7VM84ASPOUBPFNXHMJGkU6qL0ThQFtH1GiXCQlrvvuwbxsQhSM
FX3f5yk9Oxzih77yxfrKG5kfQ583ApBh5SY5ll9NXQBNUQP9JIi9cuk75IiDENtl
022dzbkKuXovjQRQMeYBdNxd0UKYA8LjPpBjiILiW0jfBbstLg1ELiMTIGztGVNJ
Njog2ga9oKxkpstlC5cOUXSrPeW0jzxhlvTWyWx10CUXN3hErTkhKx6kR8t4shQG
+/KhByiabE/JLW3j8EBDwM6abG0kJ9nz2kfNwIRixn5SgkCXJws1L90eFQnzc0WJ
hquo8U+WrZjYWJbQ0IM1vyEmsa/vV1+grIIMMc+LcebMnWKNof0WIIf8yQit8A0E
CesGP7h0gTMuoyXxmqOy+M0PvfhEeinwqV2V1xfLWn0WcdWNm5wBfUdVVbLWNgo3
VkypcWnF6fUg4sZnBx8r5Sr8JqkXNmsSsxba1GHg9Ox8KnsfSw5aS2XtIHHG3nUg
yO5vZJb8kHTDboBD2DLodCTUdp6MMvLv68W9Gigi90p8NRSYpRxKX+yZd2/5DLt2
OTvcIReg5h5bZAOyC0ya6mYJxhrW1dIS6LT3Hnta1pC72jXLoXfDKzgapBAOBAvT
7qFJZEGlGBzyvcP39dLveRkJe9VVk8Ff43Smeankd6MD7wWa66f+ClCJDU4OI4rO
5U545btrqmYFXXLkMpMPXlfe7QAofEGtZl+xBrMIYbNnaPMINFH1jQRyhHhYKPCv
SjgbeZM8gMUe/gCRDcYjVkuAqGmw01AwgcJnKxH4I6ZGjIcI5L2i0FIg/ia0vyuB
kV6FNKdXgjAbipTwyg5ZzgqHqwah0Pr90gqx1tN8hu8LVqhvzTRrLa3hHLX8vEPq
Fgd0Ef3rNwPIJ5pgJ4TsYH5WfG2ZDaTRy5fG/O5i0+BBsDgAmiZZvApPeIRd03Y2
/Xpe0w28zwKFPGgMDJTuT1uqvKDeyhm/Ef6sfB3POlK7lDhznP0jCl2yhFITC8SK
cBj3nTDvA0SbU8jwbI6gG1uv+mgY+AqV/xVZ131keSiGTENq3L6yPSJRA435/YYK
a/k18lyr/Xhmnog1vzKc/TlfKLvf+hMHkYtkOW4gQrbomSMNUPCXHenQtkUHBsq6
rpl5uj4v36tGGVB1uCLWZlC3I9/3sIeCdARV3U6Zg6td37r/6JW9tuUvuzVidiX/
PpuPHLhFMfboJTZlaOzw6G1QqrzyyZBY0Cfd9BomV3ux8gqytOGsnlzrDuplcp63
cN+4AbIn6Sn14iLr5Ystwp/U3YaOEssgAl37wKN2TH6awq0MCJuJMk5xgBzMyqPb
wqnP//We8DJ3gF07c4kjvbl9ac+qur94quyeDCK6DuU64x4uP8H8Op+UmrD2lzyq
la3lEqcfWdMG0TXaJ2N3geQ1FgK6hqCtUL2DVaoWTscndoSNJPBM7/X0lz8P+6S2
26z/JUDKXIgVROwLVRmaC52in9fLs9Bh4MXOWq8NP/seCfKZEjm8SyFe5IPOhY3y
EKO3gEpTKU2MqdkW70vtqT58kVKOB8WEjdOEv3C1+gtMxc16MqqYp2PuBIGQW8vc
WpLGegcGyZVF1fzT2tQBLTnvJ985B+lip6N2MNqy0JEiR3SHr+4Yg6i+7//tPRES
mceNg+8yyCqmK/mHfah0UbmgSTTrd5NGMIP85+zHFdEyXH1IoUqjHv4tjuoB/4Nz
2KoNcLUHLg3CGK7mNxjELAyH9R6v5YmMjQTDy+fnt70btfud9SeXWf7JIPTQ4LRC
KC8JT0/wOdBdZoEQ9y018+MBUasUkJ998Y+fFH7vLM6qz1K3zpOsNYBEUu2hkWDf
XXjjyj21P3y+i6tzF9/se/TEHEyrXMMkoODA/d/Jlepz4w3bDG6vdSG8WzTOsEff
7dHLvzakdL3fDmjqzOT0gYeFkBdSjfulyR8Oc4fXMNpgs8S9qYTpX4C6gYqv8NFU
fLK7bQZnvztnOHr9vgbwPwOmBEeOmgeA1YzFCf/6xBljxHdmqs7C1VoWt+oTrojE
Eo+9CnnFwGTM64m4WdivKWKFyRUJGgAfm2HZEyo6ZRnjbTn5sAYFlMet9UsaKoAC
ZJh/4rBSztpDFmdjAMEgoyTZBlnZhUYjo/EYeDoHcAbBjivupVOqOX6I2AL7SvXk
4PfzYrEuhvGmu6OG2EZuIYHv5s3Xil4tzf1YWEWAvq/reL8aM+4CAM+wAfBseMdN
fDFVym3MSu4EqUXfNAaQPtjCBdDGRiZ2a7qAR/eJKO4So5xsmNHFbYp8+l24TBjC
npBULPKyeTyOueIbNzObN/+AJ6uhHe10MyiGeTvXBpqFW8IoyE/sHxP9byGwkUsD
jPYzw5SUuPWB9EZf4gaYb5125LPjDiIRG/byNK39qmdlU7BU55WMpeVIHJ3hhqgF
KStgWkTEgllI3/LeDR0SVrSOwpi1iW7RQ479B0vyH4O25T5B19PMR7Lx4awVhyWV
8Q2pLT3dASleKHbkJPKbgTHPT307cjmmPzDhAmtdL/MEJ0m7MRq4I/j7wkXH0T+d
gnIl3gLDrfTMi7GcJz0B912Fh0mkFXHg94MuMFDXgM4CNe2T3C4fKWfWZOJL5BB/
l+3/8kZ9wdD5RWWVkzaWSx0KFGjBrNOOk6odsW8u3ER2A0baaLZw2J+NySmGMG+H
PzoCvL0swRu+CZ4sesOIh9lY94y8hYZuLaM/S2VdrimL7UuvcaqiDKT0QKBS5NfG
f7onKFh70kEZkx3DqK965a+2lXwjkHriiodSVLLamm71JlUFBLzaFZ0i05/ORx5L
SlJBONKDUw/f3NUrH3vvA7eh7odN9CBKSLH9Q1AMpvAe6h/jcwp8LoSVZCV3edKd
v5zWbsLZ1gXEzcUwlWMGcUCdFHE3R5actFf0wQWn+Mbdsl3ZSdP/+B5cfdi+lu1X
8ZRao6FWQsHFLjxSLG4NL01h18D9YsoXIRXtQSdgKnWf2dVwi/ZXARuOLuy6wAF4
RlnZJMqtHPDHkb/tMsULGya6hwKbEgZigSh/xFGsGTV4L2L4aIHk2x0TN4Q4htC4
dgkAGY8PeWHsmIicXXO16iyj4/qbNK3t4DpJd/dfsWHlGfVPlLhtEU952NjSuwLY
5fUntg5fXT9h6Og4zQfQoKInTsNRbcDqgXaNiejjd0lLoeoqaSZEc2qBPcpDsQ1v
khQ1WMmzsPMD2jJdXQrsUfinJLkzm0dJ6SUkxH0y1zQXTjRDz13wEQdLw1VOP9mY
Y8V2+7EKeT2teIg9rLdHOuNA8HSuHDjq/pAhmBS3IswFC3L3R8o0lXYvpBgZ0s/Q
jOx2mEMoRGedM5ZctGc4oi+Rsf/Ydznd20N/dk2n51T0a2ahDU/jUO1N2py4+Czp
w3SlMdj34GuS6TOpk+LXR/Fx6pgG20srY8eZG949vg7vLk2Aojh55PHmlAQglyPE
RYwtNZhE1X5MM9N//NuCeqrilDaHQFR0HV2LAZsan7Qaam+Pkm9gi8+B50h8h5/2
SjQYLBksOUGc+DOuu7+QM8wbMO1xBZfOJ6UpRiaZhy03wJGEZBfFFeV1AUZjfr6E
+sYFe9fysVx/dQSsLmoRLOoRr9+XnEWt3NA39LBxCA/dvK9OoiqWgxvgxIGEh6tn
sgP+rCn1MIGqYh2Zcr7oic3B9zKqstxqtvhYmWmzEcgocM3kQByE00wR05KJ68LZ
FDwkSyDbENJYbiVkQOJGAVDAOTh0HUGRXn3RaNie+In82j/GK0Q7cTY/l4/Zq9kE
Wp5IvjX0AI2HhyIvNLDO5C7MByS50NqbDGB6ND4amX8aG2k0YmBz8z4ROpblxJvD
WzYUz090ajt2eEYmgsa+o5tANUymDUMfguc+VtOUwU73ow3VIlKv6IncNjruI6AY
p3Z0FCwntpJC0yiwPzp5esGNCsEzRRWJimlkbXlY0Ql9nRgAgPDUXiVfVHEyIqnw
ib8CzYGyQu1GlafJdxsDHEejsLbevoohjaQtRdlN+3fq0HqFrvZUkxahyKkzEZKj
pNV/0fjSGOWxvXgMY4uVuQAeJwyBst+oAkHlsVAH+nrFCP9CGhHguot/1eJVCucx
zuxsNe4dqui8r0E95PRM4oiG0YR0zu4i9MlVLc4V8tZseEZIsS4TvnGRt4ObZ+uK
tRNtY32KIkkvCihVJHzjYh2U0V802L/v2fL6a0v5yNe6ZyD2YqW6EwJSulwROOOi
v0Z2XS0U01Er/fSJhLWDTS7Yv0EUt49OTM3TB5ck9k+6/IdmLkbB7zjAReMzVX68
Kt+dosQSNQKrk2wKIjFsFYWWOoxdD82isxS4m+BH82TzBtJ+b5OD3kCuOaeInUD6
/6KL6qJeurMUUH9KbDmmzo4KCIlsH9V+uSPqtd8s4QV/8ZIAj/lK0XZVVS8sVQZ7
stmMCcvaPYoAUAUWSK3zKxykIvynvHyciAuZxcnSJcUbXiF+VRRgJ0DgOwBn8Gpa
osa2O7uPJVTNdMlq6hVK7cnctUxyguYzZO0RUPeMNJTcQ9eGDl98gME1ZkqBixzw
2iT3LnT2gKcraBxYHaM2M1MccGxfwBh8pccTspkZsBM+8+lG9b2RZpnSeaNANJqt
w1exne+9DnOGkPCeCuM4Hn1xF0rHB96/HPaSN7QUouy3LJZlxdqmbWeUJuIzQ/g2
Qg80ubs6FW1Fa0sT7mCErpJUGsu8Qr17jm8KRlDab1/3sJ5s1bEXFugho/lpJi0w
2cONgdlQ0aAKj+4F9ax8KiKTwoOZBbTtAPAtRZAenWpYo4ROsi2kskZpd824PBdM
sQzQbOXC7qe0xWY7l9gvIeNlZJcUVllMSz7l8rU7pChmbGHZwFtvVUo7COUgw/c9
lwpbdhJE5QFySiY8uBkl+KpZy/sOyrxk4hBUg7Dgc3RXjcJE5c8WCCdKzsRlSwH3
9sKpTN/I32mhUufOtgOlMGpXP9Vs4GKJqW5I61Ksqn9e2ha70zwjRpsnSGkcHhLy
MxGg2s3u1PJ2ZALqmMcEifs45kh6EDkz6TvddZb643wdnVRaIxAhbibebDDSpQjK
SwhHpHE8SGHCHfTtbBWII95qtcYALOjPjR+xJE/DKJ9I/rsAI/QhDKQ/n1butxxF
xqC64DM3nIxmegG9tSUhN6xQWQmYwhG/mceygqqnvaggpCCUKi+ne9yDv/KizZaH
7t3aeIaDSKsLzLV1u5R2N2OmBrpfqJrUZDfjt9eqdz/oboS9K/m0yZzEgLNHT0b2
c8HzRWkFoGhphngHFDUQpkJ2yrCAIM7m5gN1pfEFv8mMsIoU8dkuDcIuUVp/yxqO
lVCxdpw3lc54IT+SBrAEul2n76zYO32W+9ES6edIk6Hf2yG4s+kvqf4/tK7+xt3o
NF20eUqATUc0oC55vcx6Vvyxxppc2aqArkOT97/NP68PYgVcXbGZLxhRebBGtXtS
lIcxnAxDvrk6hbsqiUmRwwTj9LN055R5YDDRbLcz7NnjSPE96wIAM5Om2fOSQhpt
p3fD8nyIlBAjGW6y0uriSYTfSroWmFpEk/AKsKkJ2KJhbncM7H3WPzsB8SCgwABy
51SZgdxJs6jlKKb5abXgbLHDo+dRG+sFHd63ezwYIC9iLSPWF0Ml4xtjozlhGDAg
z/12zjOJpl0/UsEDkLojDFOSCOP5m3fttP0DwGxaBlh2sBFSQLRDIKnkkmPZNB2A
rbBIxKgDH1YVsTqR8fTaOyqNpcAlV1xrUEkQeo3Kvc0fCqgKfLNBEO9F70rZd+YC
MAnu9B7/3iJCK+NMoSZXw81ChSU0+9gpS0BUXvuOAqPDo15m1iwZjQFqyGXJvi+7
fVHoYd/kLn+OtVxXHA/K0pFAQqGeZK0n4Yzp4XWuAXT6f3dEO96o5wXh0N//bkCp
RAa/XquFs8Gr7gj/RY+G0RT6a9wAga5fSrGtW3RPaCZOUI7KOco8tC53yCqInuig
rd7v8uAJD2wXwJoMTMJsvG0YuilGNhnICy/iu47dCb6uHAFAzbTPQWPK14thHQLv
Oh8czaQc+QRBU5H8sGui2j8wEq5GdqJNyhag9/g5SSz5F3cHDVlRO4q10X8QYuQy
aYyTPSKG/3SeCK4ypg6vbSuZRKsMmJAsKuWBjhSFERb4NM32HmCAeK8Qxd0PAm7p
mkleJI6/NftESIIOgUFcpR8gPKU66LLDgtEPs16J9NQmv2zfFIuU38KVAgFL6RLK
jbtdiMRDXZjPgxMQ9sKUujuTxNrL1lLpXGYPCK1Ktw5zi4VTLlF0mAaUyhfS2VYx
wvO+DTkUtosQQdfaDpyp6Px9Qgi5/uDhuqYM1rvBPPwP28u/8+GzC3jeY+PgPRpr
YSs3mp/WcGIEtxfowqAGUH/hrIbQRqVNv0iw0iq2BB1uuN6vacbIbyawuqfWFJ54
QiCV34eFdEQwsuT77qxXz6unwfAGB64gwG3KXvFOG3/op1tlpBkyzwZszMy8KMsy
xKUlRkaTbvzQNjqN5pde+91xlErVWuuON08FevcMXg3GhMzZBsMMcJKrWnI+7kgE
39In/28qgGdrC0KEUr4Loq+WJiJVRmLMnbJ06F94qwKMd+K4DCinFTDEMc3FzEuV
dzw4MARiAk3+pdTt6HA5YcS30JjJcz5Kl3P1XTDKCWxSFE6peiZ8/a1DrPiRUkGY
kc9R/ULaD0zhJDHKcoVrX2f7qvDP4Yi32IEl2q/WeGj2zFLKggESiUDQsfRlc/AB
PJxP/xjq4LU6IPDMv9Dms2cGGKEkYGTtoOvBDQoavTrkaO1wSGnvYo2Y7gCH4bKl
5y7jC7Sv9UXzxEY5W69CTXervnvlXs62VUD9k2joz9hLbCqsgI8TuBiSqMcBYez1
7Y7ajsxy6jHNjReTRQOmaak5V+CqUAeICGriIkCX9HzMPU8vLthJn/DcIa5kKhoV
B+RbhUlfWL2XmYuc304CBBoGeB/qc9PytopZQz0z4dgWR+TLuG4P8a7RJHCAXJJ5
vpputjvgaYRnx3tIddLdtFpykSFduTdgZxzy6W9BySlTkMWx8EaOhscMyvB1ibSE
hfNRGXIVLKN+2S+XjWnsWPI1Yiu2KZahfEMlE1twQqu1EmPYc0BVsRZhl5UqQvVf
5lrCIooKf7YXWCEz5dL11JqvopJwQ3DuvnFi1GeIga6eZnhXewy/aljfxuPAj9vq
2ev6bMgpIuNPSG3kgv2acbU9Ws4y9aA32CGrbIBtYbDZWF3H/hNgMxS+KGHhcFEA
w+e3iuXOll3MUZBOuaZfLdjP1uCS+eTh26erhebDRqACPleaBV4rFdxa2otWDpEJ
rdB362YD+upWLijkMUn3swlc5lF5m6RL6qWvn/sscOxxYbfjSq9xrEYQcr/tbaVO
ODIMswMpOpjvGq4WKIRVKF9NiJIdFq8xZXhJ81mVSM5S3ZX9uEYI60lRcSK14gFX
oS1HacRvkWokZqqAgR0hFwdStaLiRDlNeP0ltim75im1MKOVrS3/7mfivfV7HgSY
QSFjm7c53Q0LYMukd5Oa9Sjnto4qXjPeLaSWVDkQiniDWh6M9e9cfJHQEayVD2ob
+vYn33MDUquHNS/0ZFGMORZZX9SVB/PYur12mEauNQxhBD3xXAliUb7aTdZug6Ne
krQTPXv2v2VP0oYMkPDe1CEe/HFCaipZAR1WkawI3m0QUAJrvQj2PXaiS9vF/Dql
UAZKgEeFWR4wqT5Ec1FLsW2GzQ3RUOrRjaqQjv+dmPoYZp9v+kI+C2Rx3lLev9Oc
8UwH28ILRTJNvJU5zNvLgqxzzdalgD2HXqy0Wpe9lsnRXmm6DX3q9uCa2XneCv0o
fLyj4ecJ92C85Yt7kXnbjZu+8I/ATaqRjm7HtDamnCKGJTwRtqvMubiljaCmHFSo
v9gxzhXMoxEPt+hvkByxS6lVRa8KewGU2WGa09+yTq6eStZzGV3f60yl/TcV7A19
5fU2yRO7lte0S8zrsBfKpiofRF06BQkYRTz4AzBK87YVpWizqqqjpRkL+ZZAXn1d
l0p7UbHmGizBo9wyEZseyG74BX6nHjwHMp25yUL8jOnaEkvlaMmD0EELGyYTxhqL
sZwNdS2K2/g47ZC9phRmegf8rqLf2cM9wnEgA1/8b5jbQXJISxDDfVZrTwBGjcR/
19kWh0rchK1KAiu8fHFEo35CpLt0I3sTgLKoR1OhSUl2om0sQS5wqQ6v1otsM3OD
m/1pZNNztyyZeCG34KRLxg3y2o20lzSX+yf2dGFIA/8vdQ+KOdD5YsGQJGDCzLTw
5D2jqnrHnUmyfyqljuabtvyT+r1vfcds13E8nF9+qlBr4/xPJ4HjR5fnS9ENYmHU
D9c0/SIV18RQ7Sl6UR1smmHvXmqD4afv/i8i5dZPjr8NzCxBqKYGCGp8lBhhpy18
Uwn/1tKtdCMvfNjcpngtTRBxHdgI60PUz6J8z0U27zqnf6SMuotTviERucSkETDO
T2Y1yr7hZ5LwKCafbPiCgU2uZ7gAPNJakeCVTxmVxPJ6P9LTESiLSRoxELC6Q0Ok
OZgtwuZqqXtXDUbl7b8OAv242HaDyhNeeXILQvqB/XsPImzTZFX24lkkDLBo+Me0
bl2t5bMfOWh1ilwYTwVA5eaaAe3T6KWRDlbNLN6pAPw0XZeuzUvhgorGAaUcfmUN
sA8hy6BqmCxBMtLF5jneZvgAPzi6PK3GCbVTPBEdQzzwQu1+vVgaMNViKr66v3tZ
P9Y/nnUp5/rX4srRYMq1DsVR29JUyqrqnr2C4Vl5cCgj4m0ejdRnRTesTo999Mz4
kYwLM0G87JUqZaRgxYcnbFouBRQsvy7XcrRp8kEq+PANDTPg5kF9Hq/81FPc2fU0
Jr9IqBSzv06t4ChlN7+gLqe/M0AQehGPb7iWaAs892z6LovqlG7HjoKSXSoL43QZ
tGjjj8XYcV075+mrM3sXPiEUgMZk45Rca9LNwoILytjF6qaYM6oFgrTSG5eaE9ie
uXcgtG3ZC4tEkgJf1hyK+ss8ArG3xGH6YxR7/BzK91JA5ULHKF2uL25RSHGyPa4I
/vlOPFze+MAa6LX47Ct1Pn915lBlNih6+23uhhba1cK2bNwVk6JMlEBZABOhrF2u
PwkNfjVMbx8/eM5RveoVoZgxejBTl6PxgOoenc2Jll7+rJDUVyVf620wYtL1nSZ8
VaBm5hHxvvIkhvr6BlFpkaVCwd8GdGYP4RAXke8uZjNqIjTSQiw9l5TCG7At0vcf
Y8GF58MXaafXm7TD5gyDMsn3ll2ZV2dWjvMubBRKclGPjONnLlWBVWxxQ1AUU/2y
rFiJR1pbAmnXoiT85JveZ9Z7gmEKuHI48wgYPEBTiHQuKOZmHkxGS9xJvuNMyyCA
r/XmYyJRCwHb+pIaAwgUcUZwFuhsiMZNUx7EH7iIjgsteY8OGXMSMKb5uWhrZOO3
2SqFKm1hHRaoA7dXovtML3Ljf0js3r3KNujUPKs6uGC8hhHgRAnIBAWfj8GfiQnx
II+lMtiQMDf1REZyJEexB44RaaRje4BGaXwhqivSvdUNnSdkk1I0G2CI6trPe92J
0dhwUqIEvYfw9/EQoPQ3fp63Xtg0Iq6rNfUcDDfoSnC8wHnLN2QZ8y7ldQWyhA7I
i+k4zXqX6fM6h97+4VlxW6FNFQxj8imBb9JOU0muphBkSxVR522BplDXAp0O3o14
YU9NQU42nHgzy/4H4rc+wvOhprMdhWaq7dVLUtMOS5m3O2TriZwr5Sfiisi5DqLg
hiWOOlgyrAn9pffcOjVKDJayj34i5mU2ZHsdez9tfIWSyqnGWsv/+ned1EWSPhXs
mHEXu1JuPPGJgoKZquwXUSypdCHERZfRVnRrYk3vdGehmhQl/xVGOAorB3ZaeXEV
P3Vk4HuyHxOEMqJk76b2cfcYI4wkLpoV+wO0epMZ4f+3An7Fk30GIsMPM7iF6kwt
QyJ1i/phdaxWgEe/7kHHAjZ/nHyVWPHmJVr+eq5ey7v9Pb5yhFIdJpYpMMOgubFc
vJJWmBSq07j3LhcPUKNrrnUii9xedQ6OdUrJvaQZkcvjUDo/CsKYE1lvqXyL1zKy
wjM3oQHD7OhUveiK+ob9iv7lJ0zK5hsGHZFVvgRWR85yF1XirB6Xj7OOFaqZ8uxz
jiEDuqwvv8q4CXmgPyhl4/zjPM1GWWnBu279elq+QpH21Mrc0/qzwoIhXoAyFmZw
rB2dMxczChF/pLrl+UUY4a2Q6rAmP5c2vjQYmvuawyR/B+CFZhOzJd1X9yOKqNgQ
xkg+xVXee7vvyVWTURFk+UckRDYkZhzxpQPPZpgDLUyrS9nfZLgl973EDnqX6ZvH
QUnb/mjtg7lp4lbY2ffZpwGuNr40qIZ1QB7S3PPjLUJz5PAYTmW/Air1TolGXpKs
Z15A750bTE584XJ0GFcajMzspIS0hWv7SiEdHy8CeIkXrKSBDfMpiCLtFYvoyI9M
9geQfymyJT8ntOZ+RrS+6OkBqZ/B2pGaV65GwWanzSr9RCs1kVgXP1frKclxEw4m
t3Zx+UYBk0j6dQ8y6ynoo0ojrHYJBciUROMmg9XGeS7yM444FseqqknvLVsyMZg7
mE3equIJm55tHdWqCMlvKxSS/5otqtmY/2OfazGdO3NZ5ldXblDZ3gY1tlMD9g+X
lRUyvykWSkgYzE0QUfE5qMS5Yp8PgsGTuB56tubHcsKuxU7iCNdeG3YWelfoVuLo
Gz2AwiSpS6/u0YLa4ekEBWzfjG+fmf1HBZw6IIKMJ9GERWoQGDc7uSVBuA900nGQ
SK/l7HTV+BlqXHONHwBeifPWs0hGYiC/DOW13Bha3Snp35oaBw79jv4aKrtVykww
idospJaoLZd0vyaIRhFoSScJ1fy0UGQtElxAfHrS9sOUjyujZ+upcAI8Jq+Xr1cH
kAZIEAF+2Wh0OeYey69ZTp/GAxAqxfkeLNBHV2dXWI7BsY+FzrHL3u+QDKJJzPIA
fgXlHiGH3yGzpMywOnbr/NlY7MJHQV8VmycNapDGW/nWaVAKGshcfGkMmuJU63nk
+b/L8O9GWhYxoIniugbvV8OlVkZXHoGOvXgp5tCdDFRAR9+4GclXw0NOgPVj77yh
86CdiQQd6MCTjEvKzznz9j+vGOIM1eo3l6y662MwnRUWuI4g1LReyAjFZd9v/Tey
NnMaucEteg2MO/lxARRPAp3UvdUXDkviIB37KxyOCxJXQVs8alYML49KTFFo75wl
AQKDaQI0fD2x6tNmSXydD0SDyiPndH5Mv7X7dqqwR/OI4JX7dz7vdcbQh+Z25q00
O0YakGcutT7SuJwvWjHMW1rA1nLi84TLrZ9DjHYTk0+m0NICk3YBS8ZibyPDCnvO
1vt+K/cU19HQwWovdZjcCj2RBPswtrX00L8V6HN5zO5a6HWmLcbgaggl3CB0wbOZ
vmhtOlms6zS/xh0WnEBNH0ST4x1nrrJt/K7taG2x3Z5nByOBOlsTN2B7QuiHS1m6
CsifPsqdY4lMikdLGnItvLwPA3aJCH60vG6vw2WniOS6YATW6SpGhZ7IDDz9UW7R
/cHzROFgP8WZwP4LhmcxWa6cyt2pxZcyYW2/vpMAEisxC0POSwYVwDXddCEiyrpG
XD8nYaEuEcqXK+Q4NWyRkaLJ1JneTgQTok3orfb8JnXWNusYtjKWSj1/O+ScNJLo
0yiw+p8FwAtDfbubaTHoIzGdBLcNZvvMyvC3sfnji+zPy5bmuPpT+eyd19piunkt
GhOWrj5uZU50CI31XE8WuG3iDfRSxkOdCMdfSVDdwxefTTKuazg/5VrlQsEYrTdm
uAPEzNSobUBodc7Gv7LkErtBGRaytxFonLi3KD4TkrXpbLDjgcdzrRrbLlJKLiHw
0Wvi9G4MN6JIPhw7KVDUMMjrzocfJBZZjgyyQIVWQeIsh/CDToItKE6BfeKUwpfT
BCysK9UOpSK7tzu65+LNZqy7/7mHdL/tpXiNxLMdPF60mkrO7MtNsWo6Dbc75SRr
CfEbGzrWb3ipgGXuWsGMLMA8hEBUIpvr/DUJEuOM8GcK1r7Rus0IkhwDr/d1plPD
acYYqXxaVoRiS6ExbJ/8f5WH3y/LXhSZ/B5RTnV5iYiLafpmqsoSShwMwFdQImy0
HLiFaNVOk/Rdz0HPC9iHfBafy24VYeLVwbc+zQFHnUvayQxCLxiODtq2Fc8gunHy
vCHHthYnees7UTS8YQOZNju1H6PR7T1dfzuKWbbYdx+5LdyF03QPR53imRle1Wzg
eHPfFnzliP5GipAwXtrqqBfWgfAttD7X0Gt0R/N62Vo+bg6/+K0T1J/zZRHIb/NW
c8GAymgAgOfTh5tYpNG0R6Z1MGBOrQcNOGsWEnl5Q3/RcCyK5ilqkiaEyVlNuWYa
7WqWLsNeie160Tf5URh4v9CZrY002kCWRWRXQ8Ehhl0gjau00xXJ1XA1u3irvwYh
k3Q2j7hBMXdj2cFWrDiSJ0kXBm/rvio0VsZTykC4kY6AAseSClKxtp0DmtFXExGO
9wJLrZYD4ylvbj3AjEE8KdcvMUmFgkgGxyzqYwRcoQXEiG/t0yvAywxqpvjP/glN
pR+rBXJ4vRogkeu8iuW3kLysNxqdN2JFdOGmt/7wqyKzn/Of5O4fmmKlGJ2tIZxi
E34KJ7EXrBz6+FWOVkMXbFWTPFySFxP8vhsrfVuPe2BheWh3jQkELLCsv6G6G73l
+mzWjtuRettUCsWfVtn2jsFsT865UAQivVIctKFeu4iuKGGVFtmc8vYzQxmKIW58
v8BMfZfwf4UrOTTYP25FsvwYm4esDMmDGm9xzvS96tNMS1tpXdbtqwbvUpEPkyvl
sO0HyGHolvtNBgMofagtiAlB21PC2dDdRg2RW5Ksyn2LH32LvncM2HRl8FEnNO0M
/zTvNquAFtZ7to+R+A3WpLj6nF6/sBVcH6iWEg4TKehx4B2jj7zsuxJIrhy+XXCv
fvC4Ks9/qRBHK0RLm76OtHynn1wfPkWqdTFn6PMfdovaGUowoyPzhGuBstgLpqlD
SY+ExP5EgzuKj2KLBPPBJr/5dj6iRcsF8Qz0S9fxveIc0jvy2+TEsypzomkTo48S
qZLH034/gILyM/KM6jSkf8HTSWbqZwhO1Qz2i/F6IrE2upuX21dKQ+ZO1sHktECO
5kS20AbylZK1dfskFoZGtT/kahQQAphE0qBYfutN8fk71R4VkUwb+BhQiCO4SxiR
U2gKjLQWvjtuUz3I4ZC+gLNunoOMkB+Et74mh02vRKH4uc6Ju47QHiEPdeQtOvzm
ldV3tLJgjV+doXgupf08CghkrqGtX8UW6aIwzBTHq/iAInBomDESrT5LaGkaVnRt
ngQyOypaDpMOn/WL/TKHqSoZ0hlzpbVOHzyeommQmh6Kny35WbhCdb+t+waNLFjN
7Cag6Cyd9QaDFmBUhrDWCaysimlVdCKKUkk41ulPjgt0TSR+T4uKbIBzuSMGQXED
dCa9KX8JrQX5gpbNhiX4bqgle7QtIeR2Ht84B8iN/xzkCDPJO8ObifkwsKHzqUzs
66ZYMjAbHxCkC9f8EIPT9Ls+H6Z35A2DzgScF69Wc55D+eBNwWgAIH5KERTNBTrm
OQJpZZcmF2FebQ93hJVjFNYWgbgInQbPJLebtJgMLhodHuEbKuNdtLz1qc3PF9OY
SJ5p5JugD4y53cGWvRob//fTk5l0IHPDdHRi7d+P/7BsvBnI08ovhTxpLS8ZdxEB
sviPqzz/fZZYMIVAopE5dQqVMn+Ms9Q7u/O8a5K3GOMCUer7NoPvWkLmI7k5SCCs
kr1/cKcP5rJtxIX4i8eq3WLkJieHH/VaTQkVE0lcr8qrsZGOPt1WZlezL5U+v2d/
YQmRTsZg81VagV2bjl1HXMAzm3JifppB74lzpbN7dW7DIjvNpXiOpUlRkxtTrpvp
f6BVt+wjABERJd5lIAD7anGnf8shg7GG8i9ikSx9z2q/9Y/qcfWO/PlCxo7qZAY6
T5/AUFfhaTZ5vSPc/y1IkHQbhmTVppd6aVe5o7dVc8xbaYB+LnWnxEScTGY5UCoy
e1TpeUPss1mgG0v/gDct9UH3isUyI6QRjt7cy4pZcXyVHBBmmpn+k7Kra2LgRN6h
URdc6HdYAJi3xfJLCsU/hJymRAH/9heu0CO9OEBnUiIYI3POMOWiDMAHAFOK5oCL
yoFDpZ2dySkoFAdqS3ADRBlQa4G4vf3kMKRvgT5Vu+eHdTyqBeiTfScH1m3++HBx
bVipdSsdzUPHOHbD0/UYjuEY4SkJbeUZVX3satuUjBaPZcr1AZH0Acn/bJqModNi
aGo3JfIaeUfULiQVMnuWP2Uyvs286IcgRNXW6w5DMS0AWl8mYDeO9ZcE7oS3SghG
+kNIvkn3Md0CgF30tm1Vb4W9JTIkqk/DE3nIUgi4ylSDBXODonZ9nGFpPyhrdhqP
t7NPswlMPovH3Xhpiv7oUna1V9dtr9bVKpEfqOJXvdanb86jhuuNrg78xLy3RWNL
QxeDZkmRkCmbn8yTItLQ3a7pXVImIHuv6xprjaTq5sSKYBjgpuVJWrIW6/bgCRpe
cnDXmNFZzDShPE0HknLnwmyHs7mKCi34smL8l4Tzkmss+vSSjea2S2JNTmebljYW
Ebe1wu1RwRqe/urJIRrxx9zuLz4Vf6HV3p26QNCD5mEmXdx40DkJUxG6LwWRQlvZ
roK38ZDnBpDj2RwKqQnvlM+psJ7YCKfus+xdIAo0iRC93w33v+0OwDGXke4Rzv7K
nHm8yKBRdW/dDl99UESnyE0DlabI1ZJiixVtn/FDvC4xetHA3RSdelSXG/4FyDYm
2oh6DJtJH0oyjtVnPaggBWKEDfjAazge/los9MAycqX70AXt799FwXTKrCpM8WJb
qtqSsu6MuGiiAKyaqcRoTN63ROlZ7TCsMB7hUlyzA+vPi+wWiwHlPSWclWAFIDvW
tU/2e2W3l3Cc7WSlYOPmxiZrNyXJ1PTIVVFyMGVgcpFHpJS94DOqxZiGtjwyZg3G
+AbK9v9yzKXCJbOQ4RAadGyhuT8ekDLXxWe5zsa77RcCfD4krCyIzhDZ1cV6LoRa
HAUf1vS64ESjycAV7yq2gUsFd031DlTpzERglIB6u7G71TDOiVveZLycL4fjr2pJ
9+rWG3I7mWtkAfj1qB3V8UjzwuW34nVnj8WbLDZxIRSns2vMsHERz4p43c6V/uK3
zgfE0SrbkdY6ACr5HKQcDwQgzV4h/YnKops5SNJX/EmqB6wK0QtgiecK3IvTDNWR
Wb6K4B81jihvIpSNaXaeSKhDweRXqerrsB7qMwEHrGNDzIoPxmJgsl+bo0c4M57o
0ASqg4wYftuUonxuuHwUhcsRUtxkeWWQ2hTtj1KMPLfdyCJl0sHfp1o1eFNc4JVL
PvoA3FxSTvsJhTEn1LMA4jDnmMbnsKTVC7jgZ2Yfg3nGq6c9oXTF9qqPsZRao2pJ
YoHySSTApjzrV5hWgGhoQ83Xf3H1g1rxIaAfQhWsFLzfFFQGI6Ki3hQ+yoFZe1j6
gUkjUD6jBZkNMSOxc8QtsYzC7LEhNCJVxEgK/eEC0a/B/FfadWk1w55GW7JB4mZ9
v5LvVQRWfFWRpYwhmTnwbqcQ4iUn9M07IxXRt4Pov5ChM733UoESY92OttRRYPzX
QqZ1Drglbl9nAYUIv4scC1QN5yzNuUj81IgmZfYIzl5gIzwhEQNZAE8M1mY0tEQ4
IE4wIv+nSkX9J4TjYxQdMq2qhvcslJzUvg5L/NWDyaKtfoC44+Y2U9v55DEc3PNu
+J6/hSiHMV+JmSPzw8UDZwa6lXBTNPoiwHvElyD8P9Phs2js6rlbCwVhzLY7VQ3x
DJczzbNfdf+mB4UCw/L0CySeSlKdmV56Q2seRQjqcCCgWuVs5n8vEK7iJrb5RvZJ
po2H+dYZiG/bxBamFy+IejEHzGgN6XrlO2ONsk8fMhlLZm80DpDJLtHZG3sDDJ8g
/qA2JBTSVnNKaukIxMTGsdh55CYF83tamz8xhwaosWtwkd+wA9HGI+6mDx56eFhX
Lt/yrJqZhiYU7kaRy2a3XakGxwUZraLWhWcMOnxPu4DtU5WCgasjOwyG3JgEpH/V
c2e+sLwM/rX7Bv4W911pimmliV8ZCb2DG+gcX0I3BQRjSiaSWVOX9WE34omAmXkf
zCE8by4N9mpgP32YGA6r6+bKp0ndDkqngI4v70hr0zzxzMV/Sfk3619TNZ5YodrU
LB0TSv6YtxfWTbANtzeCuBsp53u7cvA7RSsQj9H4+aa5UgXPzJl2baIemDLkTgF4
rMIRV7FdKAemgFIwqMgPm3qOh93s7BJDAY/SXu8W/9xPc2jSsXHlqqhVsi28Z5EZ
mfrb/PnrD6zYU5kmWEh55HmW+7unpXm6gI+sv0Ii+m14/W17Yicaav2cVG1BmDUa
Wg0nNY7qlr0aLILOFsuOuCcZ63TxqXh2oJ9J2+suWFY371++xqghoGleQ2WxyHUQ
67rjNkpSUdyPULRIRS1v9bM0R9sYpab0frdPB+YAuRhKv75pjXmrad02LqLNV81g
hgFnrB9PGKK1O6Rr8lqCudyUqRZjz4vPRtN5OH0wcOwctPE0ShaQYNCljHWnjSix
YxtdWyymYheg8EL/7cfcu1Gy+UU6luM9uLx7+upPVGevtqvj5v5GopW2ckW2jj9C
GkUu2f9A/Ze9jZdv6KTMv5UXfh8cu2jdHiUhbQw1NTieK5wu49YvMs3FJzSSV7AP
JsOqUpyTnunP/nXkW78CCQXbwmIJbYZCZ5IQ8AJ9wDZW1BcwWnRvJRGeXxGVeuk0
2B+NCrWoARiwQLYktHyR0YIE74omeUBSvazkcyHRY/Ih5WKY2gvo7StV8zIJHosb
lUiLZT1dLSbuX8hoxjZTfn3lU/BwbPW+duKC+DZDx3RvkBS1Nf8SDHgSEzBtfpcG
z7Q6aV2+aAfKJUUB8jJ6WUfMPBLKJhqHz/gKW11ar5Dd4FUDEl7JzfMrL5XCgfEq
kuFm/AdnpnuQheP3Xaw+fCB+3sphzaTUCMm3Gpm00VJZUGEqD9ZRk0l8lULwr0T4
2rfhAeiPrITAEeG1he7dDp0w9dI6mP7wP64V11NBAJLZtV3EAU8pEz0katMFADpH
k3A0dkMtmGBDppP1E1OvA/FBfTgMiHpMROdktqLn/ot435UjD6QuOtAucS6JfLcX
5U3B4RDQNkXimX6yMBX++ehzCn4w8CtbK72IKoUX5btdt/fL1kFS//V51NRe7lnL
ZxBsYNFJPvOUxsWXONwjMiclHXRn128aDepB0i5hYFBDVmeQ+lgom50HCdtiOm9O
3TrYr9coeYIR0+79jSOkiMaLWfqjGvFR0erzMYHxpCRk/52Ms+5XIZUVFqva4v3j
qAChoeWnyzowGawmlji12vVFhDR9sWqHO0dYaly8N/sp7FGwp9HIq0f2oSVfezh+
wNr7Oay5zvtekACsHYhS1nZOwXEBkWhQ+48O5mUcyUsxUENnnFuX3zHXKuq3kI58
3Rpi2pIPSzR8R7N96kbi9izImCpjm2foKty7W2OvJPyQzu1kPU27hSzrQdE9TZws
o5OZYAZUszd8BxuwnsYqZ+Z3DJVvqglnxUiT6GdHtRdsozSv7cDBCJkoFwi2B5Ay
uyHRXf4fcPdWvAC7y6PbJO17asBqA4sfvgphmRe2VrS0vC0ihUCPCnyo9+BWAEqW
dOj2wCSNt4WNm7b0/RjZlF94ydL7HI/H4dUS7QsVAi7vJUAEuvxsCrLwAFt1nznT
l0QuWJw/0SLWNPDnj+ts18Sch4NNBXSokdWok9wi9d0tcG92M42KjPxS9giiN+KS
edYMGkxIzdqo/R8yQU+wjxf3Ukecv9My18BYWD7JUN1qIa2pMeYV61pw5yWk6CG0
YKOuohJDoGj7HIr/Bwbtt+UO4himShDdSqjfEK6vWH8R0e5Amtybr7IpIfcqYUC6
C3t7dgoU5QfvEdIrDz5cs1D2ZvP1KWKsWy6Vd+SSIanT/hkfkC6BdPKZ4vyFbAfn
nljomi4MVv+bk0H4elU9C8DKoVrqk4DmWJGamU/ZvD91hQq7weqypoaqgRaaMnk6
BuDNfOk/yLM5KQ95zWiuYOJgd6dYkrcFF/FJ8y21CeaN7si/i4T8lrGEHyu68kXr
SSo3YOZbUcgziip/D9Ha1jgpwqeZjxjVjmj4zZiR5D+60xNDQ08n6JQ2bzpiFs5c
SAaraJqkyYZrZ0yJSqTxPVvgeBik/OJwu8mzPU0b0J5vHhRb8Kq1eeXiLRYOL23I
Ig7w0muVgqgUR2rAABHYvTtI959XMafHqso+aCtwUR9lAWwLL62KfhO0emWkwXWb
VBFP42yTQehgjfxC+2zhKjIblIoKpCOaJmPGhX7SzTkV+X4gUG7gjkyOJ0aTAMOi
9kmrtYLmbh2qld3czvYN9cv8obJ5pVZD9/D1lOc6PnG1pZnLgia32rSYSlNLE+nT
6g4Te/2RwC5O2KJrJJE2Ib3nW+jstYUO/VupcGXTglxoO4s0DH3x75P3yQh28kL6
TEqJJUi/MAr+yq1tOwkrSeZgM27F9SRwz8edYMiiag8jd+mj7iWlM4tS/oyD57Dn
W6Eh01sO2Va5BXPFOhEJRC4587e4uKyyveFTM9csed443VLrnmBOqk/r5VubFbHA
4i1CAR8k4T7zPBEPFql/CWNjHSKsmoDykSFhy+JWT+GCcRlqr7nZWA4farHJbqAc
jywTpK9w5KkpyOi4xC83VjN+gzVHwTGX3MnePND0+MpZ6PlQqRnnaZE0kt42lgNF
HSA4dJvNc/06xtALCjpowoUxtuAqSr/doYRVsfp8LN1HAZMPw5Nc74hTvKMJrGyf
ztT5iAxu8zNOAOUAdDM6iiUXWdOFqzrvvftgSJ8PzQN2xaNATuJcpu6DBf1wouDk
Ui/dYHfgkOQzaa+gRtdzm3gyH89Tx3ncVjNdPDmGK4g50MDiTg71SP75OxUkR8wX
2HpDEdBkj7VIRt8+vPn2JNJsK8+VibxTYFC6HqX6oksGkUw1161iCYr/vAGqsl78
nikSLNFrLG1npmRUvYtJRhuf1ZD1PWSkSommP4+cHwkFuGXP0zXm8DsOnRMRc15W
RPgdocqwrwhBQwCgbLxEFWlz1aNN753df5vLO8v/R65oqv+qTp4iM20NEtFFXXQt
W0WQ3MTvrnvalIejHrXTSrC1HtvoPZHQhGflBZ3SCmJeFCCPb910gbFuPOXhgIgm
YSelfFXO/CPr393TzbPYWwTPFrG8xmY1UHPwCX7KFm8eSxvHT6haxzysKn+DJDQ7
IYvxMOXvZBwSzAbfvlEIchpbCC0RCpRfhks37k+L+vYY2K9DOOJvM5j5Tuq0FLOq
Ejo9tmLGML2xgU/7SpJvsCxOUbIlkrUD7Bho3UMu5/8j5TqNWVkEMOY7aWNJkyHU
x/dVNiYXx4UBVVJL5nimCeogYYCMMZiGomu5pufOERQi6+QL2SSaTUeUP7rG7ypJ
N7zCKSWuvSq/CqJwks7yEFxjzsvDgM7j0AK0Et4V6Zz25ghW58BpfcB4Opmz31CV
Phmu2tFvAv47XkbeNSJX1wZTuFBJrRPlBIlVhnKIal1FCWn3mO+EJKNvV/kbKSl+
YWkF1pozbBygtyu7uSzQMzAaY3CQrjg3rrxjYSb3ATF57sTEOcfjkq2nQ3El5nuE
4QXakoPNwfkGWyl8/fyT/DuHnIr/2fpMfHVEDxsdzxQPX/wQeAu2hBumHByW/0se
LpuhNoG73wzscIxb6WU41h2oGBKQY1DoL89O2y2rRfZGSKTlv3HxC2kk6fhyf2v7
5azwIrDey2T6wMqTUtXbnhtoqrnUKtItFme1mFNOnk/PiZGSApf7Ga7BbE++VtSb
rPkmTTYzfSA0LuwYNiBK7uu/JN5yguhBaoRkS0YSj2I5pTR7F1O+83i4c7HVUeCX
K1u8AISTQxv9eV48g5C4VfoXxbGlhkEN0U4M2vE8IxTsWomx3nnq79GB3zrVRbRk
0HqnfH3EgabxYqiaH4ORAVsm8E7K+kXvCrk3POm+jZIf71cwN18RBYTrb8zZM4Jo
/kT2LMYLPlSmdfOPZH2KW8LCoUE+SQKy6+UGD7sAfuCTcE2winKfhXw++chtnryM
C67yzg5Sf+UM/qhFdNsaf0O51XTAKDOdgnKXWr1fCKubG4h5GKwzCUIgqPRtwx1R
3uWTjspNn8g37FS5qyog7oQNx+R20kqZ3/2iVaLNKqqi3mcuz3YeEhZ1OgmehfRI
BG2WScOVtznLEkLZc5rZWCBiW0j9n1LEloL5LO8R8BUSEyHznk5gSuLzQFThNpVN
hoFDwjQXS/61ffeftaLsii2J3FfpRnSjFAkjzzFOvQH36KuVTmL5RX+RpRpOqFRn
rxsSgdzomUvfMnK84jzWXava9CtXlFYBCo+shZzZBLB1Zu3Cy5R+7kwgML6iEQTF
DgXP2ripVUwSMxgNv4yo4KxbaOqC8oXitCez7VMVmWuvfPnW++XqlYq0sI455fqn
fMXToO057+PkwH91OuF6+Up/+U2hq5U2PFW7LmY3GbWV0mqDkxmfLfMyre/0T1pu
7FJti6qsfztwy29LAuvvQvdVU9fYhrEPsJ1QFKqvzZLG6VaF57yYT1gFgUnMGn00
anWiRCt3ydHxneXJ6CXH0+JrhGmxq65NesYPXpBbGi8gdgedbhEOu9NUMoRajqr9
RrOZ5ZXcz1X5qHB//ojxe3L3cnW4dC1DLIBDM22Y/x/IWdE9qmk0v6XE9kVIlyVI
SgRJwAhUNQc2hiEXWUlzmLFBAqtsIpA93TfNbAx44eRHQpFxoQ157guTGaerWRCY
rTGTjXuMT1j7aBWTWJoPhUPK4f0YN4mCwrS25Svz7R3zzeDTjqgLFQFUBzXJUBf2
TJJa+ktaQft6rgX030d3scc0CnjFqFTTtOdpKOhSszeo94AsQNSgWlEysTw+2h5c
A8P6uyRzPssQnwQ+7vpCWnXrx/GERQjKA8L/BllS2v+8LNGdIjvmex9FGZZ+33sb
OJNouAsU7iiuCZ1NzJcfFBlJ24NI0Qm2JnZlsXl9bmIkbVDbPcc6Wxjb9HgvI36D
8mM463ei8bB4vyh+sL++JNkTk6NCe9k3F6qYjBjdnGA+IeZJ3ZQo+TK10jw4dVC+
4ewk4os337wbJba/p7xjEzwpyg2M5pxLQvc25Y4yBtPdg99+dfxr4/Bd/ABInCXL
YH3bRa4ZN47hoysA95Ku8YEIZH3w0D2Kmvu9irQIUTvS+zKFJxy1nk4lDnzp4HKw
bUtAfwr2Ca8WmRbLuYKdX8wUzAvXUn9ojS06Zn6SRto3oC9l9K9fqMCaWrjCxFHs
wZBwFQeTVZvnXxkaIjP1EIYcJfeClE+znv8RWrpUJIakv7Gy6QjfXDZSz7okGbmD
HgPhKETsbZyhkOp0dzHHQjXmHZngqCX+MEizaMKsSAcqCr/cKYaIeHQk/CS8PdI9
vSNtDVPhyyictY7ORviP8KOBkecTX04CavEikEr22hbA3salgHm6Lsn5c8phl24K
czoLsptxDPLe6uvEKyXtIt0UhqpmOQ3QDBreZARck/q3hr/M5zGzeP5TqlvnvVMN
hi3rKO5CkDVdMzsW9nC20Yovzp9Pu0YyA+zZnxif6SZZ33L5Jf/4JTqXSf/aBwIj
DJBtKYHwqJtA40MU86556g4ASRCTtrideLR4QoxbrZdUH0zmXjg/CRDwB3aFH/uv
7YGHEGmOJXzfztd6nnf7B9kGrRXnf72qMt9mRoCp1CLbb31xSR//Xw6GY00+QmHB
ulKouB0D2GvYPwzPQ3yhXqlyTZJiW7DKu6RlGZFUe/59MJ/ZRQnM5UhBzYchi6nv
GLip15GXRCCAS8+nTDyWSu6S/jQlLm5E8FgzTm9BQAqutXvuDORi7M8FD4gsU5m0
Vo7CvCiuLm9SDYlah6lt0G/q940pYvVM4WsDBaw6Qk2e9Jptld/b3YZtKmSC7wS8
rTHoykJugz0HsjoyuorGZugegbFzWhm+u34pl4gtgO4YoGKV/ma8FixkuOGokUvf
/8rbG5ZSgwr1QdHnTJCmSy0fAriCVSE7045lQeTJWGo0Fxy1vUQBOaBcsUhssIr4
6NQGOHs2FIxqsiOP4gV7vJeZA1P3zaW7jobMpd+5tV4sjZ85ZQrTSIb1wgcJubbh
X2nTHpkctwYKtyy8veeMBwYicyLRmwkjAc4fTDT8115t1wkrf+MpveoZOCJLq9I2
DshItZb2saj7hUJnyxyD21mm3F3fIzeAJQQ2Bw4YzvtNy9mDFrjbuSHCevevPZte
DX+us6zpZBa+dkqwRCi5+m65yynfm7Ake8nYcExB5GzXjFbNBQR0A0UQd+3iZvPz
zMyeIKbjXk2+g2vBGG3T304IvVm3PQdQj7zIxobShNpJ5og1BcO8kxjUMg3l4O72
a2KENRKsd2houscr0oDrLGzobhrcO3ieBYBlFw104nm43dqv7RjxeJJ9uVP21jrE
QdTjTjYS0VLNbT1my+C1Dit6aheBFFNR3NlQ3OtMU3tXgY+/MJagRX1gI2JrndnC
O4IurkTPTxudCI9WEm3iH5SEM4dA6bFHYop7QAiCIfjvBPghV6Q+y13SLo8yQYuF
8blDnI6/nbSvUer9uEKuLoTRYTegb70YxcG4j1odzU3L56Wc02t/5EKnxH8/cFsy
59S/WPnG1slpSWjzBu0aHIhC8Ykc/9vC5hlabzCL5g0D0JzDEaFQ1t2UwnY3l75F
XZXimUOiUgdJQCWEm9+TgFqmkk2u81/8/cd7yKNaRApi2nGnCx++PII/glYYRjNQ
CA1hPor+37VBtuXoWxGDqdAzHFgMXePJxhwt1f+z7DLobZAQa+JaKJFwTVhENRmx
tFG8NKbP0J48+z931mx0Qwml6JJ/Mt5OXOwULO0hr1uGVNV7kzfZwoGp/6PY5hNG
iYOknpiJaO1QhOvbR9xmhzTPV8ux89RYufrQET4BxAob3zFHtuXnP9pmfrp3JWKJ
/7wo+7fFWlYZMK8T+0rUIB7eA7m0JSC3gqXJ6Ws4texnqyLHJyvC5eSPVsmVcG4c
PEYHmfqu+Q6fBeCG4BL1D7PJN5KYNf1JJw4H0jWWFg92UnJCkInFWMt4rBmc2elv
ZARL47d0NtpDIjAql/BKaz50vNwv0MB+OVzGIVhNXbw=
`protect end_protected
