-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
DddHZHwglNZnWXgXUockdmbfkklhBlX5Nlo7sAUXhkTG12MQY6rt7gj+VH/Sj6KLSdHnR2jQKwwI
ZOOcC9ZY9ozNdqGC1zOrKarNWvqJIc4i6LHJRgjpWtGw/798Sj11qtJN0YkuFoqBmDDxx2dtGJQm
6GTWDb15mVLBlWi7rB4Ov9PYehUpy6BKcDWmGXj4XJprfk/j+8z4BJ+Zb1Fvmm8dGlHfx+F6P9/x
6ZVNDe/Js9oKoFOQVJ4LvWf7eZfFeaMu+AmHfylzqdfg6oX79ecBELnl9ksKLDwECkO/1UdX9Pm/
5Gr5sPOu2JFRiRECibcTohlwT/L2L42c7O4Lfw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4400)
`protect data_block
pTHLl3iXcyd5//bQU05LDgPPdUCoLNjPai+X4fZbX7gVgfnE7/HrTMIjEYYiF9H7HVHyQHK3HVzG
fpHHuBaoizENDS5kNmMRig+Ak95P9gY4SYbjDITcG4WuejLHxL5CwtwagFWNBzCVu0FcfgBPzB5L
EdIpIjUtFGlz5uf0i6aaYXpUUzM9IDHEVg+DsaICTjB4Ou2gmySDHIycZohHEjuUYVLRt+OD1gig
o5DpwoxCHimNQO0PSytxsTL/UiHQRMCptNhqDdxf//HFHQsIOXkN/kU2Y4pxLDlmakNj1jBKuu73
MtOZG+giwqF0xEv9y3UVVMTKyJMiYObl/02h2cr/TR6OtVbcRE5PeLJZpAggEchAPThPrmD1BnLO
5QjUL+f7cx+teeQ47sc2JTbrxgfnfhpBhOYDkBEObOn3C6D+oSY2DpgnBw/rcfICfVzKLcbEPGFo
GC9phfpfRR3JZ0qkUODvQFg97qlCSo4/9iFSZVYnbBefiqhxRa2NJ59va3sSaiPx0H6M1S17z1a4
m40bhVF1bdc75kobIgT9/Io/CAuJJHVjAo5Bcyc9J3gg5JqhYiBxAAJEIT97VB0UlcIvcvWOrm5f
by8sNyRel1fnCEvaam9orU1Sl6Kwyz6+d2tUmF3RGkHow7ZPgtCnAeYCMaqp0/+OM4HvBnYricDL
j+F1lwDKlUYXieiFQkWx5lfIVNxbqX0r6HTlx4ywvKhaWTsvyGJ3gEZbyIjBa+/2wgimYdO4aSsD
oeXiIIQQEhR9uEqUyf440OBRLngXkrMHd/YwNvq48BlhmNCvCsICNlLNVtn9pz9/2AMQqBvjAvBl
qw8YqYus4MmZtuZWpRN32WKVPS+DMWCe5vucp0U0/Yoc/xsECKgCqFr0htZmyQFV0eVjZLlu48rh
RKR4oyKaGC9I7Loka2dGlME07ej9YhUr4s6NS2++YP/g6IPSMOx6pg+132kmIh8ENZznPaoe+ECD
Prla9uDf6afvpP/IAzc5ezU8BMc4s602/yRwdnmU9T/AKZZ/R9ilhL2dIQ2BBJCfCbvS6Yl5kEGT
OO+GOeB3GToI1/Q/JAviQfibyS92uSJsvcNn9VDkAcCpxk52q8m65Ya/fKTyiiwgTRuK33qorezM
AmCadnb37NyZE/hAq9R+G89TLgWNgMJB7aUOjLN/tDZMNDOjwvbT9nvgh6WkzY4AYCIUKMLiqEnP
Y5TDeaP0xebpogOijzJhj/UtdNJGmZ4mJXSNHGRzMNJ4WyMY808O9juqad5yu+DHCz75xT9S9aEo
EVE3RNNsNMRf73+QExRNINLQxPqIC72/7SU23RsNTrYBX5uAlIYMaWHrR/Txv4UpQHllkIuIBF62
pHIsfFGm8ZJSf51k2S0Yef9pmb8Hrc8Y0/CyJRLnDL0gg0PXbys9e+1eoKT94G8d5/K3e/WbjVxI
8R0IjclkQ/2xdxunWIDrevFUQolpwcfEkzTvDJqgs56Bq/4kiaO0KgERT6Un6zrL2rR50aPRvIwA
owoJHRkIVyrxGj2DerWRfCwqZewh098818Gin1nYlWO42Wznv8eL+Iceowa1ejLdcYSA7JEjTeRr
TPFrvSqXaHHZilCeAbxVa3rNgerOgJdZWeoEzzf33OlKzSN4jIKJKtzUvcmwGG8UcnTum9UJiJUq
Q2lwiFN1i6DOHICoWoTeCuos87pLLPDYeV1suq3TxycwFT0MPGfNkam60LR+jJM7Nhd7A2H9sCC1
HH1NCRn8Ixt/AHGJ6fNM0BZZJ1ReTAPDJloylJlW1ZM/0+F2ofHBpsWOjgPCVderVfKLHQCUX4gG
mkvy8bVg0H6rYIO1WbrpIdaoBN8OJ4/riOWLBZ4lDutXr6xUfErJm+1LHeWQjXfE0ImjHTIagnBe
AgH7k2pjJyzm9guKndtHtGHbnzpcdAaKKx7j5RUdRfynjjgWgYoNB08k0YSx8mpuH4eHXVkmhHmV
EjV2qgVfPMqM9wUkHvKQp16wZzDTceF9JXizOBjyIbKKpZj9mOENiFwOTyePyYDF0hwyKVnjwNqr
lPHKn+GADLaUPNdPZPEM0nbd2aSM3jz1ALNei1b9EtXxwyNLc0SkZbchYkpjHXCYFEZu4lHyhZoP
y4cwF0P1YhN4EVgg4cUbut5E1STlXBWhCL/6n8bPpDNgsGIR7E2DS4WzxycAKdTUr7bhK6UcJ2Ze
1X34nvEevpzRCY+YN3+os6kBcqlliNmkndrqGqWqitP0oQQAFcQnntEMkPkqKMEOrCvYMTlvlgEb
4O9SGvidWzARn63LhlPpJKQBZ7RkNH84DdEN/VqAu7f9ud/snht0CLk/9sb4IOrMAHtyAXDST8sV
CagNSUVgMxRI89PbcXO+ezlDg04H++syckTI2TNs1ZUkwaXwlvZn3Ux9NjtX6DCwxzkvSTCrXt3K
AvsKYdcM1zsbXHj22es7rxbtkv5Ib+RiEr9Fi7j1fmgC25x4OpH8TfmF5q2CE6RhsUiMwMFoTP0R
wqvRw6t0U36myIciKo1a6PFnf48OErpQF8m3VC4nuli4kO2fg1OSEUEjRfXDbfca5q0ofJf8peeK
sN0pKZgDeLkA1+yRDZJTep7iycljuyU54dI++0b+pRSuMIY3JS2tHwJfcJQwygUtW/6Km13MX5V/
vxyNbLj/FgAJIET7eCYP1TxL9SDVrpgic06beD5M5KEFY4p89iAAbzNV0t3XA0OxYPbrnHuqwmoR
OuNuTC5tQ6vSq2c15Tjft/7+zTMbLr2Etp//ERU/hB4hrinDG9FJkj5dU2aIqnBYo+yHg/669C5G
w0Ql4r4vsLogJsSbuTgzMmID1nz5w7IBXT0CTJtE0IVyxCHz3LnnCk8HFOFkknN3rBJrRGcVA6VI
yAWj/W4MAtE1RcJhBB1/d4Xx9RYE56RPTfyp0mpVqkU4gjPJGVUzx2cpFXcXkR3kZRF63L5RWMeK
uERIhFY86gHnS8RnZXmE9b5senz92TxCZ5oh6Fov1Rj2gphgFC8G9A263u3lWSfEniLl5oZ/7lhp
E+T6IGoIFG+bX3tiHh8Z0ccC2N+zJ83P0bItyFS6lHDYTWXMN7Eta/n+V9AZ81gws6S4CKNWrgki
MEhvdD1+4k5x/CmZZ4POIvKDsgO2lQudFl+ZV2Ia5gdIX+b99WyGREMkkQki+xGA5sypmLVRjMwY
ekcm6SznGgesrIT9BS+BdqgdyIuys+XeplV8AjVIB2CWlG/cy5POm8hoA6N6QiCcE1Ubp/cBt22C
D2m7+sU3CFYZvirOI4rUMfcIVusZvMB223X1Vl5ZSh3fAxsjtKJ/WobcxRaLXuhI5ue3KK3ula60
uj++JNU7tJUdaoCmo7/tmb29hKxaVEWX3WDKM1MH5YctqEin/B9a6pYdXPYgwdW+a7O0Mf/lAWRp
qYZbHFp0U9v67GL0AYQnbzTYXcV7tu44XhJMQA0b5sRJStkXgK2EWelxxRKnE7tq3G2u+trvQm7N
VmJkwOR9nuTNrZkSwFPGv2TZcX7cezsZfALJBzTPNt9Wf+FbXrvu/9luudXvxqqT2iltOaMLEvrk
QI7CugZhdkc5zz1iawAWnHs4ncc2GyEWY/XFK0fPHuPGuJVmhjC+HDDSlrTI8wQNdomw32V8VTNN
ry2dbBUNiAGSe/YN5aNzo7Nt2Yi+lD3i0x7QHCGUNCEHJG870cU715litzf5Y6fu1Lizk/Ml7Hlg
7PUH4/FVFOr/YzcguG0NcRiSIEMyOiDmh/ZyIlWfAy2kCP5KG3l0mRp7ebuUQAw1v7qglgVcL5Oh
vSsifOKTgZtwlua68rzE+Z+IHrHc8oJnTtSJQay8FNx7cWnCGKEpq+NJPL2cFGGBiuGOFQYW1CiP
AFQSnznLX+nGF9P16rFVbYfzhkpeOAl9duto7Kn4pfKWD4PMq61TT9NcKkr2hXAmSRNadaK+bj1U
qHNcexY+/HwpaUxvaU1Lf44Lm/RuXl1db6eeukbz9weTV6GeMzGlNW6/38XI/krkxGymjbcPZdGE
e/9OgHCr4NvPOKoxwZtamJttyegirFmzWKChmQnsb7gi5UV9N1I2rBe8hsmV4ewiC7umzY+MFqDA
xb93BQ/NHXvwksH0VLX0jMPyhZL3AnG/1ubkVNeDJA5Rq95aNYN4hK/CgjMqBzz9WHasKvjes7sN
S4CcWxksN4Kagw0yqsY4WI5nqFF2t5OhMHecQAiasAKrwh9bpZ/kpFZeiY5fdDK32Im1kxDN99L8
xKr4vFHnhJdEyRiI4a0fAL3UuYZY3Rb1tGLNxlBV2GySkM3o28CV9CjuRnveiNRIolQZBJL8ZAa0
n6H7Esxz+99+l0qbg8o2gKqqxaH5JOyw5w/A0nRV3E435vcqw6psh3s2w6OrIOWipk5fG8BUzN1E
BSzBOJXvG+gjY4+oMFSwfcYYVlOsfIzJSzCO3cFpNJKkkRkllyHbnPA9Hj6Dwze9C3S+z4nKA2jm
zfhLSalI5ykkU8qqd63uvoLRECFQRmfQWoRLxwTgCyqEXJxB0rbUJd/F/x3WMHMvf+Jgi1Oh4psy
0ZOyPXl/8f9fprBS3QofMVMk0nfuMOcKNdPVI+pRStPA9UAQHyVFzFMValL6GlFJhicFsQZFjDEE
J6tvypins/5X3FEevQcNau8ZoysxyRetnvlbE4qyIPIWcTBBxvRxFxii/DpY7IoT1eb+CsYScem7
mXr4x5HhS1KN1UpcTd7vPo0dJId3KBPfKuHz3jqUs/OxFGpxXn6K+WPgT/LxYEEumRJ5zcwI5e22
Q0doB+dNOnyRbQdlvP3rr2mvMbDQaVmYV5a7yK/vL3ZO/LXdIDBEOM7BnFIltEc27ftaWBjZBXO+
HPsLTG3YF/z5q78zdwKQZjfLID6MuLaJ2/aDDPsKSmR9gDadabuumFmvnEdmOsAvV3mfq3aVigvt
mXjA12a+XHPfJN3H93exPnRAF9fI7iwlz2AlUUMEQQ77KpScRrtkh5flafJDy4w54dHh+RxfsDFZ
AU85YPbDLSnKWl11avM7ZtnKFvy69cZ+i66/JlLjVh6ZmIJUrbpYwLBEvWkChHGu976yLVSYF+OX
MioX10td+EoIZ/uj769kWwzfTGDo3YN9Gy3KNo69OClwb8SMc00AXSQQcV8vffWReEdbNgchZsEk
H9mokNP35CmkM0J6Xu5RimQIql6QVgMENMjAYE56IpC0lBUCig05evl8I0tilSblGDVZkYR80hVM
74MVb0ONkAI7aTL3zIZQT5B8JdkXdMAQdALxOM1C/eVSyVlLnN1/lMbNeLxuuhMFqL4rm4jARruF
XDe8C+EvG2yzzgbITqxyDikrKcoD5PUKXm5hnB+R3hbRzZqlGpWwWkHuHB7n9BahvTMUAFHOQqyq
KZwxehqL5D9JGoGPMv6G1+C69wORKIK5zxUOuI0hlFQRAhy7WNc+53fhJmgznEv2i0Kj/Hyff9vl
KQv9Uc4c0r5sGp9B3uZmmU07jjuQafH/RLlnko9F0Q6HMp609jQFW0q6BIM4CqyzyaDnNUcWhxBU
fZcOQmNNip1a2qVU5cwdGmSEoyqBNt2tVPK/BsZ+ESUFpljib568Q2lZTDz7q+ePKRSXnACAZlIt
5TuUN9xP9LlR/zdLqfzRW6MCOjAIzcAvrZIVJgEeq5qdMrkuGe/T/HnLfkExk9CfwdpFZAobWnWe
Izj6x9QQA5vQAJwOtrtzuzkDXFn93ofnsKDilcSCh26LL1I5IojLLho4YOmwr+ZnV44vPGInU5ps
LguiyCpLI2AfUTOROpL0BtutjsPufbo5sXTrqJ62StJCliQEOp6GeId9SvV44KTMT/Aonp+I2W8a
vKSk8e5vg/ugrTY=
`protect end_protected
