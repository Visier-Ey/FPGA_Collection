-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
QcyHfNMVvmPGXI6h5hpw85CNUue6s8vXIZ2iKQfJey7Ufv0Qif6VYLs6xQ1aINTZ
9GQz5TskI3OV49BRGqFTlD4AQvwsW7OJgubs1UGpKs3UiWQS1NR+HP+OA0HDbBqn
NvHRLEWhpGefe1/YGDIh+LwxfjC+FOw9IaLpC2AOYfM=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 24685)

`protect DATA_BLOCK
kPdUu/QGu7CqUCS07Js4Hh5zP1JUmqP9dSf2DjAuNlWbdyl1jl6BuGFQ3GtpAObA
iOoZ6TZiCH2gSpC3htx4A5NK3xUsgukAXtUreqi7OrDBDLhwI0oZixxJPkjAD//N
DR385MQG9DLR+oRB9EJ61CUYH8FqOuCVwAoqN4ybrBl116QQikeOav59lb7+X1ZM
DLi23PoN5alGxeKkClsHGxLruic0ZOz76AJXI0PXJwAB5vyVH2Uot4yVyElUdhH4
HZwD8OE1+gTV3d+37/bSOVodmcsyWlu6oqpOvUVOwT1uFIKVn5WcfE6UhT6hoa8M
sFs+uc1LwNwFN+aRe0ZplevawQoj9jkE3i4feoKoPn0hYu8V+2aO0oMie1oWoRRG
DgjcQ+VnJXGn4EKftCcle59f6YG/NGbh/AUYa+53P6Cc703KVkmNQnatU59ITC6F
aPx0r2/6uOosxN5QEBHKM/lJ9F/oeH6ZNTfmiYM6bVQ7yM31Kto6Pp8LZDQZh6vo
KL+l9D7WKXAwJW01+rtTaGcVASWKEc7X7S0t9TOiGMO6kD4ryegazeuC4cfp57mL
aE1AN5ZcXQ8FVwWYfQrZJCX8mNNApkj8xE0c0Tv1NQmCgRXq1aYo/EbuWKxBHy25
4lAW8394wL0MmFbBaLnlY3cmgGggvJ2HxLcy5fgXICp/W+QocSibMu/9HtvwrCsp
MwGSwEEFWeRUb+uIvKZsyabglFk3V1NNO+ttgDagjkiTAjqtWpOxpVmruFTYqjGc
V+21BEkDlUB/WyAHGjaz5SBrGBiIHiYBlmYaEQK/ITFEENEzJZSaxw1Nvds2gPZ0
DqKj/4vhs18U4TRDe8PK7xU6tOBzEPooxCYO7Yw/8RswlBxabXX35mJYXB4ajMtp
3K5Voz7YhZTJCPuQXygz3L2aNntsJMkNk0OASnEEpjcN/LTx4MQUGRTcu0RoKOju
SUPgMnCbofqiYEclieEqLUHafcdGcR9na8undAH1opirD54NdEkG9ubQ8OHx5jTL
ueM8k0DYjkN3hG+h5ZGvHFcWpzn3lYpyGaKLuxpTvUbWonjtxafnQdKTO+HWODwb
0gqrJ2cOCj7dE8+ZUG+cbPY0PtauyOi/wRLxvGZc86a9SQoTaWsGe5enbu+a6zh1
6q7Y7Vsmc5eyeMR2A7xWJaEGCf7EHd9rDyyCahdNJo2E6p6bSOAHto7rWu4m2eHA
77RD+MskTKHWIVg0/wPBv61eaF6NyB/JpBT7CpzqX9Zxb01uJnnVVR+emtmX+f4/
boMrHHGH9XWDwShvz/D0+ae/6MCqJpBxRjAjXAgy3Nbslnr1A/phZDwmt9sEFrVo
snYXSh413+c4RofVsXxcEzHzEzhWE83uaueV19UXtMoJYwhQHGJa5gGGGGQ20DOZ
HugxEW9hkEhhht/+KGVTFjYnWZVV1t2SxVgTFwPRClRfmb/XsXwSt2LzSRYkgIUU
GfkbwUayvtX6fCjVuGyam2bdr6zvaQ2T+FDUhY/pxl6bmrnGhTiOPtAhNC8pJgWS
yv8hAf4X+kL4a9Lu3/3JsrtOLhLkF2RNRO5C5mfPsmRgcZ7eaqxWdNQDMFWFrXqB
3UC8dLeVQdlO5nVXvNkx8nn+RoZv0ZVey4DIkQUMt8681mI+M5hi0mSKji05aOnS
AFam1G84lfxsQLigJe8eidgRLVfLwr0vS2GyZoGGIZxI4qyyOrMxAg9pQdD5YLK4
43jJJ4z/uboMX8PrDMeUgqETa2Wsb8nrZyrIq/j3g+gsJhyvaEjvOFI/+SaKPbP8
AdI77Pd7dcbKbPd7lrNXUXcF+jG259gY4viI40Uy54ofgMD+XLjsPGPeJM+j3YUW
WI6KNDTliRNJqxqBwbh2V95Mu4UswnLGB4DUgO2jNgHJ0MiEYLtYw+HEPHtUaHMS
fpNu155RRIaark557sTHrMiMxv1Tzv6Q4NMdhcjgTEF4GFo9jOzeriQx1Qpjobsv
OcEVpoK3fMLFGZBKGuK7BFteQLLAjDVnYYSxyOtyq4NXapnDraN4w41w2AB/OXMw
2x5gRHv8Np8vbay8QvALJKmm/U/0ndej0W2dXouCa2pcLjA1X4UPvaKbSh6Lc8Eo
mSqCjc0Nybt41QsWuVwFPSw2UJyojvIXH/GWSf6wfpLnGLIjpqGioHTxRJJT1A4K
ChHSgo7/rY+dHUjcO9eENFdRqKqXBuv1uA4K348VfHt4IxNz76Tou/YSVIFxPTUo
bskZCN+zzz2rmCnBnqbz1MmhQ3m+FseyelNg0UpsXnU4lXLv5qYrQTpVwCZQpnPP
+dCqIiYZGXdWJPn2TDUhxjwdhmTY4/C04TieP3YBFJLUJgWMJUE0+HHJ+REfGhQI
y0UU4H8cdnCQUdlfhp6PuF/Q3xKY4PKrQj50bG/l5SvmdedYsbbByqLUKSfIo1Hm
aKxs1HiFbatykhBVKVkvry1JyjY6JeqGd8Tt86TrmV5Fnsaj6tZxAq4/vaSd7ZVE
pzs2cD9BpevFXVwzsMWteYTw3jD+jl0OeQ9HbVrLIUP1euIh/AMXIhbzJgVPU3kk
u4OTXR5neVcyQTU81t2EgChBL3hp89zcriWLDZdvxTmWlJAE+DQdXLYzyFd+oJm6
S9kWvYYzmWOaAoU+jLJwz9MUXFgs0+YF2sylJMzebpk0G7DbSYG5TU/mxfj0R7qb
Ma/7UunZPmTA3AwDORJrzXbeyy9n69rLakLQkYZP/TMp3psYLEIeYXDDqXvW7OT8
auYXyF/9FhNQnCT0IvKKs+T1gQ5v38wPinzeC7VIM0BMI8WdiJys5nRELzOBqu3l
BtQZai2sTbvzU/eMB6xfHqNVV8yYzb6CvIfNSPEeoHEa3Fmxkcn3peRat9DJdztn
qhbifCUZg4BILRqi8fl2OnYBO1NrsR6iuX0eBAYIpCOHTmVVoQykqbSp22RIqKRs
x0jPqXOJUs5Wg3azxMYiaYgstU76zsRWbhREj1IvmxWgfFGXZWdcDwYXU4Ooo2G8
T2cex4+bXPyHaE1yC1FD1FSPxdgLssrZvSxqb50brFW/ZICrS66EdjqPNbZbEdqH
Qa7YP9gFBolyvdQ2SW1xDEGGG6a3BH+Pd5R36QY/vcO4M5+ZiyRRZD8Gw9gkeTf/
GP2+TJUMutRd04JV2HjN35t+MKmzw4ER1ZOABcWCcxOWn7BA15OdpOrgEuaOVPPr
w58apaLiS+XKCeX24g63HR7ENlfPmCB48vNyLQB2i7F2O8kGXVemneSOe9oGdBfF
QFHcAshrXbutzxRa3w4Y1to/x13Qo2INdipqGNR/9wEtIY6wYVtUpOD1cJ95Tezy
c/HyLA5GZZbzID+JpGuDZ4xnoccQDu7HCEwU4a4NWg5bogLvba06VnpA6wDsv444
a9rR+N4ntvT96ldAznRUf6h+/WRIwR1HbkYkCVaEahZdU7yIubDAOTL/5q0Zygy/
/dBvrXnQdokqkLk0zSU4muE/VaYVjzNXznpenX6DIR7XQIqtqMQ6wVpQStcAgW4D
WazCTTrsZn///aZ0SqMfMkb/Kjd0jnZZpzGpl15EE8vUaaaiKDJQEHpEdgV17gfC
3zAf5DabxnpntXBgnZSKCtD0NmMoNYs7/J6L93xRvaSqel7fE1PfBDIQ716DXAbt
0hUkByS70AaN3OQ5f/nwWmXI84A7I273BojRTDkCb4/nWQ/AgEK721l28d9IdPrr
vzKRIRLeJs9r7NMEC1jXqQDpSNEk1zLzYRreJ1Qw+vGkDJ6EgUS824jZkzc4pTx+
rFsO8LNu8KDjPKRxFfa+I4nr4tGC1jmplUe00ByL9MY1XgJhqxf3cWC0JL1RwfcC
FfBw8WhIrgDsG3U+AcHyCMBjQsqPJOz2dkdbljVB1/goisvjr/LIw5KwotORrr2n
2cKisWNQgSzHU+lHqadW86ddwgkpCDy19xc+b0aLIDqz1uojgnYk0f8Gg/Eu2oc8
G4X7EY/g56wEIKhkWioCKciLpXAobGRCORrJ1vzOHWW0YoxoVxffWwat+XxvJgtG
/8QKEN7gl31BdPBJp/OhhBN1NnC0OEDCasPz+240CHP6NJOfBOAsmLHAlZUIGwYs
VyGylLAl3gGLsQnr1JOffLCsS6948WbiFr4uIWqiMDRRWwMgzqOEoFlLqAa+mgq5
Ju4DkfuOIEDMc+5OMIEiNQlSHTPjWFzmQPvz0fefDrLisQ/ZMwWYedHOee7rHIxE
+mC+AFuRJU09O0qcPQbb5Ji3hLqC5eaKs61peQyC4dJWiNCUMEjGtbgfroc5tM26
4gVV45py1Ooo1Uw/pvy8Emlo5NF795K0J6WcD/MndUUtUbnUQF2yqOGrHGB/7kfU
wZAxqliIKakdMHtW7TEnoC4E+x/MccBoJHGtDSGV/ER2qWLYLkfXYmjYZ0b0+5ss
6PCGn0d17aQgrIdv3/MUHk4pf2ddqiGIt6PQyR44RvOxl4nvPt46nZhH6TW5QSyq
0WsrtW+uTRhP2tYB4/xP71zCR38gQeHxq7o+vWpiMK7JTgUYMuWnUZRkhfuG3yCO
PCMjRn7lNBppUoS/3+0PTDvptU6bNQ1QMK4Y65dXjHBrBcuYxzMH8vvrk2EZVvMj
Zogs62McQZQX2gk0Gru0FX7F4xxk1DSE1E27QQJdGdRoTNCOIxASt0/G7kos5Sso
//iqiEelCTQOIOjXy4jIwIbQV09N9JCCjBfW714A4bzRzAvekGTqqe9tadodnFKc
NqtffL1V7ohgezwGR0P4H6i4II8pi3uQZ4ebRRt1yy0u1qQQqKI5cIrkIpqv8VYl
/HQKK1iGuHVmrtseOo/aEXYlsmKoHxrCfFwV2RPMazpsQiLT3utKgQTPJFu0eFpR
+gz+wElLbqPDkZAzug8jPfsUkx3m/5tXOhmbsWJvuTqeaFi5ELubKVDQMgoUk0rs
Xjh3EliGZ88eq8kSiFuvvKLOqUpc6/Dz3ltMrpqGP01gUkVd73x54tUSmvoWRiHE
ZjXUVNdDuMfzIdh7kzyVO6BBVQUvoILXdB5xGkA1jtMG0jDiMpoNVyzXekhbITWX
Pszab5qf90ohllJyquYDvyrtbj93jEerQ6iNb0m2SqvE6lBunJQrZoC5cMJBUwqC
ZQA3dqWpwFzUZfpKXO4TOLe/99lm1CFFB+a5Sg+Wm09vRAbLfyblIqGnpkhGg+N+
BlDWkBZLn0DJ2sax688V52aXf6QaL6SXfHNxwUnVgoNrhNYEUymlHPnsuVDKrZjr
P7T0+nUwyw44Jugnvtnuz71fGw97rQY/E4ZWF3NJwJzZPQAIwcytd/HLI4VO950X
T81Vdt43r99e3LmlJRVn4XVICgP3eVBWusAYe9oQXdMUExoDMqRBWnxHHq9p/N6q
pdpeguR91PUg3fbw+wjfSs2oDAbiEWOosQaEebSV7a8bPbK4FcsOwWxdBJulP6/X
mljhV2KvlqWNQ6mcN2PLiVjn41bR1z7J+gZjERcE5JBQPOJShzv8Pr+m4R7tXcVs
o8eQWeAoXggI9MLW4N7FvF+6oPG8PqyxKjTAUXorg/Ur6uZ9EQQgCRZSRUS5iHbA
CRVBrfIY4/TbTmJ6wmsh83dNPAp18bWMACrO/stVgMFNhr7iBZIUWJ6MI82Tmj+o
aEMQKbzyhDAjakDY8GpnWeiIzRvXfLuk8w2bTPcor5c6nMW+G9fYlio9QafUyv+n
4Xuj+8dapxsP17a6oELS7UUJwHx720wSX4pFvDzzVAL2KEUUFvq0CQ/6Iqe8I3T6
ytnbiY8klAjWG0aLg9YhZWBOna9CcheDQucz2D5r6TAbjUqIdtKk01TW4duL3Btz
1SMS3rku03744Vs+DK6bai6zP5nhhoBzVmRRMDperzAOEJ7mGX5F5JRToX++vT2e
pKiB1q0YMHQYc75vy2ZR1Y3q+VwS1b1Wb1FHM4V5qebcgfBr/ZcP5xRPcs0lVFUB
8/a/OsxevaoShYy+MjRFOs2ejrtEHfCPww2jxp6T94mMII2xGKIugCavNJ933Gv/
FxORuqFN6ryZsWEWkzPtbDeIKkrF3XDGAQNDLD/d3cQJh1DSIawfoKIVawwmXmFf
33VFhSgq231ku5wcVbruavnkBi1z0NhbB5QxgItA/T0y13tkjjP1ae5lSTul0bT8
PVJzyDm+7fho2cXYBI7w5ekTokg+FT5QZifeUjBq+EYb4q2gkkRNyc/9LiTnLX8k
h1jBQ1QbG0PXSwoaj5uE0lvM8ypEeRkF9Cj6uSiDLsAIB1R0jLLp6vMEOuKAS1ar
3KOZQHT9NJEpTpsCGQ9v4YdnXjt+CudimxZ8a2RQYKaOaLNypEj4u8stuhqZWAl6
4a3A34KQsldhPxN3sQM8xfDGOMzdfwD2BANwvpsbAxCX890V0rOD0r3BxpJXy+a6
Ra/pUPpUpvr4uvIzN283b27ByUmOm9tL9YGc8sGx8S9gfXTFclzmCsIt3ZILC5X2
QZTNUSXzlpFoauAAzHO/2H+Hu4gn340lJbPRiEbibq76uddMI0/EsmWR8qOq6sl8
lUwRue7V2JZNkItNdD6i2JDO65+wsp//9Lf3ECJjiYPWgO4Qa5ugAedbfcCbArYl
3A+Aje6627+GKdwkyz/+2tXhXg1LJGWR0U2EOvduX/fo7DCKPuYqA1hGB9xsT2Zf
saDEgU/4TLiGcrNo6x0yOizg8BSUadWyN/tLUYo51Jtlcj+CnhCqKqkPOaO91s5Z
8/rcnE5NemAlTEzs08gW6UFKfUwN56oEZEbp+ztx9txXRkA3BEW7bDJdNGU5EILg
i+H0N0WmVHAV3hf2BjDdBMsFAWcSbnVWsO50Jaa57iU/ctEpZdgnuVyCwGkk0TEv
JxAe2aE6rQKpxPxlGvfPrlXiLnBQjfOkjpGEpqSbTI7RY9gPziIB7+/v4So4z3ih
GNQEG0oAgLCItRHIE3Edym5EtaA4qlYec0O8KEOOj2IESRsixtOspV28DcHN3kgh
LEQEhYvu7+oy0LwXEvJFmcjtYmndADVEL4btkjCHnv4SiQCQN5l6bnU7dn71d75d
F0/S8lWUT2cEd2qezjfXJkB6jnXj/WOpgfHyrJ37snHKBHokaI4aD368nMj7sn62
laZ+fcSoM/tEJsFlPTYomDgw69kmQXY9whtFVbqirx1eydFVBZz7MBZZp3SsMEva
zu5eNDamMqr0k/zuVz5ynor1lEOKmG8cpq6XNjo5tndMSK7o6ajNITJGQCB96IhI
CoOH0yZQ77F2Cv/bTAOowijBc0BJ/xwfcqGqEbRSLdV1ER3aHsBWDs6shFcwK2kO
qp33cKxKq7XF5kH95cIfYgaA/6UKMXWj7BX4TRvQDeWKdNd+en7e4UeFXxDZZ3ma
Qy/QIFuGOA6g1m+jIbbh9sVx106ALLCT848LpV+wTEKUs11DJdKePJ9sCE7s5Mfo
7//lH9rDJpfoKMoxtu5+szVGaKdodmvkdgVpCydFFBGpHfU+cxw4Vw7xfHtaQPVN
h8hAIm3DWDw7Ds3vSwLFGXpIoRjRlekpKRx2+Wd8Thm4pRhDhoOQ+Wi+DfKRnSa6
1seB7nOcP+Fz0Tzh1uPWyhAhl9BXQi/X7zCFMObsRivYBtmvxG13W6cYr21hbS0j
s/mwjCxNBb5XufibCkjFU4eCWghnfHM5eKnvtf/OgMaJTSQcZhPqwH6VFq+Ho59Z
E0V9B6D5g8Cocz4smAk6Od7t6m+26GAtK0Y44olS7XqkCplEPSIj8ZmwwmpaYihM
3sP4qjg+VVm4xrn6bI33ta2joqP65c1AcrEtNY3z5pqkTfGimjreUwhq6pkmlgy8
GFc/2mew4u1362b15cFWS/KQ6kw1IGxIa0HiFSCoL10/XtAJCem+gQTNCjMI9Q69
w2sYTFiJflr3MTdEteqbSsvr/IQ02RRvrNieZKREjz40brK8fhgs1KLpWJvBRZy7
zFj+avJF49ccd50ra0opN2EeUUU1q48nCIGXrhJ5VmYpZ3hN83QXjxpTkeyiFnW1
cs+88g71d6tpErZzVM6JeVcW9Cx3IszUcs505ln5xDnnRhQZELmOYULLex8kEvqn
5iugSUSBfe1Ujbye+sWUIA0uVfXLfQdMVkaK9UNIG/9CI1ICqk1UT+ANFaMFuxkW
kjviUOduAP//Uq4+9TcNyGaD9PkLorGKKpG/EdRJ2iNNzA0pYf5+WdKe+88vOrw3
y+FDrJq4e1aSHQXSabZ7rIDygjnfFY0N3lcLPsUrbV322BR/rSStqUqJHAxT1PCe
E12osdN+yL9frDizX0ih3Y4UNhtdecEXQsEGc4AZrTom4bKjWEmw7I+/+zbdJj5u
eUxQMiGoQrIhobIvM1Zx7Hzjy7HDZMazoRFvn6G/LeCpAObx5znZB4Rsu824omvI
rWDQLnYov03cJDgoJKJzRkX4FwdGs6JQkrnGYanZzvKdBJ9jZd5ZvYy8D4qMLdzY
zF2tCV2YMROBX1m88VdmRPZgkXw5xGOarNs2qHG7i+4tUlUVxyFTpH3C/M0o/J82
Y0t5lbkgxWPL/q8238IM09QXzcvUhftCicJEsTqfpcARNls52/+kVOzruokH/jwU
zHinAWUATcg95scOdzLO3tT++Wg1V+gh4uNtAQN7EuWN4UrSwQIcyE67djUpif5/
hljZYfNJz3T/Zx0h2zrXvzmgwDj71HdF8uvPtme57+19JqJt36kenobYa4rv8OJ+
zzJYD3cPQ38EGBJT0h0Si2GkbKSSRIdw72iXt4Bi9UpjormVg9RGuRoh2v9d3KAd
v5X2LlU2lFKO9NuXX4OYoTugfFY4J2cwXktbU+77xyCnxVSPnWAQHxBJ/CAfYky3
MTH8rpcT6viDBAxTVe1QJjFkyrQmCgvnTSFonLtGxuhhnYtExse1A59mf34PnCua
r/3LbKXKfp0m/sq9roRF718BlDElNEi8iHoLZFeNUHw7FSIsXQXFH2BzD5pE7sE/
5R6z0mC0dno6yHeaepmiEP392M3NXd8yFs5tRWwwbQQhifaYUKv+LJO3rNr1rKJg
RNQMDlc2hwsPp9wCEjjJ+kn27HTmMDeATzAqTuNEKMuqZ978ziQkitOd4mRriMj8
auxWEmp6B5cRcz+ZbMIauy2r3UigKy5cclLIpU7J5n7vUnsXFtvYIXgEJ5jlN165
+Q3weT06uDBrEsKxZwKos9yX6x0p8il/1NPSNW7FBDm7h3zlRWtVECMu7sblYpb0
jUrAkS7uitu+KmLr8Yi0ZjcNGlAo1obV/APlU/buvzNIBxVbEupZYRZGBUSxfm86
6shB+aXC+Vk/XucFeOQP92MeUH3r19hIenfDhCY7RUZr76SNHWk3GBk3B7F513p3
DP4eLvvKrfNQBX2c3+YIzZGew4CdC1I4YZlKpOZEpGgUEKeFVUPOKm6lgaj5fcbA
H7RPUe2yYs+cBMO5hP1OaSMe6V897C8QjJR5gkHZYWgjjpWHgt9Vgbyjla1bH4Vj
5Ybyq1BW2lZq/4Urv4ZstYtaF14lo99WKilD80of328HBPvHGlDFT5CyyO83mimn
U8eQkXVJ/8m+ZAItFF0M/dQDXZ6tGHpRqABy5aoy58g8Nkxutoj7eXLzG2VxXR/n
jeGr9kW4+5IboEdMGVsU3zjWC1PwPQIOoTacs6woIssA8fwMJEtr8coD7YxlxhaX
ZEkpoE5zHrqdHv0zwCmE3ZBANBHj0DRUIJjZoKah6ZdpsowyQeMyiSiOeekrOYPR
RBla1jppp6fKNafM3IjTuLAvpBRL2G2gP5AvWKJHT2R6BgMGjI5mCR6J+0pMmLnm
kX2592OUseeBIql3VLjRcQMnGFSqRsO0iRGAbPNoQezQR1fYggsa1jcAXn1bVL6F
879zOs92/JoccnY6wRBnVDrIMRUcIm6iSXefuPlgl3bgj4+1SzMeTx7z0FTIZ/+C
PAF+gEFWPTaHAANFesrbOddw/V+4qQ3YSFCUg3ciSkfckRY/tDUqSfcPhy0Tfanh
GlMETKlm6/rMAVT1L/XEOQeU0Abqee0/SGjeDykikJ8F4cH76vnFKJgUcarLseYq
mPUOPg2fIoxQRBJHVB0CnbAGXme4UXULsruqVBrKwUCst96HUPsYcI8Cmw90mkN9
p3Lpq8B34XU9JxIHKxegNAa0qMHPwgTB3iuIipndCy7VQKVmAEIlzXsCTznNxqGx
0nxyVKz3PrZWpQDL31J+Py+8dxp+xyePWEE4TCzRROXidiG4174lUyn+rnp1Nii9
3xO6VCkhU/lkSuk6wSnRcgrRPnyYMFe3zBZkRLYCiyl1b1qKF1qhzd7TZ47ce5S7
9Rd+WonH9E+dM2IuJ+DGxnHqhjzke9zAgNNUYMkVYGCjqfjXx3OT6lBKLzlnTr4l
noPGX5/ZRsGEtimdLQaT8ZdXpdBLeoFuLMQwKIUHscdKe8eX7Sg7czZXMiuke96X
O0LhVOJ9Vw373P7s9GBKwX6Temq/6cDPbpSgDS4w7u8YG2Re5cySYCOG5JC786JY
r2I8l/X6LmxM++Uho9Z6loJ/mFWAYkWUudUGgAi1el0wzu0JOQnWIdK2EnSJW/Q3
3AtlMj5hVZ26Q4l7XbZn4HRvCZfYiE7919+RdCGDMtjlbp7dxmjfHqWZqYQjvNGX
mQsqCNsYFHhE42B32WmODXDpYTOTyZh520diT5Sfhj0OJ9YEQvqtte3ogLEzfw7x
UpRM9Iv6T4Qgdoc9g23g+qQ09wF6sbqmcdCmn+QYXOMGsiTdhY3F+8PF1bxJPcPa
HadZimy9uALfhVJEFgcYu+ZiDaSj7jafomny3xvocO2K+3I8YWnrhBKT2Abx8XZA
JK8naQRS0sd/jKpaD6jyYWUm3HdHliX5zgo9TCS1gksTvGYn66tK4/9c2C81j9jF
7dYlveP7abbcKWrtYJEU8/Ubwu7zqY3RCfxdB1bgsYG1YZhlDaZXHoEZ2+QW1jav
qlWvaCSafgUyX07ss3baTpZ68RjHg4O7EPurQt5SN9qMgdjeQsKP06wJKE7773D3
GSbukTNXhTs7t8ys3T2q35XPTyQ29hwWJ28V9q/ewN8xSm/0ZHwlLzIG2ox9RRf4
sPNdKoDwMkbpGqtNhphitJVnzgk+nv6RgZ0aPuTOAOHzk36ajPRp/YtK9RIb6UW9
ZD24XviFU04LnyYbS2DOoit4Mq+BIAP9aISkwnAvpCZK5CxIl1+bJgs9SjW/gOb0
5OsjIXxW6e5H8J/q7bmAqG5zxyuCaMVzAHWjdKAGVqpWMFPahxkz2Hsv5+/X9OIe
KvK5UnAdHCkh2sV3Ycz2Px3F2ls3cOOn3o39a2HlOILZzFFe4T/f8Jaz05GaJ772
qMPD6s14gmgoUrj0J5PjuESeBKd9HHdgiQBQ8VE61Tqg6y4UcpVD/SG7v9GH0o6e
kik3Y8TtEodMqXhEe7mtslYG2Gi/ctcepJ6qa5DUInRtipKl0lqVC4U5hjZwS6vX
SAjYIr0cioO2izz8ZNZRd7UQF3sieK9NTYm0coeuORQZSR5ggFfB64Pm356E6VwP
YgpyBZ5N+SsbncDRkSMjWkmQV0+L6J8RFpBOc1AVPHuzKzl91irHelhS2zmx0Dxl
5GqGeyJTqMtoGmOipnuKH0mpWnfR31KCu7YzFT12bZ1vMDhsCmj2so3Vrgj3EjWn
TgMswQ5883tF6U8uP6vbCKXsgmeztl7o3DT8FqKcI4rKZPs2x1/9XUQ82Pau8xHY
p5ysKZh5wOrzxTX8MP4qr61LOPlkeNCbmULQjOFcdenITYJeUvKtH4E2HOSc2WSU
LFXkYZkOUVHG4qY0AFU8t8gxpyrumaSt5baR9IG1FLhzXxNphe9MZaADXB+EcK7E
w5mH9cTABxVNX6s9Z+NrZ5S+38/ZcQLNAhSujGLTIGxoJYJ31COF9B+EuV2Lv2lq
AWgxUqezi7usHc+goVjWN2XqrF94kp0fdRS9+f+2pGivtewkl6QTY02apUX2jxkk
2Zpo7qUdMqQ+ptjJ4aK314zImmpEzkZwgn6T/DkADUc1Ldu+XidO5omfegsHoU9s
EUfC9RbnLUTLlMfskk6InD+b4Jkhrh1miPL55S94x6zKcS0PTP55ibkz1J42ZZlW
sxKdAVMRaf19mD0V/7+XuNfGZVOhAlh4F7z8y2U9nKtYROb8rmG9ETrZDJhrnLRb
n2ZiOyN1DbBgPsrOTes1yCJgx97N++Nrl5121rUB7LtMmqxnJ3EPBpMzRvJAbrpG
BGb2OqC79FGh/uzisT826vPoDrRtZVa7I1hqioo9/csMd2AksgYlKFmiiw//4zDy
x7T3dwDz1Nj7avIxe56UlYIwF2BBrZWICEIIjL3wxIJjQMKjHHJSgvAtftX0H0Pb
a44+sfX7+ntqlCLZXDhZiNDwOE+jLM4wBQ+++YEs7Shc8bCN0EkIYCiv8LD7CKXo
LxTruIvo32lQfYcs4zp5+yuAfazaeMV239RwAI9uJG//rXfz3Ikjl3ZliuK7xHyf
dZyJel/1woyv9LrOdYljKKQBBexiTeWMdxQLZzOn3UyqEkvLhinln3KJbjcpbvd0
+BcaHPIsecdAglvKyeVJJ5N465aqkKYCu35buROwSeUKmWZTbxDakT5e0Lx4rdQZ
wP4M0zicF74qCO5RbsDqRrZG+uaPVE0AMT8LRbDlrgrdWPXowvGGameOj1b0FW6L
17gVZKrYjb1bayPVyYJ40iIF+jfj5hD9T1weg2SWIIt3tnYTYkWvpWYOgeY5YjRg
gXnil4714sWpm+Uh7I+TXoQFrYDJLPQFGnCx9QEzSgDtzAqyYovR90MP8048ER6J
R9J/ZUJc9eMTs4s7H1k4B9H3OiRXMGX93Jq86W8E91VkxcsJrA1SS/mIBfEMpWMw
j0fGxF4M3SZHVzyWr469uJr3D6rtjI4x+hK2Vp6/vTob51x8EKHimdsY/TnYK/Io
xV7NawGcJyC45pQsIcSwH2q7Se1f7hy/zjSx3Dhv5ntrvn0hBgF71PEMFF3+EcMd
iw6T3Yi0yv+8wq1ysbmV65Jwujh8fCwdsEQ+WErbQxmV74pFoGtGzlV3Hsh1RQHY
tGZ5MFhciDtmyZmAZxoTWhJowJY1ZlPCduGvT8r097cERxe25+sLY6G39/S55xf4
sC0hWuR8Kw6fmdrwtBLhzq0/x092gXKvykJj1LVd2BALBq7fHNNgWpNAvyiSMNDG
I/MCQYPYuQFrqDO7ZO3sDEoOcCklvf6FJAPlf1CBwUXNPNSijZSYrGtwwEQP4aj6
xsMWr5kRdheMknqpGxcVEGhVmOwct4pfIN6AW0tPzHglVYmXzjCywKQDj7gjY09b
YfhpdAjGgMGiALyz8EqXe+gtQl5ld4HXSZboey5mmgW7UcMUsI6D4bSpvoSp/Chm
voKb563Un9emRZa3bE+xVQgKXnRyGgYFm/xLFa8+ImMpQdobVm5Q45hAktY+foEI
ChmcWVM6VtPpm6lRAp7I9MNpMV4Wxq8atAFrNGAuX74zAm/9i7/5gDNOUiKMz1rH
N08KjlsKLY2Xot+tWkyrkE7CO09DxAVAwK6qhTuLHESd3+vvvZYpsiL8uy0FzJgP
9Iue/sp4Z5xTVzFGPdGOfv+MANYmBeLC0U8otPGLaLBM3ZKgvWqULjCSG8rvnac3
tL3V143p28+qwgI0dJI+TsUNF02GArqjPLOSxe6M7rLsNgxSRFezUAxEQlLGabfa
jnWOV3sxVCpyMl4hwF89OslaeNFS7qj87K7HjimCH5yKqgYuZ6rcw2xomdPJDzkV
DjYPJ/2BcSUFkTFonLgLnKAND5llH2/1PRSQMdDG4TMQurTUaw8+4ybMpLeOo1u+
mwTzNQ/YjFHjwWLEKvvpRWgKohFiWbfZwjlRxtyiJQ6y8o9/7qsznxkwdh/3qM7t
NCOhHq7c9gOt02N67Oi82WxZlYPFhD6O2dNpoL/9vYRc+DaEE8IdQV0DIwu1zewC
NTX8EUeD5M6I5bH4KMBEGqa1IAJ+9glqcXmb+I+fqLJtFRbKGxVkIY8xEhPYEGuX
6zo8BGrTwGW/oiu19mWQwt/A/evFTTj6AD9Vc8nkjopnc2S59ypOCg5ukycawOLg
OO9WzF8KIja5UeSICdqgJbO6q1sUisWQoCuj1F4Ck69wNFsHzJBBnDUhWvbjCRZI
sfg2CSHiJATigsCPP/zCaNbXSooEaYnvMX4w+L8LIJBNRzsirUBaX6TthU06Bqea
fx53zp5faBcYjM0tcUXRv5OmeYeMm9jIvDxtat9T7HAPEzSLQDBnHNs/nGpT6zwM
IrLeNVut4jK9wosj2ZW2NszJLyEk2EaMiXU9SDxiV7CPY4bRxnCZFuUGKiOBmbJg
c4FVRcfTCkf0k5XjNLLDDIsJY0Z9lhCjHWR214hQA3MyW9wRFhy384MSG+jI8VeD
jxYmn29f6sm0E11kXhT0Y/E0Z8VbPA1wuZ70sKqMaIkGyKziy5rtQRR0qeXCWmOG
E5iOg0eLva1uLBqV5enGvBsMQRMtiFhBvMYGcRlwURn/L27natfLpTIidyJMPU9r
Vqgh6ENQc4H1HuYjD2KxE6Hd+U0Rq2T793ndTdoZzldMZNPDJ8N4970HpkwiwNGJ
+MaYbJCjhqX++KewLXe8pXNWUq3BGCVlGrFOH0NBWimLXpQsH/bUI/eedkcKzMV7
OK6AfiY2CkWobGt611UjUEQf8NzSVRSlA8gwZlnMORfreoU+zE7zB3+Ast5ih1B6
7z0EWujq8ER/ZMKRtqL3zbJ9vdj+7xpvqd9qU5122B0kBF5YBUmMQVHN8oVfC+wg
D+TBO/sS43P0g1ECBnc1uDiyCQ9wKKXq63Dh5gPcySz48or/vUDGP9+iHmj0Otf8
LY5e5phg6JWpmg7zqxu7+7ClM25yu9mY2EAukbHa9fkSWF9aLq6hkpZndvXiIodt
o8aewXmgbmDMACr9Zwo1uTntgaB4exb9kaV40irY7Qenwkh7tumBI92PprOgn0xa
U/lEcdh4AWpg/7u44Z4wf1FIe4r6Cft6Kn0mO95XXXLNARe24MM/b3LyoKJnWmxh
BUjUPE1bvs7/ukMPVFrZ16Ek2oFULngaGAj8xgboRGj+lyhmBYPElrVOpk75ob+V
PSDJm7iupvGYyHi0pvUoLOxlkW/Hhppo8Q231deYiYx0CChT8DVK/mb9kzXo5jFh
LUh2WNhFRWomEAPNzTeOpxSMm0AsCAhrkw0A7ZtM4OpCzH61ODHvfkAFxMXQqugA
0oT7LYSgVES5AEu5asa2HPqWAnx533i0MR+lERiHPIzgz+GgcZDFv5gHmHeueMF/
fM9ZfaMH/3f7bzk6F36JyGFw3d8EiklIKM+139RrFNMZ2aZLQ04GQYdAheYvEkjL
nd8nLMNA2WrT57cHJlMbd1vTsNnU4AZEpuaCrzjDaYMCGMevKB7eBSePwIHctfZH
xKAtsansSxbYrHjcn9PKK/V+eL+DkdVBSR6Qml10PvMGzT4fN4s1ZEvMxOm64RjQ
UGNBSM+5De61dJlFt+M7iz2hatvDN9pK0nzvIl0SlL1OcnUSFtDHazYt9lYFsQYg
aaMifXwIGbplV2FE5gkcLW5+Ow/pIw4gS5mmTgfrM1svVK2uAX9A6Rb7DrO+J8mk
MdW9Sg8jc7HWTfhsjsIIIn1XBBk+IqW6kb0Rm4ND30i4JE/AbtNF0NQ7c8BbTOLH
tRb6iJacHW911cmlLOWXdUqc/09TXw3qSnGa5pk2h1H+Wo07V7noESNWqEcCpeLu
FGjSyKpxufVScZrHVcnzcaZgKHHPTmJjK+MteElsxa/7No6y0dv1LXu51fQKNI41
aQ2WXEs7eMjBjRk0OskudXRoUtCaR3k7QqHP/xzgE5YlxuFGmlQLy6p3NZ279qeU
3mDu+q622yVgdMuDcy/NwOFHl6DdRpfLOElQdAfiWyAym8qoDC2CPwaDIwkedsGH
4+ppZo+50zobW+vRF4ZqqY7xd08Y4K+GJy+wNurhAh1HdNQEWbEhYTVUBM/rSsv0
3yTBWBNNImB+0ZJeF9tD5shYJJQ9dLzmjUd/5OXkPidm5hX3Eb/nQXpCBT7SB/aV
3fIpXI0PQIE8wecrKDvXi+ap23/cfo97b5lKKi8RXm9Ebb5NGUuZPgpe9i5WdFxO
v7u/ACCjARBVUfYqFvrWGplfnxcBS/M6ElPSz1jrvY8I9VZWh1pD2NQMhT6jAvcK
2C8BEJjho+ol1HtTkBX+5ngk7p5ax9QZc1nS3O9GdNY1d9mWzAyrH2FAqtMDlH8Z
nR0u1yFV4bOkdGb8kFOk+RRx+qO31kIoYyRcWIC7Al8MXFEev8h4BY+mQKClbkIV
dfM1WVM25Qp2uI2KCLLwnQFH1Hz22GOSlRPmk4OXPxJe0WUJxlgJxAMZU6XVCzc0
/iYVQ9FjBln0cyxcgVycwZhlZxbyX9ME4U7Y87Dy/fuG8qVl+S5A89ce6aG7RLV7
QyHdPwqHb5G6/0MaEIvFXV/GkJpqKtEgDgPyzsrQef6bGGNAH/o/DjqjANo9ZVH0
/AcKrnxmfnCR2pz6xe3igun4mBGwRlakXrkXqUgRks5dgp0jv2J5RU0EaMkPq61K
C3rqNApgklfOBtZpz1vv1xYnw8Y+Ex7q95l+Brz9gdJTPwSiK4+AMP5n7DYIpwVh
0WbVCKA5XnAtRXalEVU9hyGeIYLFsXtYsT07SlLag5p1RCN08SZP3Zw3llrtErv+
8ZpG7cNugKyT9W7IfX/mVe+wrUczJPJiwuBQ/SHP9HgETzjI0//gdZLFtU+oyxxE
YSUg1Khnj68yGyrYVMyBeT8S+SJndQFYLpsAESn3s2CRpiO1eRz5ROkHmgpRH1wD
j460dgbdLzbf/uG9mSIxZtpGYWKM1iyZ4bqTZofTPYkhMX6FKqUomDuyhs8i88yR
Ue5SNbPbpO1mgESO1f54ic1oGyMstQZM+xhJ6+VBMwvwVf3h8LUk3d4Qq8IGrTq8
JL/yNKbP0LJi5wi2WEivRNAUmRavizh9dNKL7fV3JqwFkJ5NkYrQ/U/Bb2BT0Ywe
YvEitTK89k7uBZW/kVEkJS60M4jE+WfQi5FE5w9PuR6ft4AahC+cONtOWwA2jqiY
Xx3IcpEJ+YQJ8uprrvzdSEDA/CXvUywNsNW2lSFxgEoMLCuipDil7f4IWhDBrxJT
brpTFU4OdYzADFGRN1KVS3CZ0bVRdEntyCJ/vV3e4EU7mmiC4gmBEC/n9NIhdV4I
xPn9w9lV0gGAuY0nr2AhxXl16OUJ7mp33ztWwMIkWzA6ZuqrhGF13QIqYKzfctVL
5cJ2j14NAsCluDgFYSL0IerkGiL5u16bcRj5UDU9mHqdc4Fcrm+OlQ13sGKmc/Sq
erSgmWRJ5sPQh/qCpGhjobcNA5Mx8uTgkvymIeY8RAXOGvvjKH4Opsg4iBM39H3d
UxYyalNtExjR7M/AuhEunFIJoW75uOvCwtHwGVB/vo/iIhkzTLWSf/iY3Te4iRYr
5OZL2lQfSHTomjtIo7qY313AbhxaC/uOeoLC+Wz+mgOZvvLUMo01Rc3aqTrK6wd6
0f+bRHRRWb8OFca3hvz5Y0ILsydXAuNbc6+64E1VuUHLqx+ysbBg7xIQiXx9eJcq
ZqrQ/Eey9uiJzwNICITBP3IiIq19jdPpZWEs68hiLPo5+BFV7/Gq3ayiU1tlpUgV
1A7ne7WXr6C60XHcT5d16qnrRYezsAofDhLfidZLz3cyWqrfUl0yKpPqW4K6iKq0
e+nXMfqo2NzcQT+m7VHuPf58oeLKhMgdiGKd4E5xUS6ZpnCACW6uJXkyhCq2gz7F
eM4zz/BoI+xIrj8+D8mxkZ5OgiH657fkORuokFbTkmcrCqEoAmNcbWufGfWX348j
F6tt7eYspbYlnaPBvO1D2Wsu55XJhXi0tTgTsfMZHLT3UiLNeFfF9RRm58HafEtu
sK94Qfz/17zzV0byzNVjJylQebkCJFzt7tZcoDl6ht42lOXsZpgLUmt6IaZme2dG
If4p/jFQ4Ky0SkyMC74KHGF0sm2bSIZK8By8bbVaRRwe2wyTyXEPE0agbdRSe7Q3
cAe46N0AnKuYR4F31/7OYYQNB+EQyCUhqavDmC2DQTQJehgnugPXnWhesl0Cel7C
z8qlYHi4Ze+IQGxLdIo9Dtt01snkC2DlaGBtsQ3cTd4cRpIJzGDxQnjayY1LnL9K
2UkvZLNMSz5Z01fN76h3Ln+EsKvHGrCq9f8R/w08WD1K+JMKoEcPwNHGAru39cFI
Y40lWEoBBZOrxQ7EuIe2QRzdhRCc0o/BVwqZmhzkiaCXm7tgNL1aRIgcq/pTR46y
JyWFv2CnlEBfFy7jjeqlJ4/pUybC4PK5FP2MJyqQfBoBXy7ywDimBdAWyQgfmecY
tcQnJMPWruO82nTB84ssADEJLZ3pJY93XOO+WiowTv7AbAOeKU35u9tF8JgwHZWU
98O/EkF4vUkS4fi9UDJEKrhE/shc+I3iVRKF7tp1WlwXFIeI4PGto7qk+o0wQRqq
xI4qVqHAaF/fgUnEVEULeoKbPdOHridOzwvAwmmDwMzqDOGKC3He2IuKEHmPjfWc
GmIc3xGcgOM1+/2vuG0TJ1uRD/90m9/8isBr5LOXmq5JoefCWq68IWqrR1q1CsP+
0icGAtlV/sbw+7AuXTt3RYRlpXPKIf8RU4u1rLcUZj2LezEibakO5YI4OwlJuz2Y
CMthy9rOmYNPtWYirQDUGDUpbelWHdMzlhPFjLhYtk0Sg8Mu0/fqIgxIZNccKI4m
NfPNTKLzCkaRjJMs2xw/gWMrQ96l/9pLTcq0jdawKeQF3SOxyGo92VwhWnp/JvOO
sLmw/6UQn3PPRnCiN0hqbKeh428as9Oc+RB5TXXJub7CGEc1Gw0Ui2qC/RzwG9dz
iEvzgiWg77tFC/+SVKd4dxGeQ4oUIPIbXdfUa2PLtdivy0A/I8172+4Brivk6FrR
kCoQ+I9eTtrYLa+pweV38xW0NZQxKZ9UQUaD7T1+RThFBTs3dgbK8YXH/cGxqXcb
cq5dYuPYogVyVxwG/nSiY+9MczzEGcUNkA4hVnZ7n48UDV19LVXF3X/gI/qXGRgw
TUQuxLUYmHAFvrrmnW6cbq2+axvxihhzVP/DGL/EGZSPaC7jRf36HXtlEo/ZngT0
PLVwLbx98mPzo6WP3mXed9Owl8qDQ45iY202A1vbGVxw9XgDNDbcygygF3GJCzta
ca1LVFf0NzbOc5cHOLK0W5Vdv1ot+IoqSmZJGbSkJajL+E2BK4Y8wqHozWf2MtFV
jOfJRy9883DxPomeeIsSnbDNYTdTi72KH8/M03eXTi17g7qe96bi9g+Fa1FJtsJw
2zuavZ5zUtSKHr4I6Hr4eIblB4pqQk2QUSA16UZSnzvrBoMMLHY6xsXIiaOOrKiQ
JjAHkoOaDLkOgEW1oP2OKqv5FB8NHotA+4Ncu3D1MNgrAUUoPkqDRfYSjVfXrvr+
6RcF1PVtcto3W9yD8KVaC/fdyy47UhUkRZU0T8XhRp/UpnIBrXbqpI6D9FcUrtGk
IbLcLQNDsSNYb9A9ntPm246miFetrsuB3YLk+/K7xIYfJ2MIL5ywEYILE9bfu0kE
qX0z3bxyLB9GDaBOpBoDk2F89tHUYDYyohjNZ8FLrehdNuKww0NBN1DH+NvVEHEX
lsjv7A5dW4HWbfqDnEn90jSkRNiyMG/fot0UGgi3ZZ5jicghvDhsJsmVtXhm/U2t
C17GD+ezwEQsvQJOQx+mv0J2h0hUviLJQtkvh6s9NSsVOcaXnmWH17Tyznn2h4xH
TuIbGdtwpl7vEjeHZibxfgLEZqeyiEVYT53Ip5syvaGX/VFfCe3KCiOId8fVRecu
kMJ5WcYjwyWPkLdGMKHZUTy8FUtsXx1BuTp3tOIXIPEGKBUMp+w1Ijx/ruqqVKVw
EqLYiMX4+CbpsSXLS1Mxlq37KCGjdo1L6q0YtBEKOqGrLu4P+/KRstOrHAC2x9Xo
QDGjiNsf5QXfPKLOgnj3Bz3o2oCSGWk17B8P2hSeHvl1zKF8MY84OJyxIEitPnXO
c79sZzHED54uYJI/i3vPSvba6jPzmQBfRCOefimNn6yqxK6WT+XbW5fP+LjZwMXT
g9KbCBxTTS645B+P5dCSoYbqUtJZ97q9Tubvx6WP9n2OxZCdfbLXMRt3Ct5d3iGP
ORTK1ET1PfYbbf4+4qwJEJV/bj9xtlfbi3BkheWzJKppPyGPl74B3xfCGP56u+er
6fov1oeqa7ETXCpRo3TJEB2D6PLvdsBwQyUqSyUwOsQbTj7SBdzZWQ8R6AlacEo/
fHkIPqr6WuVEwMaYgi1AcR17JqT5OiJ8C4c6u3xALemLATEkUEeQeFbRAc1Ss/ic
3gItbnslPIR4fXV8+hYx9L62oAMmZLLQGlQWxHMUBrcx0A7JEpzT7sgR0hSqqh86
oayl/xE/D3aiChZ6fUPTQvUHEZ680E5JwA2buqN4AN52ElIP8/KiTqIZgUJuON1b
EM76/luFqp3G2CJY+/iOSlXbmr6fhnn/omPZV1xqea1doQJ6oFO/ztShtkFD4lwx
g/4sV9Oef7peq/ZVXcKJGD9IGxVca8qVroL948Jx8aTWCV3XLcCM6QvHWUn/j6st
w8HJdq62Zkn2Xpo5b0tlgBs4hLIYRO4QrdlYdJPtP0Q3NWzhqY2P8ROf5zEf2hqp
VeQHuKc4KfNlGircAps9D3izq7/De19Wv6Jo/eau5utls28TEg2LCw3ht3YakbME
KazrehoB99bCPPZaZ+sHOpqCjq9Dz+WkmioCOKbwnApu1VRJyngDmapwMF+kcTXn
kLRLRNBSR1kbNf6Pqejh/Vl9OBm+OjOZ6xapt7AZOXO3dBR53QczTqNIFW1ClXSi
MWVO3fED4M9jJ3HQKlPQhhthz7uOQOFGMXdx6gEsZPL+xzasmJrIKitX4Eqq9Bpo
VqcEJLFj+cB8sDJFhlf7vTfDnQPQkCJvYNwiSnSjoNOIhE45ARgMchRJqGZ7xK6a
CXxLffu9YVycTyBuPf9vXwt6J8n028VfKHCEgkx83RBLwPiDlJwUuoDi2MxsfWWm
s0lz+ig6fnQR97p4GtH3CZSwkUCTooZwuidiiqM/oc2a5klMNVh1wf4C8dDvFwIL
PSEmR8CqOSlbnf6m6y8NU5XKI62hu+mLC1hOyZ6jmzZXKWt1+v5Z5zrNzfRZ4wZU
+93NZaLz9z2rKAIdDeruV1JvfoVZcTF4BUpRmEQRnxJqtVZYLxCIa+CSBeP5xsiH
gxMhBo12neKmTU2uxyWCQIijDQ0iVbTjrOHrsX3cTTremgGSoqm+6FWktphz5Nlk
jASWwiX/vEEFmcZ7NoVUBLn5ZeD9nLKtSonqtAE3ik9jekGwJ4FA7jCV1hda3paO
TtY3i3v/fWzmnX7DmAyuNh3ZkMhvtk0ljKayJJ+jOwcPIdih6bdVPD8JsgClgwp2
xhhexsarbly6Ogr5PPeODawt143lPR+d/B9x4VPGp30qR1OkHJXSbv6+AVC9IAQv
VfLkIIk8UtWqomTTtKcO4LrYWDL29MsnzjKrDPN9fLlHCGjcZE55WHooT6Xwuxsd
+fzdNmhH0RTglgqtBC73lTSTOKS7rZGcQAtOx9bN0YLxNRmyQ++XbmJeShOFvJ/M
KRIBMVWFKcNOvLDKenAAwDngWFNj1Jl3dI/I/6ptgmUTFzgYNJ+XEtAX153DqI0F
l5W/gnftAkAW4spu7+/e8+SHM3YM51hahmbuzpMXsQVb0blrXQc80UDkH/AwOtWy
B0B46wHpYWzkjnzKXK9TSnP7pKX+pt2sxXfxkWZWydpUFbxKPmfsmt/Db4E/FPaZ
rdACsnnB/Zf/ARxY54N6vAq7n+hWfnCVTpObL+Hz9Z24Lsra+hzsHjycTrtvZn3o
9YEziV9GdQa4PVll3RH6uoigpCeb+/myCE1O3kLgsFp6nTUhrQAFN2jYuTs3sTCH
dG680hfFzKhJWFXA5XcSLn4iklUiV9rDPe15dMJk9oXfZysck/+GFkDGLFgRoQm6
Qa7juQwFHkq283z/AUFDfKP+1Hl3kzUOi0NhTpVc1UvlLs4NvYKKyaMmlYU08hXF
n2oAuwZ4uj6GxqoaKvqpsNtxHkqE4k+3M2Dg5y6Vr9aeiltVFKZ1JMK6ga8J6rX/
B+RI/8tx8jlq7kwS0PRnnz2hLfrkoWSSuR/Ev47TL5xk5w1xCZmZCyajfSPY+ZL6
1Z6oL3DczZ6w/+he3tlAIteYDwpAwC9Zj7MxN+i5L1BldJ+C8K28jMVE4nXo7nMk
J/G4qMz1FsOqrGAcjvO0qo23JnhXsB2a9sFiYr1Kq9YKtP2G32r/M97lsGeK1nmI
Q01//VKuVXUI1ce7wkgsXgO/gl2+LTZ/kuifngA+t/bb0lwQKfilqe/dhMIO0/iG
FA99W26tunSLy3m6w2tTRKKOVOt6Az8Xg/S4AJzEaB/pC8yjvmIjz3nlWImyHOj2
/uCWkbTCdSrBvkt28JtC6Ed1yqkkl06greCSbPl3FgZDkFtCoDPNl6Q6MC6MaszR
vllW6NnSGQ727vrdEr38pXZmCxxEOeQdHMEohA7xApJrty+7vUsPiqlHRyoi0Xqw
3cIZYyd7xkn9QYm4546zbbLSDBJK/0epq9oB3aTqVJqg0tC27EC6BrBw7rjHsUKO
mmo354Eo7zu/ay0xr0/rf8adGopvMNmXY/TXWXo92hgkpqpoKBBEXNnEfEtaDcFw
++EFXJ6rTc1Jwu9tvKoU4azP+hu29YQnFO6WvNR9ra4kYhco/XeK7DPhK74IboNF
yJjlwtC9gmurc7ULTgpAlLkuhjH+cTzUQwq9j2DXdOr3YeWEj5VPV3P8rs2+qHnI
ATEd8piDYOkgU5rgthSX9y025facNbpvZftcBoQPTqCW/Mekj5z4iKDzA/KOVM7F
TzVOfkpLHV80bTRJK6fV2eB4fJe6XHGs6bdkYSJn9OPr53HSMkjZqcHT+L1KxfVa
cI/yGPuJyN5a1TFMIXHtUxp9mBv1N9d6nUSVgsnRWvob4VHV2tg8x0M0Z30Jn3eV
SYR2rJBjEP2DR7wGEDiR+pscFEZ9oA9dWOX1rRDtOG3V3e6/OlyOazgwROHZneb8
Jp9zC3f8gRjEYIW0eCQo82s0uN1NtWdHNaIer5H+fBqNXR0O4RI9VGG8kGqTLQwq
oeY2y+F/gz3lwrM4XXuvK6DXNf8PwS/l6yPbAUbRnFtureeMbb9wPwjLgmb79/qK
CkLDhza+Dr6bsQRIdB6oXz+fhFobaoY8/m3dhFma0cQzmypj0bvN98PSUVqPo+pA
kidRJ4p8+0+BlXif1KfR0RbmWCdY0fvNGXkfJsbi1R3xUYQ8XKs7IflFNAaRnIDj
Ff3gxFnH0bOZvVJO/haxT8r9ag208xFQJVzHuypctqmHz727IJwQMq2fv3Dom9on
mMRD6/w4FfE98fe9DbfRKmN5OQrznk0XN02oaLo4MyqCE0pAGipIXrsj7E8m4mgG
LUnxONLL3/bfu4fIvgV9TY4ZfmVp6Qv7FKs9vB5Dvyw2fEhWadkKTgNixAOHxX9X
Nifq0g3fEQaxHHcQZYHnJcQoBuyLHg6tL5KFkXbz/pjdBbYSkKQJVTw1oBIRBcys
n7+uv9z2e4gPhyVWp5G/6BaVcCT2Wg3SlnbHXOU+MD+jTHxB+gW8Uulva95CyaaT
Nyq09UQKvJ215BDCr+pL6wVb0S8+N5ylGsRePsedqEOKgJCFH5CA/Ri1vb+iM0Ud
zquNDgO9wfMqrheX5zow048eAjcBMlMxg90j/fYRWRsl82iOjojvNkNrhXgdJM4i
Cxx9T+Sm+JS4c0OxG4KIyDfwYGKwaePY85IOdUctVmcGhIyx0VmPCMXDkjdcw6LJ
QFCzVSCHKPfySxLDt8oNEny9jYRGm3n6Kg7834xlXpU7C6F4qR/4l3WrQV1xZs+3
38hBB2m+LUvNXa2WWq3O+QLBmY0ziCJREof4bKTiI2hS/RznoXKnYvBNgkDK3Q0Y
fY8NT7YxcGC6kzSHA2ReSYIdajyyXoijKBVphbfdzzmHa3+HPSG+M9/5V94tothK
+idGGdghnkJ0VSybwpsBBR6PBJ8PvjcHsS7+8dFgrJ14mUl8pkj0cKyZpZHkA/Je
RtVub0u5IFSqUR6pNuEbTONAt6w5YFBg5q0YR2DOHOq1Phyn2CtTu1KpepYDTXIi
n/nNI9AnvTulkl4PzACoz6MS+g2xChpVZmsLl+s6wxhyhsy1gGZ9FnqOIixPZbHh
dGJOPClnvnKPHAAQ4LNyV1GIW2hO4mBwkMQVCZx27ehWUWwEhBJDxzfd/M0dhq91
QpuupZBQNzRrgaMBkoBViwhjaVWb3F1vVOYUKDvXsxhLWtiVtir7ThxkAJ9lPJVd
XwTrPoQYxBsFEY3EcQ/0+aG7s4MN24IgRLYJIdgkmwyru+Dr6TmUNza+S6kMLXGM
lqd84nCrfLLSSdqmYeyZWcFiG442oamCUSiJFm+3R0zjttVRa6fHLUzJVc5kfsWd
pAooF09iHZoqebIgSNcm4BG96jalQrvm2W72dIYE7YHRMgpMi+kCPSi3XS4mkEzX
N3gpCloXHUd4Yx6FhFWJLlFe2eplKCRG0Y8SSBguNle6T218D9mV5G3aNyd6gT2w
MfbD/mhFWAz4iZSPbUzbED8tr7xfh2DEEce9wsFdSSvLt7dtqVn6EV+mlvXtJz9Q
2c//qCUA71/1YGdtK+dk/wNJ8yy0YJJs1Pb5h8ffYNOmOGj15migiIsbxzwrYaxD
WiFxnhq8GJHbQMinerF0DIblFGyU/AshlShyUeWpvO44Xhl9+jGe9UYXcZaBrseB
W+/faL8FTujLS9D9pjzEH0C7fyB2P90HnOBen4f1AMCvasAuMKAktO/hRdmnCRRF
k6bRmAtShlNFxjYEjf2dZCspbYE7y3WMIKi/D2nSXQxsMFHSwNsy7d+syL1KyFPy
+YIPIokePKUipyU9ZwrIemsPNJTXxKo1xu3ZYSPyiBA08CjsQyLNTdbUhogs4RX4
3sJJyJiVgYNYLLmWGhr9uhOL2A46Ihh8QhwFfXkKk1rs6hHNadcgFaWWCD0a/cz2
4jgH4z76CU1Qf/52IsUdeuryUma1h2TQm78igeK2AkCy+v4kNSF1vjpRR+JSx7/9
uXJ88ZJ7YFs08LoTgzM8jdA93WIwhTXaDLtsQuD64+ZedQ1kLyih2eokLyx4kr2s
u1f0NFhmss7ITA7cxZzq2awN3htWMzj5WpOpFPhhIJbxc4yzKNmOzmfanyCZ6yLT
xHuH3kWOgyqcWVyvLI4HoQlVotmeiBJWSAnQIBFeaepfL9NEKlVtXoHdPGZ8M+rP
lxjhCimrtxB76PzTJRkerBXkQCVao1ep7lXg6aIhDwS2EUQUzNj6Da5TIGPzijlm
Q/L7HQVpvq9u6yV0e/dDAeX02T/ahaUQ7Tife6TMeukZgQiDaTnvdUiEIgKk2Bi/
6Sk+qeUUhMy7KE9SjH9+CZRIJ4nxW8DvOSw6VRuNfNoWB0Aocz8iHe/J9INGrww7
I5YSmocApOz/9u56PBluN0bVZOFu0WaOKus7yf1mpl02W/utKQxcRMSm7TU0CVnP
22LDsETGS8jpMKnxlu8XK8NzxqZy+7RE8H2sdnsIX1zSFTs7OzxaZGBh+k/6bIHk
2M0nOJcctLpV3FJYUIVYlxTrM4ftQChhzk8w2B//u69ebEfwjqeFan7o3fOIsrQ3
Na+39tbxzGzPm67yX4HG0U1jtHZne6GWJ70JlNyjb6CztusxlVyWFVigX//x66Vi
e6LpkhtPXEpXJvL9qoPgc1Hq4KG/EFVl5Im3p8Dt6vKvI0W7nzW2cYUB3OV5gulh
oHuH42gvcATaUXEZNdbUOh5Ko/IstYleynH1Z4hcUjHEwwn3ZC06g7D7Yw5OfE0L
cv5N3Gh3SUJFFPfScmEtsiVCo2cxuS5974n7WM6zIFCIj74Lzx1vi5I07fek9fTM
VszUeSEe1XGiryvsDV0/F6ZIEmJDwrOH4Cvj1T6ob2yTfcOyHwtMfVchHp3/USiE
8jsa5Yo3EFlc9xpfHc6RWGwCLjC68DxaMaH9bI1/97yQPrjXaGvA/cXIaH49B/e9
pZvyiQaGc3vYcKQ3CveM3mvOkz/MluaCm1GMM0PPwZGoCOhDlzYS3fomzTqTumte
TgG5iqAnYSmoWvYDXt/1waizPh9MacQqTSvyVISh4tMKfZiYnZ3yvZQooysshl82
YT4ROnvg8h8uDQLvj28FoAGiv22ywW82D5/kOekgH4WkFqIUGGtptvV8GhQvZzgF
2FtV547cUzeC+QTxQM7Nr+g+M3RI2/GDsZ5zaj+A3AWNzx1nztgkSFLOVUJietjM
hIPx1kDnJ9HpmdY2BX0hfRnVXoE0X86QY887ZdiYVccYFRB36XW2oOQL5R3AtC2M
IHkREmdNACeafmVni1nyNso2NzeWjwjHrK4ZvMRYAZXr2EUhmnPsXpldS+xScTLe
7OIVAE1T0niMufPP1DuYSgVXMVXnrOBQD7Myn+OxYCrxoRhKc0dfjmfLXdBgZ51Y
GMT80I3TkEfOTGedxO2ELeiaH7RMEfzzttGN2UO6tGyo9Vq48/uEjhQVzy1jjYdt
/y0XhHK8Ip+5H1QWFn8XU75DIKWBekoCGazu92ioK0LDnGlaWP2h59H9NPpSPhp8
lJV2zQf++fJgv66Ejhm4t9iCZ716RKrbWBtkU+rDjIR0E0fQrJ0cKQ6FBVE/Vyjq
9pkFrc6TmP2fkjgHnaPbPO4KAhfWQ+fIO1LvHpWEDPKAMFv45EuxkRCzmpoe4Mr4
gbeN0H4MeTCuPe9FZC6yF6iDACfgqMRzCEVcMTCxlSGPpMdSnuSfFsYAdWTVQVjA
C/4mR6WeOvNeZ0iX98jKlisS1xT/4T8DqI64R2QaYRfLRdj75fxwyLiwImyGWyr+
QKuWKI+FzdVS0g8VmmRKzKhRznGgr78CWafx7WW76NdRrcEZld7A6m9a8va3Vqtd
NXCCwK8F+ZINb2fRUSWyKlhHQrTMbrtTUt14phskV6wX0KyTgj30oQbQkg92tbpm
cMnFpjQKzXxPo0e4ToFovunGQUAZ6bhajeGUlHpyGCUJgDrJLwqViL+uS/YOIvnJ
aienM11pO8mhu5SP96W6pXWn7SrasIGGBrgNlwnsbKfuu7NJAYkLGXQe7ICl6vtc
kTvd3666/oE3V2bKR6D3m8QgkJM6mRwOI+3ddtE6LeS4Hp9A5d7ujcpMx0jHCTfH
x2sIn5j10M/iCsqI1W9VLEHZf3U0p30XdTgClaCyxJl2ICamHXolFQ000DWlbQYF
FLNwrqo6noWM7NZArdIU7iOH2W9V7JxcR1jfNZSrHxHcvul/MmoyT+U3uHQzvv+3
S2b38lyMtRXgMZipINS+H+vyoraGIxjde5uxc8XWKp9s5BPx2p7/dPA3l105pVQ6
0c3UAyPrTG9vuozYjqmLiX+vuP/XJu9tpAP3tnidxyhhCiK8QX3CvuOYHsHfgDxR
SuKx1LQS9u0PjLJ+ESTJDAufNlyes1F2hcNuaELiNjzCdVRjEu6dBiniJuCvErxQ
0xYF08J1I3bP8qhcNGphROIMn/qNaGfALNG41e3fJPJeRfJblBW/ZKEeV9Yod5xo
yJZ5nqNkADNKNRTNojIvZAEmjudTo5de1vwLobsERa1yxfvqhb0t2INSI6KnkXne
kpx2xppBSl+ciSy9cFlYDF88tiQUdUS6B0giqhPfgFv0lBk7cnCCH/gr6MglOZlO
7EiM3FZ9QV18D/ScaIk3Gp8Fx99Ny8eXMcF+jYBstpiFGAqEq4x75MOzfOSb2Zm+
dIzIeMVzuk3qXT6RhZJ0z01ZJ7eNNgobVMNC19W1X+cPLbtkbJTY0nMemblkbuMK
ArNqSu4xexI/zjMpBASSFWCcHspUqW/x4LQKG3q8sTlaRPba8BA3TT3TTwAGxP0m
fnAT0Gie5Ok2qBDKoiOmwFkT75SA7i1Ya4S5Y4OeWRBfK6gjgo6q1vaeymW25/Zp
e3XiXIeCXKeBWSXEJkhaOEkLUpwVeiB/bK2UNTmV9JY7LzrapLcIrYL+aBue+w9A
6R1gP0++tkBphcur7Gg+iqB+8vTkyyYP9amHlXALjCPb7HzwJt1VXStz///eP3vI
OPQv15xMs1ml+4uqSrv8yOVNAlp6h1B+/tkKzI2zKknUvrif+kyOjNXr9MwZli6V
nupF4fYTN0A9BKIa09LNzoSGF51Gx2q0CihR6PTkaUDiLq4giV3LkCFDwRU7Vg2Z
Cqmap2QqiAx32wdelwPpwOX3U71n4zc46gMWspQJGk4ikEnfieOCL6E7oWZNqoGN
XQSUrTOJ3/QlXOIYKRq42X5hHlH960hHYvRK01KK5D/3gOyTZw3eHIbVTqhhYcLb
U1a2noB/yrRDi33E2Q5DPqREDglO4AQulWHqHssUxKsQld1WMPhcDtbHrqSWAXIw
+oPPzOx1c913frrq/mAekxpRm73Lw3tsHPdUAOXSMY4HQZ/CZt6UtWOcELI+Vp6i
f/dWCBjK/Luud7cbuhYvkzWu/ENYWKh9bXioDj9kp2tusDcYGI0k0buP0Y+7+MIB
LxdLJ8/n7751fe5PHG8h60LXIZOCB5sCmVVvvM25Wtn4EIlzy96fl16WwTLpuU7g
onYVgCkDe8NruKZJCCskr8NVstJaJ9sLwsiYLW1hId89B1xvfap2c0eclq3MV6sf
9Cpprzz+jfT4xMOk7AMb6DmIH36JTWJOYUAsLDaI5mPW8BPqnyKVomFLMJa8hEvk
qTJvzqNbNUI8Ejs+waYdgDfjTXIMl9HSUN9er52wMr2AHZZ1sOUUQsr57jtsAcOo
ogvU+6k6B3O0dm2CtOBvk8Ns7EOmuqJjQ5iWgSB3+fRLJmqL7yi1VnkcbZwoUmUC
My1erWjSvOYUSNoAmscrtzJ0aQ7NJSsubuwEZm93RYqGMEnoCmA9zBd4GEO1Ad3a
aldIZ1icSeG0MRigndncTom5j+aHJFBoyJi4IukpaxFcihhuELQDMBjPdv33bWah
hseQF/63TD7R78idQDbdOjO4Mjyfl8Go7vDVhclqjgdE7Mo8eTPxaTU0rrv0THxf
hk6zshuVN9E5zlCCcaQxQQ7nVKa6YSWjSOVGr28DSGKiLcqHk949ExUJHAZ2TZ2a
ny6ERIPX1+/JVnfnB5MMo+M7zAQuzQe23b1U9uZxXC7zou+srLVZENCiYetvEvgZ
vBCF4ZalmOhH3HL3plqTEZQE3AusSUmKPVIUf45V0PvzVbcJ1hVlX9Go3M0ABDXq
7jUyGlCrzWSu076tcdzUY4chOWslLR5et9rOFPKGJrnq7WmZLzo+wgTgnYELBI3H
kqKTNFSHXf24jU0xaGNJyFWg44buWgHegJJtWczdt6aquSKNM4ClsNGcao3pwv8d
g/PKyVdXuwjkiqTxg73W9VjmAyR5BO0vQUvJi9wj5qFm4BKTCq/uEz/qa5ea2+Zp
FDa3YXxNJMGnaEwDipsLGLi2fYTujrPAJebI+5Lpw/+des9F58EuXjTjeaY7Zz54
2ulbFtwRA28rgWUvbD598uU6Tk4XS30hYI4PsWmdDhT2phdYpNx7tssbaLKmGneb
Rg6BHLLOPKtMLoZqEWnWH8+YN823yfQF+2SZsOdyeu9PVW8onpanWBW7PqmT8s8V
AaMRsuQBz6U0WNHbILVP7jcr9Bn9MOSKWccZxEXRwQohufj9nWZV36NTWqXPbxfW
pdfPeYGdYLt3oOW6uM8W3O7zVmjRGYMypeCrvVkC3XzYFu1EZA8diZ4bSIZEAZ9t
QUOe9U5CI4itOwKX+IGDNXYBfD5WE46bUS/oVIclclznO/G/uow4B9D20uviG5w6
04kTULdzOgo01XNVAnJrlOW5pe5cMUQdMhUENO/ecXhbBwLxrFCgrzspXOLdkjk5
voJdD8ujXvsufhC+MMNA7qEW+rblOb4pTxB2AkBn3BXGizPKK6KAhaesNROA7Ehl
M5y90jqM3Wwak+JXAn8rNz1idBrrfHfMPR1iDrY3OD0BwHvkJ1QQUjcTPtsq40YO
NGKITfKvOWGnOZcULyyhPoea5PShKAjKrKZtt/Ps6grGuYKq7gpOhY6DKhdkQynj
IkVfhT4VXoBQSKW1CkGcpSjeI71SUpj8AgnV8a878aBY/kd3HACEJ1CFwCQHgduQ
iAI8HSn3aQMjdQCSFbi1A+4E06Kh6FmEvvaYXEYLxcnyaS5PbtI4E1KQT2xcVacX
ak/5vqbhw9qH9v2QATGD+powycl4S4/9zzVTQ41UHklVyos0TQgJKfOskBINR/gk
lSSTQF214Jri57P6VdxEwZiE6WdYv6cd9iyXIjKulPJ5E1S/w1H+BC3XYpxDhU/i
s5zajZr3MpHhfLliobG+5yUwBrkBCj/El8ZSKrcy2/3U8P6gje0DMs/+rWtSnHmk
1o0iE/joGU63KMo5bQHjBfqwA+iOQZf86AKNvBg1NZ+6lhG4JRPn0zecgASVdmKl
xvQgHGYLksrJKZv6zrkrAxHFqK+N67D26R8NuJjcEyPTnEmUz2GWw3bq3lTEn3JN
DUqxg+cgp9hhTOT/wI83PL9k0n5ijZu4s6PYTeFS/gtnQhfReJhE8daPBHYWH3DK
rISl8b92+pbV9uI7jrdqmaGV0pvkiuxNS/VAQCOTUueme1NLnqQGWRzJlKaIy7kV
NQgt3cHJA/UDXvKk/w8EtSV2FQJ/wlDwumhomybidyseg1MzSMkfdALI+AvGkMLa
+G51D6LkktGPD0ZxXvDZaqY3d6bj5dVQl6g5TuSWYLK+owWhMxgMpS/IsiWTxKl5
CqpXBVnTfX0RnH5104l8dFyRmQJTNvIUt5/q3H+/4NBCXKUtXx4ll8CsvHdbUfjt
wPv4faU/QePGegcTItCmiK/NjQg7cCHn3IMvplZbDZ/AsL3+r1fesRlx/hIG9Dkp
7oZLWF6ICG21171MP+PnnFw0qkJWkrjRgIJC6BerKTMHPTfC6RAPB9Cr4i3wY+Qe
qVl/PGheHsR9lAI5lJKjZ/sUAg31zruErD5Z7mWBWyB+b+d2bdXLikZI5FxiA79Q
NxGoi9X4oqeot2LPl0ZcyiDiZHBgLdE8qMe1tUarvcsPgZV+JxwDC27aPXXDymy2
UWQVM+2rUtK3UMoJAjmNj/w9k0jTeLY5u8TrUXpBs8PsHqCVXxCXFgBz7ra6l1RJ
R23vbfcJ8z8IAm+Pr9RtbKKyXNlAInAlx9vdjb2OgQ9wHVujd5C6LHaZ2nvDs9SH
Lsnr1JD8OVqzOQfxYAzt58YCNqYc1PUdk3DUH2oq4wffslz8bvz2N1DxJOKg1zos
Whdy0wIwnMSEohwtCgolHLLlqaZgwczl4q5LRn8pN+8tgODjiYWPqmTiegGdDuPI
tK577m7FXUzmU/7jQ7FQyyL4ul3789E91fClUsyGL3ePa+b2tpJZ7LPmhdAjB8Uh
JLieCGzrqBESBZ2dVB2yj+gLm+zlGvZwyNrRSDs2FGKkcHsxnnGlZYD0ltZKcDmC
nVS15hs46abiUnvUYDm/29OFLvY79JntQdSjYjNkiq22Syir6K5g9nihTtfD7f+h
rFtltVsQ8CQ+dHRJ3fKhOWJwTDl9uLYSvjbKNLArF1MvBQfPwcIK5aKtng32tdgm
0HklCmVu1IhHCQzOJkUE8r5xwZHG50yo4kwHfF+1qYNKUDpAfNV0e1jXXF7z+GPt
aKR1tWvzRTmnn0g9Q2tmMAfAS2dc09KEw/L4VtHwrGKK20WMrDXKMhGdVJ7/cYh2
cHFo+2uo2r++RKzV2nNq5AXRos5AEgB4hwUpRdrRYuKS45R4mPGn+0wFZ6+J3Inw
7CqIMW+2HbjSXL+43gB1p+AWKjVu/YO5AFT9v2KJvZUYlfS3StcnwMECiyQ38a/z
j7oCJp//atcD89l9HaPZK4a86/hoMece4czirIlRd4pxshDLlms+DlVSlaYqyXeT
M0y13Co+ZNiCDYgt1BvqYASYwlqX9muiq5lPTiQ22PvdaCzkC0bYoH3z6T8UnmHm
Qh0hFBEooJ+smPqKgaoqjQhLmcq+PNMMNt2k1hGIoYBVudWf2aqtmqxXQHnfF0M5
osTKOrVB4TkG0C9KUU/+BE0cjyE6BKYREpEgdEy6gXVcNk6i4f50zIwq/GwFF+XQ
oEnGlckrGlSRKnafQf9RPYkriKZSFLyfbBmFKFChWzZKIE2cOzjQPONKzm35TBrB
B69tfr+fkFLKxMo6AQNTRixY1fiUUko5SDPC+PisbbM1tb+HLSRUKCI0aE8y8bWj
Zt0YygK4J5PmuJ6QSeGLXYOkN4UquB3JT/Uj7N9OgWWstfqZHRrS9tc2spWw0vCF
FSlcAJhEK2qWhSBXdbSoCGc97LbjiB/blvX3jOlImwMhonpqH58LC/H+2yYSoNAb
tU/pFDI8LZNam+EdO8iLZR+G+dMHVm8l2bvBG6VRG/RIyTYwFYfLFaxJqa6Eib2Q
/j9nwk4YwnYLpvVCerT17udgCmS/Xqtsj1LMSsyORtjrxoyYeuKcqarOQ6BMEZXW
uGhwgJe4sBUjH89QMfUNyRIBeuT8GN0Jf9T13qj7dqFnxVk2cBD7zDTkWW0NtUu6
ODAK/ZmKaepyAF+d4U6tYyk2gGySIGzju059CJaE1oi3STQOd+xC1dfZPK9yBN72
mca9Ocj4JcQOMcZgmLCDNsYzlFyHRi/dP5bNYmnFmNCPco+kYkvuCClYpFUICrbL
7qq4fSm2N5ORZWBgoRBM5fKZ20Sz7dnlAACRcUR2cTLUmCRMCnMW943aqQS4DixR
nXdBnm2RCBSs5sKAZBlkc2wtR+HiIzUS/NQDdk7k07bvJ19D1IDLI6O+LD68yWGz
d+6+5s6syizVMYD4x8MdIRtazF2Z3t0Zm9d9GkUVKbI=
`protect END_PROTECTED