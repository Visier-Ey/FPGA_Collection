-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
--pragma protect begin_protected
--pragma protect encrypt_agent="NCPROTECT"
--pragma protect encrypt_agent_info="Encrypted using API"
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
--pragma protect key_method=RSA
--pragma protect key_block
Cpx1zDCKQUZr66a3Ql9n5UK6gqesp6JR65nBqTQe39LISQaCfut6P2gnnMHrHNK1
BOHRNqUMTcKoNkkeg9Hzc4BWKJEsxuEEIb9FcaOaCwgBlAonzBz9AGcTm4a02AV3
1qJR2B++OcbF0R/9s+m5QtyPGtCsaVbak66yf+K/7w9bVw9j6IJUPnThZhyUqdCe
48V0Z4u23OVnXBm9B/ohSdY7CEWhBB0gXS6k+iPsh8ZN9O22d0I2cBg0334ZT8lT
NbVLSMzF7ITAT8REtkQ9eVdsZTwHylRXSyebFkZ5LTyMEDESOeIfR5K+EzBSPrMm
+f+Ii26jiSsOSXf2jXikSQ==
--pragma protect end_key_block
--pragma protect digest_block
zf2ulZupggmOzocr6tDs00IbkMU=
--pragma protect end_digest_block
--pragma protect data_block
R595Icfui3/c5o8BUBqDwn0Asei4FL4mwQaCDvw7aQbE+G6KGtRAaxHl6u87uCtt
1ljhvtXW0Pn/vZmbcxQtyWHwjD1aM36FoJvgLbZLD1NYKkdOGYNZhozbrNy2ZmL0
jUg04OpsRgQHdW75wdY9xK2TcFnA5/hzcB4BjhAf0xqe2bVb+E1bjiZ3pMhvqjQ/
cnapoLDIt2yYdFiRG6Hjf567D09Qp/OIuQoCweJiJmlM5eXe9Zj+mz6O41+PYWFt
d8QvepaH+8GPq+0LKBQ5ERrYnzahUOtRlP75j5wuLWFd25GBvOJ3rt1bBV6av1nl
kgFfZSwndFEIXr6zu8h8P4Du/WQyQYhBuos3NTUkMRiadUcIHsC3plQQ02iBs6rE
bFykHnB0U3sOkmrHbnjAGZWfsvveAEpZXi3rV2BbOYKYdpmjtf2J5fZev25JPJXT
fg3HhaS0N8kPMolS6JFKebV2He57GtHZxAqpuEYVuTcQn4Pvq2mbXYW3N45JIjO0
pGFEDfj1YDiAF5JM9C7228Q6ZJfG4fHYAOt+FEklhcRlwJnlER7drlHGp1IO6s/2
wdFRjzd4MTXR0HlwTaEpQfv1pf4PexyF8jhOqJqol2l8WeK2uCTsiW0g/0hE+26P
wA/QTlasNMK4zu47QxgK36jwdpLEwqBgIZAF9ONCE1YodeaTsofLQXao7JpnWaR6
SARQ3HnNTyTrUV7bR6L/VJPceFePShTYihl99kfZ+zexlL5i6cOUpSZ1FZV3uuSD
yfdhLepFf9C0KFwplFRGqppUMtw46YkBU/lpq5xKCemJ3DPaHARkPdBMTXKfC7aj
NIQYfr/nYxdF/kaAqxPlH40KC9YJOvUcaNmSpyAp4Ites5b8AFcoX0b+Rkrv1Xz7
h9lcpYCGx98lkrgpYYd1a3bXZl0B667iLgMAHIez08qDYYI6Xwp2P/QY+glqFxDB
RRu34h1h9S5SP5ug9IwRBZs4gWtV3ihy3rGaVmJYqc7ct5L0l4/C7N6YHSsWxP+d
2DitDjvNzk+WZEpDpJQUVB+AYWmRYUKN4DG5hiu8oTF8sK9q4aR22XrX18+jFKqH
OVan6qm2DkydIZe8MMKAg1qspTokUsQj/sBsNtL1KRXY2xvm8EobR+8qLjmLczKG
OU9PaDItK19Aohz01qhPPkwd/Sj+8E1qC+nMyfEB1ywBU5qQhUg21CTlnT6+qIdX
Jb5kN7TgeC27DyvHhk+4L2gQp3ZU6xLYEcG4XCRxOFTGaN0mYWAOVTZ/x8txWcNe
8egWFlctdae9vx73RmqXXGv7CiFMDQepNcO5vkdQPJ3Y5xhYPJ3NTyPhVSoWVAAs
i1lPICrgW7QJCxhAC5susJMLVk/9NCiX9DewQWiVm6uV/XiiwPv9wrhK0ptu7+6d
1CFoRlAGbnO7ipUX+wFVzjViU/ZpduYT5OkZbI0fVMHza50Jfg3kDSogRPkItZ3F
KiuOohjpjY6rmPovbsGm7YevSkMaxW3gcPtK1yq8XDxe80jQX4EnZ9j949p9pN9N
lmina6mz04WIUrKQN83z7libaDN3KEgZN401431fBsAqFC9o3nB1FmYS/zn5jzqO
dByaLVs6g4UIuwhsU/+xGxhvwGy8gBByZO+P9fMMYSD2Lgiu/cWhOlITvUEs+wIh
4j3Vmg04an3YDMox3RQvPrirADt3yT+PzYpMXHXhwqp+VTS2KF3SPaLSE45hm/1K
+4jjEZ9GCE002OnO6iWmlTbW/b6ESce8QcTw9WG/9YNnHsKaZrLhzgw0qaxLy80f
xYz/mZnTxicF29vyEikpAVLWxjbKJ6FTPRv3pI+0cpPvEFsEyyCWouZ7twY0/I+T
MFiZzh2u8unVF3QNxOv6LQIbKjkiRCU/8uLQamcTQEtYkfK+ZOAQiGUkYqXi0JLq
MiOHO94ZElWVblACFBIMwBfUyKAlBwll5LYMbl4ap8eow9z/ZcGGdYlUf3ZMz8OB
Gey+aviUqgHBBjHQdbj66RtykwcUaXZXA6mdHNNFDipidO26EuWn87AAtPqTURQ3
8brKpYhSZttgqYbklx8RembgDNRu15SE6iwRtkIg6q0/XGq4K9YpAIwjhom+aUsh
jjZn4ieZn2hDi5In+Cz/QL1Gy9E0pfC+UDTVmkygTXIss2c1XAOLuV0rZI1lUjoE
09vaNoiwlYVjdfcXxjYegVlUpBhWK/9AwvxL4Z23e+QSsFmnj+ZV5c8euKFj2Un1
m3H4jKquox8CWIQ95dKn40HruqCZ14gavnTMMsJAhPEFZPXr+JFT4ONZr/YBbBLv
4AEhXLjZDywLfbQY1M9mX8uo7QOzIcrLI+nwrwngS+NnMK/VeClHoXQU7Rocgg+m
IbRkXHhsMzbUo9OsH6ktArKltvzc4q14KAoiHc6c8EUjUaZ256hDUn/11h8gSoI4
nC9PL9Sx5AwncCu3R2mB5HVLt3kgj+42NTpZY0Q3fD8FF8KeEsPm3HIjQvnAA9Ty
QcQ4G2Ju4365LKSiBWz2+Pzp3Y2XSM65BNdWR1ch+Pe+fkoNyeSgnYQ+7IhX84t+
SSmvGCCK8aMWLtirtxwd8ty0GE/3HbOhIO9GzdlEgrfKnOXTG2IxnoPtrwpPTxn1
P1uTnLlAwWT89AQvM0lOAigc6zPJMwzI5/i3HZUASMS6uoSTtsQqFT7RCYQJmjKj
xAxh/2n9wQAPe9cKbEO5gaFPnkBnxRqKlevARBRFIc179yEOKoGpaqjttSd8L+XF
EbqBwjFb7sTMCnM0iQ0OGZy6X6SrFPzbQIx6wFFKlNjXXm9u0vE9fWukkJzm+Wz+
a4c2xZBDc9xr5swAmNV1v5pI9KB8HBv8J4A/TlDBzOoduCFUT26QxzvBoK9Gtz3+
BjFvI6Vj5RYh5ZzJ9B+8K25opTtJS710REovllE3iPnB6TnVTKYA1/GXjb9s3rT0
5IucB5oE+3SOnr/sUMOZFtxrqBozFzmMsGrKgxORdLt1Drvy54Q4tgUaOcJ4b7PB
29rJjFR4OlVpau4CaOaKoJUN5OmeaApraY/SelT74HQ2JBqGlCpfTFcOmuJ/PzUw
UZC9RO7aEZNxQ90nTRgQ/vqj02OmXp13ynRuvuM+g+SIFWXo5BeLpRwJEDXM/KOR
XHBy8ogUCPFhV/UH9jd7nxZJrTjwIRa2YZqgfe7ZOi0/U99AziPmcUq8arupRSxe
JqoMcXDSPFmju7zZOyivY5XH6W4DUPNGSSzJN8+0jFtmuf9QCHJh/CrVXUhWxfzW
jbVRYVutC2E/eWJeOIdsWrtHeEoaFceaETVAnuTFSi4iGLO5dxX1izxejNXZkyDV
Eds1ZXlrVeJjohVIDBfvbwJ7fGN35vLMy/Ahb4Tm61oAabxWtS+fkGCIRIdEeb1J
0Z73XDxvoy+Bn6cZjWRBUodwNdjwYnkQN0S/acu3gtkrpoGrJJXkNCNO32C9dowC
SKoWp25T7RfBVD10Huyk9J6S2thH36plkC9GxzmERS0vrnhm7CJzz+MWmqao22Id
xx/afvth1/a/4EMEp48CJ5sudT7g52nA0S9mA3eUffY92sIrJ/8C2vcaGKqOh5y/
rTG2pwWkZyXN3K2/v2wYOECB5GPIk8LN8F45xRCs4B2g5YmLWgZLdRjaUGtpP0lN
S02CRQDTIVF09aGTr6xkTQzTjRMtau2pJjz60qc35QWqjGvl5hevbnkdqge3Q/+P
nobUuPnrBXfC3w7U0dKoY6rQxBmgAf6t+U3YcfqTR5cmZpHU0CA3Wg2k9LdemHoA
Kap9Km/FsDXceZMksbOx4835SD20Be9egAoj+qM3vu8RAg5Wh9Ocko7E6iHtsj2H
x61xXG6YiBCSAtfonY/RxgIxxK8s2Rcd1jHijX7WgoRDyCm+/nRICit8DlLvASKn
HmC6osFewJZYIx/SdE1VucJ2mVKfLgtqMiDXp4ZUEkZA/7/U8LsbGGaH/n4/sESe
gfHEE/GDC2Otwblu/8k9mmxNFkr+7Bs/7JEt+Z0hbzz8vAODbwwZU0hStrJa/ZuV
QMMx/U00CAW5kcrdCYclzn/GBFFfdFCx4qWpJ5PeUJaAaQu/gOJc4lFDAENy5G45
yF0qkazMRw88DmV0YGdv0/tpWpeBC0A1Xwz/mqYjmdTwUHIUiQyG/dpMFW2Gst4a
mXQVuB7eBsPS4iEPtKNCCkHSqQHAYHrDoxJL9srnny0kGVMj4qBF3DFSDxzdtHB1
gSWGJGWyw0cl7o66A7Io2BzY6n34cd3iVb8IYkQxHbXXyEB8YvzkXxeIiJSzf7CX
A48RqYj9L9dqCJVaW6mu20EKLV/vainRgoAURTifkTHp5KOze2eDrtxpnsCB/ZNs
wAgzmZ1LCA1BIa9DqgYtpi9L5isHOeAgPSZ1EZqdzDUeJ+zwEsz68FqCiCLwHMoO
lEs3c6nXfmOBYqKLw3jOQwoLTJUtxrl9EI/Iju6ZhGOfb2vBrYN8k0aYzuomkbb2
cyc/AGR5RFY2kAaX0W41+39xY1AhpMiS7l1/Ps9sPVV5gDP3Xqfo6tKgAdv7oOER
xeIQ7UbvElapTtFHTjwBlfhr5m8xPlbEm6YmsRZbk5CC4G3T2XTCOBo4yI8AqcNi
nSAnnFf5DVEK+mbf/5Ms6QJv6dpZrRHsCvvxdHqhLyQfcRbE5EnHIowqDAI+7KFp
DIWPql8xru6e8LHDFKjfd9kV0fz20Sk6w1DxTDPQg1BO8WKIVbSiqEg6E2JuZrFY
LkO9pMrzbQx663RqFGE2GozIdPrRHnC2YHdlb0lfLYoxTFai+DhhWukNxcpRZuC1
WBCEoqCc1Fi2hYwO1HPZolwjY3gtx/FeB/0KLyiMZAm29+d0BNgpzEaoB441FuIk
1JFgppppI6Rqn/chaVYemNyRHVeNq/x1p2hywxQc/Sa4wv5ROfGqboSFkuQUSTw6
nKPq34Q35vYm+SvYK/hIpHumTneBaCc0Jx4bacDU15eEVzgT/Ne5CQ0n3Y+u9GGT
YeIKD2j8T2NXvjCSrZuSG4PBThw8wjOrpS+NzKrGzQbmCxDGHHxpir4kyeVb7hOD
k9n/K3aGqqjxJK28/oiIQ5C16B8/cTP8qZt63i+vGavxMwmAyy+S6ye9a2F7d8Wm
+16JL5Hgg0pucRbdbzM0chhhVC79bjLGVAALcA7wsszBQ3f1K1sNAREwSTnzlhMl
TqchY6CCQSfJ0+iYNtUpzcLEwLYVrNcPfM110xZ+oqd87fMNJ9xB4YtTJHrPvpZ4
O6xlVhqqKSvb2HPjS3QXyYkncpxU9QrW/Mnj9BLG9Q1KgJjFTO+Fw4NELJTJYOiU
M/xD99waOf35g5a4tLu7BYwRBbhiYSMF1I1YtnOQIh0XUWvGAeKiJpSpeEg3xHp+
JNjVuZ5NHK1hKAXucZMvSGAf9Ec6c2F75sfdC7uu5yzzqP1c0qleunJdk7Sdvc5o
viFZHO3d2z0z1wPnLe8TD+Q+fx0cQ2VaEzt6J8JiLSxoIq5TnBfw6oVgEhVYAqXq
7gmSCTMF0PUBLMIzZc/8FKozALhfOOdiFqWYJZEK5C23S2cicUDnG4gxjVwOMvZk
8ZVUS0VtA1WpqRjESpT3Y+Bfm8jxQnOhQ3bKUd94YJpWKZzp1F4BzWsitbIBqlNl
SwyScOcFK38sj0iS+Os23y4Ij7sOS9PyQ0axLb1L94ainPuyvMUon7X/4DKq5KuK
jJnMdrXgfc9EWH4A5dy6A2QqAoyGC6Jir5facmvDsXGG8OdkkpZ9PCCRY5sVnA28
WNB1fQ/ksuJ+F2fOv43wpSI1RKLr2hX9QYVDG6QlvD91e09YL9loCq0rtNrNROvF
DO4ca9VcqHDtKZeNBUrBAGKtonWyPdn0zjjtwpy5fhLJmtEBkKBW+U8WFhsiuLZL
0UbSHfRcU2eYBiMSX+Iqokds0M9+82md531RhTi8OZ8z+JPru8PqC+TUqnCM6mQb
LH73idpSTDQyBPhrgI2c14HsGg1pVSCuelJoU/GLFN42+ICl1zaXt0ehZAYFXkLN
faLCbPlJ3DLl6gIlkXcT04cBrDO0vmu6b1I418j8R2AVIR8h8JycEZ/0xWaGoY7s
C1XzA8oEUH1F1B2FfOrPWbyiiyJq8Eg3AKNmx2snGaPYUHl2vjldegrFHpbeDXD9
g2bU8h002OiNv6WB72OI0o92ExOsOFsPdnwJ1PClncpV0IdrYvFAoTORy/7wjQoR
0gjG3+Owvxpbvf1IHtNYFznRvGwP/uNSL9kSZfsFMAwlK2tVyzz3sJwA6mDNrdMn
XU6nf6Q6NfPEBwlhtXNmOZitMoQz30r+zyXaxhHFD98jtzjuSGxTuueQO7LggBnI
sqMnlhFsGNxju2bdNrWkfi8ZZO8W7EC6/hme2gK/DdC6ZFyix4sS+/iJA41o00bL
/QaR3vazkQRmD+to9cVlbKPqXyj+LO4jI4URQhmIws9xqsr/TeVlsfu7zFU56B+j
g3K7f8SWZLCNWX7sNPvXmTjRL1u7rP1u8Axl1LjmcGJVIcdwHzELCKmdrax0PXkK
MvRx97lu8NH+/SWj/6d1AEStDZQ7RB3JDx3IwAh7b8LN1i0uE12dWI1ONggPM7ac
R9BJrn/Zt+iOBWrC+Gtmc12CTIMFn2lYeZHi0zkQgxDCDM2/ZXLtghCFsPI2NZWP
Z1eXs+5S7+qZN4xZk7XL1z6xSvDTd8kfm/HvGt9vfos7P71OKW4nZoheD//isTqT
+SmZPh4HZw0IXLeJma3GiiSa1QzcCq+QveX7lnNEfi7rD93umhM24vgpYDfv6Exr
NTUw2zj3D3sMOFvabuFtFcuOpOYjUs19rMk0XBFK/2dFwWbFBLwUjjZZkYFQwT1J
wpcGuuX/oQKGU2OUzOn1NoY510QOaBJY0BooAdGyIrammojpqM0c1qRQBhmh7HOb
ZJ7sn84O3kCu6FHjUDBmKEmS2jA9WwNG/WXoPpNAZYBhvQ/uQxIV/tLm2nj06CVX
L/r34EYBd3w2kANkou5MTB9FrNK2wIP5KN1xd/x7fF4ttZdmsO5TdD32SzN6kJrw
x/5nEubXyKkmnM60ZgbAEBOJhj/cLqM58zBWH9WV4sL4ADQFB7c5kuSlqpZp1Rqa
BwydMcmq+8hxKCoL+ykqGSL2LS1Bs+dvnTT+6uhRjB2EZxiN6eOJE87QKxfBOXUz
phMTed7ipvzUf7ffhEfuXHbhrIkZakrBZuNv7OkEPKJtsR4JzWdl4KVz1yfxYj5O
2E5kb8MmNSo0vgLx29xS5USFBwZk6tSMHEnTi5/Z/4xy6+KKYbslmAR5eu1z1+WN
mMPzdOmUNbU51N1h75iOrtOuFSeiZqiFfvswOVhHDf9PNX4NrRdQxE3vlqH1SS1A
aMrM6P8H8ivk8YrU86yyT7YxqmTL9jSDgvmmgvd6LYXjlpqqEe93OTY/u2OFhv79
eoylac6jAlLX0SMhP40s4bgrIFv44Z0aGZE4VvBXB8fg8cwxKq9pVayfxBWrkf30
/p73lXTkBuyx5YLEv6lXjMArVqFQ2pBxy1onzP1xLaJTddDrQEsEULHouPJ2zr8h
szlqlvEWk2wHS/7L04LtgA7F9Ci8pEvPSpI0XhcXVVwzrX7adlxiUpHYwLu9Cg/I
aZoHtovasOjBhHlgHtc/bEIgAxRESgXfK69kaF0FsGdaGJ+FeXi7P1xTtyTaaMRi
zs/aMesV4sKySncSorQ9IZBWTntMUNFYj9YrxdmOLpOd9QbW6Mxj7JU8YegWAV00
EpzP/z01nR4TCmjhWcdt7inLTWoS8x4bvxxAroBKbPsmseb6SGIb+DQ3q28+QjWr
FnQBSwvfkKfRUVKNDIJS7yHT19JUrcXcmGHuE64syvwe4jOjZFDXh2zDEByqRChd
dvJcauC6aWjBiBIRhc0Scuaw9xOQ4lo/BXDNBkLv5n2MnySYO+RMP95vtTdOy6Rh
Xaf611yOi3C5im3EQsW/VwYTkN+bA+ve1pX34381t7HydjGoTsKcH4dnHm1k2E10
XryVZPOXDoVhs0y8hfGcmbLtkICbBA+DQZSVuO/1n3JjGlgMS9YVLoBhpfRHVIM/
kvazAbueNpJUWHmZE0WCk/KUIKLEKPhNKgGNoUOV9yNbo91O+gSRiXPI65S8HP9d
ZRcDk88hHYc4QIakYilCVfzceO3r9RIFhQIT43NVGkT4hHub1NYx0QraTVJcfhW/
LW6bMbRbhNX05VFFxwLGiQenwUZy81xXe7Wg7w2EycSBkYqJ17AY7CoS54QB9jsB
cjNaSWhYRQkXxOxh49sBopt8wJCX3Wt8SqftIzy10kQJ9O6TsmOHLPOKBJzYoz0C
1+Xu63o7Ynm8fGOLJxneycYseY4oOma4EceZpmWXBxzdw+MYBYqxi0/HSXgUZjXQ
1dtOJc6TEn5WUhNg20d8UGl2QWT69GJGyA2O97DlHJ+BWgw2hlwP4SeC2GbEsN7X
eLBbQBphBhe7jNtgeYisnKQdftHxsJO6kLE7mPAMPBcW2ZzehFrobGfLxoJh3EUp
ZjQ1+qz+tMV4Rc8VbByRDiffBREKU3hPt5g2Pv8jsWzQxmUFoicod9k4Npn6+G+c
ZUjsem3xDmKfvtH5cy5MEedZSZcbFuWsuoBfIBBYiZ/9fQxh8H6q3QNi6G/ZI0eo
CqPwCWb8jN+X9gsHFe6Nx/cLgoZk9y3pYBFA5OG2nx41VNNSpVQgHnO7HUysXzXS
+eaectDgqai7XyDKK1xRebDr+jxI9xn0Jm6ytRP2SDKwb+JbghVc1sxo+DbIuEFS
--pragma protect end_data_block
--pragma protect digest_block
1i2fle0OgQwnmYcQZpPTCQU7ISQ=
--pragma protect end_digest_block
--pragma protect end_protected
