-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
LN6aIpEVyp54rCQ7obzEQsoDqv4FhnYut6cTI8sLfievVS5vT/OneU8mT6p8y3aSnU72Ejp/qE9d
Rahv9Ia/E+Ew6+bWS0JQg9NiWuH9YD+tiC8lE8bmvX7FuUIq0M0kNXojxX2HkbXvemcMCyMRB3uZ
Hgxj9xnJ5fZDFQbrEe1zcxkopqvTIORQSoMUYl8IurWwrbubp95EmVvPu77p395GmzOiiSv9+43m
Hhvz+DEX/kVMRCZ4Sv9GctqFkE1RSFUl2g6Y/rxC3Wh9uvyZUKD55ykQf5tp1kgN+5vvqD8y0GJU
GQHZzitIZzkaIM3sjrrr4QJ4+03Qg6CHFQ3KJw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 11552)
`protect data_block
e0/swfQ0kgOnJiSDWfJPPYROkkHe5R+4Mljap/1pgNA9RyfG+RCCdBLBHcGLcv3BTa/YRNB/9dbs
q7F6lSraPcUxbSP58w9z3hhm3BpriDmO5I5eM3BTFVYBIMtZjt78UpnPLW5La+M09h5nhk0Y13o3
3SJpXJ7GnhvEnVaE4O9jygDQqJtTWpl3jSEgP+v2cJoCbjxOfJcsKSxP9/V2E5JsO7amHD3vwgYu
XGz0TfgxXo3MoNdKwpTm1uwfB9sjy//tCBYJ1D8mvr2ZdSPGzyzreX5dh/Zc82msnoA1soW7iLxH
Qlmoz2++XkkKzSoHhkLb6n++Mhq+bnjy8kqIG3B48JarEKKKhATdQOy+hOPLZypakxI+V7Gald4i
GzxK8a2HHCv+SvGuAyW3Ozv/e1EOxmIPaL/TZ1fgvmDDQZGoXJJc34ErzjbeDQsZZUI+x4JDT8m7
CAbavUnOgBUkDrF9ABhIiaAJwwfGRWtxnhmWG79gX3VYyJCFAYUxMNCKkGOb4R9mAOmHxn2QHyib
q29ZSnCl/RIyiyPnuiSlkCxpCrI8nbc0DkaQLbmN0kRUjqN1IAb4DfyJWamD9SeUUkP4tXlT35Cj
f87G14CoSj+vNhJKSudEmNat94Q/dkJ88iIjlWekAhLi9auYzwQ8bY6HuhVITxINb4Uct9vAmy6T
VvW2c9z0kScLkog0WM48WfneoMHJD8wWP5qyAkVm4X3tJLsVdoCYFyxx6DiuE15pT5lnOOyVZxMj
0Ku5uU4LRUOqWFAe+TNdBA82L/Z5lpuTf997AxZyudI7SvwYwIbYQ9NFQlxpbYJeHJ7YN5hG8Xlj
pHjCfa2ETj7Dp7Fw70p8zAffy7jQZ1DDhrs8R16+ripDfVd6WJHXV68hGBOnj71/DaeN8FBzdJLj
4CbpVcISFLhNRAk16PfLIfczpQiK2wqQp5gRUN1xMAnAXrEYe8eefkBYwCAUGdH7aWF/CCgU5hbA
rH/eActa2jUqS8tbcfJhhT1TPCuYgL/TPul94Cypcra57534mD3WqTAVoPzTtP865o15NM3av4Vp
WcnudnLKvmqnzStrEnk6yBVr/XAUvdm5IT4KVvsMaAzVPTHqXpExEM300ZkjwIPgz0W9AbkOBGMP
yXgpYhUuCUqpdjQ37tSpu/Pw9t7UwtfbUx0nrOkpzkTgqgJJC8eIn/MsPRuvpBwuple9AcOs1K5S
/4nRKCOd+9aJwxwMS3Rbqga/OGVZ6VZaSoKZBU96IxH2Qm/Qcfuo32vF4KtSjx620nrKd27BWtZe
ctWIAMCcy/STaARZSm0d7sYEHvO5MNGmeWZG5mOt2Ykl9SczyCUsddzZ5EITLs94eGdvVKYpfGAU
UuCq3xC9qi1vMelcKI4vlhVYlpoxx43M+beDsp2bwrxXuUwdSfHSZkUxjofhHzXlCyc9Z9GBr6pv
MXvL8HxlnAUJ2T/ydJDX6zfXt/wrUVxQLwjDrb2jn6kXLzPZQvoRDpr5TRunfs2oPuIXAw8cAtMV
07JkcbdXqHi4w+lOHMWenp/c0aU7fkROlIKKcKKqmnrnkz9X4HLvizF44urqG5dmwoqcMe8U9urA
q3T6qut5XGqL5p1+v/gil6XyqQcYQziEcwTLN064qwarvm13jsOyFZg/wyhPSb6yo2n5pbjEo+DK
idohJHLHjXXraxorJ1FtHvXux/0kRc802CeeXUM42dyWJdysyzQtXHoRT56IuZbpl38DR4lYmJvR
KLiL+kvRi9DACctUYqGjHVSt4CjGqa7ssbHEQYf0aamT1b9wq53jThVMGk4mqZ6Jgmf0PMZ/q2xI
lXmrZ3XNgfjpNS6V4bvKSWdXd0cjEQSy6KkkkBu6NDmx678cy2kRl2IV3O1x5TmGIEvmiPYdgbj0
EDDiAdc+wiqI3yCwoTDWVMrmkochlaZNcxDt+HYq63rEq9wqsi3uS494aJJpIpC/fSqm3H/B+xzS
G0C401+xNrw/1FqNpnxelX7Bl0tgd0kT0d4zUZ1PknECcMnCdexW/2P2txEseA+lXPNQAl4U6YmC
I8rhbvEhGf8Vgz4B2Y/pZSw2FnSIPLEpabspGXMctLCTgQzmr/Ra45D6HA2pd4yr4WAanIpTq38N
PnxPoAugpu7EcdqEnlNVkRDZvPiiOtAGqnkBg6e0IdzB4B0XuL2q4LsjuZ0KWmU+7A3Xnswfo3Ze
B8p5bsCf5O4ddYnvIoIugQJoxaBvxaqlqRdIkeKW7ZmLQnrhPOiZKDS6lE8ZKJgLP62bVKh89ZDv
XPALu7UMfw1V3TTjafmDiPtB/rwBKbbj2EEGCiW8tSXkxFEZtxQXjMUgGaq6+nji9ThQSYbKTcbZ
RQDAAgi8quNYLK0MbEzrPdMuM+GWJ/It2d39Axjz/1iAj7zV+0TGI2vfXRhDgRoVy/P4x6JDgWM3
FSbr3L//EleWZcFOTYXfisElYRneRpp9VESone/5bvVP9aO3oq1h3yX2W9cJ9ljk2STHPWC2E7WH
YFdMPUFqwJBZhxDLmgeXWrrL20veC8bGEkOPDF+s0wragZhLpDLUxesxMTGmjToL6HjSBQoHj1PC
rq0k6sfGzu8cmHqFNM48I2LduWMmDY6DumPri5xv70xxIxO1f/24Tr8eB9suXZNsdfS7H74TfGdC
KpO95xKyPYJB++GVlGWrhyPz7bz3Bejh1WExVoHBWqbvC8djPZasR/lk94x/e1C6kxVmp5PJGwQZ
A+nho97lVHesFUJuhO5ntKo8L7SJXRF7ZaC6NvofyvPZcga6TEH7mS948PKlQ2K08Vitg/4vspbh
xPJe2l80pdhZgiqSpoqMppoiHhgU7bNS4X/yl0xJbB+VK2WorazWiEpUMhG4ER6hr/CTK097RbIK
BT7entTRsS+sjVPWSOJs8uUJBv8KvSTTv5Iieq853Iyrkmpvv+xXwHd/9fVKpW46HoMR2SbbPez7
veiEF5TR4TRhSCwGPHLgfzcq1AdCQ4zZw9fU8dviZcKgSmJAjPIhYlm1/2ThSrG7sDxAHK8S8MOd
Lq+stclfn918xZBHrv9ze71/diqa1bKWLQk9jpdO+W4bzaaj48LYiKOZ+A2V2fU1i4b7HJKemiiM
5u1OmodF23em/qABDbK9XuKnu2KfqbhCC8T1pqBtjYyBNf/yKVfT1leDZ+mYVE2MoZmzqQap6wbI
kT+JINxcH2W241dTRd8r7wpfBfPN2eMvYz0j+vYH1R5kOS1Rl5tWAbrmxopiNgZogmklIhBzjRMj
r49xfgmx6SveR/c0v+RxqA7NZDH2FfzU+mfRTQwU1dpAx9XhwpbEKp8+Wlfss05bEO55jXpuF5zs
Svqo6WFc+FX4erbUb9MjaBkijVCCKkBqty81Vkkvl7l3KhhkKXWzWWSJ5WBFkKEgLKM+t4rH+z8B
vIXUNUn2969T8zkP7L++Bew7Afk06ypnNJB/M9Ii6xrKrgul8sjNB+T/nBYIEdEgCV3RppJH+cAm
W//0lArc+GzNg5vFEcMJmLJkXfjch/7aHwPwhCs/EMY2xnLlg6p95a+BZf9hqiFM+MbWFV2sNQcz
T1awjoc0kCQiaFIS1sbejF6dAGuKOJDjtFYlGygoPWHzods/Fe8ENgfYg538qKQ1iv83Y71S/mCY
QMaUN7CaZiFQzKMsW4m2ZAIIq7TW5z+4I23uJUF7rw+DgrH3hokdNZPS7hX8VwaVDeLjFUaW/PsS
gQk4OD7XWbR91SIJj9KeDx7/UUQ3eWUs9FIzHqG5qOtQCT2hQulI0O0yPwgnPzcXGCdAlclxmhQh
lrmV4/cnxQcqbGlZK2iDszXG4jCZVDdB4DVCzXvxBAdCnoYzmVGxc/wdBuEwpgf+NYR056+aC+xS
JgxwIhPT8oQp05TKuGfbEMeMImz5eGRUyB1MAr9SvnI1QJlKOY810eVT/u1ru/cdnjmHY9VGImYV
SiDawopnjCT3gL+CTQ5SmiVo07hW//JdKXASmbrMLubB946+QUm8E9+sKfDyeVrPPpi55aiFxTuJ
KYf7UraCfAyxXDa3wdS1zMriwgm+LxJNXamz3i/7EhV5E2wCdg+SylA4qbdGGJEOPeLRCfeYLtMv
N4bbEi/Y0FPXll53zHIqk9jgYsZKPM0yyNYyWLydzNlEWyripUVk213bDEGs7Fa+jNl6L2X74i+O
39oFeUZbqHZq50OivFldSihJiV6ITBfeFWqZYVJuEqaGa6YxqFN2M+CBIgMUyri9DBK2nkV0h28u
K7/AipPsPBlH81I42lyui6nqN7QbdHVcrqAmiKfA2+O+UqhQVMoQEcVb4YgXrJRZ0yulAXRpv7PJ
KQXM0OvmwWBABPM+T4Uc/wdWGVhhEbeQnK746hSh947xkZXnTLZIzxrzvOajX1JyubTM75zUm9oW
O1G8kLLUDHBLps5fqgMhLZV/CoxZNEPso8KVP6fE6xxmwi7JXbmB6wyW2orSuijaridjEDNICqqh
cDcBcHmtT8yvQMGfCakgrPLXpS+f3JAWqbDa9BXrRn91wREjOJa5DPKd5SA7hpqRNg4dg/mpqu3Y
WGlQQV+FnDcwbOE58p9kspxBG7GFjPhY5uDMRdSQBm+3aVSCf1YvMgHr1pAjpCrCqg8tPZW5NPq2
WsLmkUVjfzqH3cx2Tq50RyjvYE2AC0BodwZZYpLf0fcmMUY8jGLRpF8M+sj1HJaBiACDgbIGKWgK
CoyqGojXLa/9L5acYR7B3bkHDMYyTObou6Unr6NsgBH6r8FQYsX1O8junFoND1Sazgyz9qNhjXiy
IlhPS1fmzQHEUcQLmOtnpSkM4tp9sUP6dH3reZ523uGBKnxEmGz7vmzDC0hdbL0XMP4BIpKrS8PS
/vCqtajL6PnTKkqeqenM7VBddv3G4rVOtoG+0YlZ6+/furtZYwa9hi9iU0ar/Se9t/gccGWLP75o
bFUfYExNohVkGjUuXuH0OKUgMZP3ivzKWNPFQtNx+UL9etrGF4arAooKpjc7HfzLAzlAPovDBfH2
70ccFYVcgX4orwE0gkFPA+iXk4StmISx0H33k6lzZe/Do1ZMiK9O1zBpxPoVcpUGdyQq3c24MeS1
R08f2/K8n5BI9FEoN2jfvKkmLWsdzpjGiJx95Ka9ksolwKCJR0dkmzw3K7t+xuJq5r67kRUM2Aa3
lV1/gn1M9a5/bkB8HGsK8voxLLqfH4HhdgIo3+GF+tDsQ64FCPwDZHiS4Gnq5E7DGPC6GnPayIxt
KlJHBqtFkHYPz7MPi4eDyui57R2V7g9j7I2r+9j2ztYppOh2Q1ysN/YrXfAaZifkoqU1DEozWXoh
g1YgPmQJQhYmhrpyrdkkOErK/YwPVOKmK4Qw9prOy99HnmFt5k0hDitXubzK59UKxru6vNIPadbe
QsjQeX6izmyhSomRHNntLTzdoF9+CLoR2maAH7AlkQQk8BP3QzcAGn8cvdgSBNrJWKEqiNiM1Zhv
ytBBZlKDq/HNfVEtpqUTWXSU6KslMs4GA8btkY7UXwxcW3GJcUk0HkHidHq4btN5Yqgq6rsBoGR7
zgmM5XybPywSPMxCbJ111KDv2VqYE6Rs8656tropCxFGznRcY7GSG29BpowuXoyVkJsKINsKb5F4
D1MMjXxBDfqu9Dm9E/aInC71EuX1TPg3UEArnPT1XZn6c+tIKUP3w6SKQNh1/lfD2PMVQFoxv74d
gyXVtiRJVwkXbd0Tg+a05rReJ966TUNlGtXB++pzlQakR/VbIf6Ob4aNfDMkyQCemGqK/Y2rtcyS
aWDZAt8dMsXn1tDoX5x/BxUu0Jy4ykc+jUVxvhiHXy3Rzp2Xt5239ZdLz5cHSZ2xPCU+kiHq8dDr
3XVJb9H+xSMUqXRCDw02DiW/dsyS7WQAYtUpXCrMbjmlTOAAsdySmR2nDRqsWP0AIoLY2yc8gSf/
hv439j2hJCgXK7Kp/Nl1ZqMlklsgbwSA2yont6CcxscgOlxd2QY31AAievGPAHPVKWjjwYw3nb/S
eqQtyCWD1elrIIq1dDMTqhjdkhrqy0V5FYcz7VaG9/ZbShc6WGRZsBexY8WL1F4Q9NUjPAvt28Bm
bun7RfhF/NgCOfSVMNHExjH8/S35HjgHWCNTr2HxEF+VeJ2wBFEhOHR77CoQY1GZ7IMUJKoFFMHT
B5N5HzExPKc9z5W7luWg6VB9BRnUuJyCcYNtO3+3KPm835MKG/bg+85pp9J/5wbAcGA1gFOp/nHV
Ltffhabd0hfAm2/zk1wtcW9IiJn9p+Ht1lVeTl/ygUWyMzN9NTgOGR/zFuLQoKkFNuRrbkw+hPdM
qnTln5sbVD/Yg1WLUnFZx9if8gADFUrfCgl27qSs99qRdQxyyDoLr+WMNPTw3wJrCa5U4vZhfiM0
JhyLXxMvZz0IKElvbWvCBrJ6dQmcQrUOON577aMt/RmwMQ7eY4LWEMIv4nOQX82d6Fh92zAf81fc
a1erxfAfl6AWD+sD9Mda8z+3qCN4HKUM3/U+b1Y6pIi/tzSp7kyAZIQcJ0kVRDV49xrfOd+ds0Pn
VYVnZ8WVTSdxfJj6Sc3OmWE40IdVRvHZP3gkWuDYmXPvu6zOfkgS3MXgZ6DLazXB8MoRqBy8Ljkn
Bmreg2TzETOgju6lZsVRoX6JJc60WGE/x+Oc2WPmYRxyFmagaF3IvFC2kMX+vK5U/skruyP1sZwv
O/7EORZIGUjtLFPWERCslney3NjfeShl8BhD4ubysONzrmAfQmnbzl6DI4klY2CFIaNUVVOMhRV0
iZbjR3BmlrDybYUkq4S+OvLG6WeAejOh6yAx17sVHbLhDSyBgs3RLe/LuL1nuVeAmDzD5H8g2KNK
Zq+klf+TVvjChLroD/kjVpX0fjcfj9n9oU7hFREEq8iCtyqc3ieNriWv1+NQ7rYqz2zOCcZlGHQ1
lcMJvmJeuBMybT2dNarmowIEeIsyvIvt1vrR6hCSppC0qZ5z2fk8kWiLIXo3Our0eAbuRDSkflnm
wk+dtyRkNGjsd2hsB/A/o9sAy5RQNF+ShJzklf/x6iAP/30xWsHXaC/O/LEprkmw0GOlcvXGl6y5
dbjW9h7kqLND1C8ewtsTWTxN5Mw2A9ecyLNBAO463ZXBjkpf9uquo+X/t4YzMd7zdjxzSXf9tvzT
caX1GRvgtJ3G/+5dukFoNCpemWd8iGEdJEzqKc3Jo5I/DJbtl+Sm5CFcmn7/r4xYYoLPgtDjjyI9
24OL31oz/jRKBGFd9155USTOVPpzg89vDByO7GxUczM3pCCjTQliEwoEefLIYPXd8lxtbhp3OmB7
sOUkUhfvLe4VDAwfqywQqLqU/WbM5Gc8D8sUK6Q/MZxCOpDHX7X08BaaBWzF94q+y30BcC5lz2Ml
2qJ/tOgEK9bKaE4skwkf5dIXFF4BA+5iiVRmU7Wd5lk++Nfjk/UZZknZL3kLhzNUjNWoPhBYDPII
L7kFuiBU/LVtoeeU7g0UOMCMvUBRfTeh/wqqXjMM5nLZ6nqFIqei2oZtQJyHMNKIBGpWsfBzPiMx
BYp49NpWbOCTB4AFXVZlg6m9zh34Q8zVPt/JlPFGKNvEM8rWgXpm7gdKr8I+PUH6CUaRer0uqJlW
EWDZ6XxVcKVGruS/5P1Qcet+4UTLfetdPO6CAxl6GHnm6jqXVcABstVsFkf7GwCv5aOboGeZ8TgK
o3+HjN2naHqn3XBM+eFwHABg5BCh6pz3Ms2iTq4VxfHgXUOrVQePT6D/soGbkQ2WjYl4B062H7vs
4PXxf03GWgQQ2vBx5Ni5SlO8/dxRpYemnbgOpyx7BXaJZoKJXQCmT6mKMGaSR9qqKdXHgv03L1b3
wqxT1VyOzOs7n4CbueMNJOWn/UcgOGHDgKh0ysYNgIDVF4jGIaWAso0geTYqhqYXeRTJQHMixpNY
gpL7Z7hUrLvVnHdGukozlrb/riYYm7/sAH3KUUFXbidZCw35ZR5hX7UyxEHkUUEfpf8jxWZWH2om
/8hTPjXgWRb+gsKQaEhVZTm3EmG4cGka4WJsL1vKBoOyUWpxEEALo50xVvUmg/cR5d432oXn7FUT
njUvMIQ1WMf72+x/wjLx38Ke2igiPC1+PKExG10VHSUSSGYJpWblJtncF4iyqYrCCTlWRHR0OXoH
pSPHSJeH69l0xPHtOG/u1ngoc+rGLlHbl+08QOfm1Vky/p9X1CG4m/fWdfU2x0pCR0RJNmEHq9Ib
BdTwrBZE0//Dz4eF2RQ0j0cM6bvJksBIvLEI8UfjRcBSbkHnY8n7BjZHWmHo3F6uyPdAbapILv3j
D6WWc7LaPWOx6I1pVKPr+rv22klGmzyEAGWHEYMiod2CbtyD5/tjYD5igMe0s3StRCdQevOtvFor
2834c7TbCzqXd/nvCZPjNP4CaDvsnI/k60Pj9bBYb094zIyC7+L0MwFuJe5iFP/M0iYnlfIxXO9t
z436r60UOsn8P8nuHDT9D0Ll0laseG9hQ+YDfQTfbBYdAMjlXUOxeMEijfVUYOK9EfPmBvxqlQAg
4xG3nNV2MR1RejQ9GeOupYIQPZ5GRKIg2PUvIw1F9a9SGTyXIWs61DjkzqOS5PeLJaee4IRM0KYG
+WB88Hd7+TbuMqo5rgE8WpghAoWgHxuYvm6iHAvwgITU4dfu9hATzuvDctowbEPEDqZ16Fu5tg7x
Z+agVDUEGWI9C/yvWWaViGJYMIXrQw8naO+w/DIGGvu1d9rkkY06MqilLkEFxy0X73aNODAEkh52
7mwDDfTsCK9pnUiQTIf3G/dMbbac2nvrC0IOMRiKY0YHN8teZLYg6n7jirbEfliUvu+yA4bGnQvq
BpKKlak1fvxMb//Xt7sAgEh7Xxd76PKK2OydpQZAN3FoDOb9ZNSpwPWlRooSc36bogLVf5ePQsP9
rEsDEGquHEX9LotBwA6iymzOnosdSLjzHDBFcGQzNpFTalZzcMhQVPtLHueVgsWW5PF+RRlbLlKP
U/t8HeJTlzQ6vXFIjGpVD+62HmA0MFWVT0VwJYd2zViWd85KzSC/D0JtaLNtWqBB6FDelQ9CZ7gu
mS98nycW8enNRaXR+wnyfpMYfUTPv9v1BXMrJptvsZD8SKJibXdNTAgPtMUszvL/oWCGr5TGuerV
f8wsfS+XDXsbrgIjOAssSsyiWyZEbcLHEijzNUdC/X5Bi23tFUCQvO4HXY/if67i6QZwnU88xewq
z+Q3IHHTYwkKg3lmc1ru4oO3306cVzuOu6ahBOmJciao3sGh+thdgRXGLZTq5FxZabQOvQGNHVXC
bxXYTcUraTsrIYlS2ZByemBK53Gh2TGmHDtN6AtPH/UG7KLPkoah2e5N4DnYGo5FMfljQdClJ0+z
vDnaDrdju34jC+AWAzMyyBmkwmRhIc9GgbTaI3YG65PhMO/Rg/QY6Vl9QbOtu4qgAMLfsNaJG3Ok
1s8dFJb8xbbPeXhqlITyHgmJ0yr7tly3X9zaoUFoQoJa8cmtkzWu6WWnOysslmrAqXVkGWH4ejkn
xvMMy8dz+Q0RzYjUHt2LyJHxoF2uNxSi9McvXrt0njMGINDDH5ypEFHi+ApAp2dxDD96b3S2IuB3
LfkWDcyd5cBSG+S45AyzgH9OTDYux5IBqW6SqXq8a7OuszHrAQgouEqlQTmn66hAn7p/FcutC6or
6nbprqLr24tCuRWC0dCdfBa8sYf4FAg++h7f2/U0krjvVoduoq4A68fpwCjaheYy8Xp2/Elg3fjt
TDYTD5T3wlpcMhzWW5iKbUswbrfImF4EC+W2+3hzvxRqzuOVkD7QVbfb0Fo6p/fwnjsT5xq2t6FP
rqJw1xqc2QNN71M8x0t02HyEA6NWIJhVSts9yvCTX6uyAdK/IQgf8gHytnHPf5WOetdeqNesViuQ
sbzTNGE3kM0bv25GiUoyWIRnN+TUuIYubf0woupLbaBv946ooDP1+GLcKZy9alHDvlwHRR31jIZZ
aZmTt2BH0mUe8KtWRi3jp9xI/c04yvQBvRZRQRZlokvzACBbJYqLtXjCWQmaYUif2BcoDk8KddxQ
ZOsYxlHntVAQndBiKSqrzPT7m2dKeDvpQl5j2wk/Zxs5v2ysFhQ3Am1DiyqvHmlPMugvTr6HXKpR
DdBh+VWX1H8EylfhEDtAsgdPnWMQJigTwOd6rzaeaZ7OvgexGyirbJNLotvs/tCqUev38GiXlEDU
+KZRa6ixhHbzZAjIEi5Rid3lWlQu/TG1ZM2t/BKcbSEL4jkFS1o4IBgD+FXG5cSWuciZZkQbclza
yYkRJD3lETsl6qPmc5bft906hTKOjoo+KdAGAP0xHVJfprfpK+RpLjJn7lkHBFgnFIA91/rYJ3C0
zCDXyVmlyVSf6Jjau2gjIer1v8GhulBlJbN9vsptAI34ENdBvFcIL5CLJUR9SFEZc2wjQhuGuqMg
0y2FSfmJGGInzuLsiSwbvI4Mg0fZdporBaHmd2CkwV1wlb0z3+fKeiyly//M0ozSGV5qBuuEXN4F
FHjCFY5YuhV50B/urrIUq8aXaKZ5GvLzxeigYR5Kbekp8cSjGc23fKjEQKCWVMa42flsX4fhIhGQ
7Wn3ybYz0re5hZPxxDit2CE4G9KnwjA91MuO5i9BBxyyD7EI9R2tFblD7KOxDzZgEG447cBAx8iU
7UpjsR1+jRnJLQSwWIE4gFdo1nYSBUzUAvCmo3F4Almv20ssveSV2vN+/543XjLV2mXqewvdh2v1
d8uf0vqgfBtjiPfkKHK99TuO8RusePg19b8RbVyLNRyF/BTMn2Lz/bAfIucM5bF0CAlPcTwBUBca
tyrleERIESkRE0AbpFBBuXkXz8kdYd9bPF0cJIIQhBjUQxRjqyoG9n7WL1ssh6SRKubgs/qsJUqP
ZOKPU7Mp4TKvmOJMat0dTGRZ3uXiGbsLypdmr+c0olW9BDYtHpmEQFhB2xAcExfUBUGNLygyvJQi
WHSKFpFASlfd0N0Hbynrz6Mu5DZRdDB5hPVoy5SKC1+Y9TSm5FSMRalbuYZB4c3Hn3JaAV0rzEwl
dPMe32BBttQQYoTW3MNaSEFJAeprfXqZgr6uuU98TQmZd9coD3mmYjwLEbhExhpMK3oD9r+J6ALS
rWVq+8E/Q2mW/nud/hx54oFdLUXDhmu9rznEWryUxa5jNB/o8NQw4s7F1LdztHFdfGwn7SnTJ7du
igxJXH03zJMsQR5iGSjohg362C19qaZdHP7KDHlPPrMJveAZA93Hhqg5IhiIZGT5CMZgxpygfYhV
5vCjeHihzli+HgB3jC0Glt9mdVCuunMyEMjmMj6pnm/sbFJCIbhQY1WQo5F2j0jTtbKUMtYPoa93
w+tEjMMSkbe9Se+UN/Sj+sqreZDa+Pqr8uYIJCFQHCMTMRCTpQ+EFUBgb7ff9H0xrBFfjbOqrGKy
qjkuX4GIljONbzYV8XOGS7bGYWR3q/NpU+krtk585ZCQWJNLU9mwHoweK69sehOSZeY1Y9ZHSm1h
BPzPvgDX9NIPZ/e8b85zqyLdrX6UFfbSa14WpO8UdQk5U63joDMV2aoLyPMpBcOLOY0z9DH+OPtQ
C/Gr/mfKslbpGTPqlR9WL9a9bA1XppWu8ywE91qf74ydkFK1+q0wboRjz/g0tPI70DlUfxedkasV
rZDSxH0neRCHuFjNHue+U0AogjS9bSHnvcQbYXQwf6smQQENfrGoYWbjTrNyiLyN1wqOzaG50/mf
F6GxPZ965vjRUqX+sLTtJzn6/Jolm7pgIUYwzuuzbZA/FzR3R+/COb6mQ94HpWSp3sJIU6P3g0D6
B6Fp6vR60XPdXDCu+jOjihALrTzTdDhOMUn3T3L/A+wpeTDwfLCumtlursPVWLy3upjhA7M9XW/1
8Qc3vF74QiCWVyIE+dxCPYAyz0tFMIfvgun9n0xTaddh4iSzBHhNO/uBT9+bQMCckwWyzgB3Nm9F
+LIOCtUu/PZawankeLQuWewVMzVaH4xvdO852ZhKc/BOG4wSCuw0Y+U0aYCOzj6WW7UwsXf7ebzQ
EoCkcoTwi63J2LPaYvToN90Y1c3U4fYOBVBukM3c0mgs7yFrCzz5jY7i40Zp9WQr0/3g2ZF/OgnM
g00A+8qDvMoF3tzAAQr4bggxQSoCmhu1x2iGnwZNRlMT/twweADaTWrPthWImx6h//IjB56CAUwm
PWwRxC6l1iiFHAxyTDo3PX+AO5Ncc7QiYuUX/2ZHgk7DfeJ+yG4yqRRvirgyBpcnJVmyZADBWc9w
z+z/twimXA+5mhtvYED+hunZTwqKvhUPvYlgcLPfg8o8HaRIsl2CTtWi8DUW/kSlOl/eeNjsh6Gs
/TGC+yajewp0CnT1DA+27eg+hT8me16LvjkfYaHYvIrYi4T1u20WT6oOJByjLDqoEbuNS2qyd+KH
Cg1/DrzVnMGozER13kVaPf0romX/mtlvZOLmAF6LaLlfeM/4juB3t4jE97hJF3XSxohZSvLVK7TS
yHvK1XVwRgcdJjYFw6Zq4WnZpZKY0LE5Qy+JGW/xl4QRdi0Qfyz/fvXMB9NfvFW83h6OPBf4T1hi
AuxwFmyPE1MGK6/5mAn71AcQbQnv9d0bLSGEYKK6N5qz5Joog0x5cb/V8855YBHc5vfLrK2JEcGm
Wd7G6/S6ghuKNos5NDhSvC9PyASKXFLyVcMzHovPTm9r3jM4CoImuDIQn5n0GmbLvQ2kdSXMCtEr
YLXoXuvRVp6VRbmWsgSLX9oJteBqnyrjeYAqphDAmjLEu4jtGmCr4ufCv6s5Qqf3Dd4HwJoU0Pd2
SJIOr2wUEGNPEUfmdhPzVW7hxl43YdMVqWTfCGdeJXVDNdL/Ma9lBsD5FF+WUAFWVj6WePr8xd1Y
MhnmqAPuqpP5AkvtEfJZEVPBzuDeZrUsFGGLFgyFUH7qfS4OnnjUrclS6qTWdcaypbKFmL6DnL9q
6Rsu/ZI8oRAi8U7PJZgZwalKP0bGin8vW8EJZW5B5MrN9l8RT3DvzY4lECsxg6BPB5wVpZ+Sf9J5
GN2bkC3j0B2G+z0z2f8pN6PoG9duWr3FeWmICptdH9oh+mFeqLgAO6m0k5VWKpbHRRYoHfhgdnvv
1Iui0AlG2SgAJRichOPJtiQqTD6wDWJ72K/NoYsAwx5Keyiqsh0bLp8hAsOKeYcHrYentBDFhd+u
z8k3DKHb5mmz8qZHGCfSHvbq9HsBKNLi+Jf8KXPbmSiLOTrD1uw1TirxVEZFsoVw3L6bod0c/2yb
0IB0pNBbXdEavxIP8FRJ6akn3gdM8lGZWCfsOgUL3z0NSEfn6YCO55LuH1Kg76lECA2odwPgIWzI
23mwJLxA24gfP/tORqdkyxq9EICMJmpnusFow4yezxAjE/VYqaxJ9Qt3r0Essbu3HYETIMDJJ1gi
a3+i6KJV4KvinRE2Z+d01H4wQPI2lnZikolFeoyTRPScoWgWuBZjSyFnmVJIhMiQtkoUt6aZoRPo
tQBw1gRsG4ER1AXVBwyyeUprMQPNUCjpBiFutXJbeVEYsW8NW3+qUn9BPRR5RSbdjSNUZab2ht5B
Cd5q/q4bcKgjNkpz0o4mARhEw0UhVv9akRJU+UvV5pSt6cefm45LFehBgYKhKxnT3lVZoDk8Mdm4
EHw7HpLGaUXuqhK0bdfvpDwjpgqpGDjfdGXSYtVnySQWf9G4us5olhOajwW8wxJc8UZq5ynpPuLY
H/oD1Sp6ll6yZND17s+T2Tz0MVSeh4uD2Z8XPTu6y60wEYSQBXVPWU56arj/wwcuMvfbz6Xc/BVd
tRbkR3+cQ11XIcWJafAvl0D3lqX73SGKYo/ItPCPVUT8Rm/URtC9nwNP6vvAUajmVKydm84fK+kN
hWsWy4/cUAvXR999sutRrSxybuynNUxs6RP2XFOUAQlTkE9mEOWGQJM8Kt/H/yVYu86FPtKWTFvm
MilpWYFtEOuxA/EOZzsei/vzST6I2BwRmUYYIRloEu9/UyWB5tADiW2q+pxJVkG/1c6Ea6dLEzro
tmWiOy/oR7VBs99rDLp9eh4rFEndSzVCq1Kk3yRDwhOVhEjz8eWKA8Cb1+C0U3he4AjZ7J9de/l7
V2FfEzVLOd0oic2kcvVQbDK66esItcjaxKqEUDVvU2nnIsE9/UL9BHBMrdr7c7pOU9JYXS5xMXCR
H5F0V/44IjCE8JO5d6Tkk1Rjfpq1mEe7xVQfwbfaNl7jYwKA3BSb0YkIO05vbFXZDr+Rvx8ML0Nv
aYmlgAwoFi3wP63ivO++5MTXhtAelQDBLhef3SspSj6IVebkXVFWe70j4WGQLIyQoDGqM9iSC6t3
K/wlHGmG0edXWbo4oFjpsxfRt7563ReoeA1a6QNVeuDg7RQrbI95sohFVyHORL/GNwX4I9VqQXNV
AkhpqYt5XWfYpR85DAsiRiIBKTUFvCn8Q7Ai8+er8cggPX8BmfxSak/utDcp4OQXN/ga8G17qQ6q
kuDL5//FIgH51/bhf1QS+AXZE9dTTMLRyFDnv8Ac7KTl9NpOCYQE1MC77RljXXEcTc1AJSmXel1J
mHQHV01lHGLSi4Km86Io4BldvDgug+xArfRj/ZYCV6TnssgtezvN68fKa9vJNtj2AIKsLuALep2t
1QAqKO2XzlQTT4wnmeMg6mjBbS08cZPKURvTqLW2lEZlMufwDKsKv5U2H6+lg7R1lq1oJEzOA93S
FZdd8B0B/BdQOw790CKXv6RcJ3PeBZuU4FhOKgGJ27dfuFzHMcloVHylspEq2ogknMjeNeBspykd
oGSavriygrEM9W/Hnn9IeBrgZ7LkuYXPZDvN6eU2Bao43HV2Ju3V9vvlW0G1NVAMQYQdiALj0irc
w62nTD7q+MFP3tI8iGjmVSziXxyYvmzhtSo7Q7W50SpuMAUGqFV6W0bmiYZ5pJnyY9UGsMmIXIL5
E9pdLaAO/o/o489Upcy1oLy6NKNsDS/kYoH+RNPRRZG7sTQ7cwapflHL+ogN0N5wSA43iTQ7jOST
4ybx/Dvw3bFI69OTqnmfDK3v5A8g2pLbaMDXBnDhmV0Ustm28YBulvnWpVgTTlkBfDwFSp4/jB2/
QY8/j2ipFQCmwDuoBbDt+s0BLEqyKbiKWeaGSmBe0XWEWODDSWlyZ/184Jb3Yo5zhgK0dqkGILa/
w8sjI0KZkbVazy9Hh9NWozkDl103M3ZdzqPW/BvnXAXvUzX2/E7VpSHs1vrFl8IO5f14C0Ulvgxw
KlEq9Bg5Kvqhlv7smLGnQHrBGTCd1H5NkfcAw9NwyS/7p7FqTFJ7PE5mB8iuW9ntU2HA1h/wnEQu
ZY0J+4taUMPZpbryJHnNZZhrxXEW5rjjstxNrxmu0jgVw8kkTjGRczTL9Bc12mAyvk921033qQwF
Nz1XRvYtzAU38JZWyCEstBlXKj6r4O77NieNXtmk71uqNy+/zYk=
`protect end_protected
