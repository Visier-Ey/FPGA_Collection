-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
KZIdeiUpUufOpW5fsVmDLiva31WgHNwCgZbbBsTVxuFB54anuBgFHPzplqykYPfQ
CtcjdQxLXPdVS1YjKwrPhRcKR6589f8jftCaK6sc8SlkvIWS0lQa6Q7sLy9bpuYI
2TFI69vF/d7KpLZ8JBdbDmRk18ItSY65NEIQCUfZg9s=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 4653)

`protect DATA_BLOCK
4/3300LMXevI2gTEdHWh92AI68w3eE/9+8mrnZeT/JlziyqG8kqBa3B9klfXseov
GA26O3yH0b7W6qi5ZxN2Uybg5AaLNVQtW8Oi4J+L6mnDtI4MiAKf4LquiKW3mLxE
qEonKYMhQ68kVtPGE9b/6i2rg+nPIbEJNGOSakdY5ngEWWs8XTuKQlNSPihsUwLt
pzGQSY1mI+ntEOVDv0QeJH5zd/JOuCweGt3tNk3q48CtV9tlTunx+6r5ttQtdv06
T6svRyre2vfSufGNj67nqVXpzIM7ZLHmS8FrBG5M0KgvUATvFykzXrLzluzqlwaF
3BSqq0QX9Jmzv2cU+pL4PYmTkvQXi8Vy/h5fUab6+q9ZqSVaSUVaOzjgxiA4Prc6
aqXtns1uNnxp3VMA6+16fTGkzljeS6yYad72/creixp8p7J+4dtfMtxwhvMcV+kF
DBKdAIZTvzVZc+llqlbWgkvR+lNJLlWJpg++aNd8HKTcXg9J9hMh7muD09oEcdym
SCV6B0v8GtlSTizIOfRhrZTsi3uignX+AbSf/8eL10TZxkaE7eip8l8Q0ESak9Ui
Uy4QK1GVvqXbjIaIZv+tHROc2o1yLCV3dIxqn4Id9MugavlZ4MEpGLogdsr7flU8
Dx+dYAPIrjmkmBvqG5XToRIkPYlhUq1cCfKKPsint5bSDnoDc0ajdunEhpQGJ0EL
9RyNh1S+mthLQ8d+0/GJbQKJJgqRvEl9B858T70dGTyw10qRPGRGkI7q7NBTfRkx
GwesbH1gGxlRE9E1gduP6gXFiKYI05CVGPL4G+cT8cmtKs2YSuN1QU8e91UfnMN1
/icqRp6ERB1lnCJ6OJC6Sk5W+kPjbqh8Xq5tyZcppxCtVIail4YY7Ph/CHz3ahBF
2bI98CD5OQ8w5HZ3JYoIrylyRSDAACHpIiBB7+TCtjAmzRHl3KxyBQURFH5NyQCy
U9Da3ADFuN+5IqZzpmx3JBqHP2x0fUS0eHcRzWrGLUJtPW2JytqEtYJFOAVrCUDO
WdGr48fM7maDXuwGWT2LYJdeYI4mZklCyjGfIfMm4Eshn90kOgE36Y0MP2Gg6SNA
IiwVvjfLXaG3q15ZzSQsrL2q3gfJyPjWFOjPbtnSI/nVSa0ECooKw4u9VfGBqU1H
X0UaRC7PlJzu6FgqpgGGHoXOcv9uLv538ivKbXd7/5YsmkbTmpNuWWRtR3qJsNVU
G37GTgum4HV0HxNVQt3XBOm/MhjOttIGSXpYzxYZIZH1Slkgw4UNY3DbXlKw4COy
ZcuvjQO6OTBlKooslMKM433WcwaL+V8ZOiH8etSerXJLodim2u7xRgCP0bT2YJax
o6DQy+JLHuzqcsZZt4KEI2xEbX0PMO+obmONKOPk/cJGYhsmQsI8+1oy26Z0Yrbm
PbWt8RrvXx9uasVY8dsKdRnHRCtVkmwlZ9eMTBYMM3lpp77e8VirSilw9wUHuJQX
rHY8Be8+yWsCphayWBPb6eDcTZOZDymAfuklTKb5SU0baaVNW8BM4Eef4qUfdyrj
884Inrbvh48vVfZTPaNyCrAe/sdmj46FoYsiwKSDGiasfK3DiHP8bxR+8gU2SLjU
jbMwgOOg9CUdvr0Zirea1mDulruiqj6ZC/2i+D8opTul9jbObi8IaoUkNCrpMoHf
QVAkyug0bB19f5plFdk6MDJl7jlg4rqBwTgOVqLGjx9HbiXitwV0DOdJjn9VNNoA
yAu3Y9eFee4Ul/cvbezHmxHxoFaVbvG0ighDKQbouipL7bP74JmsqMJIvBiq/boR
FItX7Rw6/2v96gncjDIyE+xyX2KqS5q+c6ivI8QKBdQipngJnDaBqEtjxeit9CMg
u3GOucxArpExUZjVsZQSK6hP0Gs+Z6xme+aDAwE33uRb3fZ0Su7116mmDiElRoDS
UeWkNSeXpKUmDIkCHRoNIIJal9wycuzGGUG17YTJ8tuPHvjoyMyzyholNthC8+LP
c+MatpaxOuxRweAzqJK48SkwKqrq8Cjx6dem3HoiEbOpEtkolWYWZwaOqjnqZyCq
jMehXhRGb2prjn7BkxKsm/tNSOrWQtAsYfZ/AKX+VRdagakfni+lUz0S3DkQoHDQ
msO0sUWNVzTW/mrinu8x7wL8FrRaLLuLasKy8/EqlpLUD5nTKqAvyZB8+5ZNJ1LP
whybRLC0NRoXiu/rCdsgZC/09TXs8RvQzeBOl0EQ6HTBHD/so3lcmbuhLS98MI4u
ZDDUoYHsAk90ZrvSIF9HIM2skWy1K93SceZrRBA0ZvQ+MZ59Kmu807DMUdXyPilu
+04jMi41o6TBkG6rTB+lG5M1qDIEeqlwCXBtHOtH4V1hEye/bwXRo6/1CXFaLCFp
t4CZLH/dPFybz8nI59KNCbkp9iGTwtKHs0DnsnbBbgQwkLYc7ZDB03meNaqVwJOf
iS+wk0WrleZAeFkH1Pgo9FKqjbx0u9+86WuHaq37oITsIKjQ/jtfwKObFt15ctKx
hvzA3bQTJSXQRymQ2Jg0HQZ1138GFX6DgpNcikNpufD5/Vv1B2+OoINxiASjG76A
JSm/3w3m61qejoOWsZJKNjUyHqxyLlaJQB42LqbqGd6pw9NPxm38RHvMcQQy9uDk
OFfWtn0HUktAgIDvo2ESEXP0lnMzuqhn7d0PMR2BWuELuPruoku34VEcT+h39gd2
AoXOBjuE4ztKkPmeOO+cQnfv5I+SMXJSjrs3t3Ylqxnnd8v914YlB96/lb46BDOp
4ZKclLg9oemrexhVmJu3UDiQIlBTRvyeVmmj7Kb5WwL2lCMdgSdyPFln2uPtN0qD
3DfWD6wGYozFlrTw15kL8l8FpsbsaXqA/ZgNZ1iHbFdlpk9tQokEft+Y0xNc2sY3
kUx4QlgGBfjujPp2n3HopPfkZVyos7uwHfm5FYaewqetm19SLQgqvYsJ/nQqYkzu
6wCORQybz5YynA5WI8KCDqP+QCqyCU5qZVXC3pNZvfINHUuOk0z2OSRs1WVMKSKY
KfBRFJ2XpwHMAXYREMXM/aqfgrJiix2Xb1rllfY2phv6oNq1gHvh3GKgTzuN9ANu
oieLMth76YZllp8cxjzdi5addYxORe8iWHtWXExGPxIsTM/5joJr6dbyzuJZGF/Y
DKbqNjCXSXQ+axwFPNKj+Ts9vhWqKeVnh9nf8e0wAqAdjRgAk1vJjJjiSkt1/8UC
tyAj1h5LIbpCctdgj0ZYO7f8iH5qDkuu1tIVtIoROA4BC0CShXbkrdLYdfIEVj8O
IHF8i8KG/HrD7wBucJr8PYgKk9KiYtx+oOWBVbMzilbcY7KTjib3okij/a+cbMrE
LYurnPoRVBP2yA/bRdC9ijOIG17/aCuzc1sAhzO8/IskWnm9YoM8fBmE8BRpcK2A
To/0j1ssfxsNk6/dphyosyK0V5ncj3dDRwMadOtGk1tjs0VfjY0X6+qNR0omL3Ii
cSfGUQCSHvMbp3UwYvQ/uugvKh39w22WheWqStDvl3kjRRIPuX95R4TWpJ2rcY1y
mZLUX31MxL6/SwMD/EM8miQ1qmpaHO1qfznc3PFlKUPa0idBZiraywaZ5TwZbcuM
3tN2LWhoZwn87YrzWIwdrQrqZejtGq+7N+PhlD2LEnAYPEtEz63qhux57tIyhIFe
10mAifA411UI2WILui2KKmlOWD1NXsAAhCWM9XIWJou4PQjiRW3nyj03X8dhZCqu
N9H5y2LnjLTM3xhVkWz94bUR1IiEstpEoLpwGhu3y/4JWjg9ZkisOa+6wfVGWfLA
5AjBTX0cvflp/KNEEEA+y4sYxZMsjsV25zv4dMxKonwrG4KHYSo1JcySbN6JphZ4
DoVFNJcZ6KQkNEP1XeWrhXahpsXHb9jmizWfljy2Ah1Aa1JTLjS/qbZogTFnZM+n
7KnOii0wPJQcPufVBMNosfquCCJM+YH8+SwcqW2H3qiXMPqhQYKTHqKLIe8qklxS
yevcMj00sdUosh/fF7OKnoskuGfoIHOpqKAMAzcLPM7DZYDDiqmrz6EY+85iqlw6
TOgiz0XCh96ntg4oUzXLqm3szVNk2g3hY+cm2r1Eo+3TuwMbn0rb69BYV1+uN1Z3
MhtQQMkDmOjUygfydasG1ZbmIc+CxbcwZowwXVBDo7sZio0Rxm7p6R4GlvGO8irG
T0k0ZZBI9hrkH/VfpOExEzZYRPT8TOXV5Y566qbKLAFk98+2oGpW4rJgetFkVOcN
O+zojDzelOirWAkgqqd1dh2BxdHoWcbCgyZSZIeU+FIL+EN/brQT6dQXPzEoa/Vu
PIQ6oYnzLbtM32Juwtz9MgR2pnA1PLDcp2KPq2x+3ujZqNP2UvRaq7JelqAH3lFw
7jnsJxvnKhgyd5PukjBIuXMhW6T2udjbb9j0nDr8nIuI9RbP6yXsGFZjZf9hSnDv
MOdxlyLpP+bSGxe6GI1Saa4mSQfbarBSejipqiO9KlbIzk6vtwIhzv8s+cysxoIt
4HbBqttFESu6/AtR7qoBOeJlmwusI8losgLh7ou954MekDypljmlfyk7s4/YX+xd
bvaZul5JYCWVM22jQ5NFhp5aN5UG/9d1eH+1q3Gd7zoqssD3RMe/HH6ruhM9R0OT
wqLfuQ+EBMXGK5C1OvwNY1j7JSOfV+Q2I5sxM7n25WijBZPS5ZoQVep9DJuo7cbi
WIDaFK5Bq/m5va2Rv7MK94hqv+gRwLE7naVcT8tAz3DXtEGMp700vOWZme61ogyX
dYAnHXX72ONzYjkqrBMo+kKVl+KnhKH1wdqtnORQmLEGqPKx5EC+ZdZtSZt2oV+A
irSOQhCJzeaucdS8wjxG9QsOHusHGw62X+KNJPmjzzvOSEyxjmXPzcTp16A4m2SH
AoZD0U/KbcsMqt6X/TF1o1MujdVrf8SjAkYN9/ztAkuweaqSSuxYopykf2K7Q4UZ
hA7qhGpwg9nO/U3TXQuk5ZIWmkCJAvaoNu8ddEVRyi7i1KEp2gNPq5SchXZdojuQ
50gA9coP+jCfYPNzxJO1uBdllHVGcjAouG8BtqIzZ2NvZdERmsTaYDvQC21swshm
NJ4+VPr8g+2WQXfS8thCwYbHqeRfJ+ERSJduTM4RquY6cILboaRLQNOCNWhIQjJq
jeg+Hj1drLalGyGfY7qSJrEMb0HpYxvDYmiBw5y54G+WqGwOoo/N4f/1lzUj9HJn
wkzCAJA2DPAHW13KrxHmX0dzG0o4hXUdCBTO6qJHjlUiuutO5CQPlHnACReqJ4y5
4boSN0mnnhYGeJwK8f41nFXsh02/gR+hOP0DeZ8WhqDIMcC8NGOpYMQ8701AL55Q
f6GUFa01kYOErrfLP3iGejq/Ukh54hya3HzDOE9nYfDjqqDUkj9O5JODofQjmFmb
FNw2LHBGBl45TVuFemy9dHDx2SrmpHAfNyb+yPZj9WNuOUAnreXexpiMV8riWiYI
R5vW+aeZyP/bZ/wLCi+ZoWjCEMtsEVsFzIa65qIXUCcZMWUnT8GOQmlc6xX1yu+T
ZgYV0czDiXf0hVrLfWp58d8MKk7dE7MjigePcvPVOmkf0kGpejWRBFw9ocABy/Zp
Tf6q2VRjiYuIVH9LMiVvJv9Ukscd9bShj4bYWKP5IZLhXmaDZDuaZfY3N52MUbiT
iQLsNvuxrBIpXocRtuMyH4jY5ZZt37QVL1SMh3eOewVJZl+DFVGgWRZa84o+SH8P
Sa88fyKsvTnebqcnk+Shj9i4G2UlllQPkmoYicLV+rTwsJW4fBTc46abGiqYzPqi
/Cjg/CiEWNJ9DoZDQhBJRuTApYIcIA7WMNI32QEoyMlz2fAN2p4lNdx9CCKdovt2
BO5VIEkW3Sw8QlFxBe8FFvFq1qoeGC0p8YgQtC+myztYvQ+2mP1tw18mXM5ndvl4
JUGdcIfn9R8YaADmQ2YMIReZ4y13mqtMJrktXZyMtp5NH7BOpPH2YqbdbTecRAk0
uIjEg9hZKUqK4DLQq9HZsX6HXxo4e7ukBSeBsGLPQ3Y6S/ZGPVC4PfdLlY7aix7k
zcp5vTwf63sqn/8+iM85PgtD2S6BBbFC6AXmdn7xK6idSxoqO467vLkxSdnlv8K8
0ZFaavCh/BQpHk+6Ac5tLaHcQ4W9eTww8RJSaMR90gGQw4JsfPdlQBDx/0gI2xlV
r5BdkwgbOyu8ePRdKVs5CCuBNRTCcRanVhYycyL5V5gF64cLLK9BZhsOdrHsoM0r
xOBXotmG4cEHah5sNxvaww==
`protect END_PROTECTED