-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "N-2017.12-SP2-4 -- Oct 23, 2018"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
lH1RlaXvXZI7ctQfVcezxtSBsuhgIpluezOiYDUAsVSWLaHMSc59QEsvWU2Buvc+
OzMrMdrauBvuSwQkTmRNM0pL8Ka1jThLXB789kdyWxZJnGeF1LKTgWsEs1OZ+ikV
KuAsph9NVkMmE8BPQZu/xwoYMUfsx9h/BOJ2WeL56G4=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 27776)
`protect data_block
OFXxxm+T0lkk7mDG0PFl4aDZyba0xkbEoys0AQQWgY+CBVbuQ8/d3vsWEBHMvJY5
1WJCUpLPU/0hO2isWOHZtApQj0jaeZ+/gdxKPjerVOrE41DfmRhzq/nbqDSD86ts
xfUwqmBLPDIJGsEzPo0ZP41xcmp5WXbAdRummVE2eVzKJcBnYMLyFnVLEmhx4zHX
KtGZFBJ7y64AslNhwPATwHUXMdmFEyCKsXB0XiyEKou1VBx2K+vn7Zg91mmP/m5r
WNzcI4RNrjOfY1ZKNFpHuxd19kwT3fs9DvdG1NMrB1mSmTDpX/pTPPJxWhHxZbs0
u3RJ9leQeqITzKkyjRR3nIjs/nG4CI3QDgT36CWPAeSnNt2eaHdXPOwg0pFAszZK
EEElY0YIolUGgEbvEZryyssjpUuRz8Dy9wPRKCax19zAwwLlhhFiI3ajiv00xZPF
bpVGuJe3li6MaDL3WIg3h1JFhDXn+tdekF1FvloeyYONdfYPusHnRrzJArey8CNN
0u897qIVyUHdrzcLfE2dAxQKk9QxuhBO2jTprwCDG/o++DC4MlqYJ310dydY20Kj
6XpGJ4xRReyFyIVjgv5Gi779tAb2QvHV0blAhHwSZ8LY/OkmLkfG/wN0kDLXbTxU
5qxEnguiYQIdh6Qkbu33cjGDqQ4x7xJeTen2kYOrJzk++ra3EgOplR8M4yFD2WE3
BCRisNR30O7WfL1CqMm/V/aeLHwn+dIanRa/hOsf2nj10Y1OjqJaz3QpejYa9XqQ
t9MN/3YtLfZd5mBy32lRtxORhPRqwJtpkr6fjTDafdY/KDPUvGkTBpLqOJlQ0NIj
2tl+ThUm7sBifDDLLhYoM2V8AYYE0ntPNqmDcHxvqk8KBrtXi/Dj2u/1d2tkJu+Z
tzjWyInlyBWCesAkgaysTyZ/ZXkZfeh2bXTKHUUvNPrVPoGzDKjRHFdl7DTNIWl9
Hd0rftmrLyeBQmyFwK01h1lVks3mUgTJiL2rldbq2dKy0S4sqNt8Vhft1lN7JIT/
LoY8wV0uBKrMKlO/USzR0nhg+kQTdrXNvBpVmfnSQW7XKKTKwQikWnqbUKGdzKyM
IvbD407zBmeSlh/B++iE0DWY6qYRxKtS2qry7SLOeMqJfew0lmtSP2AKgWSEOVGE
Ow06KecMkt4WGPPhUgivvYzZUpvgisLv3CNV1SySMCzJ+2HJF43GtDwtqSX/bOAC
5uzes3UUYABA8WniLcn2b82KzPOM8oDtvNxCL07q8LYirG7t6UT2dNTNVvwja/7H
4BsgwEtMBwxIrWfaKO1sopXIU1qUBweNnZnd5dyp/CQan751XVFtenoq/m8Yg7HZ
RQw/T0VrY1XRIJNZWD+Q7RHRu3nyZzDAiM2vjlsH0dFaJSle/okcTUd/95B+nk5v
UaBMl2fxVr8FnQ83W0if9k0/ViA988rewbrJPq6HQvEFQZxy0e21nEAqTOZIW4BP
ATKaLZ9qeuCBSCV/ZzjGlc2EqwGb0xOpwGPp/s/Ms4/b4NHuPpzKmkx5HhbSjTx7
+r/IZfGNAN40aP3wl0XYt5SVs79lZA0SmcrXKHNvMID6qfqgxinJtDwzN5k+KNgM
mpbap89MhOUadZ1IQJno9NSuh/4mN5CXSGUzRBqWaHv1Bq17yJHILcPz1XgvYdXv
vu2zZnEev8mBPjEkJ0Sd2uN5BOtuBsEObP8mS2l/uE6oIpQrp2/aa8+8KDaHgYsM
bb7qwrSjnwgVXoSAAH/bCz14TK+KfEZXE1BMVx6IyaMhEgggNgYWta1mxzo8FMOV
cEx9BZZaCd0UJvHDxvlATnH5B/YCjofLam1NpK8WAdLIG/CSHCTNcF3Iz216uAoW
sA2rsrilgTf1TmEIZxWDjGkyvAYvkBBoSvaoaXRnSDHxobJQ80UvdetEumV0L3IL
ndoJ/lhYKvsI8s3P4ujqzK0aF2ElL0E8N6iJdjKGojWjqfLo9a09de8y5NIvbkKv
q7SYH4tTMEHIAz7ZoPQQS7qjid388dbjRhzAA5+CSvZq3W12x17l/bQ/crKLnYPR
Gwoou+Q/ZEQr5Dskf6cXhD/faFCOkafTeZvqnpqWPVB0DzE1yJyzVvw/ourkGyzQ
A8MAHd0z54yOwPxp1B3+Pli1gLqxgTQq/nXWiC4zE+QNmO8f6gp7NmPyUBLfCpVq
SrsJc80ACw47PV2bH65+N6C1SY/TeQfMGriR28IPbxJCE6FFAoy652w6fwzt6ZZe
88vuZSZR9Ocxaxa226nMpepxjnNBxCAFA06uZSHrmiCBNPdabaiY9F4ysn83I2oD
1yeYy4uDPaGAMQQgZDkZOiNMg8BcCiTZQFiqPwJHaJmVeuIQg0rkD73pbgGdCmzl
purFCE6ZJQnsgzW3+5JlRJ4Iwi1P3lBfYLrGCBZ5hH3kpfVCLJU4Jr24xiGKab6l
QzYsw2GYlIrIHPFxRQrWxlvqCjQ/U9zqTbYsBGFYTOaKsUh8pNXzoStyyZ2RODal
1+wMIETfbbdycUiiaeywGdyn20DKUrSljog2xEPk6/6cGxg6c2f9Mp6OnB0euxIF
kyZv1/+cagaLgtIMgDL9kWz55vnTSSocXttFQBBpERGjt6qJiQ/Iy/iG16G0RzKk
f9hUOGsRPzKwFjMOucAI4QUmB08N6sNRFTopS0eHnD5WNqWc0fBQlGud1KMNZt2x
wuq65yxxnE1IfLVa2oH+z4e++Go/YNEHByxK7WZwrToWYfsdMDNqHX40IsMgCgw1
c+MMI9Cr+ZDDypm1YJksNNBINsGyP8zCFIHDWUd392iXRGOokV+dWVLZuwm3Cfkh
vIHDGMDNQXrik2bvLOa9P2WD0t28gLvqDWB/+zcSLsETGvapAis1mESgPnyCmGql
NlDgzRqTjwgsV+z7ESyPj9aFoNvPe8XxscmZ9TBucfmMghWAZuVbAWe+kRI7ra8w
M22qelsBw/uULWnWZy28eVeNAlou1Fu1AMmBZS5y1t7wsEzGhlHd1mbK+5MxtNwB
Jy2F9BFnpQKiiccdxjucPqgIXiHFbbZQznXW1vosuGL1+ulBhvt25JZEYBJzzsPy
NOtO/yynThqfH6dytZ+/w/sC2R1NbtTshyNfR9Eff7bo5Fn3cVX+X5I8LG/w9jBb
KHu3guBSgkAqP8p3yY0VcOKMFAUreKT71ASTq8zG83DLcdKlgVIv1kOp9aZhP2Os
Q65D6VTnuOrZjS9J0fRFTjmFFR46iku9wOqHJvhcjYvNFiS4CfhYKJoHYYkFtHUJ
GQFmXcpLUFsZNm5VqGi6fu61A+BRQw0xC/jXGI0DPp1NoyuM9bwzphM5KDZyZ8Pq
xgeuRD/eIrH1tAXpNBVv81F0G5eduex22hnkaOx8bEbi0Qc9OC83pQLl4K5cfvAD
O1uPfhQZsUxNp03TFqoJLTLTaVvyCdGnt3m8jp92Iiq25AKjFggzltwsT0DCxeRl
8EwFU02b1BDPSuS/2xwuRn6ny5NrH48TYjFEQoPNUH39mlxldsD9q7JbK65PaEwF
qj1as7h1o2SNZVB5BXx9to3TLCZ1hJR77xx8ATS4h9cWEKkev8ltxLMQb8HqhXRw
Zhp6NRaaznaoey/g4v9v5QwplphX9td59Dqm1s5jALkA2a7QMQq9u9/4pwZKLDtA
t+g4DDp1KaLCmMA8RjEUGQxK9wLo+WZpL/pcrahY24HsrW5jK0YCrSHwRsmukOMX
diX54kRl+C//2LJc3QgJLmTUsQwZLz0BWNjBUn4H3S/Ft/Yjx+tDKoKESUmgweBh
sbNN2EhOmpPT654ASi709LYiq1zy6H6FeINeHx65UqSA6kr7GxfTa9mL5QUgmsp1
j0hh0QT+uUXqs4omq04MWd6eAhHTV4BCGeZJKvVnLop1MQj4b9ByzVHTbrbjVyLr
6VU2/c2K8lz5UeyyI2zrpC7D4uBR0OL4sp/m4cdOlJW0ZSdbQSU7hA3m7KiMxSj6
hlsfw07ZNkmV/2VE8g6JZ1lSRtUZX7ZnhxULaHKLnyh8j9C5IBoufWfSDL7SQAJf
ULpo0Y6iZIvDeIArB44wjFOwfkJIUkAgU+Jgc04+1C2aS8QbGc0MdJq4vqZOsM31
svYhQzy/ie2nW2OPVOXZHWIvdVCZ9PwNNmPlyzTJr4LJmhpQPsjDAgW3weNCDQ2j
5PvTENbbpwP8MsIytwZvfTCJ1E+TbmRReAXJJewNBIIpIkDJy1c/PK7Y1JWiNT7f
qsKPUv8K9/1GXROajFEfDvgIvbZP5y6FaEwNwmaWSKv3do9fLDmedhxL6Yt/CDgs
9XtMqwxEEWSE2J+Kop+lwwPD+qubcoawfoP1p3wINZb1l+HQZ4OZk1ogK3yrt3YX
dMLN9h4oh1GJ3eo4Zr1qyOE9855Cgxidzhoe2C1uXs1W1+TtK5tFaVrX4tZHxFgm
o1YXsipu28gKzNx/26KgQQI2c6MsyiQLJSpmU9ukQ4eVdSt8xwqb1lqrnzeaLdyL
TzkYrYIczv+wNqnqndLVAtzDjkwsfQNMM8d1PdFOWMQBqCJDPhr/oT+Hr45UGEHe
/4QfbfZT39UiVLVu8KHYu9IdJzlX/IEzenVIFFj7QerGwWvpBCEdq1WbJNtKAkpf
VGT0y7mwFASocrHd+5csQ5T9mWDlsqTlt7PkBK79OHffnGx0+Mf7K2l2oUeJBJtD
0rTQu94RROvQs/b0Kek5+opruIOXki8DypfxBgHuD0jZ3EZFgM10wt0iEDeNje+y
DdvtUjR83AkXe7f0oLkbWSZyuxe9QCwGFYIqwWw05P8S1lizEbZyj1X09CAto02d
2ffbRHKJ7jPEBHDZRRbxj7bpWXrv2osz/dQRho12no+VQu3Y4MkZUFkreFnrZSjv
0mH3dSvwkPsMXqB30qERvOOAMHvDOFyWFGNQ7+zuxF9aXhHkIYoUVx3g39LsEThB
tj7fO3BK5KVVUiqrk0zJuQySluoGMOHPLd5CpgPTDhNpuzanS/uC2Nr6OtxQ6qY9
YohobLERc2CnKDx+Oy/cLkWPwcExps6qv6cijJ+Hbac6EzB4y4dP1vxTGQbwwfjh
L/uKii3YgvfQmkn2rv/mAbGr6Bpuq4ZoeGVZOs/C/0oOKsgo3fxR/awqTLkDvJkl
E7DEAQfrJj4ZNNonXEiWIa0gfxmH0cRPFpJxTwxiPJtANG1nlHKp/Nhv+xhbBWOz
GBIQ2G5DysqjyRPtSgs8fnyNhQqYPPB6CYgNhaTa2oFtHjqylRTCMS9OsoA2dAIR
TSASeSu7Qmb7h7v2oXJej3Yw1orUD1Tn1QIQyvwUwb6HImbCCKfzvlMf0L9hQixH
YRffYXwjg1I5Ysi5j9L0V1ccSS70ROFzFZ8tfNZF3is9AiyeojVMtxuyqnkX7omJ
0Ua5eFIO8b/enffIT8NfTrdRapDbGXcoixS9g7BNasyKiljovp7spWxhBD+RoEZS
8QBOA4A9mURImukoyjRSMJ4T5HfCwOBwzBTsnkPMyOpxVaVN/OgpArtfrZsFnp1M
qZn0G8ppkSBSt9xZwYELCmsorYNQeWG+T4V2bxYUMEldYftCGBtwWtYl/WZZBUa0
3p96ctK2XsanyhpyZ+FISUed+MGEYGqGjp8gPBFmmo9oSHfRRN3NNMDQ4AZXdM/T
NIwaTdKdlaiwxvJGe7oBz+DWNW2HVSx/lqj837LS9PMYJF3+Y97gG1YWa+KXCfpE
37zd/bCiaa7yIbx2Li57Lw06SygeQa0VOhG0VR1QqdXeH7TXyU9er+KlJ9prSrtw
/xjXFpu7d0qHSJZwbgE/fJlAhAUGZ93HmNDR1TJzU2sWl2mjJLAPyNwFHeW2nPRC
J7ohgr+QCteeFyE2Qj3DipjgiyJpWnd7QU4cWqKMnDgEnpvc7u3NAsm8oso3AaFH
QKCKgvx5SEb7TraaQjffSjRvdxzkRMpg5SmH+dJpdUsNqzdDDInwylz3R2lRWp3/
4BbSqO3aXZwAbHC0Ao7UPjcw+JdS4sYvyz9cPubnOFqCtIRpHC7rxMhjwX5cC5MH
PHlWFT8rKQSmu+Lm86QzhGh8B3yDog1GrWq/gdxSS5l1NaI5vRRBT+x0dD7Ctyir
bio7JhzyVsk80eodl7fQl1mdBOoJD7Vd/z881g7Y7ApbFbNAbQGScmOEncDBGiU4
xf4Wzl6cd9L+gTjwpbkgWXhSRV265MbJUm7Pi2jLD5ucG2lXVjphjPs3W8ATc1xZ
YkqM9aXIUuzyLZtJFb8458P304oOFlfV7vX4jlTo2nWTXiFMUJcuqY0NJjFfP2Ou
10feGHEYhf0IZO7yfjOtzXuhsELyj51HbrNE9ZCkeE8ETIL82o+iUawQgHpdNMiJ
zl6RVdA1HGXT1PX5JDy40zDX0lWaBMrgw36NFLMr5kKszPJrWNiA/64iYAHbaa2u
/laBLUkeMLuTKws0IiplFVEwIvJinxtwICXUwyWvJ5Wr97W1NP29E3vwJ7dIUwnD
xw8H2y0ZVN+uYWs9eRgZC6Wbb2nB+JClcsH0mCGq/HvEObjn2cx2X2QvNRLX3QSk
nJgA7nYy67ePMCW0e6dSdw80B8zHqVZwEIKCjdeHVnFRla/WouB6dRGcammqsmWK
hDX6p01fpymRDfJNBP5AEmI8Gv0w0prg5GvH3q5XLn4pohfi33zKvKjpcnjuGAOE
lPWlTF9hkSXdLPggIAvasuyeU6dQQ+G0gMdOgUVvtJ/lVPJdmUafSX1vx8OqYjoM
gd6DdgNxe5RyrdeY6P5AK4kARrlspXdTowEV2LYDLK9UfRg7MAsSPalp7UzjanGE
kCbwiAs+X0LnfbvUKReCUM+dl4eLxkXUzFxYfTFe2Okr1zXPG2DgdH5D52V5fSGA
j2kZdfGZfb7rSloSUVcsutN58w/Iwj+mLz2cRSHw6oWpPmJTiALNtQC+q+LqAO1X
xi9aSzUQDA3scEFdhK3lVivqS8GfIKYeqNgFKX0tG+PRtymlO8gH7BJKtyuSwx3X
hHW/OnzMmzzHYMjL7SHqQdCx7iw5C2ldrHXNbekI8tVnoZhIIGhI5YZ8k1y+4jeF
lA++L+IhddjW4Gkx9JEooFq+bCzGnOh6Sw7pZ19KtFHhysTAi90HmWQcoplmXlrs
fSkIN92BdaMf/7+izuS8achXVKEHlwwNxZTw9uGwIzmItjfTzvii7xeh1Kt8CJay
MuIrkLUluPC+8Ny+2rKVK5gowSJ1fPAwROtHkanFAPI0svrjoQpNoIfcGrxS5gYD
WlAjQ+HerjqPGGUbPusmT7zcPmNQ1GFF9D79jLc8PAyYaVVqm73cBcURMxvsVEoM
Oq/SKQUSeWAWKq4GVnVTq46YMzkKgokVIFbuU2jcJM/74CsX0i3/MSzIjDScKT8b
2ooWj6byql2ZL0xGXB30df82hafep6OePBHzhHo1+yHh7hdwY08HLLomM0UUAfcW
zQS9qAg98Zv4p9X2O43gNu9kNMxKDm6ouEIkbs5qOdWm8BdUxT8p1amxoGNg6bQ2
UY0uJDxpaCHp0xMqkiOUl/2RuoN0gKcGiLB8OHiAoo3XDji6YSkgUzmsDQJ/bK1c
BS7vaUuk8Fnll3J2hD+RWCij7epVOqtINJYmsdEcmlPDFVqJLenKVjsHgCKXGgea
QKaRRo6RU+Xi1D44EFEIDowEhnv8LgMfSKcWrtFlEoUyXevSlwBtmL6Ab5rkXO/P
SEipvnBZ9umaQPCpeXRP8HwC53rhu00WBR6VnVEuNmP/YqG6Y5ivJo/FTB8eZSFd
tgFeKvVJzZ6m2IBD5BF9AUjyRUSAf/5GgW2MHKsFh0ihetV0i0B/qeB6a7KoLdV6
p5g6ME8p+PZO8QAd4PtZaQfrNsIP8Byu74KNYVC6dxOFuEuPqICjMhjD7ZDdrtYP
48CaxoNNgUvimw83t5SSOI46Q9F9D12yzdtveAFg7j1n4+aSae+nwpgXCkF1bpX6
Ha6V4heiQIE0BAirosn/aYhrDCao9/9+6j6FxqwReJT6jXkYfwqXsx9xsZ2t74/A
uuqe2zqfglwdtZaz61mpmpWl3Rw0RsG+thMy1w7wgERz/ff3lJonJRvWEB8TC8ta
Z3C5/Rb4pWgV/NO6ECdzD2j0SW78VsIPUS1PYsDZnV8Et5lAPTwauFD2xKImTLf6
6THMaB2DaSN0PtpVXC1W354oVlEAgvHDefokzdALGhlCmjKC7jAmmm7EOW64I3fz
aiAXKptK5Vqit1geQlBn1rW4lBOZLgHna5ia+MDqS25/vn2ArOO28ydl4ujEgRXD
8p1mWixx7pKuMvhY9E5g3ZqIVQYwQCyhYi6ujlYxoLrNTj0C3QIvoBmAlIvK8cBB
mWhUPVB400flYXCsTBCvHOrA4AfnLNNpsSMEHXwkjt4Ilg27L4eJL2IE/mACskz3
OacQqE8PZifalCXrxAG6KngHPEy4+HpRnHTOYHy0aOf72wp52vWxVxrolm1UsstH
zCvkgBWScnnV8aiWPSjzRg4tDfzt2+cIfIfGZOZDILwNAtKOY0PqDhfJw+gBXt0Y
MlY0kZpQO+BXxjX8AI//dRPGewgJvl6y2S3Z7xfoIWqLKDGJ+LagQyVcy5WxW44W
rQmAVW2iEw8ULrdZkWP+5Y1JKw8iLfezsLZZetGDbFMhm2xAGz+EGoYL+Tsp/fqD
+i1LnG8ItQQarEglvMocXxB6kQPMAmO6D2WgLoew2cS3NwzpXpMGTbM5Rzv9zV3D
Ilq4cUpPFUzFzZhbEQzFjh7/LWkX1a1lTpdVflNUL4seuWkWBnjnNJMhSGbUQPUs
R8aOLXk8/9p1qIbsyv8znQaG4Zc5Fv0mmUOKrSqEZRvP89+JmVLpf3HoflPpWUcl
RZPvD6PMWYzRV5ttMz53LWK+qNMqvNhLtBcKEyk6obZzqd1ajc2tzMds6GTwxlWA
gUbc108y91VvFpVXSOQiv9gyswdBSi/RpxtuwYE7OT/xT2ekTUq3dGgpmVEXnsmi
/Y0IZ8rsCOL5fY2CM5UWFQQKGMiBQC8YpEn4meMJuXA+wduOlOCAzbu0KIWk+qBQ
0KF4NSJ1qi/bdvBFfNQqwpOhOsyJCLQBiJHJTc2cuJL8YaAxOQrLQKOsJrLcrUhf
zGFDOYDALIHyw6jBZzYOK0qhsfptX9NO8k+wQJSEjr47CpuDj1zDqCWZnUQAYLh2
ntX9N2xa7MTS4e/BFXMKbiDi/gBWu87mPiiwu3Q4vAIGFyZf+LqXOpdvkPSh/3n1
z2JRhXSxt4jrv6ujpkf1sjUt3RcxnLlHjvRz0RNXx+hCHFA6xAMjFX3JKKPft+Kj
6FJTUwHx0KjHzfy0fzDorvYih7rccPXf/6+ud7qMGZyaSUewBY56lt0rp57HXXU9
AKfQpKkSdge6/FVKvUmwDPU26ajaZrQkxwM0zYnIkDJvJprtdtl7d6yzJIkDCBo7
Cxcs1lX5FXctGy2cJJryoMIAqeegr6ubLIP2hbKuBtPegw4vkGymLu/tcCDkYNSD
Taqmt5s6MBV5zkHlfqBKxkjtT+GGrGRd5cApcWJJVibXL5EhCYSMUUpY+KRBSjAz
EILBJZOPQ+CGd2pD+j8dCcTD+NbumhAgkvGpL7Jgo1FaWe+lDAJsJaIIKsFs+I/v
8ZMQAPuqt80prsk8WYf2Lp1CPLj68FUUg2keF8ECTq+2UCm6yzFXPZFJZCjn+fGE
oXHAMrHFmSEmzUqSV7pNxfxHUg2W7lLra93vjpA2MZ5FRzO8YqwBSWOJcP7OSkkn
Oo0LVWsiXgiXXZfbfrrM99IJ9Lo5ZffWF76Tj/f7iRjTxKtkxIy2FZWBmAymKnbq
QWTk1BSfagRJwFKrAnyuV8jsEGifib40e5oATbwGIaJ5Ri7WJ7rIG3lns9P8pjTf
9kjqr1/Dp+4naQV5T7dw/QHRmHDEcn1seYxJpkYQCg12qP/2+fZBnc8WWAgrQ4RZ
ecBxW4tTCuP4eNVaZCCFMDOZHn+OuHdGCNPFMB59Rt4eyx+OCDlUURQ/Flr6E9zl
in96f6xKGqx9vwW9Ar9TQT+kMR4e4Q3p5gx7wV1GQNscyqRnlxN0f/8Jpzzy3i93
mC2au5VlhRirgk+2veFUktr7yU8oXBkoAmVNwc8QpiGlUuyiXHkbKZru1UQ654sR
HdHK2Pif/+cAqNkjNPoAqsqvUupl/434qzH2TSRn/z27WxA7/8aD97TqncZhPD+E
SMOaPLys/PjEntpfkY6/Mwew0J6Wua7ON/R6zOD5r5ByMblUV/cgd1h4fGkCuq5k
D1bj/0nMxEPpOyxmU6tUWP/6La5rdFLDEvkx4VgxCeQb1aGad8YfiiHwF0taTUFC
woMeO8FIgsMx/986xwYXJR8NJ4m4mSOOgR9J7xiOMqizTaCcsY8dfBvrm1GYj8jm
jbkmsemm6CQG2suOdkQXjZg8NlD+Agc47czl94yRoVSdu0NJSM5Lpdtuks0E2OZc
kbMigYVJSqX41X0AmYLKdsLlcJTQV6IlqzViQ6AgcWnxY8+f89YQQZ7I2SJ3g5q0
MXDjSC84BXRuBCwLS/7KkDEJaMkZOxrn8+5Hue8zL0tAWHfIgaNfMOXK/Ixmn2tq
D0P5ThNYP6yVl5AZv7UdBU4e0QvRk2MS5/MPTi+bYcHQ55dpaf5K+F3pp/GlCLG8
JlElwWTBh23QhCKJjUp4EXbpTKNKbN86ZUrm47eE/evgrc8SQiozfBeMZg2K2Mlb
xtchfWUIjGgHzWHmsPIN9PIiqzSeON7YOphlW39mbFSBW/KUNZuq3TVlo5NPXIHs
WDNmwQUtidOg8Xm/QvYRGQU7dvnScrnaDL5M+6AB55UZbtAX29E8D2A7v3IHfGil
TLJznnaMWVKWi9eglAtqinRQtDTuTNuGPoqDiR4DNhFLKZVA9dbOyVM6001Vm10w
AYm9hy12JNcWVjLGdO1ftihsLLpayEEoKHQGotyu46yKYTzoKO6sQjLzf5RqwV2b
KvJW/Ql/6eLNtpMR/ilrGJdq8bCXYo4DGYijCHwqqjw3Py2rnMfzQeeHIGc8THj+
Wq3OvOkSC4E9R8LNmNwGLzsWoL0avndqLzFQ+QO7qM+saeDcgA8lcS7I9KQG9mRj
Gvg2YHnIgWaRQvj4oWnAD4GzthtUgZq//cPZKp/zH0IwxindYcXxdOpNCMp7ez5f
7Xz8S39zxyYAFBCjGPLytKboezgbNQM9UQ6nxuiLJ/C5ziYm9+/QT+DmN8OV1BO3
eXC2bIzHIdsT3saX3empchsNMT6JdF/NgV/eDF31R+yw1d3Xh8RbOWz53OXupZN0
xDg0OSPYcM/f0J2FtdmWlLAu0MuJI5/RgVRQJAVdbzfQzLjMTUv2l9OOWQa/wjBx
ctw6VaznyrWqDqp4tCycMnwP34ppy+WCwIEKPo5Cc5GXWpgQAxNA8V+d7jd/my8A
gQ5cB7h9UInJ7O1RhWsCVAcH3C5T4PRJMqPC1fuPFTzjkEm6QR5SS8YDQF3K3bkj
ckLkh4BgZ9vPGCitg/PHp4c1KKeeWclF0qrSXFrNfBF+lAoRHGXn6b//Jig2Po6b
48HrMaFYX+DIB7loDJuF94tpI2Xqi+2R/e5yq+bOG1UfrogQBZ0Y0QCJb6CjqZ4q
7HkkscHR+OpzLcbxupochB2Mgy31y1YEHJewbYD5pXXpsBCHUVJCOCs/HojqNBFu
noWHPDc9rnzSHoL3xhKW0OwjM+XPANhAIePHzPNvLYvcMNsovLcu4yJg6l/UvOIN
RDuWdpyXaeQtbfknmZEhAYlAUPT6VT3YmD/ghx+WFRvtewaA4SlMpiCMzWusCuF1
BReTJ6I37NBefm/YyNgz8ga96S9CT889pXkHSv/PZd95J9fMxltYcrF9/CQav/sN
bKaSdK8huVYErFHmSGRWofSUgC4OzXa0SiitlZk2RodAI5Z2HgA14PJ8R/Vb7OmO
kLIJ7tyYeSctztluNUWFqOp6AB6cL+gbGzd6VFOxNio6q3LtOjbvzoT+THAC2ctC
DBhZVpBA2hWr/1Bjif490WtooB43O9m6k3MlH49jRiaE0Y/wkFRWjOm0NjYPefgZ
FaH3e7QYhKrVRiNSY0tI+W0EcS8t4/3utRD4qse6pkG3qhfnl/lLudQTtofcrjGh
OlPQF/TLRioZ1ZRey/nYVuqEr++aVDvNMyiGN01g4F/rYZj7LLH4sHZqQblOx+2o
5fDehsTIqVBlNl4xP7hLB/3p7mfiqO7Mu5qCkT7nzmXwn0v92G8msxUu9L7s1xlR
pLLNAzxmmSkFrzNrylqw5B1qRWcCkWvF19YJ0hU+qwYKAKI7NQUCnUSd4UqlmbHy
AJO0H+SMScVZWbcA+gv9qVGhgq5uQYKiou7jYmr7S655uMSbH3YD8ptllzkvpydT
q1XAlUyQlCrVoLcWJB83mtAFg0WHSRSvwAPS+rEOXU1Jm6DyxQwjQHboPZI+xNfc
s/jnqrt9jcYDmXAgOMlK9AN8kH/uxyLBSHo+kE6BuIglxkOmbQnRaCQ/Fc7aCxVY
DGniXiVPWhnWqd6krLgxWyj4Ug8jGbcWyaD6uC813jpVNqPztP86jFaWmcI7VHGB
1yxaWKnASeJNNyAKywEyU/3hRDL4OhqdnZOJtetcQtUKXwpJFvqyV4A5HLtP0DgK
28wHkR3j0NP6AwvW0/CbvEstEoqJ61p4jIw6nRTDg3E7JJ82NDtgKX+lxTGHpO8O
rnXxVSFFgmDw1i3nABBVwhceIBbbXCcyAIioyFWqMEtS0/AtQJSetFpqKpq3l0h8
otOJO+CZ1ymaN/4bpzEkwlBwK9O8Tw0W/WwNoYbyLFZRdkEZtNnR3mFNR3H/LqH7
5BAxWl7e0Pd68WU3Xp62m/RYJm6++9urUnN+Df7z2RYY5YRz7JJT2rofVIwGUBea
xpplUp63tOYIp0v7HQeTRN2qfoPiJedueyU9DKscml84NuuDqjiOqySWTeSqwESn
ZRj7vMjxE+6PQW++YWWebotvXhzG+i6QRE/kv4OqKRSuea4DyyVJ7Ac8mRzugiWL
A6jlo4PxEofeQyF2JCsqj2Qm6GzZp8xhp5eLMVYkI9iQ2KEmPfEaYec3C1WHkvx1
EczE9oFVRKktcXPfj0/3qH7DQDtkWRGV/xvtN9gho6Ms9RkrDnpbD7hB1jZz/uMH
LE7WoOvnppKak7trfJb49Rgm4TnLLpzYr8aFpjJxc3SxtIHnBU0eJVUbAk06ckE6
PyLZJyFZCCGeusNWoWqq/l4o9jFbQHdGZHDhdAjQ65MjlNAvB8cFD7X2keVoX1Cs
rf9p+K0JDbIU4l4y3dvs7+rwoG8AhiofF19wfX8PClAkJumWsBOzDButzYigJjqb
l3YifWIL2OYfmK2CZ3UMTsJC9x15CDMkQeQyFW4E6/b65tYIGov5tRdd4XgEvCg2
iMAECrnM4a3NtkXl+zEO3CNfx8Z3TQBV7lcLxB0udlp7mEEYU+hmXFymb/KwSPW3
zjezvdNmKp51Z4ooZSgh7BsMNW8sRfKoi0Jh/k9av+c/78sNvHgf+4sjZbIjPDBt
3L1tKrBUicUxcGVcxPAASCsKnLmUc821X4vNIMKDMbHzijIAjXHqSbmJa4+q4F9F
9GNcg6Lk200g+Sj4HJOlRDRtGRKjm3ZG98yyGw7C9JcPY5yNAdP5oVr+5RgReORM
FCTn/ZCfltIGwIY4s+GHAYdLBQr/9ewyv5UYSu2aqFCH+lT/pVaP4uXUBGuuDGYn
So0NtzcPEMKPtFbbLjyxOib4mpalG31xOO/aAQ1WS57RcCuo3eSVdoQRAVHPb4eL
8mv8sfnRZMF1PweyXM/r1METnv3eIKxyoo3/Pl0dwfr28nKeks7ydecWRx+Y9Rd+
hBGPCNuE7XqdtwQJZuoVC1JufsL8/mk9ndlUhf6VL94/+HYKy7WhVxPU8wNug0ze
BKI8Yfzz8LwNle7YYTVBdy0Rs3pEmJtAuPYYAmviMqmZaH3zMx7XjTLE7CascisV
w5IZMPcaExP2GCsZT1JzcDs1y5ykUiEp3W4iX4EefW7sc+16lR2cGGaIlloNUjvP
xn3WbvtynDgIJ3jAey1CpBzhj1zq+XIuSNkH5F2S25PhoSUpQTRzQHsN4qADdQYa
29uV1lrmBglFeNdlIC0Iw9YGKEPmX/darXHW62NMFoeXsJu3ywNK0Doz+t/oH5rZ
cvsdqhM0YarJyhX9tD5iObVDanhnVJ8Z7Npxk48KpQ5HVC22RV8m9Qt6ZkefsXtq
sGkNJ/HPAiR8FQhKXhugxHbzdzEUupGSfMLA9u2XkGDFAMw3P1qwZqOad2rz96Np
4aU3dvg+LPRp7xaKH/EJmz79hvEroy4ySxFPcLwYXWdCAQUSW8ea9Aw0VQQlHsCk
7QR0yRkNs5K3qv/JBpiD4Py+TefGsUMar895TKWmtJu1nYU3HeWGi86xg8H51LGf
N23Np18tMCPRZ/X/ceGYzBg4lZ6e8xjE7pgz1E21DgpJfgSXkqT/9DO9YA/1QY34
HrxPQwVoHItvKBU8NdAQlfi4UiAZl8/WPrk15Tl35dW9AgOyVAAAvQ9PAkm0cen3
FbdOwbPK0PAp024DZrp/Y68h5qVcBhRLYGLsFD/iz/wc/nmSTpxhOq3pISJXsQ3r
RSlfSZYyV/S6QGm1/voesbU6u/g89iMWPXZy3pNOWED4HYCNNofzDkLM9bWDgelr
PlCDTtRoGXLixwOsPIw0GjePeI7Ceu/ZgP5W2ST0SQJYcU56FhogPdYzseo5UVmL
bDZB2gijf/GuX6fkH0SXYlXPU5jGd5r+jtggArm4GPoDA6tYjQ6oqGTOOlMyz6dR
khR7Z4kF47YgclW79NOrSHuRQ1UxgTpbHXFx1l2axNGn949zrP3FeWGZR3VpxOA4
wPbFu6WMNu5Wow9JlXg64b1Qarn68y6qRa3vLTQ2Sj/fs7iAEJouaJBDwMaeMb6V
LfOWATCc7WvNEcBZ4kIrcUapTCxxAl1KfgndKaHOySfnCv9EJj59hSwVpQrfS/Zu
4rDfgLaK3NqsZA3sezs+pKXEblhu2AxAyF5+G5GyNlNNdA05PurhdVh1hggW771g
uHRncqoJ58OSmXn6lhEmGG9/wKkEdxb9eiKVsvrvMmU+/CDIxnb429omLDfe9X0x
bZyqk1an6jB4q+qzn6NHg7Uu4tyK6iAEY0+c9+2LqJh3v/lY/KTAa6sYdEbA7H0k
i4JAL3ct5A/3gRivk+2GxovjBu+PWC3XvOvm53IvUjqFvl65BEKFFR/gQQT/d6xI
qjBD1IyRWmX6YI+7ePRdj2WmYPdcS2PuUCR8MtXjy4CB80qI5tWIgiTq5by6Q/7m
rzDjZ4l9/EHaNt6HPy4/P8hFIfKXOjkr6IovMIrff1dVH3O0PBLp6JPuUZcKmUqO
RN2gQqhJokS4InQWMPyc5GQ3PnO2VCMO099h4+elkQK+hzj38yPg3WK4XbKwvniA
bURrrDmx9lhuxnC/MwRPz9KzvoTRTAxjWfo3QYVrYRzvXgzHD9hJg/ejhnl9PulE
CgM8t/KEAHGTEofJ+LevsO5/UOxEKdZ5mjGGWoTcNmXhb7pj2K++Q6xw8r1ez1QA
tPhg1m3VFw4g5OskVBZSHXY6LPwLJUYaJ2aCO4pHatL+n/X+zpxVK+VaeNJIY890
MRPHPERdjFiDwEK5uDknvKZqwXA29Y/pbrjxoI8O3iIaoQVNc+6SSZu21Gco29Oz
aRNvUgk+YXGPC8Psgkbnu8aJ52A7yMRrEg66eYA94+S+r5YQ133B9ee3DGKGnSM6
+KWqNoQSD5HGGNKRI3Kps/3DWgu6Yi3cO7b0wi6d8eBvgxi4rxvaSJdO++zWMDQ0
C3RePLzcr5pNFcmwNlJTScqgevZjWGFo7EDCDBOl2amHTSgnRB+h9EcwdMm8yP6D
x48MuPiNxX2r2xiGC8vNxf5E/oQtG9m4i7J5BkJL6HPnOt47umqY7n3OuLT3Y63k
nTQQIQGRYLLNhPBWNTKo8T0i6oPDxZCgi4wIuSEy8beWUhM1Rb/Cihs11scFxuIR
W2gLNwaWYwl9xKB4X7NUQbNm6N5rF19+GjzPWa1QtJABKjJaNQQOmGWl34Lzhm0Z
bJt8hIG13vrn1SdBQR/yLCoVmO6xvgFGWSjFQTKPlKja9xKi7YIZPRN/diL5OpGN
cwBQmDbmVtxWToSfv8Ln2S3yJC3LUSMYXnMFe1arHRa2S8YsRf8LCXWqL897qvHT
LgLxGfEok+EgKtBHaidSonJImcY8t7YOJCXjAFbmRHLKz8p6XJV/NDusikyqZxdi
BZax2kmXkRZnwzANjLcob5hCYZZkp6FUp2Jlrm9DISJLjG+jo3GQIb55wusQbmYR
lN3hFIsTAqXA05dH0UKsOxm2wgZAh2SDOyUEnB6q8RvncIDwy9DJYDIk9r6HXXPN
/wy0hMRvF3/j1dfwSfapsDlAIW8avUPL/6njaa3BbFA3yKMgaQsHXz1KzqK1wnTI
xpW44iUT4katcflRCYVsgeyfWhor7dZp0QEBjimMdAnZYWycDhw0PpC5NDstCOUf
Yz4/OKDCQY4yCYE7VgMRGDxro7XrkXnroC1dmPUW4YfTVSiWqlbSIvp1XXQj/PuU
CCJnYzZLIq4QUK65koaK4RwwkDIfG9xlYTRr9iii8Dfx676Fdi3xLO8AAE9Y5cdc
GO+Gdfq4vmmq5+f5Wq/dSsM9lZaO0jRxYLfI0x4rJ5JNtkbtzs3pWDI0R277l5TZ
zHJgbLIF5Gm3j2vEgHgjW7Cq+I/SEhnN+2eYaTTc4May/JTJ0xCKlBbehQRNbxvE
EkNGizEzAry1pLM/OIOxlTM8qAmDKxVPeh7rFMj7+qJVe95gvBd9N1+BqU1rnuiA
lqenAlSreM8lu9wlhdqinl4Fy3ySWCrWokXfFvpdd9vbhPXbArHonuOsyWnrzdYZ
qM99Z3L6BO0k5bB8Tb4+0bldS/QqwJckgNy5rWvOOSFk6lP8/HnSqTAnH2OVN9co
F7ohKiOgiSZW32LoeB8vOsgifnfdAApWVaYSvJGqLcibUdugAbqwXmaAMqaO9D4H
gIcv5v5fd3zG546X4cmhN1ZyEiDYJrOjnY2GQo/Kq0anvzBe4xOmjlyGODjbqfvj
FKyhm7xJG68Lm09fei7Lk2TqoYkG0bQ4ccOkLGu3902UEoPmHVznPZ1wgl/zl18c
xWf7M0QSI0VAba5cZacZjVtvn0t27X2ZtiYePR6SDIQ8c5rhePzcZS8iKC4hZ1hO
3kxaE1DCbf3MLGtyk9Bh32QPswcQd+nury3jVlCh4FyPlPxvY1CEs36k9TSKT7yn
/C+DLMhcR2gzGq9CDfUSKzuMG2KlpHzbTXplMhsiDeeJVl/Fchkpl5IuIvKKIb5U
KGU0FWzwjF90KQAEx8mqes90ILT2Ym3EJQxF+32zEScQ5Hc1Hvo5EkW0g+MymHPz
HcWnwmcvdhS4rlbU2Rm0ggYH6XjYyjuyJcqvV3NeyyARGgai7Scl3wyw4NwC5rE3
n5hhdE1Svim5kyYtKpUVYqiG02LERoWP4gpeSJFo0onq90b+aCrn2dP2vn5eylat
We0LyKpYckwOtTqnfYOuiqGxzHHigKJ2FjoepwCD3RJOwD6kTlqaaKMoIIwL4tRt
4ZhPKxKt1MvTIJCPPHa4b4XWc0i8nijPhELa8tiG/I3xCO0qfUOUBS+rWRf58vqw
ch6c+cGcKvu3loBX549dfnjkz1jjvdcjSCQNUa7KNwQs5GN4RTQvNENAwsy1Ziox
jkL4XTP81BZhCV/LGhsNoLIorEJD6LOItthJRHCLPlYCoSJZnPO9FU6pm8IiCkmS
xdlbGfIYR/D/uSsuY/6vqTJJhf/5YgZNt/5GeHXdcWROnY/X/2FpaIg61fz8dtZW
Nd89jV77jAi+M2OmQANHrEChEvasYlD7JXaErRo+YV9LZ0zyUeF46XJy/2P7JSgf
xA9GNJn18W+PMLXL/vsLAxSYMsyZpczQPS9tK91UpLAnKBMFvKidjRxrM+Z6zs6f
MKXhQ3CWNcaprsj+D9i2FeJau1YGeeK5gho4yrE00/8HMekjJA8mqfsDF/7D2EJE
J3+CshCbMvWzTV/uyj995JBlEGvD67d/EaRGpvHXn+Kf8zCWCZJQq4EvsTLM0cXd
E9cBTLwWGf21pOZjx8W111NfYkmwprgS3bq7W4QVcs0bKe3yNuUNPAAGnCdDiWd2
907LzDdgJwN4zRL5z8RzOGDo38yPlU1XnJ6qIdWaCiW1JrcoxIdFXBLfD+MQWC/J
ExGocG1Mc4vqTWtIhbAfBemsBehqCn/LZIHDwLoE63lQEmmHf31r4nxd1/ZvzrEs
fAPs4FERrlNXnYC/z1bh63jVl2cC8qEpMWvNu51wmEcwIXpFmz/pikPvUOEUbMmK
bfJUTEhz7MmanDJp82n4g1NG9Spx0A+9nkdD1m4xRt2NkzliTdBtcwpLQNAEVkWD
JaRS9pU2pGDvVV9NMMRuY+qHmk9Q9blE0wm3wBsCy+AjBQaJFCmZqOmI/OBDj2+y
rtcc8oMCGvYeidFYV+HArKnLFQP+8hFCB1H53BL8tEdrpUTOQtlRo4QyZLGTQ+zo
7JrxmI8VNvHLzDA/3KMU3X9jQY8lqjcuMqYOTUVPgYvZsTM5nlLykWrbQSIcFBd7
HnDRGKqCwR7mvUzuJWLXv7Me7ozIFg0wqigUL0ws9Ulvn6dZ6pkgUUPLqnXiHh+R
RMUPEOHVTZhMSs3G9MBvcKh9OpH0DipD0b42Xb1TdZLBrvCbZeK6Mtdv/sFiHwHP
9aSpxUDGLt794kyeyntHa7i1bCtPm/pBvrksUxtbP/r4wGTX4GvQGgpEEZhftjaV
HGuj2YvtxrtuO/sCHRizZiO3zEANEHuvZ0OhnDaC7IRs6U/rI/3TaWZUfA/Oe7js
3FnM+HMLuJiUN14n4Dk6aZDkd64YgmbOlV0rfbmqmLTc0Ld0t3hDvvz9DMPie8oZ
rR+CBtPHLGb/Z6xatXefDSQW+XPy7LIls9X30a0l0vIPQF8eBDQBu3P0bWbEdhNO
adKJeG6yzL4BCfPR1JnpMYcjGLzCEG4PiQsljoHe1uQhrFB0hPxvhCIegSrIs2Yw
OhNu0t76pLNwWXWy3H5tdrJJhZJrxThZg72AUqoEN593oFoQO6KpLzwQO1yUiAe8
ayysax0lIKicGvwdprkry0WIw7HdahxCJD3TTT93/NF/9YEfCo98qD/0hAzQ495y
95sgKFaN2pf2aPCZCzmNQzLxPJn3ZRAc4F17LQNN0rKvATgIePWkdHEzJzS1qWL6
6d43WFPDDkE4YMxR84vawyu+oWfk1NTEfsFXzq6pZwiJwBKBEq/B4IsMKXHdtk1U
dJdGJn6jLzhFlxdvO4vzFbXPLRAN7/ETQFxPajua9VFt+QgeyteQPitQtLwiZqqz
jXor32JRJBIOCFqu7hJOiLLe6iPc8gtkjcfHI4K/LL2aretnD+pYr/2VkMFFt3QA
ThMupckEkhZXcMshLoIi/PmHsu/wNcU7IoKnE0i/KlJpxZwmEiGWe2olUcuKgdOS
umFUv/ozge3yuZa7pDDDH+x2RkhAS0VQxM8HIV5WY29TV5paMXVy+bgb20koP60Z
GQZwBdkdYs33Hgx/GJwSooKgQyx5Lr5pz9omaGgPweXzmmnpspMTjZcqHQjXMcVD
Tnfx2hFPGXKLYmO66ezuqnRXF3dUbLeAq7Lr+yVad8SaZp5EsOcEjrrXHlZcpIlo
Lsj7bZk4/0jCllWANsOBfRiYgnPnsxrgk8ejVG6K6q60tRo3qoPYMqfBeFOnVAjz
emzVawzoo33T65iM/8fOXqh9poLjohvhsNlm7dOIW2iK9w3XHh5OFDyyPrf6Euyi
Xwr48Jz6hwik4+b4jC52ls/6SvlYot51WTnb//oXcFSrXG8v6uu4KYjVKIZ/9JXc
L2ELfSnEVXFP3Fp2nBvdW8u6oRC4I/HzhlDgPJ4kUhokzgMdM/thGtV7j5358A28
BOxX3v8LjazCDUjR8rfsD220sYOnqxI/URdRo4i28bu4cutAtsXmAzj/tRSlISmO
4aj2ZaZ9sltqWRas7GPte4q2H04NaI7v22BRDx/c+T0z6KLqDQ9M7Ou79L7c5l+W
RE396ED3dd2N1K9Kjh2gbtcOEraebA4uGwFLhgg3QFyJqsUIk+4Mnk1S669YiFI6
bEWWdGpkZZkyuVXCMGaLtRNClMSI3d6RHs9HGNvaDQX0Sqf46C0QyqsIOaFgbkFx
Fc7iMb/EvU6PpIIiZG0595pfLZQCD70kSFMdYW/YKTEMnr5TgaYCyaLLgOpcKGTA
Xy6205M1HnhQIVkg/7HxHf623RF6nus7IJ7pIEldOvx2k3k58PuJNZL+fLq1LVQL
pnkhipP0ibdz8zpdolrdOGTaV5dwg84XWlpF80NrX9QsA0kK0iWP1vCs2Dnrmjg+
spSVc7Mg70ye2ss2b59+3NTazXWFYwTFEHHVN2RJGC2uFRliBtxksjT6Q52IVa3x
JiOpJOEvH3qUBx6GK9gme/UE6/4bD9QGGK2G+4f+ICxqVn7dVawKEzO+WoeKUnU9
3Y3ZXjSJM0ZlsDbz0Wr5LdT6Q2WwpjzNVX+4zq1DQ9GznVCpgddUjnoFhaoWg646
cC/TrMpYKUYgt26vS6mfyy0eYJ2p1BQTg25Cd0rrfjw09sOLj4s9KBDVJjkwTUGg
+/ko7U/IQVYICUoIAqBbW1Rwus722AlcXlJQTF5YPh4RD/zcqDo6jSPhz0/MknN0
8HEJQyloMgzXqZUkBNwEaB1gH1+ID7b323oB3x1L971gl5oXoy2KZEvl3Fiq9FrK
AJXfvvrkYP09Fulzpfwk+lAoF3GFFfIStfCY2O7uUUAbBQ7JMoampp59eMmQPoPh
IthkMG7NnAHXrSNBxZvPgJpf6F9jytYOJRv5e3UZqMkm6PDvNyRV0FI3WP9Q6uBv
SN4Fh6aHwap/jolDMqPj/Ra4ZOr7vP2iOUtCBny36/zfy1K0lfuqPxu35wtK3ci+
OcCwpgQ4QTlaJEAuSLF8QWjOqKYYPmrlGKxfLvbWlAw29u0tjYAnUvam5VmEowkU
54mpBvgjgI+XtltiJu1Y/XJ0qFpnSFMFEiNpgobNFFev8IU/n7IaB3QWeLi1iEUE
r/SV0CTKjrsNkWSSTBHyd+HdGwvetrcaiZjbfWd3sDDnBmz+4ayXWdIdUlAC+Nx2
fV5uA7RlP98FSaogMeLyLdxe3tpP5JBby6b0IoNorSu5D9Qtrx6SNDPQnq0Gq4vU
XYdbO01IwO6t0C72g051A5+yJP6XhKPvXXOcx9WYjFS5RSN6IqbjoFl25VOsQp+D
wd2ov51PKrqF6SO3DwqhpRDgHOoUHPP2QXSAapJfuVmuIjoBJvhtBCHmtQoRrYyA
yajPEuidDAagIiqpTCTGyYVWM3wDLCad72a/PLf3X9KeYjq6wVPGFxd59893CuBd
/eIZz6A2cJc+zY+apWvoTj+92OJE0skE15KcM5G4hogUdbRm+P1DMCZAXrJyToWC
0g8pBZDZ3VqN9PsnlFZHhMTHFA1ShDtTuNk3QlVpuU+ox0V5tql0pFeC3YDirVjh
qW76a3zVXYNKinkOk8/oJQ/wyiy+Y6y+KyQxAOxgJrpNXAUmvP8v+IYzVHjWdc54
ptRTbHq/2J9mczTHifrEYMa67x9+0VdHJjBU5HFK0ptxRSI8LA75nMLtGxqUskck
1F7BZK56GbJxU+Qq/CLhHfDX1sUCEoJPC5iKT1UmVtuAgekbsFSXCA7jPrJAPDNj
Jh8/+q+XFXEdMf+xDigCF3e5Ms2Kc+gHSrKaFf2IP+CXcZg17lhg1XZ/tzUYZEmL
BF2FkaPNnEWA3ob/FJtVp0puA20uFWN2WSBJd6OONlJcPbRxobABYR5l9kSWozzJ
87PKko6m7T55FtK0ILkAeV156ZMUxpJQIFMDgKL05td+awIKPuJVu95ie53mDFJ5
79GaVP1Kfhm5Hv9BAE5dDpt2NTSttFAAdZfOceByBz62s6sg9Gjg1eRclMXe3wVm
086mby/OxQgq0DjnxkjKEU/YhI2hRMPFQl2hP5zAH9E72KcJWOhmycF/Fab16iX4
PBJMUlDteE6kaI3L+eysve+oNEDOb9Vm0Ia2TGkWVl/dfEOMEkz7JVN6FIsAmSuG
goBvm+adEIk6qJTix33YuQdhVqW3sTRfWDXUF+8bsJAz6OFTCH/uDs5pEHb+N1Y1
Vr0dq10/8pv1nbfjDCVf7W2ZTqJxI8P4LOiOPT1l6B1VPqR76UVpPyZt88SJ9pvr
QIKaSW5MqHlRv5fedDekd2QNSDdX/YbZhxRYLeTguJKKRdPggFX02mzzWBCWhc8T
312a9OVFsbMntslvHoTN9HOTgHbq4E9gls2U6vo2XolUnY8tv+1wZVZyAuyD4hb9
KYwxANcNXjnMiRTww6ePrPdOIDlwRDgCsfFrt/ntNNAz+n+C5fb5LlLSiFdcgqPd
8g2z/tT+EREPHEU9mAwMJ/m0WA3Ng6c7N36xINNwYmM2hxBrd1AOhPreNrLFyDDv
/x8BqMSY/j+HaHH/y7tczL9MmTM2Ow87eegHgZdTRjlI+fow4iIRZQCZHwWiLO6j
7tf0btwMWzvbAG986IZkQWKOG0DGCNHbtr8LrKO6D7z0LXlHnfh2JmHRPqLcHaYw
pZm43RSl6/sgWRfcnLYkKH1BDd6qLOWxymnMiGoJ9TCzDCd63JxbiAQpn7l6W2+m
Ne66fZz+3IX1irk/PtwBDxxduoRa5ZVcWa9FQ1MiXD7AHrUFzd9halZNuHQCnBPd
xdlNi7Aca9MBC5zFXLVPXvohTqEQCNxQ9N0LVdrp8Ki6qqVcysIa2mS1JACUWSxD
ZeOSKi0sgXPvQcKcsQHeNh0QcmuaZ9hQgTYpxueC6J+9IxWmUq0lO45sm7Zqioy9
irPVtTUhqtW7jiNYavw6d2pkl0acCzkWHgEV223orOKnrrY52q+5wnB79p/NMJLy
RiUjnsa337UxtSGrdtxlgJRH7KCFGNzJeYDNwhxIvR+vSlz/EMBM7w/UyTF+8Qua
bVhUwGOZdLr92UTbMokcWa5k1jc8ixGymmF+exYjSeO2F003aeZ9cfQasbCiWDWa
5u1DociJSloGdnM0sOvU2vP2NHPyqooSNMwcRYT3q0s4+5dXsWBaykOqN7U16dE4
CaezTWBW0UmalpXFTeaKRr/FuG3nkuIKoW23hdTFtLA2bQV25sRuTlnP7ml7b4wj
ZCJi1RRophf80NzeF/bKpnGYenlT68WvOsvcwkygBrBm850A0BtTKGJdjDtIlRJa
zCEL0UcUO1LqHB1Bde/jWpC2DWFlYtOiNkFYP2X7Dpy8kwgnStVLiTveYcLdyVBf
s9YUeteV1keIVBfaq99xSVX4DsEEQjv51/TQPimRY+oEHbdbLGpogLxFtu9KPSSQ
vWR6w6Br+ok1GoCITEUxoJC6uxuRvnGwHxolKuMf9EPEN3+mGLfBrZnD111vwsKS
2eyt4tIy4wY2gUK37Pi6oIHmjLK+H1ZhtULXmxgjxLcOG5JP1FTP84T7jopWWDkM
Bgd4F0CKabcwdH4qRec9c5Rkj8/ygtssWNbh6wgDcdu70eGHynq07j857SXM2pjb
4VZHLPKLs2CNQEvkgLveUMG3SAIC2MTj1g2EIwEelIRTIC+vb2lXF85NAo+AtfBX
8p9CTozE+7PguXRgI3JFpU6J67s3Da5U5CYUGGLScokWElLrsRZdev5nkS/XmLDS
15VRnfxWpSV8P83SZRamufcnPdU9RTlPbaXMq+iAO86yymXpNp1SEmTHbPPhPQiA
Yi65uPVazf5SHfkTG8RwR5bEf/BoC00n3Knv488EAEq35FjbWy5L4DztgOpvuaq7
McAblPB9qrdlNmugGm3Z0xNjkeJMESIIekNckeU05jm5Rmxl562rpklMKTJFVQkm
TQ6couBX5rguq2xGG+06UyMqtNkXYm56ekEeJ+u8XKZNb5sXGzDNxv4RMWwyMSOO
uuoByvTRJGnC3dw6ZJLjxUMr67rdhshHk5x1TUHLMUS2q/NbeJmojSPm61R/77CK
LxSTa4UZWiczHogSlQMCobbVn5QAWnz0bWylWtC1AdhAsaeXSW48l1Z6viz2nqFq
tOlihsqu1lyU3xNEveWA2RHJElhziW4Akg1dD/2WEotkHcBJ2c6QnCwr50tg1+rw
EdL+UeGa29B4a3HIysnYoFIFB35Y+m1A58BqERex/t/8T9OReqo7vH6L4PFG3WtM
JntAMxw6trOkwYje9HdKx4uusWoIQbuWKHsnpP8lsm0f0+YM/E4xHLZtDumQV/sg
I0cMUMwWDo6x1D7TNL9l4PExcH86P38k9F1p/9aW81RAsGYqmk+RJKF3/YAWGb/Q
tgUlekkTMNf+wuTzMTVbs3uWkNIlbT1LShpKCQK3+6Z7UWTwLW8NyLlo78KH8ILk
Hze46/+ge4I7NjXz0N4ay9hkPF3ieQZEi1SIsCis3FDgUyKjGWlqdJh1Nawa+c5C
GmuvOFKvs1zsjXJR+lLFIqrOQWmYS4HsD1yH82e1S0QChzRFDjja0TryzoBTghqv
NlhrQ/dUnnF49sglW+HUg4qX8EXqz90+5+VCtukHkvnmqthUuuAyxMMtgIUYwvrK
8kV8mvSnejR//Hyng8yaf+gQZSGpWnpVmf7M4kR+Yec5JDJoXr8rv1XDqckgDKdV
/CFt9HQRqL9RfM4nevwWMSOmrARFTD5pFIsZaPWhIEissu0o/mYQg80/GAmudD84
IcKhJx3rNlSj4o9w1kDgHQgtAsPug5M818d6LaKa6Kn9qSAon/D7q9Ujb+WNV8TZ
CS1bkPky6I2UQPf4xE/gqlhOKrIaNyJcKQPOLiw6k9meCjTOA1AvYM8r0QlS0A05
yGfiLDF165v7+A+nUrOJln/sLKR+RTuznzObpBUP2uG4VmKF4tIbda6tciGAqqSg
o4IIUzmmLyLoh7SKQ2POLy4RfDU+TRd5i0vln2riZGRuu1uqOdQHEQpwxAyTawND
gjNzsVLq48woZ4RVh1E8IV8L+Wc/Ruwa/BnAu8MDJHcTlXXvK5FAlOq5r1hhB9Og
+618Qyt4eUAa7STxDw51/3SC3Eqf8IhM1s87ffjuPtaSkuCfl8d0Ooh2iP8ORMu8
STCpBaYJPcShDAW5crdYiKGA+5EKsHX1ztbknbwwIq/kPiqL7s8q1rfK11ssJ0lR
Zq9Bv6O5TAwWBU7YOZRU5PjOKJMLvkZwJ/IgXO2876YPy4q+RANHpNwWy5UgZJ1r
yxqfewm0oca6f9JYtL8DfyNaqIYvmLdv9PQfJ+ujinIVrWWyJYjebkkCbAyalKW9
h2eQyOJaXmlivsz6bpSSncwx1gFMyYNbaUR6v6oxQCtZ7NPYQeJ7nFQO9mNC4oQm
PesB3Ccm9UC4oJ+L6rm34JojDEliwThUB5oubpd0OaIpgWF1kHBylSfoFsQgEFnz
VV7RaG+e1RMdGWZ+DiLCN5Aqlq3nElpJpSzAnfH4CIsBOopmV1n8QthkGgVZLq11
H3Yc08HTCJxtoaX7uz3XybqakdSr1NsLryp/F7ObAtAu/Fc+hTCI1vntT2EzxxfR
zZA+Rzr1ixLJNhge2+J3D9qQ5lZBCTSs9muRcUaD1+Sg8fK713mp8VqKRYJ35p2w
yI3myaPWUOhDS00qA/ChdWxCvw2jCJYrbJtHyfKL34UgnMdjiufQN3fwrlTHFLH4
ZY7955wbyo12LXKBta7qMnt6KCgbxe4y/DVUTmfucITRrXepC5LyN90bu2A+Carp
1zhnDzt03ab0IiFtHPmlPZL448CVl8xM3eUiYh1dyjxfIHGkkIDy0i64ZRVmdcXp
8XhcNujcM0z8xNTc42oqGj6k5JtiyIvnouVtt+uJb9ZP08z49qYulEn2XgR5xlff
PX0sJht4Fkuy51/X2PYtJGb0pOj7YEKgjIvDL/2m+yzlHqSwnhlpjRGF/uKU6z6b
VBwfwCQXMaUyyR0hEBoNmj502bo4Z6+yu3ghp/eel7ED19aYTODd3WR4QDa2BkMU
4J7FNpFpXUcXi56lJa54l43QRfAQDETC1i0d573ZyS+/BhB/ysMcceWVVrzPn1v/
QEDrmG7MunHqknZ1mi6cC7mhEuIzo3x5PBITEsosTDgS97ZSuM/yAZ+xtoiwsZ6n
GeJgiQx2/m9ytAGNp4hZsAvnReYmyrVLPmf8529NHUUXSGPpEL3gIZlU9EG2kK3G
oV43SZsEu5ZFJf7/zNTRaVRla61+ZneqpzKLD+N8L8UvUtZHPXLpR0XMbJJJIfl7
0HLht8pvXNk/7+7p8zY1mNjkMQ0jJ7GZZ7sR2mzoLWZT9fms6OLIf+Hk/MXnfzO8
P3PdDrPc1F9bm+bMaBxManSsdBNc/ETQp/9V5NnuvBNF+JqPO6n6lKHS3kZiHo/y
7+GEdRNFbhyfcl74i2FSaBt2uu8mZxaQ2V62aKK3FCBxTqlJsuGFHw1xbSr1hV0p
f4dru13JhJXEBFAVYTT+1tc9bMnFaXBf9K9/sPY25GrFw0jYcB1RKws3gTFmiqdy
XGvTlOUYyWg0UZBOxO0oJtG6Hu70nUlFFGbjUdWrUzMBpL/lLObeGHT3ecvCAW6M
m4UQCJQ9tpiMvHwMUF2p25AQevQWHpJkYDa3MZnzmUm94L+7W44qyBe2xX3VqKsz
1P3cbEfHVvWzcSTRemdRPAwx+8T37PYDEP6TcI0YmPoJPzW5MmXFqP8yQmiUnE4J
rZrtO7Ou+OGKwkrMionk5/UjLebKETy1SMGrVYKoJk6W0/kBPS3dJDwI5h+nEHF3
9oTzzdsB8dpy/HZ1EMEFIwDrfNDerfoZTErP2MdjfPx0MjcQdfiadhbQBNaGCt7Y
1MSExHyyWaT1rkC2Q01Ie4HBSGaHvm4d03IXaiStW0uqfGaBDdbHwi2aTyTTgeoM
qhT6VE5y09su1tN/U7zhX5n+0lx8IGLfRmVRPiMUshr2uoGEcLSExFuFaqqfLL0d
YzD4qbd+Voldirx4sV/x4/qmQILaRwvwQNfDkC5gIAjzuXLvtHVcOHjw9GgXgsuq
4CtKbEKTdr/E8+d7c3VxZXPOKhEAIoLfiMLz8IeQ1HlLO8fV4uTXYHmzQozCQl44
xe8odcs4PJU+OYNvF+ZQJxHDF22LFPFfALOOjyc1SZdMEF+ZTBX0NUPXh9wIZdb2
j0czgOdrl96DIwTkPYV369oQnmsWoWbHlr1EuXn791iu5xTWPA/mReBSR+VSJlro
4TlfkJP+30vfmUGMERqpcB2aahViPC4ah2jb+o2DOe8J2UGQ3sBfmMrO0FO6AmIv
n37jkeYjm1pd3eip+ZgKmN3T/WAqxHNnvrdv23BnDyswXDraq4D3Otc5mlDDBzy9
V4dR71C+2lZWC53wQGqjR07TXiw+Po+3QzbcIlhmPPO0KMXA0SbjENeF8LkUfNPh
XpImQZfKQQ4bj2JraKYte8jzEBUDVn69AjRJAvxS8Y9WLpOZIDe5Bmys3epX6Qka
oMOoQLxzgE5Qfo5D2UlIEvRTVYlZFRP5ErnW2AM3QwIZG2XuUSzPn07DY0bAMzFp
gaze3X5rJ48oLe32BXpV/AHZ0E2lZHjgfxU7Lml9nhHxpfof80hxfdSo3DfHcFgm
of1bTtTxJt1ZfAEdz8fhUhsfvWOiVadmWglBVpNn7y3TRKpMOfYIcNjl+ncVNz8r
D3zZ+2NealLGa0I7mdIGEvIQY/mISE9qo/i9QfidZvIhGZkBkbL00WM9FYA2Tpp4
IJG7E1gv/jlS0WLTYCBMuinLIKtP82HWKerQWZWxcglfWfvIJ8m7Y5YzTQNAUnaM
sShZOk5ALwzsAv72294naXZTaq7iqyFOZ8sgj96KUf6IE+NQuQ8X/T6Y3aVeozvz
1vuWnamcdXHTPtPabpb5NLUP3Ps0p2L0fxuPXVAig/5B3NL5OT3/FxzKjQaIct3X
9Cj4TXl+wASSg3sjJqU5JWQ5WsSwmh+L9eLkrih5+8ztj6kAMTipK3ykKk4Yrp2l
xKw0qgPCKgxCojjnmr1J3Nt525/gFLbIccJUv4wXmYCE5kzSvqVLtEDY2dLtsEQu
y/SDZIexg0Kn2MV6EHWdowyTN8QyYwb+emhshTAC5XL9q6d0Gnmhatxeu4e93oV3
QBrLzGxrAfnK6CqRQA4eHSuvZxojmPcjBxQHQT69+bbQsRxMpw98GsMJDjyEEXGx
1h9TI4TC0r6q5dICrASgsC4tPkJHYrUP94PMlqkrpExu4n1By0ggNEzRmluqtHkv
NzqD2XN18PVvlh9VUevBzyNe83K5JO2QXqIDjCEt3yjGomVhjW+L6XXL6v/1sG8r
rGl1avMtPwbxF5KxX3PjC/eFNlFHFBsnvDkHCt2plgq592cXP2EE/GK9kygg56Hi
emM/LLy/tQYkHKsMtmFyfLJc9Q2Rd12Otr7vTQ68/XQzGJmD+U80XKuTYH4Kiym/
G3z2YxU/0yx7HvQ4yRaqZ6/uBm3tKpd11eJsl0uuypdrcAN550klBHX37qgm7vAL
RvO/6S9XEmPe1d9kx5csATdUPVtfU/R/eqhVkidxvFLnULYRCwelBmmEvc8ueytB
AJ2VliR0to39q+HDSK8hRMjkZATpAKU/8/ZzYGD/M8zZY+9Qq4L4nVhuYenwM6GX
/Tb88+bq2Ob3tL+PoeEPQtZC2rptMZuu3Fh7hlQ0tAlJDyPIM16iqtdDaLyV42b3
hrcdpCEIu0Vz4HRFzeswaB7tF4mPfhAN1GAtXfV8hbJSVqGIGYaU6WKREbcUoUMy
hj4YpdLn6852gCBhEeZGP2CFGE55nePmHN3U/73cRW6K8RGZP73fe2Q7pgAEBIIv
mjB7n3+N8B2Zau3bit/0rJNBlxem9ef91L/MTRP86Cs5VCfKJmKr5JJBz6rro00f
4anmjPN5veZiNvNKS8WRPnmLtLio7eSW3J6llx8fpKEMdEUqei2cPCvlEY5C5w86
3z6qo4OWc5nUJqBKi1QWMFaYX899DZq/1dfmrOnJhr1HgGq6icPmYnAFHADsXJKE
tJPfowhI74rim00husrBfA0LdY3rpyey3o/ve1hfP+KQ1+hPmjwXfD9JYYRn5UvI
X5IfiiXDa5FCZJBEai8zXaPQFPJ4B/f3gs6Wo3LZi5JDBxVB3mKXzO9aM/uR/ake
ojyTLLlY57AyXiUvCOjKO80lxkDLxjXbJlmW77nVYgFuqt/IvKSYNLKbttPRssOU
Dbnq4i91PkJ60fSlnf8MSxYUVNivXRP/ETcNlice0IA788rENRMywou/O+nJAHjC
27hOxqCQzK+RbTz0IwLFzgcP7qAriE7M/ug+1RS9gEryLeaaIwPQx1XdAQX7nqrx
fZdwKSWVTiXObOdc3fq1X6o2BfTnL7Xxap3PpJlvS1CFmR6Exhmq+C/yhLB7nTxa
94rmhD6BFNrRZTnqwh+kSMa8NB3iRr/YScI9JMgar/vbpxNQKYDL6lem2f+I+BkE
63unb9Z5dVmtmfdWgxbnCvty0uEVSGvRlFDmEw1dy3ACwa00jocSKWvO+udu65JI
BklNeGAXOQnyLhuO6c8Ao5L0f/2Me8XjlMBGmEl1tc0/bbrIqunDIRr119bvZaGZ
hIQGztP07FLNjrTzr6EfnCAglxgCQ4w4LT2F+qnHJ+KtOVbLhyEk0VF4Tau96pV5
UpVtqiJ3coFgE/nWXVqPR9q/Z7v5KGDOYLN7MD1B/3RHdLZQCqUYKTDF3QPQIS8q
hoRa7S5WHlBCiuMGCAH9gIKtmkb3565VDoI4w6MtTtbjjZrAThVYdkmabBHJqQM/
2ZV8ZpROK/UK+M8zGZbPVyhS+Wtq7FLMscCxmbFB3n2oCHswpqEdyB09rFWvJ5p4
+vQ1jOh+Z+yGcJLtxeAjt8qg4sWnA1x+mJ/hZOycZlrl5gN0mYqdp46B4acGaHGk
eAiakTJXf9rmis1KEy6xaovFi46V5l7UcMPNfz14uZxwKtiGghDpdc1bgfaBoulB
yCmTJSPXVlUahAEtDXxXOeU7dkoB/cb0gmVVmtAsdaU/NS2x263hhVcTPDi8zEYm
U2jQFX3+HJmN+j8NhIyd399UB6dBKvavM5yC4mumiaNJkRsXtakIqOh+/sUlXtZq
SoT55dQuxW0m/o4itEXW4GM1xO/0DXEbc2iclIe7EaKNuV9ziLp1g1Up0g5pklXZ
gAEDJPegwdZOZhA/6yFP77cCDTeig/nRaq2XhcyF4lFlYNpIPF+h4Kxh0NGNy6FY
oIrZZ5S5eMi9ZC2XKIP5OK2clYtO91u92bNfq6iN4MHjoGx3yaG7WOmsU0CK2NCG
LWvS/gZt1pRpkqvdNM0c5cUO1iHbV0K+ShBm4bRdlpySX1eX930QhoIica0KZKPM
6KJLs82Xt1R3D90nOzdkUIVTjNDVfqNWsCxUrukixgRNKCP/U1qAKNjKmStsmrkW
WBdTnwnQTWfYkfoW3f8tG/Xx3Ia8ccL4fa7azLKP50eiuT3ZsRLak+odtoHyGW+t
QYKbLKiD43wCRGPnj47tWXdX4cETlAuUU6BFAM2Jz/kRsiO9LyT01I0VKB0txTv2
FJ2RW4t1tkqSa28V7H6ugN2lzp2cb59aDBsFeeD+DNZ3/K+jJ8VMbaG+ve7V5pr4
wI1uUF56MIDKrtpd3pJQyZzG727yTZR+Ohx8m4pY0oUHyhBIllWAMfFXphC3D+W2
K1tMA/Drpott5zECDzAtNbtKiKcsdFAW8Sf3lE2Wfe3ofNH7BkPNzXW4tIV/lL9F
s8PCs+Fi82rP6AAEANeojj28mV7y0RVA8PJMEKMN/hW/vd7WwLHnzpvFq4+2FD5Y
4YdPjYxPt9EBMThOZipFLF+ap40ckQquRDpOF80CXqpLlPGPoqV0y5VtTLydLrAL
1NMvkUj8zjjd5ypzsag/fYBwvTmtqhBIFPhiT+3AdXgjGjyW7zVg5h2D5fNoomcc
mcT+KxOLsM8bKYcYJVLwBs5Yk+iZ0s3IM12mt5iXuV1JTXO66KeiRJjd4vagOKJa
p5GgN/vnX4KjUSH8RJS03kg/2p3DuJ/XzkEfhxDJP4ENI7UYFIpStC9Z8hH5Gdjm
eyIA/qM81vvQB7THSyTd1pQOxV2zEmYWyA3kqF1Eqo0L0KqhCvkrOpFDHdVU7DEq
V/GUD2usx0m9XGbtiFL6UFB/UxUuyVvJjctHa9JrrD21ReWwpI6021F/uFfCnAGx
AInKFy3veK0KYk3iSDsUFCe3L5R1LyyuYKxvW9opH3+FTxQSZeoLfMOUL8igqXaD
uQ6YNApRd44P8zNYL0GhBSr4lwwqOdgnDjd8LBoO+Y4yBDzTG+NsptQMZ0kDDfq/
IN1W6rkwLMY7t8d2SAwQJTRxAHI1H7Hf/cnCcS/4WDF3YPVBbKlNVz18Q7ZjjUU5
XOPElTsTXnhcaTmcbDxrZ6VYtaeu4MGR3spIjIrQIJaz2IGNJ//kf0sE/JTW0zm6
mvlHIoZD6jOE75EidZgvpOHOfrvwtUd84SSmNMEITdIjyal2abmik+f/CBW6SRtu
OFzzIu1uxMRkxPrzXOsiorZQkd3ljo+/Y4iawqyqY3cAdlv696SOkoWT/zP/HALZ
t38kADbOVsV0zKovn2zfkQD3X+vaBucQHBuaAzR7arbGhNYlnHRFGTIofcqlLbXP
8PpVAMMB8cVBBiNoUKxsybbhEPkeFPz0vvfmj9Z4Y1dBeFfZxK2BSziWORtIfEK/
n++9NJXpJgEUYbRctej4T1MCJDbsyE9GwPkOA5ZHgGkEn9Ba0/xQhglXIp38gZ7j
D6YPg3EYpHOUQcKykn5nv1SCDo8dlcVG5FKAICg+tJtgRhGoN40J3Z4B/uhyuQGk
0Jb4WHwRTA2/AzYkQCfbmVaexYVsIaX4hQAE7Zgy1oGIfA+Av0VVXv9ReWporK1A
KfM6eqp+MNOtke9W29/6QktcmXGg2Jbg79oPJePtjO5MMjb8sCXpPxUVDM4vsE9c
miu3GU2s9fqhJByXxs0mQsr98iuKRtGzDc3DN0VHcSSeoYIZziYPFrnxGpaNr+Mb
C4VekITVkt2fie284aCMItGi2rxPG8Y+SO7MB54KGI1LbIT1TbC3HaE7Xg4fN3MH
Jis0Ym9x4SgrT5oWONyhe189kRBClNYEzpJ9+PtyNzz/uSvcgcCNrglMBvjW3fLf
AJxlk1hnfiefKLsFz5pwLSCvygrnUM2sOnbYujxxyIvMbW/6OUhrNjLw4bI0s6nH
LHUDo97YvRDA8UJ0K+6dq1Xw+EI6lXo7UYTIv4LV2fmZf64Oin/1k1LsiuyO9orG
iqbG3bEiYKlS6t/xSkase8bIKx0yv/3uNkoq7kfuLeQZXZzseYmKGLh3k+i5JLNw
STKd+l1n3+kk9+bpqR+P6gpnOiCEcUWNfGCPaIJc24/oQRIsGE7dCd30da3XJuX7
uwzM3kTCr2QmIZJeWGjpJRpeq0fy1tiUWX0dfn0TLM5unQBvo74209QEwsykohul
V2AqeDuzmywaxZ3RyYly4Jr6G3ai9UEq8jZ+tsBUTdoGByJF7S94JEUWMhZL1nTP
w2elskuPIrZZpmQr7wmdJGwQvzD/93bugsuMYk35aeWp4qaCYfEM8WyWjw7wJkp5
81rA3Cn3THvqCjzELSFNZEGVL+GVAbH7U3TOcVms1mPH5POXQA6L4JbQBH5c8YsX
vu9giRPPmVnThRWqcg80EUjH3tlSz9u3eN3Do7nOYDkT6++9371qNrzDmEvPO2pr
Iwn8C+C3N4TSBN0fWylDchqBb27qK41mj5TDQQsXg2XGmkFzJVHjBvl0kkSbj+oR
YBS0NrH0+boVxZZSqYoVUTJYV7sH/HvS1HAudTOJTXd1MAE1+0xoKAT+GADuvPW6
O1J4x0E/M4kyClZOdBNLIgf+ODSSMbK0jdxbwJjSGlppRWQpY/w7CwZiw8AnEs8r
QA+D2LNJfxzZPy/7z1tGyOdntCbYRH4hR6qMyI6aF++A7aCmPv70cKDKkX4Bl8Wm
wDC0ZtKETZEqlYofd2DWPd97rZ6WLuAJDSsNsZdX+/aEACrfOcMRQ97GhoHveXu/
XO7jUo1OjAIj3ke3ELQ0rX5egPBoCX5I/EB8cLRXaqDmSWqjMmeI+268HLH1b7aG
OmLeb5G8QvIXiJHF5RxE07P5wTzd1rdC/e3YPvylTSTc4P2F38u93f4xXti+bdTt
fjpajtp7u/9xx0dWk20oNwpYgUBhnHxrmLj6CkLUzfKMMB64X3ucznzJftwlcRXk
o4etuT5mC1hZT8oEFyxmi2Y0xwF5vI5arenHXuM3bVDthvIZxrVTf2a4P/Wh7x03
veg7GRvjiKt5FBjIQoyosMc6rjUMa1pHDPh/IvuvOS8bl6xMIi29D6z3K7ntUwf3
ebe6x8SIoQj7fjr5FMiaGZEe7l5wh1iy0LSNv/Tf9c0KA7USQdWIa0wfpwVjZ3e5
nLB2er7Gs+BBu9xASog9TqHMQAm25lBh5Fl/wr+SX6sgyMH+aCRAmFmkItSq2AD8
IqDKHTLsGQyQPsEa3JV6go3S1Mbbc2ElWwhNwea28jyPYCA5bSS6tg1bK9szWO8S
q337P4oS6ogEYe1ZBsse7Z6o4ypD2xVtVRMLmjn2MzYTyNKD+DV9Xm7y3fTes90v
iD1cZuBCiDH8oCDxATKgt9wSi1oviNSA86bm5H71jdLSqx0zqf9eKTCFJjyqP9Ez
ars6+5QP8DcK/qkyXaps2NbWCkAPR5Sva7WPO8MmpD+RIH+T3HLlkuF7wxRluU5x
MK/4XtB7czhlkC+/ilpbANRTLxEgea3z+Ax9vd10Je2aPREi+2LNqotfxBa0o1Zh
+PLrm9MjY8QIy0sXiNf1K6og4uDqCYQsO9FF6WoLgY4IFe6+nMTPfDLckKUptaTV
mNROpnUlm770QOFbb+SLlQa2b66Ac8QFyTsmBDFyxMoW6EruBPUHt1xol+ukAM0G
lbOiG8+N8J6oo0/BpSJPMztc40rSN4ikJl6fC00AoxE++twGkTwoj6S5RqLy7H8C
6EkF8P7AODK3by0Kbaw2zMDsZU/Ws3GG+KrkFgPlkhXEaU7lWvxLIrhHXLl8vFqK
Q0lkzR8fSGOK6WQcVU4PB728kJf3vDpERn2k2U85/i7wbn5SpPAPdEumWKKE2JsA
akYBnIi0BbksAbTq19wsTCRzeYyfCUNBoHuOUt558nxX9OFz74G5iamJdv9yTC2I
jOl2+f/5hkbOT3jE8ofKST4DEzny8vOapcarOPTjQ5y1bxwTjtX9m+l1I9+5yuY7
IgkJakLvPy8pfj55cLDHlnnKX69lJ3WbBJYoVv9dQ+5AkgfRjSeM5vo2UT/P3h5Y
HPEyColuthMzsBeEbiEUwYTZFZV3Hoz9nxCYmbnS+3N5jKQRKwvm5nMUhS6F4kE+
i1SgDXXSKd4FM/2H/oiUYNjLDwknlPUJcGGvmNIGr9z5eT/d3s3GWqm3e6SVNC0l
aXsyFj8nRqfR4Z0T13j6sQ3rtI26y+IDwq3qWQxa/kq1hYmF6iwIgrzeMNeUFEnk
wnxmm6DI6QKMuhX7qekYTIGvxQjmhOzmYu8VvvyvEfxDrux4Py6lxbDgl1SUd2sl
dRcv+qLu+SF4qMv6eeXqS2HxR2fDP7RX73wcSuxc8RTlX7k6jMrF//tZbovQs3k6
aLmp4Njm7FHYSN++lRY9mq2hQ1wb4NdpaqKGoC3H4Ojcvxx1XZCkP/L84i9zkReT
7XUcG47QqcecZJY8Web/KYf2avnDDv/IR8YjDlRH4ik/rsu0x9517fBTHx4qLxRX
5mqRIaw3CyYwQUwRSpKBzdjhPIlQ2si3bvoTgOs0Daumqbqb8bkqoyAwao+4YcqA
bYkRjmp1UVaEaF0NPgNPE5QOkkPzRBH5s9xDmOiZJk7yavTw0f39PT9MTEEsAWsv
qg41fCaVI8G1Yc5CTd5Dcv29YeXr3UO0zxdJWMN91dWKXqODl5jz12mKIbEviB80
bcV/CovIQxl2Lqdpe+HcKvWLDPF50VgghKp+j3qVZfBEBxSLxkzJ7KCP1kRcJYAD
d6zU/mFzHkH1INcgRpaU4WqflqjZ+FpS440RpvywEL1Y/7IHeikwyvxNK0gQDRIp
nipvMtgIkk8+Irhyh7azaFwq+kyk+USGCANQAdHBXUHt76aBJjwFRIrY+5+UIIwD
nB21Qbc4rTc+LOxUXYhiOt/dc8/84bEvzdPpBo59AsDi/zVdfy+5PX0xm002GbI9
FD6yQume+aUV2OEiXss0rbocj/6nt3KRD6Sh6inzG8/MTGMsU4KwTAyXcJR1unwV
dA9hc1lVPMnlSj0WVoI6WLmCzBRyX8XWrC/pKOoAiOLPPpOV9/3kg13+GkruAqkz
9YfzzWxeX0PRj0WCxi8xzEwzlpBs18SRKtMfAtNp4thFuX2Dhi2jQOfSzR202/U5
83LxA3XHx1SCHdVnE2/54pBM6KPG0NS0yVi7teAwBM+zbhiwO1j0Lm6VWRMgNb/C
m+0APlKse4V4PQ8VBhpBuPtkCAjJkRUmlQEkC7QiljWBW6ou/9F4hNbfWTRFAjYp
Jb4YhKOFP/f/TqQSOdOVwH3OQERImqIjD0CRU0MF08R/o9zAvOhyAJLYHRk/sRpV
T/1PVRKZQcEsIJdcdqeJkUWpdXvCTI9by6QsnSwIOpLkGaIE/XfUgqZtK7Sww/vH
9cle55L5MuBffFK1Lf/qQcF/eDohhoSpp7kp4xOv+futR99LfvGTJftkS0z6GhMs
uStG9zWlcgpgpKJgm5IcYpGViIz73HPhRDFUmeWXYV5DO9O/XKev8kAOEqRKq+fD
zPH7fHrUBNuNhNR0924zdBfAzvZY1UL8YzOrK2qvBnXdz/gRbWR8ljDVRzrJFY8B
otX4cnWYTCAZ3dLFMqvKYMv6mA7ZtapyeUjaDzlhFNjwoWmgUd4CrQmADASuilEM
t1W77V5kbQFOCNANwYK39BFdpzhgrIuy5oF/ESzW744kWHe7CbDYy3GlI4DmDntk
UI/U+JoB7fQk/xWEo3owU7SBMG2FxoeTG04dlcoaVJAQh0Z9b7/2MXWd2m6WDR1n
6RsUxC0fHBYhCOGuigHIBt+sG/CPX5503hwzubHz220DdvoSq5gqhyCJvEtU1yJC
Vzi7vzYO5wFDqJ6OIDF7hdv5kTswMhUdwH5KKvxDUFKZ6aK1DE7L2hT7y0W1SDQa
r+nYHvwpVHzteeZ9Zg/uvHiWgYOZMtZP8eaBDFCII+2BQwxK1q8ZmLCs2Zt1kvvb
01I5bNLut4YoAxv2K04TFwvZ4NLCzrWLzO4C6xpR59MlRIump/MdML4/MmQUHdGS
Ycx0eRtrUigtZqJ/tYMACq67rrRzhBzUUGh4cHwy35a3cUnIdTk8K582MxymJSDv
eiuYIqUAdH351qumAzNi4/015xJW7QtI06+cCOif09zmR4m/30kEK0NWPgzaWQZT
ZNG6gdPuem3PERqNh+3ysHCzwHqK53WJDZNYmjGkVUTdUmOkjC5dTKOuAAT5Olrz
mgEEPZHxE+Ka+YZa18xL22cCQfZ6/Vd7j3MaPlOlCjMGy5SMbSO5lpOYaqh9AwT7
QujiYaXP0BthbC+Ph59Qa24SVGYVtnM4wU1X0MRNkksynzKZGjt2uG0u/9QRhr+r
v+V+HWDT3leFy0aOK8H/LgpozOMtEFaYldI/NAFyxZEBHH77mW+vGkNVIR8Mp3Yo
4T4WfsM2udiCjmGd4seuz0U24OOxxJMIUN1excS8bkjSdgG4id9C8hO9rgF71OS1
imTRn8Y7x6hwBOobACLmZJ1eByDipfkOKmgEMd1X71ZwEoG+jbG7JVAwuOmK/jcz
73SW55jltRs3Oj5mJkdEtF9ruAfIK1kkfqmk2/sEoKX3nRu/W9mgpnaAZi+uEwQA
t+Fg/mrp5i2qQcj8nmS9HFfXwniWVMrEUCAFQnri+oD5Uw6+NMDQ4EfWzwbMEfZV
Sn3xjMnrjY/XmPVSrt/2Vr7uc26oyt3eYQMiilyOxIY=
`protect end_protected
