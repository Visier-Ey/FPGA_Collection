-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ggrOnGVMIkm+yQ9kj19IgnOldP14PT/0GEuB23waZO0ynjKysQjq/hHZL9toB7He/rVnwIvg9NqH
Y8NN80T1vfnW131hNBN8bnzuAY6VXvorJBkBXj8DNWoK8MkyLKs4gVX2ql0LS37fnffBToi8JvF5
mEzC/3y4Qm9yk4SRA01v2zuzFeZyBsjsR12/bCBDSXhMx3emTs3MgrfGHuptvRUjm3QPUrraVi32
gN0fQKJB/tFVAGmCviDuKzORNL3qg+tkWUIZwmXGK/swDpvXMnVnYs7G5a+2YvaYTqGRWnGOrv+4
ox/8x7RN1VMckQ2hhRq8TrE+f5cpUWx9C6isjA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 28016)
`protect data_block
1x6geiWstIMy8yO6dLSwjyjqf79se3+coCc6xM06GxCxW3DlvnBm96iRTz0tSAgKoVTeg1mZpbJR
JlAsbj0lgyqwnbEU+DLZWbV/ag6XPFZA9tOTNU499JxB+GyjYthrV8OLdHgsuzpeMF9OEc+eQGJW
jweNY236L2iNZd73dNAefVv/Flo7FQCtNm3jyjUlEJIWM6a1emXb/1wDa3ft2K4AmFiESxBPhYgY
IR8rxFRZ8ohjEsRaw252NbKfurgwKOQXGe+VL7OAHq2UgMZ7U5WY6r7yLwActD6/JOPcimF/XKxz
d3jAUjZtsQPAuH1myZFp2OyUZNntNESqmI1aQ2/9MsoLWcAw+Ggl0+pqK6YWBch06/uugOMt3UsW
8IVZ8HsHmrIsV5waPuNcSCEfbB2AGk8BjLQLgEyaVFVP3g75ldi8oOnYnGVpvv+sDodZ9MnsSR8H
Y0P9eJds8lVyj61dJHaZpxTBg51BxVLL0lLtJAed1f3rHLcqm07oQ9LVtoI1BrZW+l7yAttMIcCO
P8mQ5xLP5SCTgUPtO9YrGJcFR6i8KM+dLTVHiLRDeenFttbFQwiOr4+N9a1UtIP/2YcKbJdjtDzu
aGBLeFAO/p8j3s4HKQ65wlawr1P11kci9EU4KXg0tAFPIMsb6jrN9+pT7+97U4kEXvIdhA3svSEQ
4bMcXqJTzSsH41Jiss5xwoAkgO2+HKaZGjUAYhqQttpJjCwHhjbnP28pwzEtrYRKO3Ni/dgKIQ8j
Yu3gc5N4q8jqCS9lo1H/vfk+t29k0TqAhv1OFdvcUfW0JKA2wgUW/OQ334fMR0GUUG1e/xsyIFau
x2HlYC2qBqWR+c3x7zakH1SzvbzwXWSZ+8gcqz7Oqv+JT0Xt/2XTMSwYHVIj3DaQVWh2oNyn7owK
eY3ZxJfYNuf1BsRWs1W/o1qSoKPCvJEbrsaQAWMlbLuz1jOyyZ32TgSPvatPCkzmG/dHoDi9mKxm
JS+gmakmHQ12dB1oFMJN4CY8g3O+f34laZLg2ZwonpOLA4G56fboR9X3qdqoPQAPsIDMqvuUbYcx
UMHq8D1XgeDPuZdwke0g9/o9iD3X/FRXFpwlFzDM3XJRpGtZpE0kGwcqbW7r9Jd7oBi4Wv4cnWu1
OxMn5JkcTuLHGC6Xs3mPtLaJcH8yDQFG4lG0/+oq+GU6phtfwOHc5/gO5GnQc97hWQJOOvlJcwSZ
KVBfBaAJ+ZfC/ug8H/lK1IOEOEN0aeVR+Xz7q7lmczsksbGfBRWNVSHEdLHZhbDvE+HdEAnjsvQP
c1n3ZR90gQOyIkDLZorYCgLrOk3R8c1TVontOoE0qcvopjeI6EXUD+6OwmyRDIqKnrYY3zXbdPiK
VbliUlfTtXSIklmacUdx/wNL2CZxl2yRoJe2glFXvBxDoxdMgManhxxhsVzBv+H4Mi+8rfZW8kjI
XpyPjmqQobZ/up/uhuN3t6tk59AZPc9OBFkpguqIikwXpQKXcXgnwluuI4BgF/a0QZ87MEzUuU1x
J6Jml4mEurLh34eESTQ9c8sF3jj2hzAhAHECP7sVCct/1qx6dQGKSWcP51tb9DTEOuB2SCiZ0Gnd
rDSVcVa3SnwafoGsR1dUIiMEy+qzC0MtO/2xjVs91LgeirdZGVt0ZcSV7MiwmZlfH32G3CR6uwQG
p3dxn8tUwZ/ZixuV+o0A8MQbiEBAdIIaDNoDXHFdzYzg+nansaUJnrq3iHhrxs2qM9h11aj3gtBq
TgQ0zjsEI3IY7k5vURcMYvZ0wMNK4h7KHuAuqHBDjCl4pX6rFgkkG2MInO0OgKiul9NhbN11TytN
R8hTUPBvwDJS715HGc6YpNlDvpFXcDW7Ec1tdr7nCfUhxEWbGgqKHYkPNUdLkkuygDc3OnlH9Rki
Kyy33k3MZbAmymuD1NK59NAqM6VgIwDjhdKxRxP/nwVhXF59UBxUxVzhCn8aly2e3nnREkMNLwP7
qCjuQ+M3XCzgMjgrXHiN4whHW3oVEzKiTAM5it8sGWbDOIKBrVK5WATZo9M8mc5IooGTjlu6VS+w
ND6bANPV6+NJDYoFIZl6y2d6ZidbXpzB16p8aGvmBXZaukc1qeV9U0i7CAe7RunaNxDfWTKo8//A
UYw/tbv5S2+Uv4srbjaMC8t9xJNQDY9sddvKYaXRfjN/f+IEriITaPrZUXSfsxSxkKMl6Rut09sK
V575rUBNn2XVG6TbPCZEFH1Y5eclwnerx/v9BPJD8C4UrVXaFCfNw5e+XZkpWaGHzjlEKzxUfleA
kG2r0+cnXjoIsPeBAdrIyE9D1gDprFWkCUE0H/UZ3ZOEgcLpHagUkDHGyoIh2mc7uBfwKQ3fhYno
gL0UMKafKzqGRGeHwLstWDQhjWHYV72HA7r3GQMyigu+fRfrr7qWPFMdClpjD6eMuu3ZlUxEqCWi
OJ6wMnmuiF3x/KVNETSaeusMMzqjlpEUxPBaHdriqLtXsgsF7ATTxExyZwMvPTxDnW2+72/JDy/V
xkfAYShyLMQ4fe5D1rxlESjAdMh+ap8j+VkQ4wv1cpV2CW0U3OvoI8taCm9Fd1un3ydOi5uj1h+i
bJKMFD7fiTK4YjuhZPjcFKrJc5gSZ90Pww5EsK5ZxlwlXSfbVsai4Yj6qYPFRcPlsjsVL0uHs+Mn
6fxlnV8SvlQ8ZhbzZVwoKLTo3qqTA/nERwQjzcaTg5kt4aOOZQJ1CLBRBAZjFf+dEsgr0jnE0GqD
MqCyK7m1GbNekkoF4bh5SU+6jKCvWpgRMKXThMMsAketxCwhWx5RWIuTzyBPlR7LrOLtRWlaJanv
dcSsPgZ8TNt0TxjQze+jRX6E3C7hh1CGrxRtZOMaVgfpYtM4EHwZe3OENP53Afkyl9InsZyX+w93
EVnrpm2ZXeAofJ/TJqGL2TphRztfWGR5w5ZzgY5So9pyddh1JdDQg3P4xJfQ8AvTZr+z3K2ky3Wi
91iQqcYB+n8jkeTIc9WtUz4fp5gJ2ESrK8jhs4B5UFFAP6KqCEOwZUVeToANaU1Z9IHlocu9W/ju
OLp+zCO0M+O1Doln1bMv7/N453OPrIzW3MyTlktOn62CJ8cnD0wvNpHeS/vJ/3IKGbMT9fltzI++
UY5FKb7qcUsSqUvoIObSvgWJQCZIEiZ/aMZALaCv6IXHKBuievKHBtCL2lFsAwFQzUYSe+4xmUGm
21Ekp3KBjeZHi62ckp1dQ/SNxNeRxRtlUXB/neVh/LhLBdt1Xx8+GAEjFWRntclrnctSPDjcwOLr
kQSEwuCmUjpD+/0NUTaDxAMmPrPdog8x/jtjCX4kcYRi/GNnotGIEL5TGRvgXyyTKPkCiVwQLBS+
rMLCQuYIFfskTWzZ1FZ+XLG/g1tYxjx7VQ0uS7KIRnrzoNZlo1bCySYfLxNZ+bNkj5C4lQCWSW/3
liU86W9jcOLVPHIYhd6PcqLSHXRBruyuUKfNb+7yGBF5MWX/WJVNQITtlIyV09Q9fBVPTCf3JqnR
pcu0ecJisepBbML/E69mgM6LYqe2iFv0X27A/onsmTgmhFHXy7Fr7NjDsleAbu6im4CjZxmN8SS9
1CFwpEiJnvazInqiHQ3iORqAbmUlQjg8fioQHltVgrfWac0qisiV/J6ADkRZUCtzwRDzjiZcsNU3
tpfI6XyEM5TDN12IHYlHfRgc+1yw4WDonHBhnqEYGrRW/XqI0dQhrPcp2oiFfFrUyY4B3Qkwa/Km
I92Qm2Ad8JuaFTNsk5vmkjzpAYML8K8boO+XePGZDJ6+oIz0vwWiBSdsSj5zLnVTylz3oERrvQIx
jOGBdPxYFXm+quvx+Lykocf0L2XwBlcl5Bet+NQ6svFbK8+G6Sjo7U980pHfsBO041PhZcKGlVVK
YyYIiwuQPKwpY7D5V7MZUL5nUibpVUqVCzD2XqDMdhi/1O8+RI6eRyHulxtgeJ+RRgS3E3UN4p+F
DwEZpyv0HzWiqtlGKIkyJzkOWxBvkkxstmSaYjbnvMWcg2rUkqbEVBoh+/uHDGTxVzAnIEaeoA4H
cZk1iyX2aJq37gV/HjzY/nO/DCOhsuP6oC2PpCSUFHvItG3Bll6g9fX5fVc911vEaQQmv+/sDRJw
M6gVb9ONSBGxQRpnz8mIp14qnh8+Jm4eZFKHKzu7B/KeRxd0WdbSbfmpIL0sjgBm9vrfvG3psQ34
tc1MQ6hXOn1bc9d6MhTKoi+J9CDcfviUI4NpuwnwKswojqGJplp4eaR1EcxSR/ZoG1Bj4tFuEKHx
LgZr/R5oG1vKhCMkjo1d/1hWINCRdqoG1+FP+hW5SlA1bZdHLv+dl3hiKPzxqaURYnKq73P0MRbc
H039Y/F+QHltTBptCs339d6jM+1PHl/UWS/2hSNGvxfBniAhqenrGL5MZLEfdujKIv++XNGEh3yr
Ui/oBzFYgi44LqGub9b8KA2XvZAGFU41R9p0jkhwyv5VH5bbPNU0OG+bQJoWt6rxMibVJmPU3CZH
LGPFrmTIzMQ1gGqmqOr8+p4IpgdTH68tznf8KLiGIfNwnvm4Q/lf9X/7Q3hhWJe76QKJnz6q70Uw
4osSK01gqLgqenpINySSQD78PeZptq/RVBWSR+4nVJFG6cA+rkzOAjkqQYqX5Z2mUE7wxq/nj1OZ
3gJZb4zAnTfjrOAVhBng7PyttqqtPa1MycXxqiWE9OGeercxO0pvboEuLhEXbEeu3U442kd1M/+X
T+q2zv3WWPr9YtO3yVyXqloWQ5jSaQOr9DDQpbXj9c6VL6AAHu7PzmQhp0I7cHKQQFzCk2q1nfBF
cM7dWVY0vOOi1RMBy895D7ko/FvH5rLMOG9ABR4M8FO5epdMgCvG7LyZueenieG33tgYJKL+F09K
S4BbXjCiHvkvedh5NJqrEmaUAZEm1q3J0wYEolfzZ1U7D4hyzD53ravXHTtX+tbGCjvb4xidUm8T
kInNwfmMi2G+5abVD4+CLbVU4geHHwZ9VBSSYGkpkK7ravhGDnxROqC4E/Ay1CDlahj5olBHHJs+
4+6i3N/J+XFeVdu62z8bZl+h7ueBPXevl8ldUH3yXr61SlJzKwEkdvS3QRas/oWqEbtXRjtj1ORF
mdQ4zX2zD5BRxZpG0Ul3TB9wieCE8UXrMdBzLkCeKoP7PBcXot9Oo1MZS+9F1c9yxqIYaheaOIb3
rJ5eAQXLXB/RZwNg/q5D4+RFeYYNK/lZkgJhtMPpowdGKDPPKo4xvSDuaGA8nLGbAvrgJUFh4n1K
b28u8aXmPh4A77HCzggre1kstoDT7ec8kGPNAUSfQIJnF3vWoYRajWv/69lxEi1FUFm+YdZUA6JA
oNvDzyGTOavW8gyLBbnsCZD5dTgyDm1c0Gaf7KKIxsHVJZ3xu8hmfqOyTmFfKgSgyslIWenYuv+5
Y2CArngDBslgJECMb5whyPYb7MJdr+MQVdqw+IQmALt05fN83Hlv1lFj7xAZyfMdYXHOBf658xUn
8s9oQKUWms7w7ejU+HyG7nN0I47griIGEKFmyJr01wSv68OyDxqj7rLBUYQ6vNt3AwQDYmlPOEO+
lEEGqof2C+9l9xPQVpYGHoTS8XPiuPR3JPAhz85mNI6/ZjaAqzLnMek9ckHOmEVG3rKSK/YNlae4
tRupyi2OZ81qBkDPOXS2CBsH8FNvU+IS5cPqbjPak26eJONZ7B8t8gli8u/Mbdze2YXJ6NOkrwmK
RVj9BiJ+Xmsi1is4ENtHBfrh2AhxQzM/Z5zVIfvRXYEknw4OlBslho9bYOWDZbpRQtWGhc0CD/OS
1W9YpBgTJnTlqq/fW5CagMpymbFJ1UHZI+smTJHuUayKCZvlfDGBUR7c9F96H9w/zgHUq9NzpGg5
CpXrs8tYQx5Bkku7K0+PrgzFW4MmKKqsCHSJKVlDRjZHwoeKCeSiqoAWvbmpSp6Mp57Q2KUKQZ35
al4M59LL9AehgSJsAGqYcF240q8nh85nwazX8+DTWWqwQxRHxdDbJvOxYLPGHRzO7reOy8aDoHx4
BZ4bt6q2BLLLJ19fX8zRq2BemRdK7mFVxTiYFMj8jwtPmFSQM8Mwh2+l42FzYRIu9ML9qG2ey3KH
OOTVZb3wT824zh5O8K6YiRkS6GxqTgMlOhfimJ47wvlObPFq3yWpdgv3N0naQAm6aLnKNSdrb8QU
qztC6ycKzDgtCC+bYA130OzMeeXvZ2GYBuXZ4oLgeq1VzK1ZNIjDvaAT5NWwYJli8ZS/q1xsCVo6
x3SHuIC6lWPKlqWGpfqcTHCaQHtvkBp9H+PiG7JwDCDOMECK6LYBIoyDMKwukisvcCV8EYL3loLs
asdEtwtVAKfY9H2FFeSV9VpbRbNh/sasDYtfSaRt0g/ij0jPjHAByHbtvPH0d470V84JYQdgRcTK
QiE2K8n1K0bVh6jepd6vHf5B08nZAVNiBS+fal5vE2241Kp91h0lcj7BwpHqF8cu12NZ2G/uhfwR
gMSytfAs/F/sUeTBpHfsrvPimVKim6EvvTKYVK61o/TSJhd9FyAtb2nmEsYSh8qxgaVlajnzxX0M
f3IZFbPwc4CTayO5obVi2YkFJMhiL35D4/XVe5XAPnChe56+F77Z8t+VZs2TVqMzf3PTwRPy3ZXH
Jo3BwESK/Yxdz2VuSMXh8yNZEe73JQTqy2vHzSWnktMIgqAuVOgPX8kjVOVf6M8VXMH6epo152UT
mwwzg4kcLh0osNYb3WR6jK+IG0a3W6nCO0JRpKKwtR4vXeSLRa+3DxzMQlGQ0uj+F0GwiStduRE/
4l6eyvakeCtr7pWPS1xlQaZeke2QzABGlRgP29JG4rdjxTBfAUEcJJ2slFY6bxR0r0JhLvKGg1tX
Ct0reijABfGKbcd7dO2iZQB/PyU8L4oL9wGlet/2wrfe1o8cCqg1SFSo7QcP7rp90WGUwfdgcT4m
DjFzRBO0QWTMPLS9dy9X5dJGVZB0h1GxCt+iEmKdQtX6k8kpEZtk/uJP6/Gkz4Gmdv5eTwbnia+u
I0v9cF+2qnKI/rnBF5jW82jqyOoa3yWw6JWTVYW1GbX3x6fV/hCn1fWcgawjjhHKChsi1hC7z2Dy
+v3DVPTfccZJvNNDbsLrDWZEP+GcRyIrpqbLdTDjaTBFhuTfu4cpnULCuUmMPbQTy9X5uKR//l8w
addAQ7YsdmY4fciKH1ut40GdKDwr1FaxGhrHRnc1Z922av0ntGRJHAun9E/d9dT0AE6TU4zNR7Es
Xl5HnP95UTtgxd0SxSncn6uLOl4pXCcyyA/At2jAZuwUHzrcYfuE+/jSLyvKsagABt8bD+LgX8Zk
JUhQ4x5l3Af+ezYaIreczvwktNKmjPNfacNaC9q3760pkRNhNKMr9uVJToS07sD+IgfkXdpKgwfd
orsZdB0V4Z0KeR8+6pezMX9Q9DRfM3HR+ryxTByZ/7ZGrP2Q8PrjwKpgOqrvjIDqInF9Aq9TWILB
JCH1wMdR7t6/R+G+jJVk+KuiGb/gYq3VKLxaYdVU+swCFKDGnX9oQTzuYRH692+4fiXXMDrUv8Ib
lySExi0BKiR+4Edao4sOU7fY3oVSwTtDp+VJUv/6bXUXSLrXBWKiS9GxNA8v+o1cR7zmNNdrxbBN
bUD1meQdy4pohNyebVnVLqhPp6NJ8Ktlgiedw+8Dh4GzmBW7aIWp0bTHlSjpWd/+rpDRu7ybDM1Z
iJWYyYMmhmeJxewCzHUMTZGEc6rTmcMT2CRXV51ObRRg3TTcGD70Pt5WxNDixrvSAh4QNKvJIlub
s6euE/coJ0ukLlai5WRAmpn/1x3mNNi+mWvzJhiFUorXS817DP5U6oRCiUy5j5XVXbRxD3Q0wRLm
WN3aLt9k7KQxNr/JwZa8y00T1PI24bLKDjrThKX2J4YuqDQ3LKvWZJ+0mbz4N4chAGfhjeXjcPmG
UqXxB1m/IkVqZmM9JvtAFea4qMOZTU5e8UDdJN7XBIAvo6lxRoMIxZoOLnpwcR9VcnuH8V7Li1h3
fGUdACnbvs/2ratnta5MIZJQl7dzVHv6RR3D9oOmUG5wOE03lAt9vmR461O8oCAUAYVQrNX/ruNT
ERQplKR1PwqQRih5ldEqZmw9M5Qda95WZgO8LdxLZ0hUx/NQV7FCpclPD6kshkt9/AIY0OdiAKkK
n0OjjZb5HqeBUa72TKbxR77nDQe81vs8i9ju3u1Qnlvpk5tr9v8YPGut7BE9qIAZs0pac7C5iy6Q
bTf2qPwwDqgEOlLr2LAFCPXbjtV5eSZA9KAFMh6Ar8LmCTu4kNn1NFcx8OFWSZ4dTW5hs68H8MdY
qNVNQxU0vwFtIrnmO1U1kvZas8Ut6qHm8M1GB0W7h/aofzc2CXXSO3Y475U1xxpBhGv9Wdo+cmvd
N96nJAUTrgx9m8x/FETiRc1NbJfwKvEeZqD1rqu/TrkAcD4pel6h7Q8eMIad+kURnNAmum7lMcGH
B/F1VR4v7mCQsX8+6Wkau4r6QSkJiiiikw1JhMQizQUloYcc8OUMX8cq0AEhx5mp1eTwD5iLKXEW
NiFIkPQwQiu6XIEh9F0C55/V0KewUXUS69OFtsF2VX1GPY9yj+p2VnJ2r1zn5JlYf8s22bw8PjiB
fG3VCaTnLMUtcOTFUTE48AoDK75atdSyUvhU916kNe5jMxrhb1rGkW+WxpRp7641l1P6RPBhHq6X
XZP0JOMOBrFrUHtTnZ4p+O/qgFzeskhhxW2rerSki9HeERChdtxtmz/+0qdR9cBr9nhEF50pRyKJ
Wndlc4fbvANirwUo7cC8yRjf6DiTFXUlGbo0NarmhLcxVU3PJdeHES/+JbMY+9GErUAjDBn1IvQI
7Ji8bnC55Cx5TCMZgbR6ymUuepqXvA/Lj9+LEj03gh3XRGDKDQcU1Lzk2xzM8fQCAjd157hFRf7r
M+4ndkDpDuRk1MQ9vrEFEcfAiR9SwMAGiBpGfgVBpjxUUUUlWs3vB3cZrl4bV+rRM7rc1I3YSquB
ltjEmSTj+cZeCabbcVBh0LRTDbA3fK/saMAyGvpMhJIfNhGbuX4zDOacewR4oyi+gVsLCpzZD3Ad
qitm72Qd9MKFi4kxq5gk+VNVu961uAfvSIs2XCs0EohkcEmWaF/nLxMvlCqpUHfoh1kN7zu0m0bj
o8q3k78dZALC/0C/MrZ5Fy57zGUW4KYHNLdmsbK/8ef1pBwdcR+fnagF35TICQxb0WXg8uO9QMZP
1aS3Bjtel2K+I8OG32wqVSyz7fqtrRmQDCwn06V3KC468u5O6ndH3MebSrNAoWGpLIE1+piu2UFV
VOfhvB2PMxl7pKFxgGV9JDGS5SLfirOoaBTTRt6a2RAVio54v8D8HAifwQJTu0CwqD9l+uIu79oQ
ZEVp0ZCbx/yp8Q0NJGRF5x0k3c8Xz0JolZR0QXQVNglDK+g3DdgCvZevFrNbQDLtutBhUK2XvY/8
CF9PbHtvGU3zQBtOctMaYKUgmLpkW0Rpz/EV9u8c6yyd/P0DWr3fDYaxXSt+kQoZSfzyjYFYumDz
4x/tKs/dJ6aSEUDQ3uWG5F7qbj9aMUnpL33fW/k7YrYQSSGz/b4mT9x0VtbEg4OQazSwS+QmAotx
RkfGBx0OnXRQs+xf+7AJqiL2PYIQd3VqxYb5992xjeRUnp8UqflUiAWPnfXUMa0lHs0+WwapV9rq
sJU/cgWmqfRHyHtO8QGBE5YPcpA/bHAgBsZ46S+vyK3HxcdMP4T59wP74qzoE27b+tZo4Bw/5k09
B5CbUFxo3a7K0g7dzvuJQw/UCATmnp+pLTGncf7+tUx1Eh+lsmJ0Vw2c+O+4plpZ9JesKO3yQJGv
yHdcllUgga5zTE66sF6AQ9bQxGoHUScZWKk0AECHz2AxY7u2zFnuL0qRyieRFfC0hE5Yels70bz3
iggyBHxys4JIq9DaKA8ZDJPiQMUmgMXcMOaS8+8VIR6WLwaPlsqY0OV076jSMTDdm7iICbvImH3l
Cwh3Zv3uzeGZbPOIuCBY7D8Imj3UWqQoqxLr5VMLv1wen43XQ6VrZWf4ghwV9fdQYdHXk/W0GcYh
SJGRHY/iuvUI3I9FCftp+ozi8pCkeKLWcS9/WImOwfB0rF9qwHGx/uMikTM7V2Q3lrMNTXYKLwqk
SkHS3gWVmPWh3gL2ffIMELta15ezPUP6NeSbW4m/GX7+dkBxG90MWjgMLUI9bV2HcubFpDQwkV8d
A4tgBYhJqpvtGyco2Chj2x4EjoJ+vQ86PJKFCOHaPKeporYZNdPRsRJzebLdE0esQqh7dbbpr2R9
JZX35mzCqtTRf5YoK3Z5vksut4r25PEmj8L8WBNBLV9oM0wly9yNv55EgDQ/1SRYdOE3Rd8FR9IR
SOTTpNeSeNuNWcbjRWsefVggzVCiTFd61DHZMKkoQ49oifAm8TbIRFwtEbKhz1DetVxtL+dCovLv
EZl0P9pputBSNlAZHiCPeXisKxeoD2hLODxQrCcv9j5Fkq6d+TZPcbAX3nvilQ7VnO2Kxuj9MWPe
TfZpO0eoa1uNbJ2CnmhzdBI11i8jSjGcnfwcb8lEzuROBOdCPsTO0yNo+QdXdt/lAFjA/0cksCDx
Lx8MIW7UE+dzyzViC3ePX51Vh+YQHCOqrXmRpGOUg8SPjP/agBnPfGRKEidzusr295O5wE7Aox37
09coilaF9ZQ9DgixLRgihxODM+exM8vX4peZoJeHUJr83wsDm6HYh9jpNvxZXqUf+6pUg6PHjEZ5
xBUFi9/sN/ixfJZykdooSI3YIqlUPoOueVdCZHTcQHlAfWmLBP6MN1O2s1sOzVDY6LdbAdaPTOAO
DE2xx62xRJtH/FhO5QzNnUGPgWnEXQW5cVeCEM2A5FhgG80WMc5ZE8nRB26q8LSReQWuyKwpsfN9
VGO/XsMDcUsu4G4n715SAutXndXBAbiHBp80PJcNYLu8pnPQjxfKRj5LWzsRT6psNj7dLt1jQJYB
pawYDgtLDgNCxX4seBI3j63Q+xgUePofnQ2Wi/0U9NZWCR5R2zSNPoXXWX65rfXFaDl3iOk1KzBp
/JGNvaA9FyovubtctpSWDPoWNiKZE9J1r0j3FjGFPoY3xGact7eN6r4GqQJZBMH7GnFr/DG+WyPy
Ae5/vAu1b5QNH3Ge2jbxuJznE9F+3Zppn+u6ZrzteXQbSmRZyKVUBeRwX9Ti/cIsVmkVxHybouso
c8UldZ8JGGYhFDSSfMeDDBOLz7WKkZzq8XdMc/VMSFlIftiaRfrweDBXtUCrsl58J3ThVQ7YjVR6
JtzfRzEH8kD9/1QJDxsI4VN+kQm0OHlTxhUDp1naAeLyJR9Cvek+bg9MNccg/qY7SLjCvsNqjvMz
2j2znJ91XD+DU/dCxG0x0Td2SgZ/98rAjYCukQ8Hh66UtCA3xQcZhr6rSxlmavAgX5+8Qgtvh+Z+
ScXLeYHxRZmeqM6EUXEeS5bRgDjjPjAn0SQ2O6rWo0mFcyKdsOq9AQ2JkSrXZr3cxMaALw7GDOg0
W8FtVcJuBY/lMhR96JmrK1FmOhfuWVqHftEZ+88G0UY2SM4hu0Rg9htaJmvDaUJhhxJkQriAA4s3
OXPSpGcnxs7hw+wNGwCEJZajubBlHzEOGzxs1CpAEVov2vZzNBpawhpBCjDvkg5uLq7dIA/fbftj
7gKakyxs1WhOGz0qN8NAcxPggY6oJo7AsEEGJUW/Asy0Zym1ChWdUtgvoGMqEEfSAocxb2jvfnSp
0IHWWJVzpZ5++kw10+I7RkkQfiZMMqd8TN5Y2T0zgapaa7gePfDT5P6lCd08zwNZJgvxrYSRtTOx
HHGBpyYv5QKqslaZfxz6wtZQSLEzw3ioR5O6S48cBPpe9HGrRh7At9Qs3bG//EAq/srG4W595wD5
ba+PD4ll2ycuT+Sw+ykVS/AzmV9wuYIMHryzFTFgdFEmuO82zw+WfLcDpGighntoR7fWyHgLZsgy
Z/QlRNDJEmzc7zWMsUXqDV68RyL9WtCX7irIFrlpNyESbmXDhcJIFGPDGrus4ngeSUlunHI35lsC
l54ALEATIglN2INLYjDtakKGf2CBGRDfdelAawP567Gdi+lwyfog01gGx+IDG0CismfNyM3Cb82+
7ecemGL3NJNE1UYzt9fG5Z01be5UxgoMOqanyfggF6JOCFiflQ37e62eGd0BYew35AC4WHgO1A8p
mCRF0v5TO9EyFeT8GTwjmmOu9/96JTOwj2LLU1+r3mJ4h6cuc4WkMBaiJAg4Vwzw4CbQ6HQBthh2
KzWIOyG2WQlYhbPaCeaMJJCKPmrt2qAOM/v6wC9YvIV+2l1k4q8B5T/Uv7eczx9z4+mBF7Sj1kDd
DIi2D16KBeugKxC8JLp9J/qaGsAXLrXDm04FcYWO6zgRj5v9shV+BWkkhfTHAIqcCUaO/Nnzmoz8
2zPCQBpoQhMxJE2FYxOXlDLjtEvaLCYJFPauiux8TCHNJsybvCsCFTYIIkIWgPG1H9HqIFbuNUUH
w9fE7YoLknz5zprQ31rGTkzW2tylC9vkgscAF9UKa79OKu3tNGnF08sY7CIQsTgfanVgrkQ0BHx9
jI1TtO/A4OIMyyfLI3h4vYF8imZewWmfQokcDgfqh0aO4CQZkzMndZsJSoabUwLDflF67XFZUsxw
JBSCK2O6dY1UPo2p8HS2u73mkm8X4rePiA4LeFfsVUq21N5td1Kmu0E03/R3oPvl6LmooWFR5hat
jU10xk7+igZ3V1pEs/LZduJY1R9aSIH3c3pYP3mUthCloSpVRZ4A2LddOKGAZb9g9f0L/0BJVJV2
qQUYRSjQkeRhdqWliUBMo5iOO/1cDVEbD6SvCT+KxdfQZtXLVOuPR2Lrn15mLbHfvRRBaHTajDjZ
CG8wDu52mUGhQ+0sZYu6kq3SNvpzTuiFVcig0NAYp5JW2Mmxo4JtxbyGVZwUTwJ+T79yji+IwIcm
GdsjLrAEmyp2PtufwZPyQJlqhbCF9n0v1A/6w1LWl1MDWxpMqgxV+5HiP4WmB+dCclprgYyJeWBX
/+w2xKlnIcrUEymFBr1010dqKI0XN08TzK4xblgfoLs0oxn0OSscWl8DMhU6jEvj96J4uWelLRio
LKRYpC4Wj6+jrrv1GKWi29cwgoMIqRAlpVVnd/uEUnl30fU+HdENF/I4vMMfWQqDweSqf1wHtZG/
Jz7612NBxpCDS6DV6bnXHdEXSU7PF33Ze9+eBbung54AEAU9Src5wwJaHsmtnaoPOqSoZbSW0sGP
gnBnyZHsKXwjWRg9FCVBsSxIq5kFbEQKQjLrKb+wZB6JVnjtyS98gqB1Yr0ZoLHaXDsMThOqW59x
JbJx3GY8xBIEdCV5JNmHuOGypnNA6OB4gU5z+wNzqn4srIxiqC6opYkcCTMVZvbffyj/ELzMnDCB
buE5RXS4dC11IlWb0vWTaiTtadeSVjt5kjxIVdf9CTmcx+cLwfUOBV2KdhMoDVd/8X6lRJ1qy9pn
X6XRU2f2hPRxI2unxTrTbdgqXj/s2C938K2skN9PNjvTHjiCgb1UIkwW1Q0vUhNw57q6Zca1hSU7
ZpzpBPk5d4jmcnMtUj1qcpvaMGMFfAkNQQgr2gOROPs9phSVa8re5rOQSMiftll5y+YunYJumjxt
MxWxu5COzOJ6B5mtV997xCwvjcsBpxK02CW/LVlRM9xHxRqcpWH60xLtf7BTo6N9N15GPYFBBkIV
0oZGs/twL+yJIhGqE0Whepiv2tFYoc2MJjnrJg7IjGQGMTIgnOMXyevS3Q4usLgWozS1mTv4xC2w
I4ZxGf+AUyf4lVCa5HSHcFekoz1wTyx3ILxstMzqfM29eZ4uu7sd3I7mjjbXt/6vyb4dPNG9qpn2
of+S8rqjZkweOSTLrW3MAKHf2h92m5fL1C2aaNoVfuCxSmgfw0NxgkNZ+81UDM4XweuyoyhZNX8l
WXkjCQjLFAneQqNRPJipVsv+6pNrI8ZqYtvrNaBLqUjX2zqBB80Ly5oGu/VEiZ50zO6vrb0r/5Pn
PCjd6EA2V4AVpvsD2ipLX9Gutb9Vp9/iz7yLb4X6rE3sudFXNw7onwOnaqmVElJgy6F7GKzWbC6s
JS9cvhRgmcC1cvAtLLwUGnunuodEIBQlc141qQhNqHPkNYLZqXMwT0/u7QKcbqcxGS3+3d1NV4gZ
I96bZGIUeG8GVGH0eIyhCOEC9Fn2vhx9spgq/e7MktEvLzctUg5uz5ffNfTaJ+jJzj9R1+Qid+N4
16H2iloi73/onk83YnZdsoHlnTAKOS2wQQOysTgByzYuYX2gNenu8SP6ih00idmPmIYS1ZHW2dcG
r84A7qfRDkheTYLnxeRoukdrLcmzsNVmjtz3aFXhH9CdMHi+TZMQz8gnP75MYmSeGWtsiPG9aoWB
4wjWcjUk+MiSE/Fj3VgdHfDY64z/NSeuaBNRdx7qa7PdK3265twl2tb0eNY2iuuiFwWjRCyUVjoi
velb2itME8mbt7i0+fMDUrgiucQIp2gRKPl22WzysETWIGLcc6ICJWtr6Uk2BFRNFuOOsYoMb1xH
kU/aU2shkBbihgQSo3wOD1DLi8jzTn2t3VYAr/apTAUYODhYEv+3xXPMWyAS6xRNJgVpWKZY0u7X
nB3TqyIT6//7Ca/w4e5tzgjg1VF8NNBezewPESnFwq2TNEnzjkUaNYpPKfpbzJvhIcgP+DlHVvPu
DijVeb+cNqGF1Ysmam2tnu2I1153bOtYGgzwKN5ZNE7ymbs4tAErazn1pa+4Lbu/Yj7kESnTEj9u
9SsJGF8GaN5ZNAmxJWLnez7n/R0gCYU8kA/oe3fUudiUQJ1AGHKUNWevoAPBd8y7pFqXHqVqWD8Y
ZAIOoaCXKdRxXAaxMffaJgmPTbl/S+axCUcxo0y2hx+IiPzsY83LQK44AnnJ4Xv2HW/NicLp8vNJ
9H2RF60NNYKqDp4osy4Ds9qtH2ZZErSXAIWY+eY9kWxlelWKugRJmNmeMUlbvXmwF42n3VvDcS5Y
UHa9UwQn359UzzSzhBgP6AqkSBS1R8+M9C08ivRdMnFi+LzHZxQnM1/laIZqZz4CU3QcVYcS3B0e
r0/3mF6l9s/YfQC/VeLd2/hDjW0dwaFGDnCHYYhkWBR8RQBnxItRpXhrgCywDyRQwjyLS5rAB3ga
27OXo8rpmV6j/jbZCrzBYcq4RXBi9SCOeXo5nmQmuaGMJzgmw6w5y2NvPXnsq7LiOHxnkus0JN+l
lxcVo3VCsTwlSRj73YjPJosWGNg9I55zDxV0mYCku15UEv/SHzXVJ0DK1KXyLScNW8fdIDn63et6
IcuUA3gaxwRNmntB9LHTZ8V/Kkhh7Wkbed4QSsXDY3DsHweUioXrfL1c2AKRt3gtUad6vEI4UTf2
A0+GgrnWc4b9UGIUch2Zppu5tuGckYuw+hFunZeooLwmzr8iCesRGFcrzPr5S0JEuhNxvomCNYLf
nD15i1fEcCcESd9uAe9e2thnIM2i7T2S5MZLAn0Ugu1UL/sdo//sZGwp5l4uolQ1+LIuoyThbUaD
mhVNUENDM4kOscpE9bu3rYS3zkDzIB2ul5vbWPQHH8iDutuBa7EkO19HhkyqTtgeCgXZGxW87uPB
249uGDM6hQNmM4B2Dj5Q8tBq5pM6aZK7QZ5nEbhBVxFhrBE2UOjleu+8TV3ieKnaKc/L2SVyG5Nf
03gBCQjoonO+uWp5EWZEmO8t+9jWj3g/9tdwk6Oey08rXuv/vIf8+fyWCCe47bi82PvhZfxsLW8J
yC8/p+ppwM9BoAvcanaRtAg2Yer4hEvBSGL16TKo9rc47bYIOFpgWafW0y5/mH6jRQX3Yw5/QHpD
WK3rCPZu22i+2NN1XwPXCoVpvItv/uusEAs8hs6nos/FuMMTpokbJFhptc36JaTn2IiOH4hYUnPo
AESbJItrylV+7PCPq3PGoIq+MHPvV5/rYWfWyZBIRzn14OTf3+v/I7WaqfzhWn8TeQu4BQfck0ar
EueIH8yTJFfjmdpVQny1zjFEl8mKN8TNtNLx/ehK1QgwM4Glt7NOjVKCDk9P5EJuV7VhR3Yey/9A
a0VaIRrG31wM9i/hmImsmUmnkHoJyrjnrlnp4IFA2Sya+yR40z8L1rNgZHrRQuKq6agyPcBAjZNa
+iXTJ9rk1PeWN7sFMPq2ryDfwNlUAtGP26qYj+rXyRc6KzemCggQGKsYhjSAnw8mj2QwLXme7tq4
mOq1cUIUEbS6VO2s09IWZQSKhDXhzJyHSRHESKpy9RaHOtfHtEaDMotmk8bQGi7K7kZTLoFtmSN6
ABVttI0uONJMGFvuO1kNSyZcjFjIyahqZnoXLTee/VLiCyZkKx3f/LO2aEprsYLH74h5P4dfnUrD
cRDNt5OQj5C3ZKCBDQngbDzyKsqzbPHzE6IDewvFmuEMwQXq1/J5beRqGYSwK8sITcYyBwx4+8yT
gcfPOvmZD+dTKuIpQQkga8SCQgwzbrSY3LOBZNsf+/IYkirZuTa4EmN6xNcq1W0/NVtdlMsl+WVZ
xqB8M20L7IfcIUjR46pQI06jojyiVEY6GNncIWi2v9HBJDe5yvarZvftKJcJA4d0Jr0miBhzDXRG
7D0GU+Pi//bfXTbuSFJrCGpxtofct6uB8c00oFvAISlhjrkta3Fcn3i6h/IbJWGxjtSDMgbrgxH0
oYFmiO8LQ9xwACuF8C8vVDWOuEbm6gc6u4DmmsXDuTzrqYEUtJ+bKAieWYMPkmvHYdcpIz1pHzJv
Li+jne2sgAhKKOflcje97tk1smosms7rsJmOyDnFN6i62mBgAf84xqcqOLjnyec1YbjbOp8eZkmu
BlYXxEslq6Fz3eKrqZK4FfwWrk1NsouRqGY325rz9pO4Sw4CDmhd8sTMo2skqsj3pUzBq0gsykU0
9mtWt5dK6LHNtYILAu/BYoC3IZx68i1mw/sp4B3KD+OO5CLs35D3irMI6NP+lYsBAHMzl5BYYoob
UoCg74Z33UQCbEUaEt+iiHhkN+GT0jkvtr6c+6k9b1cZXWZFLK4YWBMMbRuqZOLHJ36YsHepRx/Z
z8mL9RDNWWf/uwCmV1gGjWKjmpoGFxOAtR9zAkGPyFwhD5yE2YOglO+KDInmUt0eat/duPzNQ4k2
LGJip9Dovp0wtAIP8jxQ7hNJpYWOEk88KE8m7OELGw5k3n0RqNHoTohbDPuWh4FLHSAqcAa6qPSA
Jn4qLkC5mSz5lM/vCc0TmZ+JloU+Q8eJ84AzuMrHzWiRBKgTm9NPfJGNkAY1V2+rVV+Zt4skTI05
E//1xW3ZMHQ7JTVIgSTjEOy+8uTbNEA/0mXSEimvEjRByzF/Xw0QpLZGtls2BZ3TXIqhDsTWv0t2
YpcTHhddjso6xLTGrCw8WEqFRlmQ/E8HW+Hy95sPNbMYTY6Wq1uI6o1CGHYJB+2UOp4nku4vnQ4A
pABLOXqzOkIffKTRhJQbi6ZtTvI6EhvLEm8eNGmodvvWoXugyPq+b127GygMK4HD+gZZwP6CoHPS
6sYlfjkFYKA12d06sYlckK8zvBHJA4shUbOg+y5TnMG0p5SxkApT6dRc37ft/Cfnzxo85i0D+Yik
pvyRrWvluinR7Yby8eeJIr7oYOSkRsRTF7BK9gxIBJGekI9RWwZMSWeQoAiOTyXj0hH8Vz9JR3RS
UaL6nVqeyDr9zJn4JbR+J7Oah7CROd2Yv+EgUwNELbxT2vhNTknvEUCSN8Be6gG3k2ryWXHRRJvf
2m62cOtvmsM0PV/2Daj3jvO9c7COwIm77ktGmWpVBwtfhoe1NPdTMkSL67ou3kyrYqLpSc82/hE4
+pitU6TZp9xEujjwq4AvR9vJofyC25di21+5kp1oZgDZcw3ArFj1C0Ovnls3NbLlvggFRJFKlOVV
CztEP62yKTZT29xRUwCR1n76qOr+++lj1pedLFgERWN5wt0Qwhm0K/Gzvzpy1rXxFnq1pWYLOPjc
8pYhOeVZblHfmAzWCsfPeqhU/xM+u/iKhSRf/CA3tVex18tcWB5iLVY/7ERjEtQbAC00pgv5c3Io
ygEJokG8hYLn37mtE9uPFh3DbSxSnla6wXWwPGlar0qNmyhQpoWFFDRMBXTUAvGiEYzXnC575W4K
XlXyNodvwJ7XmRqzVeUpVsftIfVTyMI08o4i9AHdI0ERt2ziC2W/DoDmy0Lq/tkUzfgvtx68xbfR
ZV4Yux0pEY60gfF4G7EIYe/PQ7XANcE+EizjPdYQWv1fKx82UCaFLUK+VpDeaa4a+SIspc9xifPh
/9q63qm2HRMdw44QldecHDOjp1Ud4JxIkD3GmomkGIYKWlebFzABrRX/25m9qq7U5CMFWeuFAnn2
LuVdidQLlq340iQR4U+3QPtZ7IgFygSWsvzZwSC7HZYQUiNNfCBA6IwPOjVde4w0TUiN4jBh9jTh
eiP4JCHPPMujn5qpz1LATJ7ETODueo9eIIJ97BQtiBu6KlfqxEIq1wz3ikQEL1v8MDaSQbRy5ZUG
bJH2/k8gk5jZ4kid3ZQyCr33aZd71dDozVI8nO0XtkEIm+eYjBDQW4jG5SHK77yqzEy4AzqWzGAP
v3inZ92ZH819PO+VPfAr01JwkzNsA6Yw+7OmnbVVgaKcRnMRX1UKCLzvQJEERcmmwMzOCILE7NOy
6GCawxLId92ag4YP9qctSWdvTg1BETpzqHiChVWZgTTe2X74BIqQizklMEyo84rOpd1Jq7+vvVJr
h7V5aOm82bTo3FVjqwDZNhSgm+eUXWVQAiJKkMJBC3Z+LvbydJvGLuLB6kxLWE6IKQdMviz0RAm3
zEbTig2sljUBp02W4AivnOBafQ3fH5ZEeKAtfGgtZm4HxxMk2WPp/RCyAK/IISLQoELh1ypVe7Wz
V1F3nplmHac0RSQpMjHtGy2qQZsqDAJJ72g3Gix8OGWHdvgk2uQ6KNjl0S8VjnVN846RH4tj3fxN
Ar4ciezkdISCQFCgHF2Eija8cjlPfzz9psyUrGZjKaa8qiRizaRVplZDlYwbo97CZoWLR+4qkBVg
ly9BdZBDMf9qwuUGnIsKCfLQxiXXxypf/WRTNIJIm/rPKVrYH3b8Kgw3AU5vKFohy1wTNx4IlMfy
+axkvBJZ30/tc5Scr7TLe6f0zqRSr/pZt59n1k3AVVgs88D/t7Sh7GGS7YwyIUCDbIR3iMwudFIm
mK4ygei8kWfDe227KtBtG+ES3iigrMQI7Lis9S84h+FYXnIvwBos32MmdT710bjUiUxzORzkSSNR
BgYS0b1zGPySgI2Vs60NQzYSGCXM9X6Rz7pumZIRrJFhrBHBZ3MDaXCD+DgvwOh3rI+tYZK0ZWcg
innSHEHZXyVylEc/vbg4Gp4W5t1jPAlk3k6x7wdZiusvFwPGosuhSdvqdrn0iGIfc8QJEXWCNBn3
JmmKDXSWLAnL0C3gSC537xwvelXLVGleGyaCxgCEqHmbeO/YwKZT1CoFrxU9K/iJUMH+EzJPrP/8
A+WY6TUvW9tmqf1k6vuq8YwROv0/0IR5f//CHHJ3bEGyjJoi708H4VJqddOr3AQzs2jlKfD/5vYk
WjE1AWdo++KJo7vlDQM5TYbn+0UizdV+SOOAfoFdiR4RpVb2/m5+hNpwTIsCRjJVQpf99uYD150O
+0oNeCk+tTAuIanJvyn0+7XH7lFXIyxzJqfFdPRShk9nkESexTrdC537uD1H9StjrFQDvMKNh5Kn
JXDiyQsICVgoI4gXGUAvhXaFBDDXzxnXD7nvMOXT74b5+APz5NXUziOBzg+ywrNa89DOfWAdhH75
dSgUMUmUAme8TQLKSwGXeauz+h0R4/WKtmuSVRlFllJ4yYwQz3DRdOrKud87xvljuYMKLXc3hdwl
7gGbHxOg5JxwqtLZx3tT9DrpWaCSQQfXfTxK8l4c0RDLzfhD0YUeYvBx+UhOyVlXklqaNk9P82eh
eucRCA3xC9Rh40MNknYdOyP7v1hAzVwxRO6+QxG03LYo9KIAgVasLj0i91tcyxmHNGmZFvaS6Yid
Ydv5hyeQoY0GpbfOKOytK3wh2j5/FGoV8GJtrx6xlQZW34v0ImStN/2DTNn8Mi6ZcReniAR+pKGU
WyFhxgs2XsBNOQHVOPR4pfaN06AZYC0+YG1kDQo1FQVsj5EJS70YWswzxUv2IJ/30lcD1PSd3i4V
74hgdx3FkMN89Qr4oNRbIiG8uh/Gp83nwc2U7SSuYgRBfays7QsNqwTI7IP9c4Z9YN3OSzRr3gyt
mIrh3jzubMYFdDmVixHDiFv0nh1AxqUfvSrKRc8sLhwiGFgyKo8bf5fEsoEnDou6IrQNeHySdpp8
iqsNL21hugXAWB2kS8JWK0dJMMfxy2LPq8owqMKgTURBwNQiq4gJIuel/S7tZdM2suiIDuFRiqqM
l8bb+FxDYNqN89Tj4WyYGeMQg8nLHtJwDkKhcF4UftiSbTV/g499D12168xcW8IO2Ra4bR0qNXAI
/+uO7NxDBndCoP9yypWSgMpa+4pC5CHBhX/IA26ypzE7jXI6rz8z3o2QqL9ziZH/0INZeFMeogaF
VKC/UNzqsUm/S5o/D+rDmnEyQxyUBDDKPwVtQOXl+pu4/3XlTjaLBi2ocSGRqhwE0hE9lWCOX2PN
t85yFxlKbbrNGwByeSThaH+6IS0LW6A3Bp8+FTzOdC3ALItgAt79+jJbm8ZwPHkRyIHsQPCPyNh7
uH/0yqrgxHtCbbTJAk9PP+Bzlme9dqeOSyqRZdiBQMq8bVbL6ZWYhS+b9gDcSvXBHAx98g2zBFgB
LdkXV6TWYbjlG/Z9u+XWr+GQEwT8EbK5U4UCZozhWU/PU5krg/dlI2OJWHvRVf8+JwnBZDpBjQh8
A3gHW0BClJ3q1fDbQMrQ4GWqlXOjk9/POYk8rf4syWQNdrpY+E4pa2awnQQup4Bqpf+6dq9Ri6mw
JwxiYhu3RFJFPDXye8jSOxriB7QrIz2neD3bmF/rW/UXaWizCVx2wNAByf243DKVCtzSExtVo4Tb
soUcwioJv4yb5m7dM7q7dTzF0uUwZen4XVpz1vA0CGY5oMDS7d5j38fWe+ZgstCNsbmnuy30O7IO
P5btKgTgMPGQCcQJZi3628nu3mDwgYctkgXgbXON2xJZFIPkxPRALuJnADpKmiRWyikUCemW6S9x
9isIyN7VN7w6Rukn5XlXkEnPabcntOXoXUGeWLPRQaxU1dVEFkj7lwzFNzwbZWPfue72t7v2s0s5
zlmRXTA4FHhCN3XmyZyn0o75XXi31eYIvkYM6shVyVT+7amFA9mo2j/Rd4I/RguALvWbKHZsdYfe
RKVA/99mME9T2vBg8mKipEZGAW56TrT6lTHrBuh21XOzbHx362AWFkLP6lqBePcFKoR7MdAVJOr7
b03rFm39AeLdpmIwTZ0n6RCtgLr5kB6pcOepww3T5zPlrHkEtvnKqNrnfB1flC+vJy7EBbXvTtP2
kFhYdDmPvNVV4mw/5VyJOdGMZQYsfN7k9zH+FiB8L2UOcC+zoPraPi/bitk3+7WhF4B6/f1CJ+Cc
HjWL+MtCbExcf8JCrjU0Lawpmy/KFgRU0jdtzVYOzltaEJxtkcYbd2jeHYG/KrGtaQrNMP7fM6D2
RIncowVofIVo3c8yeSJCy4LGY8yKeCuTaYc5n3fYuel9SN+YK+YwKMnsADJL5DFywadEogAE9CRy
6gXSQykIvkOe+Aak9sKJW5F6BDdw9WbmZ+4K/38Bh3zxcHctC9GVu9cxhlDJJZ7v+Bn1mZm2k2zU
k35KKpgyxXrQby959MPt5d/HzXWAK8RdTrXpQN+iwDUdyl6YvzvzPKhJk5j4FsKEOFQxySK1zCpp
igjOqsOmO3XCkiz7eFk65Mq4EZa7ZtAR67acEOydKHh/2gS/2jZJY5rpzherdCSSfkpNUfJE5Fdf
EfI3wrkhTddRTH2EuhLWDHswRFSqjSnCLPyovrd0cLl23ZueYAa6QSl0IwNL9q9nf169nlr9Zz0J
aTaFnau/bq7Q2wF63b4/FQTQ/hgktnuxaLw5Iu1Pt2VmDKCGIziR2PFWKihG6lk5mSjAvrWbwwcw
iHUB4bIMjij29UpvGSBtaJRcBKeDcQJrT9muDdEBeh0iPryG8wexo0ZQ5CLf/L62Wz+78zjtohEm
O3jURKN0HmQbOqHTQlNvhwnQ87LrDMqkkET9ODPw5DyZr1Wngn8MN6rAHyqe8FHk6FQ0lqfyGAs8
D+t48qUfQ2CImPR4unJviDJFpSIM3+3UlLPhVYXbAO0/o27jVXDi7eXKBcIAn9ZL95/4K3Oljf07
ZctiAopPYXXRgGV8oxzPUgQYJB0ojHPqYGlt5pIfBbZaUwflbJ0kyWioBahkvqu5N/xIqKbpzoq3
lU7JatRiXxX6ul5WBpShAjoccsjcvfZdS5WtRNnNPTGize7VyeVUoWkiIeyWDg7gbmW3wEq7XrwT
AKNE8vQ+bTA6biC4CWW4XZ4fhqkjZm9fqg2p+hlAbFoUj3nmW/+iZudKF3ciuw5pnXOFTbtej3rI
drYjtiHiW6Yw1R5+JjiC2xa/LhBaVNkQSTtxfE2BTBHMa+4KvAkEC2w4upaLd1WJT6ifnkwGeDn1
zYaJdZsFSP2LWr/H0wU42yKlV2T5L+8LwV49JCR+JyMZFlESOM4URLpuGLgLs/6+k9x/SyVieWOE
E+sukMH4//G8g+V9PLOmSLyZrxQhECF11FMAs+OIqwDRnhdpy2mrWoJIMT1qgKKKZlNC6OJsPZId
+yZthVSIoKUeH2FTGQv5yTT/fXhnVA4jMB+7L8U5AO+X1z3lOsRw5J6FgD165sDF04MjbOjAFZvo
9w9XsTYVBeQZ7L58Q1F2s0DZGAO3ODn5CdMbWsAM/63ztv+FBMf0Or8R8hIN0cVxt+DxibiTtVrT
7bgCeIwvO9UTxOefgPqOG9EAzuBT80Wl5QTXjkpnWDWI7sOwVHFozu4ZIvg2jk3ix3ywLuqx3Us5
ypLeEktFPuAIIGkxpNZsiohKR41dPU2/e8+bDa/iB7P0B3MM4r0DyirOQ3HLmETcBH13HtJlKgNf
3DiTtqQlwvKyahFSaYY7RNlrtAzadC9VZoJmMdoIvv3qPbbifDpZao8Ch7COom92Kv+9zIpk1VSP
NYwIvUNfr4IfC+WTIc+CEpY+2vjjW3wsthh8Pu7rR7dslMAWWgNV8LfMCeaesA/HS52vxkEtC88j
SOGbiiBQid0Za+pwwhVaPGn17ETf24Ydjyo971cuTgbgTZHlLtj7t9c7o45tRnr0+pqh4QDSSZQf
taJn7jQ8l321sPLuQCpz/ADggHQvLtGanbnjjFf8TGGYQvszJ+dL5W4dJyEFSobu51iefE177n4L
RHqZRAj/6jjJ1bvUGbm652eM9MjgMD1LUpEtMGX20o8YFGxngNYuXrIsrrt4nizG7D7f4KqkEJ+l
CsV/Mkh98xyCB6NcB5HD/vEBpba9FIxm1VrhmzWSGgXOAY5eOZ9HwDg9AwfR0MT3eAe+lR0kdw9C
DfAieY9pDN6YR/z/cBq8GYju4QFNiPnHsBLkry2TZJuycU9uKK7SwjVQaxO7OQI9/UEN89tqDZTY
4InHTfirs2pgxNcHZfiBlb9pSO/vWo7Si/ouQm9cPVdwlDeXnJQh/vuN9RqQTV6M+kP7SXBYgwbT
1acOlzMJ/F/PR3KhJCAS7SbMo8gLzxjN6yHtlThpGn1IwvKve3kxWy0r2WdB9Kmtr5pYryimBBGJ
70K7SxQSVZwB6WdiHuGZgr7yn54lFDJAx1FEuvrQA+ku+rY/gMZIUfd1DTnSxWLFyiBHTAnaVsGQ
o6ikjGHpYjzGTp1F7wg6KRWatyV0C/x0+IR0er2afyU5HxFZKaBs5XTxHRDZ4QDiLu+L9FBL0MNg
sMaNCiQz3sQoqvo1xgRw5t/4p/kQ1RHMu1XaTs/c/pKl4Zv/7yAfBM3nQmDbkMAXabZ7cCWT0Kqa
tP1JlqaAFsVTU3TguYp0qldgoWYjXntp5iDDzb81PX1oRKF8Sl/I1snXe1CMRWwhtkfbSNxtCyVm
j/dYv0fLm8Mhy8zoe0oimqHGWjDkE6Vp3sUpCSgL/7/jxEYBTs4IWM3AJRwf1M5NTKZrTO5D9cgT
LDAxv0QX8ESKbIJh9I3Wzx57w23mF1IHDYlcCDIooG0SkOzWoRXidjZC4ITRhU6l/QUpmbgAyGvS
1PL/kBkoTYY0ZvkohqpTvwUQIeU1VaQG+3P2Jyj8T3d9pRS7Q9/G6GXtQXAixKCVY1tczsbMZeKS
8QjyFHh065/fur1YR6Q7fu1VvqA5s9tC8GIip2JBCqKemt8VkWOIPrFNl8JWjuN4hSxOAH4/TGEU
TDbIiysz1x/eJ0GjVPKSP5Q3jr7s44PyLpkN70LalbYzFB4TbbpPrHMcO8lHu/1YlAYzkIYM7wGP
6pAuRk+lsQaIFABloqKukkVfTBHPNzcyRiiN42S36u2eRcN1cQa1NDT/kYs7knMq2QQhyB2cPFw7
KhNaP6iRaIU+7jAITE0qpyR0KpZiBISN9UMhbFyH9fQgMIFWAA0LmJdmnrygrjzgegHz67CBdbLn
RsxhOvxR9ZdrZhTaBMw+5VFBNg8WRta9SsCD5NrGqucYItwZJtKWya54uJoFCZAFxS1TwVmshlGl
g3gj7kfSmD5JTuXzn9JK53drN6UN7bM3b5SGLPMN1c33NZau5BOyLAfJConjhmCuVMUM6oWUl6pV
msi0nFj9n4xyJPUED5NJzopWlcdKt0X0A5B4W8/2IsJSvQuSgDEQdGLB63n8nRH9Tn4zZc5GlpKe
Gv8cIGweTmeZR/N5vtpLAxbZO9h+doky7rlhk/Pt6Khberi0HHpnxwRWA6qw+ntjD1xjk/kP8dRO
BY3TX88kFNRkDX4t5RtFHVUF9bHQww2XTZGGE761T0DWU+qyQkh9zKT7s+K7+8ulCk2Vl8p8fOs/
/LnZWo1F6TwhUVNPmmPEwQxlfeDvH3LV+CsYxw9hfaBv+n8IoUi+6XD838tpfFcEZ99PwEWnC3Af
0k1vY7ffJLOrxRTI0Pigde8A6jImt8mOaJhB8clRCpCZcYMikeuw2q04KM9erp6EHX5uLriiDbsO
4hLhop5cfzaPn+CnRVPMpjrSavyARkgSeG+ABN23MnF5deZrt1/Kk8Jj/BUzSZAYmM1+7P1spOL+
VPF5zUhueV1S9TqdNHUIgWPghBlzVxYUW12LZGTgTC1pVTqHVjFkW2FtbvRldbCXJKZ9rXv5Azmz
hCu8BM4jNcf/Ib+8NPQcUyDoJzlAiYjaXPyuhYzrH3ZD6ColHkdsHj7VaLbls5XXr2gganaewbfW
wKJeZZSHl5zKbAwiw1rhb2yvw7lqpkFYIZOlQmdCio+2O7iXK4KUShz171E9+2V6tJQ9bYZBq7cd
4f91pE6ExcFBXt6t4ZEK3qPrnjLleejedc9umnQ2tAbR7i+4ss1Spi/JVSpybt/VbL1N+ZDF1dqj
z9SRHLEDwF4Ofpt+YyogirnT/iDqyR9+MKbad54NMl2rYY4jAjtB1dYWq6bNGIQtcjd7b7Bak1fP
CeTY0ZlqtxzDlZ18lI2WgrUwmZzWe1pbqIL7qFh3I+TXDR73aC205Zbhx6ex5R51nqQavgGQBPAZ
JyQ2n0eu9w09xoTnEvaiv+0LSEyYCNy8X7GPyjc5MviERM0zV+3XXwnpoYuy3K0CtyNQxrov2+ZA
VZhjKeq8+H92GD23f9+HJuOXwuRPBD5bUXHkky9lIrU1jWesbxUyNQrnk8GtnrfMdJUq3F9FYR0U
1jCYf8Gc5qAS7ifebqOSX4VMkUBS7MqG2scoVU+r4JVDMfMpSa4bOQU95MoBEyyysGIrZdcK7d5Q
dySe90hyFC8hK40kS1U49yfjR8E2ZJoMgxXUmlILq147JHkC+366M/eP+RvuKg2dtIslSXtLSnoC
BCnEcPLwY/kf7cwedH38ESAiIV30SL28Dlu8oTiQCc/B0RWZfxxO3ck+/WOOnm47nLWR7j+asvR5
mqB/pk49jN/i2a3YceWcDVHV5xQL73LORFMjXpmNQA7L3MLKgHyPvy9h63mN2AYRRXaI2pa9pyMv
0XSr5l8zxw1042pZPtWOfsSu2z2uoUye5FyjXty8d4sLo5b9FkDvcRMCImPk/iTeBxl9/kwXxXo8
Ml7woEkwLAOSpixisG6ujAjAYE+X1EsyD0kZWf0ulEPAC86vsMHoXeaC+FHS7pnHiO7zNPPnZfSE
rTLOokfD2h0/LN6866j0AuUqQOV2jXozBZMhMhRb5smG02rKGmL2jObhOxZrwYM/VUPoTu/PM4W7
d0lYgWtfVWQ9CdetxK96JeIiJzsvgFWnkaaFBU0qcHxJYkx8L87z596kkiTtVFsH5n00Xigbg8Ff
MlRiQx8D3BKzN1Xn5HifZfQ+0Li4n7l69kZZOtoNg2t3wBvw2QCKBroPaJqkLkPAYzEWk3K9kAFc
h4Qvrd7AEy5mG5KI3ynnuO2khZRVgbAmfiLagrl9JfzX7Jf1yViACZnrS5c3wD/YS/ZlBrILsV9X
UUAvROQkSwKNxoI+nMVS7+SWN3Pi5oFYo/Xn4XTawLkNHQX2IQLeN9Ls3CbDMC+h1hq4Fn3abux1
gHuyFhGCXCRc+6ELFJunSh/NAZF3eO5ewc+QeIekweHZBc/5tl6CsTVo+AMiE0XhE/vaPIpxsReL
KNpRV1jJo12iKh8PIukBhHVleqde+LGFaJbkg/qXCxspW/5HpZybw18QFEcmEL0HZjpSFKYs5h9H
ZGcfi1orXa+flmmDwqTW31/JCai7+jLVKL0RQNlfHqVmerxGH+ofQRTbwI3wBqHolCqL+HxYg/SQ
Y3xslrq0hFG25UYVsb2S6fZhrXVAeiqTaQmKWpyry1iyZFHl5XzSY0FgKpZXFbXt7z6UawcJclwZ
NNw41VqwWCDSs/MsAqXzkMxb/R4BSr1jfw9/+Y3Z5jpSeKn1zmj5c3qOvmeHuyilZzZHrTevcwC+
r/lddtYZrUzNRnuLyNQ+xqfLNlqmoQbLH39dxVO1lIyvo38HgcyK6RUJ9/lm3qw58pi8pbaE5jQq
sNR2GzKBPoLtAypoBIgwSu7c4HyfrchcxUQtoRRwwIPO6UGPtkff/eI3T0g639/CtKJ6KkOh4rRH
5l1x5zmEDNIa6yMjyuAjPDqgqKgjblCy73Vy55+S/QPRpLWn+u/N8CsN0EnZBSbH8reOInFvWgkT
sip8VHLnj0CLOG203TlotSyCCd+FXM4u7H5173DRNr7uqAg2voc05RxAwcXaoiSq+sN0hiwUmeWo
yeMr/haJjK5Oj/X3EExKdIkDSFdp6StKqEwkj6LnGkWi4rsVsFWgT4aVU7+VNtfz/O4poCdbreuD
mbImgCaROh8+NmCe2x9qlrixRLfzKSmfkkU3bZa+opdXVrG0q98DGG57JZkK6ORb1isya4mnJAXc
mvAp8FX1N36iIW/cnQeILZS2PSeCEghDAezpWM1UpiTMPK43hz/2r9aq4Nr9gvWhO6wDeyj6hMuk
OtDJeY39JTmnq5tnkOtFqPLiLbX3iFvfKMnBmRNw32c51jsm6aUEbFJgQnypx8obfcpsXocU4OZC
f8ZEWrBPBOGFlp13jhJxOtIR0ZOJhIsI0hiHay5qP0Jma59q5fP/ClAjSAyfwT2p8W0NP0asAxFA
5/ZWrnVxj3UcNi+KSvjs6yTiXwo+lc5G9DrEIv7cS7IFqvzG/uk+G0umd5ihwY+Xlge3NOvt56Kj
xZ2nYxU6kGgR2FVIiZ2G8E4aN5KYwDY16/RKLy3Qh0IwAYaK7KzEOjxkohyG+lp6eo6WSvoFRt3K
pGyyQW0DhRsAiSZbcTnzTaNC6r5GAxImB126RfeM2aiCC+AUDTszeR+EC+1W8x9TrgatwWO+fLCX
bCb0zJ8Myk+qo+dQ20srhf5v3oM/V4gPK7ax/F2Z6a9w393CYwpcFxfz1JKfN0fN85WRkFj/TTGQ
T+foZi8BwlGpvf3vvgD0L5ECSYuxVawA0aj5fKbCn5oZ4h8HkksUp6VEYjdHdKxy3363k8W8YDw6
ZAr5rQrzdYN0I5FZxu7DbOR24reCzKXJCH8BbfMhPcQaHt32TRAu7yiqV6Cj91P7rJPsL0dcb6zg
CCpKvGH9y2CAqO6QiC3Ck8W1LZ53iCFm4dD9nW4DGMJMBkuthItYdRMNN6EpWeIlcEVCttQ40Ku4
88UtCtAzQ8WVDEJqRYP4vPvL251n5H2Fh6dQjspNvkwowzE8r+dlQzOgqPfQ18e2lEadtSUeZMyP
o+2w9rlTXMnqgcZ/Ivi6lhaqFvM3nST5i7mTp6CZ8xxO4fZfdDzRagHHxEi5uJpLPen+/uALwTSQ
jmXLATzv/Gt/r5ms9U3MSSnXie/N4ViNQDU3QL9q7+zBIS4Lilz32IEQWv9EsWmW2S2SQQ7M0FGD
FTKsRZoEs2XsbDFXfrrGjgDUrMVq5s91Bfy/rAMHpIUwpe5HLSfYrELxf35Vl72zMbQ48ER68hKo
L8WXFn4G3M0C4R41ep7F7NIE6Ke8tq2O/BoboAcn7VAlm6WbiDYAu0UAIhIAG3G+jXXVbzejqEJI
Bg8ux5xawFFfuZ59IYTbDhtaET7+6PRKNRL4pc096Xt6+mqEsPPCxGh9mQhCAjCIBfBuXNje6efE
16u6zzAa1Uji9++EQRpnLwi2Cx5Xiq9d4V65Ty8lNTsFWbfy/0K1smtLVOYquLXahwYYOIOsaLzF
1/sEaAiZlWdoHNiBVNir9T2RH9cgq78daOIapqHemKoGFMsoqIuC+kSWjZetfZjZhv/HeH3Yn2Dr
YhoyRAE1Uc8/3LpN+uT5RpgEY5Px4t0QU+jHPSJHMIK3X0L3byvCIVUBvdarUpM5HsVZ6ojIvSy7
gJ3NptWRjuUP7fSeh7rREgjlhBRQvaKmnDEpkzubG/8eGzhi5jg5F1fY0GoS0XzAlDQvKt7XdnNu
FAID3HK0rIMrsPKoSux6A+Xxc09+gYks0LqDmlazWM9rNC1LcTCWDVz2rP6gglrrDPkSb77TZX2A
6Ik/j5nLs7Mi4tEn+jDolgRIRgWdWFWpMzcEJfOg7d9Rv8xsrZBan4wmoYwTxh8rcZLy3/QWey4m
YZPYmx+CTujiAfidGSJR0INRxcdgWfPMTgyjqO8Ua8mhQrE3zddlRl+dE12pzQ570khpOp5FCfL5
lZGepaDBbT68Aacj4se3bgqZMr0aUEK509R1lxTHshaAskqoM22dY8JZXqMekn9T2GAxHBhAwv3a
zf0f0QcrP9axC0XpcTyb5g+BAVLu6pGh26/SUOcPl2HPHJqXFEdW+euWTb3uwyxN7Qj0Nxidw2xY
w52UNiQ6HBTzze5uS2Cjf1Yz/dhJ5jl8soYEfk8zes6TFIUTx3CMbQE9IqagXvNslkl2k7/sv6ge
QHgoMGC+q3HPeM6xZk+xHF9QqrgaHA79v1RO8M7PoQCJ8P0VdpXdY0CiUNVGRoGQdjFCMYjyxLzF
DINuHyMVoip4gCjMBz9kVAJoqNmO56Lx7LfSXg4AtdsA6VDWRd9c45MefcuhSfvDf7fx7yWxJnQV
OMvP4LR/TktgppOAbCJkfkO4tfsNEoQE+nKW1AkoRubaJ1046vm5KZXitvB6y6hQgdkojOXWuwNF
1u8dE4gyEqsLhZyYge1aR4Mv88yngn3MqMkd6ZoGvJP/LRxIzOMy2eGUPA/biLIhW47Eps1lVvxo
VYGSTbNep9ZpwRxhVoft57nK0tcfUjNwy9s0YN4coh2AQm48Rl3+wudDq0621HYzPWI4JNDRhAFW
IzdwlK2XJSxDhcCiWLQcWYJtryePvy5oqbP8S4plcog34a/fLNCPMO7xDHNdTucZoWpoefWip6Mq
il+NrHAztiGIXvs7neWFqAj0tX0fWeXLi4OwooQy7JHrSBWhjjqktyUchIdYs/SZELLmAafOFp+z
wkUAXEVDGQA0WzojZjgGMP8xyaqtArYuYmh+rpAoetSvaOSA3oPqzJ14V517f19GyLwSLBCruOmT
m12h8xvvaQ/Iq06jBs886+/uhsDw/kNGf2OvNP3+weVWCv2tjnUOvOAVhLMj1KGPC/ELj/kl71Av
ksxIV+IZRx4EiWXITZaZtyZ+UUKHZTupAUKVBt2OTiuF1AOrA8eFRgplXGpJmMfOX3gBrGufhIUC
69BS0BAuFOflJ3o5H0Oqxk8f+zeEYOk2QJ2/p/DiiXlJI5zi9tzDMOSsukE5yRbJbrc/Hb/UDyxB
HK3xs4d49Hr1FTuAYaPRnz8Y2M1Bssqp9NQoyROHnr82RSD6Ed2yc73YnquobubS0aR3CSvC+Loo
yJpehFY34t7lc6q0GnzUtTPPfE8pW9xsY/RAUSYIKpo3se6QJA2hSbjvdF7Tfaw8N6AZ3OJqVYbo
WXPzAYzbcuuxMe8vmAmHd7bvxntf0AQiYWSwCdfiYFfGHMht6M8CPeAy7X6xZhK6Qm6qHBRfM50q
kt0M11DsaKm8FA/bSIPcbttKjDSZ8rgxaVQ+BExU490sbyUpni7zN+oLGPuoo0+gOyueVBhO0V3A
1CToV6uZm3NprHQcuR87ozgUCMQPrPgZxwJrKylrv+7K2yTganayU/edyVPtOeKSufnh2xFKJgr2
NMFLTUfeF4Kl8fooNiRiPlxlqJZsO6rGut8Ajg73njaQt6qEgzN9AqZJeiFlrbIbMJdWYujUXMsp
2nPkwbYT5UhBTkk/4iWoCVlHXe6uw6SIloYBZ6/6DbBgFXRbTs/P7cWVyNlbcl5lzW97jSL7R3t8
2PXnGleA8pajjyaOpdtx5IdYTk9wY63279ZJolPwFEtqRtyvZoVejstzkcOPpZoGADYfC34KNEFl
o7Xu9ikaGC43L/Bc6mNPV6MB3YfTzBv+AOpflStJObTD1TPon+6KGTLepO17qv8kuGM6O7MxCcVR
BkonRuhLoTPVO32EP4QTnjIZm3o4wkgMVOmAU7iFcGMAKINny+FQPFtBquZ4hgZJSfZQF0T6CE0/
yH4vNNQczhpXFN2MMlwxydKFMhAz7QEnOfk5HGzHcyRJ7+on/vaGgY8RboAJb5Vkk6SNXXe4CW5b
iek5VSy6J0NAiCVRTs+xCn6qQVvIfe8A3nEj3IyAX94aZRtgRak7sf6rS9CbrhS/3MIhuhHBWX8P
y8T+nXIT15k6KVaUyiG0lShfts/6+hJQnr1dwf1gI9lywiDvsItt5vWiLY4KiU88RCUcIM/3dfLx
XnetsQP35hnLKpY60LbdKQpz+IRjcudkKf4/NA+3MtJwBtPFSwxsajq9d3r2Eo5mpYgAfjlEYzzj
GK0/DoFRFhcKSkbQKX44SRCXTZrUfG8vLpoyikJwcL3fpOKZgGdz2Cd0MzWLvmELFfclQNNHbVDu
rWmsnAJkawJnIxwgk06vqUlN5nQR2M2Pf8bNG9sXgjetJ3eHr9GCXiB7zNMxv7IhD3LNLHyhua5B
jI2wjymBrS7Xht3u+35cgNUL9mAU+Ida+ulaLk2lxBcUzGvsrJBrTSAe9tMDV9SvzmkW1IOMpLqa
nJfnGVRKwTvjNkH/C5N666eknDsxlVSkMXc8YcDbu7ZTCZAt/4/HzpWB8rdSZrd7AQgwERGdk+L6
32Ll9n1aQGozMPJvk22s9EOJPW8GmHVpoqI255OQhmpWrGqNnl6Dd6L/VbOMacdh8eCbYzZGn3Xm
IZUkAjXMytDK3/xB5RaOkj7wOaHqkLfzfExu65tcHXuOgFzI2rE/qXoA6RTPYwqbxqghk0QAhhIW
q4Xay+qHGaBOOrB0Bx3kdqrexN7xy6VkFLcFMZ/uC4znM6+v7lyN3XBj22zwSI26ZwrwyrNqTctq
3FYO58M28OXnjgsbvvhaFMBUzgS6Kb9unkNmZyVHDVKbo3kzAQSDknxRSCRT3kgJRn8A34apvokR
cDLBifBQolWgwZzCL6cTYR2vm5AJy5RHAmFIsbpT3/abb/VyQt7j76OPcBB0uKcObll8zbsQz1GX
WrgF1UtJhFgqyC8Cgr4uOhg8+LtXBTm1hVB3rpB+6j5mGGsbVFnQ8lVvYcGqHypry2qOU4QjFMUA
lkakBzkpVVzmaq9jmwuvZYorzO5++gsRiY5f38OzrVe+OwwygkqV1jp27Q4/ibIR/lfX7g/ej9IQ
iwahCEvHhdIBHGS5LhgTzd2SWsZ4UrUyUd9IEKGV3cIxnxc0vpmna6egeYqZ/0oz5zYMegHhhAc4
mYlja2u8+/IiMOhMVGbVRTWazXZLpEq1EhFI7losP8fhlqnSP77aQ1TwZLsEo1S53mMRxclfgn2r
CA5unq9jehvt2TXD5ROz77jMqThEZv6Da8ArJsCLEbB++qVOngHPrpwR417x94ROyPSCWi3+/VoJ
/K7xQzcHRv7bYZ7zeP1uSelwD36IucRsr9Z7/rbtlFiK9JLPSFTm5sitfn1Arwb/VWy/H3Bc575a
iHe4fq3/E9aTOzdLSwXZOBqAXYBryOP5NKuDUf+hh3jjE1VGxqtWRkXmvGReaxJpOTN5ShO2ed+5
lJJwkO4wsaAXQb0ouu1td5DaS42MKbsmCbwCrfC46JnqnP9z+PqfYOESEKKneRBhoIkmVb66OcaS
PCYolW7IWa9psA31iYblTg90jtajmBiCa/7EpIpkg/XPktn9WMUQY4KxaC5pi+iC6wOE6PtTK40W
3PW+H25Vkw9v1/UtSrdW8mzUmC3SdSYRmPjwb2xn+niTIe5VKoAtK3RikVEbLkb2/Lh+jHtUJjK8
/gSXlC2q9+qRzoSfRj0ZKWfvSQ2zNcX7PTEw93Jgp7Zk/nZVFz8L4hR/eXIUf7SbzRSjEORyv+Gw
RqNEg5smKo6dgfAIw8t+myhvzAzH+KkHJCw4bOmDHhHsR34wDvmIEzDqv0GintEvLglH66NW1Ymo
/Wlr1gjOjfolHyft09HWlYFTnKBA4FIpyzMomKhKtEbAZUlck/aMIosDSWwETcBhgLRrJOsfKYeu
92S3+lziVP/Ws9Gcttu8/dqx11TX0lfoDQGYG2Cp8488+UFP+bedZAQn6hRY1VZtcTOxrbqQlKxp
IInmdKG9lNoAFYNbxfR2H4T4sJOILgsncSGIJGoe1dqtKOVT6/t8J9Z7eQfXNtJHFNoGnLZCom6Z
3CAhP3y28SM2GR3z9ay5XcyyTK29QCcsZ6zgv+6SnCwAOyP/DhXNyVUH8JyxNT/tq2yvvhNrn8FH
bDS1Yktv+nl86Z6BKmytLYMkRCOgC8GOcZWmCXZyeQpnqA3/IphmvB5QddE/xqb5D2xjM2IeUAmQ
8u2umLt0hF7U8mEmVkiPAPJ6cqgkrE0KGZdDI83W+gABOpBdXIOxhCXCtUls1q8LWVV+oZybUdAc
7wTBCysE6Tvnie4JzVVcWusf2DMENqlZluRuL2cpbfjs2ldredO2Efk9mhGwthlb5dDSjzcqb417
9BnsQ+o2W3+GcXdT6ncMx83dADkglUNGjICWTFxoNXNTOO41GCJsORa33ZLGFKS2jkEqeTm2htfb
+WMXigVm7LxljoRnW+XkpxaqAdzGS3RvviRmt0sbiQzmuz3SrTPEZNckqrzyFPxnxhFSSAiqlibl
aq0TO3RQy3m9cfPatDw5iyMAj80WrlVLPXTR/VAEp7rJiCKs9DO8sxr9WwoHQpl6AhTn0Yu/x6Tl
s67N87clQHNyp+ZFoMIlE/uJYEPzKGOTLkQIrvUhoiQEx+yi+Hsd/VB0E2d+RJpsDQxqaSqB9MXK
xsJT/YluQXfnkUBpFeyyIutRuFtmDYrccA+OdN88eawY447eQD29XFWoqFFVEZU/YK2xPbo//WHi
pm4sNfa9jXe4/izusyq14NE9HAd8BCki6z1mg84YNK4enG9yXRobAhJLBzgRJKz+KEER62zF2p9i
Zz2/qkfY3sJ0SNW2k8+ipOMGLdLz1+Z3qqnvIJA1YlCkBOR8fx75yVrPv06pRlpG4kRcgQDUrtjM
7zMO/rFABidBobsLJnWYpzXFQAJfyDW6UotMxHIjOIecD0ZoBXphSJBOolIGgiCH28z4U6Q/fcfy
f1t13hmyFgUmOLSt77FgZe+dHxWBSJXHMBn3RwfVAKAD2E9Vybpfvz34Me2gIkyIMD8k+yhv831c
sNezJEXhjo1pD25QDu7LuOrxnla7zGNk6FAFWNsOy6ggmFvmw8T/IqzAW5iYrzFnZvRCVcf5n6Wr
rJAWmlbcQge20BAbYJurhI3ej+IC+y73I3KrVB8IMpYFTZYXZSd1xBba+OLET35GiPd4lq1OSjFV
dDqwe4xvHoSG7E6tsIcvSdSIyZ6Vt+BuhDn3gtBBhSXDDN1mOhITRZDND7+d2QXDJszzOrxltcJe
+VVKrVzVoyC1/yE/Apdhwcjk5nEKjemXv+mfoSMNIH98hpLdDuR8zuPg8J2S5Z670THicF4N0zqz
2hXrMLMoEACXqChOdrCw/WlaMtNcD3vmyD9UC4gpEyjywNkv+cDSyqO0P+kNSgmgbAhG3pVXjtnv
nIWmhy26gZSS17o1teCYj7MqjhQRc2J1bEu55pJwEr4L710FHGWwcxwh7wfNYPJU3oGf43MwyE0Z
/dTBJ97L5nPRZeNGaoAGeDJirl4tgy8P7XwKX48NndpcRP7KGmw1qJ/RKTzsBoXrHnjfmkugbGHP
s8ONx+SMf8VPE7WyPuAZT2xKj+iC4ghETzpWGP8eYK8rarDLVk0U57rWeX4znlTUKPcRGGE8kDJG
1Wy1ZpjkDx6FgHtGm48w2EDQwgUs/+9mLl1aMHRZe3hMBXwPV8+hhnbgfOV4Gmzl5nDzW/ufLwWr
wKHNNJ46exWMzMR8u6oaA6mRX931TtgaWXxTcIdganwcRyAUyV80PAZ4DyEt6/uVv7AMTbtvYfRS
qjHq83pUkPVv/dpaP2EWpeR1rG/ArGH21ouxMywL/YOYxBRbfpzFuCxTa5K19bqdPHUhXRIEKdcN
nuu7G83YqjviUEyCargHF2rD5yKfVM/mqCUplsi1LcwP3k0nRISAbgIk1bs7YvQtW+JsnApoo3g4
h9Q90g+5q1wr2vemrXIM3AvBce73sudwSOXk30vXLC02nQz6/SPG1mGwherSkUpF8Vaab0nCv2/e
GY4sgb70Cu244TY+c5lGKb6lrU6yk/mhGhFI5BheWnI2lg8DpQS1POEjLwu67IbCsDGlTUzwGvZK
GJunT9PBjKr2OjqdPJE5HJrdYB9S3xp8/EKFKsdZ5D+CZHOh0uAScwulNXtYXYcoaHJ73HfKs7W8
1ahy+D8SsPeuUwpZ2HR8sk2nMIR8XNkkSzc+QmDNidS+VeB9ez1lsdM313KdIKFA9r5lFHa8fhm8
VxJYPLI9P3U1oTYNp+SyOsCRrQzo8FT8p/4qAmvwo31C5w9n+u2eJP3IWG4CNjvi2OobN2UXyxIj
m0gtJ823Sx1sF+NjqX9Ays4XZ/ysmXCKrF5IXqXRP6Yr0fiTj3JSsxml6Ap5r/u8RrTi8+Z/cI78
i+ERWzUBjCZkV1Ygm+7vRrA37J6k5iiQ4vNycf4O0NXo05x9q5iAdSY9+4HxeHpytNe4YYbsYgFD
wgSDu+v2zO53S0OeQg7gkl8azAppG76UzaaeVL4x0ISE+pvDlWTkWgZBJ3SEYpSKrVHXmiFRYBtJ
P7fy7I9AUz+nfGeU15CSnIIZNNilVkX2M99yOrDZkzK1uA67krUxxaCJFaZ+3y64eteSr0a+W15p
UroGT+nyWeegzcUXVEulIskYzBcn82hC7G0altD8/NFCOkU9BFTFeH6Hl3buJ6VUfhQ3Ij/q8isZ
a9E/q4qbxgGZf1pXzUiFkPMZTL6p4C63LjOIRmfiAZMHiYQ5oWF6f2gig4kw+COnjkaIMxKS4Kea
SKpqkdU9aBJrw2I9Lcr8OmU3Kwl4MRhSjClmobFvb/QWlG2K//dmiwYdvCWmFiotRO59pCRkyUNF
xagpQeN4itPTs8qes1Rp9lIjz5mZoFxj+rK7E1a0yhPWAf4Nq2OG3GgdLaMnhTlp0I7cF8EvIhXK
BsxQLnAirwWXF6Vt8DdfMkzCU6/iWFsLBAe5WCxUNrqvw0PeQcggjBksJkIeGuVaRsq4itmi3REv
4msUb4QOkiKWwQhORFGX/NRt5kD+ZoLHEoToSMP8/j+wYNeDiCe/XE5vSVHrLS0IhVjcPQBPaV4H
2tjvBr7nNd+3ekFz8JNUMBj47TIsqn6ynMiktqxSNNdkKIsDMBd1SmVf1ERq6ptHeuJqDG4o1xmO
z8SWqxEtvDSY4CkFkd+GVwEs9oho4ToT+RVzyySXd0jgOwAIMglaxktZClzzQjfaQpWzNrRFVbhy
8c8kBCapyRNhquvaW2gqRVMhWDOpBXou5RGWoQ+glUY6/7h3nv60TbmpG7fLBWqXkwQ8HlFoemob
mSdBK1iRZC9tJNi5nHWSdzR2MXynaUhlGED92+vs0CSoyOoDaX51/vpiOaxPFhwDbUgkzx7+G1Fx
5uASgMxIYw0Y0hWajcuxi2lTJvM9r2mMyZhk89PO7dv62CJZ1Crm4jG8poYZqhjBPfgoEuzMYOE+
8df9NSusUiFCxStqB3m5FOxVr3qjRT7Rcu9XwcEV+xWJ7KFC3HG55qHGKXKReMWSKzF+wo5v/2IY
c3g9pGOfhjVjs+w9b+khc2agvyFJ+EITo7qeoN25Sb+pZU+Yqo12Acm7AZ9U1+3k5XbblB1t7IIF
ighsphZZHthfHW18OLEFmmKzBePDHUYqtaUuGXii2RrcQU6Z9pM82TSNCJuYbnnvOFrvhtGEGCoq
Pxo/YWGVnlZOzVt8BdKaY2kTeMUSECMohRpQn5T06pzzHFXifF2pmUl29qilZs2EIGQpdl97hE1h
MTisYY/UcoxPfqHX5XqZoTD6/xnhj9uZhSOweJNikjwUc5oP0MZHBawOln2lU1Vemf2769n0oxYx
ijUlnovBeumF0ZaIrqHw34GosOvj3j9kaBy9Np6p2z3PqUf17Xz7scjCzYyGwRHUsDFZsu29eSJO
RfgiYBXCzmcb/nWT1z25q/FZahEWJ/JPQVTsnzsRqs1J27FJlAbUFTlwmW4fuSKXjRSCQp9U6TFF
kT03/3WViYwR40QKzTfsMMG0B64D836RIqONFr+5Y3HwerqMLjTqQLUpUo9cPNVFu4Dfv/3rHu7O
vCKaf29SQGs4H14JU35tMc7FOXDx0FX7tfL8wtjO60/G/XT/YR0Nt7Xw4YpiT+zrSFz9/dkVAXfc
HZida5/BCd5+26YYorv7EJqEuVI759S8lGjAE6gfvEM+lcBF62+fp5VqYEXiXfNrphvQWUFvFkkv
/b4sGu14BSY+/0OAlsvmyBHCBk+1vQ/N3KZN9To=
`protect end_protected
