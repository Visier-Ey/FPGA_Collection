// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
DLwmzhsA8Yk1FQSCUEP2VsnZvuzcHDGSikzWniQnrAtIqFQvLbxrilSbCsTMdUWA
2j9CUYLTIZys24yVvExjkOOkK2MW1UXiEWlXtpP/BzIBs8rD2So27GxOjMm2spmd
CPloFLESies3uG+9YDzXGCNLlItpABHtQ0oMb+N/F1TMnGlX12OJUm73yaNVCMWK
jhsWQXCdCiadEBduwjnsAxc3iaHsUXSPZ9QCTRhiFkp86Rl5/N25IO/Zi4Gwp6xk
yC5wJ/H5tp1tDRRd0FTZvcpoTHpJpRvRfow4k88Ea0s1+e7bkbs2AcspaR+veAey
ZbCj0xMNbjRkCGzGrYJNcA==
//pragma protect end_key_block
//pragma protect digest_block
Qfm0asAEX/sUidbh4nhkzXPzBmM=
//pragma protect end_digest_block
//pragma protect data_block
XMIwpQLfuIyF/56E+Ma60rHUKUNtyzBs5NHlTYZMwyVo1u8d0ROOPlqyKO+XINPm
jUVr3mYXAbQqa+8TkK7zvCC+9KMol5TLLji6hBIB+NfKF7xTUkHe70vpNg0jkeh8
tFv7A7ACMcKiGtoitILlff3apVaqCpJO3M6n74Vkilpd4lQ2OK4NZ9wfiy7o/DeJ
lhSb917lGSJkUcJq8f31zEUK0oA7YyaAW/jYn4oMOO6wPFPHZNWZq3TsRfmrf6Ho
y2QqsursYNpDSLj8uECwD7YP/X2gZgDefvET4mRczAqYq1+P0BNLMmjpTkNp+udY
0iKaYqbizo4pu7R9NNg//aewp2X1OdCG2Ct1UDwawnPmBk12jZZ36Ii9b4NkJ8j0
fRAdIWVMXw4tOdttw20kJy/KH0BHRu5Lj6uj1bSW5aNqqXn1qXlsstCOSf17EFrm
K55hUqoRr8xWBAPk02inWIeGRy8OlddYx9AWjpDUQJd4+9OkTpqh3M7prFmKk9Me
CJjX8zFJowp38fIEztyGblmXP54CvphzCGnKsR/ak/h5965eiDOngOFpcmkeDshy
VogrC2zMz911bz8y4ySjU8lHVN3cAxjK54BkH1R9Y4p3bns+OBTBiZZsa5M3+3Xy
8g3tInoPay/gz46a0lcmSks4q5VkId0uBtVXoYjOfBWXBhKNSVAXqaEJrBnCtRjg
CCedfA7WvAILbjGXQ0HX+A/FNlGpMXPb3jfSN1Wf/ZR5EOUD2vwPPA06JZH3ylAh
z5Cms2MOGV1bkZKwaKj0DClHUsrpUD33JzkjOSXI++ePAz/KCbW7VnNEJlRCnZLr
upLvLZWf84DFA4dCJR2h2om0s1Nvkz3ITEpsj7cmQoSk4jYbeKLikyy/mz8UxA0N
ZMSiIMzy10slrIkpb9jABOm+sDv66MnC+NW5o18fcSLBnbXGtuzzBZZnxuVsHQyu
i4nkZlkA/LsvB04s3thGvCgNWXTvhjLU6GpUX7kLj5g+w6igwiWNWza7zqToquns
9V4jgcbMc3PUwLoYwprUlv0sIVgTg2HOTiEDumdPhkhXZgQvKfJpxWVqbMGQHGX6
/fSSCwrDoxbaMfGScEXAN+UJgldeQcpst+QdYoTOnhnYtHOxy+p5Sf/G0zRK9IlC
UFMr7MXzHcWFyMFFgE+IV+A6nDVVOFGQ/0aUtVtik09/dJKm1y+VxovxNkUiCie6
yuSPysUNBhipO963rhvZGvYTqVBKf0WGX1iyKDVsIN2mRnvM0PB0rY43OgTrcciH
olIyxxFCd37pBRzLtSTUqxAnmhF+DO8T5U8fz8xexrp4Z60NuzvYn88Cl1gnZW8u
sQV4pwlO23x6yRhgEj2JL/uuWwSOnXN6TUdNDYyzNLXM7NNMoaAF9MmDjbVZ375Q
9MkYINifRJHmd9tAs2ftlgZERr6l2hi8RUBQHFcKFxQlX2sMACdoUctKEOpWflVa
BGG2/rNVwZ9qBE5Ak8iNqU8EU6VkW5OSjfIoD52P3Gd6Ry9s2Bukkof9DNACQ8ht
3rRmCVABTnQywI4k9nl+dhNukpFGsvdBouxLGV7xTBVEWG9bSchXRorTqkzeWMsC
FoSYtGiRx4r+HdI+ncpbgOEM12aNtJCY4qne6m0LJ146PAxdXthlltP/uFrJ7nHY
KLwYLqIB0SIokb9i21Mw0U/Ecwuipei3i8/FLO3WD61P3Rzy8EdFMciil0hOzOlp
0IbnkvZGVKRb5aHOg8z2B/QZi9NLKDp5Bd7r2D/mXanAESUtwE+Mt0d0UibSNL+h
wzAmmci48XjRi19Rnipu1vuRBsX8B+rzZ9nnfrnwwyyux1yXRpfsf7BRPD6ErFJ2
v6JcrkGUFK6KpM+5c4mkJuXNXbeZ/19ruUu18eJm/oXnmyHppBqBwzhnH4ruBMKz
l6/T7GjoheyuNLai3kZTKdcxhY52AD8DAbbTNh9l6cesP7WTOiiVPh+gIkc9cTRy
q8rK6CBzwK2I1zZpwyGxLHainrg7bS1rUw/Rmn+yonUgBNn4ZLFAmwV4zGmWDwKl
9810w6Jc0+envgy3gmAzVX+XXTAfV0OhfejlD9Cl05EmY0bi2EwCwlzwcLsLlIfB
FhUVQH6juz7UQkTwS0goqoWXURm52pTsPzERcI93Xb3mYXeTNlFsbj2hFmsZSeb2
VNAf02R85p/KS1xDkT9I8n707D8Fhilvg7vtpJIAc5NmxbIPfh6n+z+jW5k5nIpN
5GWFST4ZQqoySXufHY72w3JnqerJx6s528Ks9uDhDrLZxcl+zcp8NWKM+Q3n2r5d
kPYR6Hp3Kcc6IdNRxiClyoJl+Soc/mhFoD1rBj7hIjt4jZCicXfnovpgXq+hvlOv
VMeqarmPJpzANBcFumbNoo746fqFnp38oU0p3b3Y8y6sAOdxMNEqq/ty93s22k0V
40V2DP2oYbPhwwyxcfXUwq3flgPFoTuS407K/peGx4W59CaOjEQ9i/j7daZqjKbn
YDiKD9p8u/iS+Mz6pJhAHMatycdh5/LYP55L0z+LJHOKVwY5aw5dxuXhDDxWGE9+
EEd6jNKr7rig5OS6AQGd3V9z/26F6jYzyp6Dqi2xQf0yyDYRlIbrnjJhMTDCHYED
D+ZYsDvma+Gi/gXBb7iKnKokEFSxIfGx3cZf8d5iamrmtRrarHA3RJrD0rdZiW8F
ZKlLwvZ2RYcTfAxZikNdJhzYxTdXX5VEahtUrTyK8+PIT9p3bZcGPtHlBNTNY6EO
kTNMVHk9QFl3QP/OyLWDFWd1AGXVVHeMklbbhey4aqnz19wf4OX9VM3cyOJu/mUm
VoCD0I+29iG5fLPLHhNVmL7xhMSR05FR9Jbs6AWhsjQB8b2PXiEN/IkySUI5Z8T6
3w9LlX5I6wbkJIQSH1vHaDtz/mdxUtDFr752p4ui+YZBP5YUWaUmB2jojFfng9N1
TWUF8IH1lpsE+zrnBTt248owzx6yOHEeQuiSL2HVyaZkahtc9oaXrWHHXXKDy+Co
ohXb1kHqUotZXwYXpJpe8x02jylOI2cCWeVDoUnaTUtQTYAauD/7UcF00DrVss/g
evtJbk6IeAJh2vFuSWWAKMkRwGGAHla1+qtfv2tpM8JAKFeuz209kBKGft8E3+3W
V+2rgozMx86Nm5ZKX/jqt7LrU8870G8U34UBmiVNBvUyewYM0/B29Ynjb8igIoGg
0bxAe/d8Oa1sGSAkfG+2XPFN0b12yrXq6qPnejb4pDUdOJuklcV8ZFshziKzRImv
/Nk3m1SsjmLHhOomT+igCmLRh5UNBVSlsB6Fy/aAqNN8NieexkQP3x0JPobstCnL
Y9o/JogpY1tMvdLMsEem9JyamjFYNdlJ+a+fqicAL7bSTVxKAKMjA5vFRKvA2iwo
CKgfutfcUVN9s09blV/h/dBryMXux3mosD0Bupno7sx/0dL6TJNmQEVcEQY8SRpG
MISoE7XkOt7V6R0RlvOmWYnNutV1fpbxEIQUy/MHtvJEoDU7UClvmwJghTrjQKJP
xNeiwY6IwvLxCfDpkSoEcF066ZArZ3UnTi0Qtj5Ab5tEWYtSsXjL7V+LjnsFBUqV
J+ncsDgwQ9i5u8VkcLt8cSWKKBzX1998wKSM7IOZyf9JZnHDbIn2YV0KYH/aH3t0
39Y68WhdLl3cdSEIwmC1L54TnGk4sFv8O0lxedKjEXO7OgRaHAaisqdAzP1v637g
zRv8hwAcyxNxN9vz4mFoWjax/Ithi8OQ/4kuhjC/f++Jo2zmjoqmFkx9eebCeHD1
1HnCz7Ewq022kULWk2JDUZNCxiWf8thpx0hkbZ7SXQcexVcQH1GlWNbFQGVMe91w
N9EKmWw9gc6dmLA878G8vrk2W3oIdPu5ETnShIXlFE7LeFIg0uxvbQyhlQngbGnC
R3r6LaRYvvDuvhGc1lwMPHNhluot4/DoiajkPJLA41E9SDRU+1T4aI535mXqpxcw
woy3g3gmgSUevO0kH2oBpgqavTiy2itMxi3mzvjlL09jazr/CYm6uUR4aSMp1Ssv
kv3K1iutenAiRHjay+z46OXdTlXZuMo+nInXtvjnIna2X9Rd4DczQQIGOfg9Toep
Yz/WAfHjT6rWzRz/G5g63MVSTSDQEo3Sz2I0p6WirldyMQO3wj+j+kST1Yo5hHj1
kgaAxenJGlz8rRK2MJLN3C6LejNePX8udgWETQCMVXH+ge7eFbqRvxNqlN63Z2Lg
1jgyAtmQjRJq9qWMpblTZL8tEjlX3XxzwO/+Dt1a0KSIUOrwLCmAczGZgAoC7+KA
dqCYARr8YF+jcNUnJ51F1PwDdNjy8FGiD+jXUERbEP2AewWneGs9YA4PU314lcTm
1R/VK1dHiWotLteQ5wGTRbMiSqdNd9MRSzRyXP7amyMXwknXL/TK6OGbWg7pSD7+
Ofi2A8jlpftv+WoSGcqI2hUyBa2T4NzAY6CQsU9cz61/AjmwT7dY0h5WOYrXGTB1
ni+m2F8fnvImM+QENyi+InCuewcgFuJV+L/OHFBj415isLkDHrdL36cMuYti3Uf5
PqMMTRZnA28keHTfRBW10zEJIGZlau72zToUmk9em6MgcLJxZohLJ20JmWfq0Aqc
nRxAAhHT3YOH4JG3oX2M75neRbN20qmiInPn15V7nYQqKfKnQDC6nWGZdcYQaLQ9
+iN1WKZobty3C4UN4XqGddibSLy6o/Aby/qYs+GrVey+CYiQrby3yHQJmSHzOVde
BrzK4+Wn+l2z+vd5YzUGNq3B1nPCTyeuZrlRBfg0EmLuB9Wq4e35GN4sWn+OZfHu
KgHxkRL5cvDBVjZYKBDojQb62bhgXL49/AIdNRVg/sN+cCtmWELdqyH/3NGnGXhA
fwWD+rj0atCUxrFcD7CZ26rvErjQBszqt3ViRjbywRCkvWpKLG9SQsxRyafM89X2
QiGznsJj7PJov3LglKL4GWj7YHwF0ybsc+GvHHwB0p6cOWsoy5H6RlMBinEPAgfb
foFG7lxpiWiKSpZqW0/Sf2ije72TuMJLhZWM3X2qYsL24Dyth+vEVAB3+P6SR3GP
vlwPgh1M76MGiMCEl7prpejNm0xp23b7aV3Gw42DqPdCKXrSLQw6rjT9D3gZ+611
I5OReKE1/6dy50foq2U638AXDBptRhZlbe6J4RE266yNwPcDnj+3W04soduROeNe
/qM4U0QNfmdAoD1ADjkdoemyHhL6OdhMutnjeywpVo6KZl/lDnflAW2kJmQbtrVQ
Pxf60TSmAkoti9dufm8l356Ii/SOyDdbDjLySquYu0NW+YuWoYoshizQStlvuyN6
6aKA+7rnc40rtWcdTwe4kzSnBwn0VtvxnLjTy1XQRLVqgKjMcNdD/9lCZVQ7pPbs
Mj1Wi/PTzFyBFmI2JZfb9sUNlsd1wAzIASxHV3MGzd3NwNrJ23LgpOUWVf7f3VpI
vlEnnBh3b51P1FsCX/Bv8S34fkeqSorVURDZw7JkkiD6UY+tuKC+FsYnbp6MNJ2s
ravliMiIH0b8jx+JlJVXqhWb6QbM5AFCR9Dvz9PS41arCu/iqV5x1+tCDPwqnjWn
LT2NsdGmz57r3KvLD7MYe579M8KlZeX0S3Kudp7VSuVF1UdjPoxl9vYzH+XDA0xO
ZLeEG5xejKSwSgCLGmamhZL28/pQMEPbg8gGvB2+0kJDdeCf/g4zXg6iiy46CQ+1
BlCyI23fIQXd+VUwx9oLBQTJOpfAQ1/feZFObSOutnaqfvQHkQaGDyteE0MdNePY
ZwmH30IW+4WbyxGkXjh54njOjPxtpaUiQpGXCWWX/d6Pw4Z/edm4ofPvSQfibbNk
MZt1tF2dZXTvHduFeLPlOOQ7dZ+rnVoafw2K0+XZiuQtjCrYsdNAv2/WoHtg62aS
mzD/Njc/VF4QphHhLCCBuGzKwxWeEVCBi75lVpfScqv77oKVu9ofQg7EEoX0ASjg
cOjXjugbIU2ZtWM5vZTs9VnWpfVY+PkE1gjdsksTtLhi3Um5HURID4fE4ELq/iHA
IW9q8H3WLxZ5I7x5GhE/uu/6V52khl4BeF4R6vaMlQFwApxDRjTxS3GEq84Fdl5K
OzX2umPaepWRyFkKV9i3wE3iBBX3jcI6SNpx6/sNNoPsquy77UvzfN8WVds3dK4E
EwhFfRP689ItnnyKuNFXtOdY3EbRyNNQdHwgaTiCkjPRIe/UBqAq7PYzXGO9Xzwz
V393mHLZu7eVJYE62lX+uEOnLmVoocPxawS2Tfv5X5n4LTtV5llaqRlwUoL9yAhq
Wra0f9QUWmiGHe7PkrURX+KgZNYjtsO7piGLcZS1kC5cTHe5Fhni3daLv8PHpG2v
aNz6YjykE0w/yyQLC8oIPRaHfElYtLMeHGnfZZ51C2h78zsVMS0GkQcQ3nPMsz55
mt92sMUIjcjKBOtcGnUiRBZASxt54ysDGkn1NFJgM4vbZWtEOJaU/LnLWiYxz6Xu
X29yA6It1KY/4kVA02PtQ5oM9DEOZZMXUcYI76SKbDqa70YKvbdWMd829GdeZ/OA
4RT2C6inIUpFm0Z+wtVkK5ove4t6q9AdOt1CxrNlUDrx9VD0kBw+py0AE0q4eDB3
HRSarcusR21OLWIRwaBwWhLQE0y1YDeQKJllz6J2jvE6g5whJPBELSQyO12pyh4u
02xJRb5C9sEQdU8Vec82uAaOpUmidzkFZH14ml4syADhAo7taUkAe/ejCfK5nXzp
tnpkVwFan/5Pc08wC/HZDgnq3yw7XCnWq37ivsMsqafSPwF5GwjLwSkrDRIY64xd
M/gejk8CuYtY8s9xN072WJBAaFiJHP7okBBKKutIMZYcjo3WpVqkpg8Vbb4y2abS
S6CI9HRtCrgV6gJRUxsx8zAGjI+5ihsTjAfmjSNQWcx4gRJGii+KT9aLRXxBL+Dj
/+jdQI2Ld4nofHMJakQgO6beED2ddOdqm2amaw8CJVhKDU9sLe7xbToBzc38w73T
98VO/mucFU0BQvMgTbXGYv0pjb9bOa5hxUGPkBhWxbWcnFWy6vjAi+jNotLxnLAa
l1NHySLo87c/4T2TIyJHo+wF7s/6dQvCvyOdaeNuCM++AryV/o6smLPMuWFaxyfX
HZHFk/JT5PCXUDTiZqaY4oWmHFeN34rqcYlFDtB32xDAaU6gMQDwK0hzVqfJfFgY
kMJw3wcCuWOuljnZdl0M6MC8arXDdOHaUMu0ftjh7Xe9rFmLcZfDQq1CXGrE41p0
ILfqoS6z+hm8lOsNUPSBrG0lZ/ehKbFY8Y5WS/X3KBxXKANlcG8dSTmr8UY8BGp5
isAQV9Wse6ifjEmxj/ZzF5AGcfQ6Rdp0CFVR8KWZrrr/0Ytln98NL9UvYC6Yubzz
DE/j26N2jc43BjDi6PlbdEBLXxFfpyRygpgU3LDTG3FEpKGnRndtYy0tq5oJpogx
IUufja8LB7s9nR2KaxePARrwTQ1JBTxsSzy1KNA2TCSfw8FHXKQCm9OHR2IZEUQ6
NMPm38NDi7x+HKMClH19jH9CzmXVs/BwZ9wqmKaHCkdEdAmp6uSJjLuvjmLfF6G2
9iEg0b8/Jgz2WlnCquBwwxieN0KXEopQ2T3f2tsEGbXqFeGtaFlQNnmunCc0r1ev
jCP/PE6OkGfXzrdljd0kWAcUH0Wv6tDI5UIK46ZlImpt3q6S8tpb/+Cs9JeOPzVn
dw7MKadW5MIexcz2C5I+rFvD2WPBYXjz8tKipWzFdny7/uJra37a9pWsVmrho80A
o6qOYWz0ZrLrwl23RM52MUj26OuLuBIvFWjyvdssV8SQerOZNTzdHhsupJhlCFQO
3bmxYl6uUQFb+O25nSYa5QLoGitdpJA4ySIU8szGGS2mgdKV+q/hETXh7+nJN9gm
NZKIbd/ykw8QRAXyQhB1mVkhwPnOyh5SOhewZ3x2xa9aFdnF3a8G4reGirwB35e9
kZBDguX3p2ijGF6F3zemqcmFWDjxw/9X1C3/+thDnYY44YaIyF23ix642/61Ka0t
GJWnRKQTykpwIYYtYq9p4/ioIySzwONd4IKIqO8ujeNmikGW5zUOP6ZHQyZKo3cx
iW6eKYV/srawJU2HRrDuKvpk5fyGAXmeSG1aHFQwCs2JcBO78tSzGCHnDIJ1vSC4
GP67NRw1B8iyKonFPaav79GRWvCTjQh2F6q5DBlrCBle9gqJqzGRV+PgxF6zR4/8
bqURXk/flBXerJrKLAugJuRgRImu7+VzsLc0b8BUOl854NB+f/NX7NtiBvFMEIm8
pmBfvwsqhK9ByJHM9csfbKLJa5stGZTNdd+1HboNMyJJVSl84xS9IrjILnlx6utb
ZZqTUEm17SSRXGQNi77aGL29d/x61TYEjnU+GIXsuMZEVeyvzQ2VTvo6/FSQ2ZnC
ZmRWtFRUC0fQQHZo16FNvwI30iXKtYPvDLvCB/kCvdbUvJNO1XatsL4gTD7wM6ys
jx0eDGRSr/2/JZYpRec6UqJorTqKnE7XnPEV2XYTTUJ5aa7DSwPYUXNNiEd2hePX
wErOlHrJgwq/A/1mmoLD04jQpGrXyCT5W8H0gQ4lZDhb3+QxFeuVSuoERTKUwc/w
8ec0O2ccMFeDBaFHeRAYDh6uavzCU+4xR4AYGzVJh66nz6HCkko/os6piLr7NO3m
laQFlh06+ln47afYbUnqQIeEVD/pPoMHkCDaKJlBRJy4sRyJgNAjqZZMAIWyAeX0
UU9JUp4ECfs+DtI25j4eBa1DPjij0h9yUJ1ZB8M0ESUtBp9+ISbaz4KlhI1bd6As
msgyho3O31tpuk9v1M8I7Sd9vweyR8j4GFTweHVD7dpaAuNmetw8Ss1lv2BdYOGf
DsmKSdGtyGLr1tTcuDU8V1y1cu2uiLWD3XAxCsSzXLQoG8C7mPwu/QkshWYn3qWE
wwTCQUFxoi6Nuv6s3T6iFO9avG3l+SatoenUDxCfU7PsghARuVbq6k0QxIuc/332
IVken0NyfCKab1UKWhhd+GFAprIip6TAMvPLB8YhNU85k5s+hghG5eYsjEn6eN8i
gnFEeGjOsicptpWrhpqZyeTxI2HiceBqoeqFNID01MLbKPIN+mE0INWq/KL9PUI9
EKNVfECj2+4ouZMpCBr3Rz0hMaW2yvtvNimC9RNbeW5QdmnlJ/PrrCBdvtTDjk+a
MuehCC8dm28rD/4xaeOqO2mcfGhMcJPd4exyMBFhrcVMppiqD0J+xWib8tNU/X/h
WOLZnVbR9UY+oB4AUvKlp6Qpy3Bg0Ub5M21IvMRTmS9lCn8cHaOfCBRpYxT3WoOy
97qQNDKTP/dp/Usr3Kmm3S65DlJVlyJdb4DrRgmY+FDOKazI+GOsXy4gxiGNpipO
0xBC4gGH0HurefkO2rEcMzU21BYbo/hfz3a/nbm+m19mJWHxbi7laz3GUCxyiWbW
GqhBhnOBcz4R66tw7iECtCs2/X+LiXPWhrKNtu05wpmG3myJrlvRgxhw9l1spadz
LVxXrjVOw61jJXcLHxyZ1jOBbxs4Y4YbM91yZC2KTfO6W8rOIXb1QgE/8yANNiJy
gg2wTYMy+UoZQc88poKX+Yn+futCaFvdaLDPig5S7BgDBsE+U8+PerWYVT/CqXj7
WVNFMwpsMk6a7s3TNbD1Kp37bMECitcpVidSTq7st/mSpMzqzi6UMmpHTCBP82Sm
fXLOoMoJa8rB/hM3lEiNn8IsID+boIY/8dCy5C+pSfwNx/z7gIll024WtevZeldn
+55G0pteTlJb6yZIL3rktDG7lWyVnWVnf1V65ka9nDg1e3VJdMg85CC7f2dJqqdt
xDFbgcwnagKiY9LeSIYnpSGRG0LmZAVw2f/f5+g+k1cZOjHzJ4DNZytNXvcEZ8Gg
guA1ZeyFocQsNs367lmbe1FRFKU63FCsle+vV9/8sv2H/ylI0flWaDPjRhNbCmsB
7wb25yb2UgpvRu/oArxM0Deptl2QVOOMPIFcInT7Lmu7clGV3/xTZ34dlh4m3WDT
1Oq3thTQfBJy4wdMDxnXlsoBy6Myb7dxHeN3w4bQ5TVuXOG+KTmizImO71V+Vxy/
0Nin6s1koIvJBlTD9yQwB8sLhbG1/K/UnZyoSSIDDzto3ij2V7XlZunE3y07zstq
aCSs5BhW7KvGhYX1EF4swU6HviSUY/MJM1WH9qKVyFLULp3z/5xN7rfPIbT+TQ3S
gIeNa1Tzvrws6RQYzymq7vnCI87ykCw4RUlZN7nsyeYiHUPgyoYE7SxcEcXgRcsq
BgwqcjuzKUho1T/+QryXkGATx3ehH5iSMMI4y3fXciS/a/CEJ9/UKAadjuGp3hly
mLUf77N9inTuCbjmQEH1UUhnILBIdS4Bt4wlE3N4Epz94b22ToRsbzVGB9nRQYsW
kamPhVmyXk7NBQADJjV9Y560PVmoQ9iy7NuaqRXQFydXpHDavEYjgejirb7nnbBg
9pKvxX/AxOrykeY43Nu2CSv1gGy+NwSqm3cD4MamTDpgfmxeTrjjjx172zkk4INh
VSb633eNhGiHdchXIRJq0Fdc3RLu7qa03HtG3np3P8eXO2b1Ty7/Ik0dTH9qfIDS
DsZ6aHnWCA41A01TX/qX6rvf5ForR8KIDj1jBTlbVX6uIfxSLyGkCCF+IGQzoiYV
Cv53LrKynQ9FVpoSpk3fArvjm1qIZX2ieWm+PDIAqppSu/s1Yeqacpd1+V2EiayP
cU36maN0f/nrt1s8IBkwZaNUozEvHI45O9GcrhnZYwMEIuf750cvV+V3tVpEi9PQ
36r8MLiobcvblhAj20/5wDwWDBbN6aQdBsEg3kcec8IS3wwSmOWGIbxbgGmg/BI3
R/sQsd9aCObL6aTiOHvi147RxYfEVgIiOYO6kFedlz/+Y7Jh6cKLmbqBmFBqdvoT
6he1gHSgFZrNCNhBNz6Hi7xd68Bbnb6bvgpdqr2W5eUQeCRdJ4JUBVYEi2nzgISy
2QpS17fZCeq5IV1pvZVE/mmXpSwMkis9uohNnw16k73Duiz9YwHtKTwxYgvY1GoC
YJjlwFvA1hVKx2wQx2r8+aodfHrrofRy+8WCNYH8UST7J0+1m8mcL4RqV+9pNowM
RxBKkFbP9OS7Elzjs9n9tr+bfcdhLDpveZ4sVtiy0bgH9BdUAwCXWZz8zbf4bdYe
mv8KJwCtXPS4Mi1huNcXwKUgBENMrxmwyQC8G/mYJW0hBeU1hxCWZ5pkLiTyw0qC
Kmv0uK/Rkptmz+n4ResLQrhl9xVz8tu5CNSNCDVhD6Eak6tWJBFUNjHhpc9D3w1Z
ytAt/NXM+Pwn953B5axZ19aJUYzE70NK8TQPfLvu0qoVvOqLkNfZAKzZdD6tsmpE
XHpuc22e5YI2JycXN9GuYdDOQxjBnwRZpwnapQtFQ/oj1OpOX6BROsbSZ/GY0cjs
N7AuSfIsO3qedbGiKySjjH73U3kYme6mD2Acbwf8g80XyA9WGoAxWO5zJxb4OKK6
1zgcqLrWnhdZgVm4bi/G9qCwaMO1Y+Uvf+PzqHqvZlqjylgMPOEFvXT3HETRRcg2
os0VGh9WJnz9/l6MVa8JkKP74To5JL5pQXJ74Mr/w4I5rDF2OhOfMyOBDRj+iykX
r9ho+kYWgwFSz31rDcA7MY69F1GWyrUr/byKF5qktXuMaRIdMfl6UFZ/M6OWhYPt
6osi+5rYvyYUXqlb+qwXY+AAxmcBYPsClICA0xTXKn+LrVT5aHJ9qHGyRKHGUus/
hAd6DbCKaPx//6MjxNisFu8SkKXxvOxE+WK6xA0PFze/OnlO4M/8f6rT/SFc8ptg
txw9xRLGhfxrPcOMTaXPAHOUfKCwN2CqsiKkl208OnmteBjPzscRCNva+PZ+Ybg9
lXrAPzzmTf14i6uniq9YEHDmWWvIbibUGsrsqP2nT8NWszn2SBZG9nZ7elscXkWf
p/NGJCoX4lIw5heaNFO29fxWfQ4vuf2bkR3O43pAKHG0Fgk1HPgf+rIlSk3ISviQ
5wxsKWxafXM/6mMIBHv9HcO74RXXcJSjPhqgU9sG0ngjt96oyzyhdFuZuKwlMCzW
Gll4YAMEoAfnrpzv6yXggtf+VU0NYyZCTOCEWb1DdlkZMI0gXdrw+sUPlXuWr6a6
4Rsb+BUsK3vGL4p4Kw0lBCSCDC1YBo8CbCM4PB0nxo6ZAMZ4lDtsYKJQ/vg07/it
Bi/voosVWLpn/LB35OUBTzGI/gOWI39+IA0kNg7VDXtWu4f3G1awk/dPQ5BiZj15
Rlml9/dlmv+fuJx4N1JNKyk6y8AWubmiHfTV4IJghAUYi5FjpTcm28jviwWKdwJu
hJEKne7lfmX2blPeoZoZo0N18VtzcNdediAWeHf5BduZMZGo7NXjkN11h/6Jv9hq
hzDGrCZ6Y2beDS++WuqVFbk7Unb57EZNKCOQZwL+F5eylZj5oQtioNAhq8Aw3bKB
rhjo+BmvZZlspy8nL4PXSMKU66hmttc5IKIrjrNBRGu1SRrD6GDcMfS/mtX1Dg0N
G7N7EJs4bGN/WQ5NC2z8o7Y+LaGSawxS+GgrC7Zm8JxW5cTIDMINfZa2mF12nr/Y
I0EjGRPqJK58BkFn5DtugM8TS8TCf4sBJ171V9f23UhLfXBJ8o6hDE8jTHzHQ6o6
rLH0zaP88HThhsTOxsPfV8k3SYr9olnoOuKuOmhd2+rjCS5ieBtHaA/6KMk7EZpo
9bT/EZy/odroSAmtx5yKGdGRIt00SkeAodzn2Cj4L6iTv1PLexu6emJOd3LRGMYY
mynRt4I4F2/k1CvQ6OMpOf2jbLYfU8q0xYogNrF2kgJAftSaP3Nci8kheVjIZpNO
z7XYQQvYeH0rTH2UbqSe7ha+/lB2YMpMgvjqwXXREPmnQV3CSDcaWdJEjSAWJEHa
0Or0gQbDCxNsnMHfvYLmLTonMaJIy6UDonBxPMXNXUU7pe2qhwiRsEbC4U2HBabF
ptONWD+Yxf6oFZPnsqwIRh1DwazmS5u8yiBz7sfbaI6oqejLQLf6MnEJKttGy8Xr
ck2Qmwh1XDniUZgqnHsHTaB5OuFjM+4B6TluDcQKxm+31dMusO3AFUEDL7pU7s3B
umdMyNrSZpSU6+a+jEIVAU4pDUN/JLGf1xqZ5chovtawSgMB3VLZZETr3hyK7m5d
5dk7vLbBp78P1WfWnkS70sgdqtKa4q5ILrhUn/gRA3G9aQOhTYkIlH6v/XRKVZXB
k+R0ZWNqqUEa/tm++voXjiFAFmOzx6gEQQZxRWSrUTAqVYGRWZ90RrwYvpxQNgMx
Knh+XOgcVsO/khSniVQZeFgclN2+uzCbBPga/FY3Fc9tYUEH/QXicD3Sln+RZYSZ
UnQxW4q5cfohRio6UWLqiocn4SLuGR2PBn/zxmX1cNdx//H/uXjVA1DXEDr4dj0H
UychEujYi6SUx609aoOzKD+HLnIZEngGcJRy2xKTz7zWehrdmnFjLHzoAU401zm9
dcN3slZnAvLxBTY8ein5apf+H0Asn95GN7K+MMvLjbmKPBk6oeO2HEALJGV89NG9
cKSIkTQhRy1mp9Z8wCGn0FhOf90R+18HwaPYQM+elSTjGGMMzzOyhp7NSyJ3Bct7
8FoDc3oDzgry2kEBoJyhL92cqi7mA86LCRSh/eqKaVbgb9+bTioD5sghqicr4uoj
QcltGfmb3Jl5higyXNM+sZZt7TE6gdUyG5l3RSd1m8hy409wk5QfOYuA9ghERWb6
/VU+YSf73ILT5JaAslLnpqUYQpYpVV2vS9gAkM5PmEOaHE+h6ourQjpQrSlvzTK/
eh26Yyrs08fiCd9GLLOVcdFIqwBJjCRulUVaDdAwZQ5wIK4f20CYSmglmRVEL40U
P31DrND9HpMYHtNVMyxJTvmu61npiNOreZO8q/aEonpOIyVJDFWE4ijNusWq9sYh
OWVOtAxbFvIlFvRdpi15yq+UIhORpK86V1c65chedv11OOkZkn7CpMvmeyITz3FJ
coYebCD+qDHgWm+nOwh5l/KCK5/CCHoR/lXzZ+f7ktVrA7gxXrunXub+ZTKSfHw9
DoLnYm5j5+vNAi48/QuY0lsNxoK8FheAUumAXlL1KHOkgfDe4OyJim4SS8uuNlZI
SzdI3dz+g2NV6yIO9C2RMepB+fMSSllLL9LbqJPGwG35RwcoVbjmPWFnYtJaS9m9
aHeu2Z+yfq28KQUr8soOyoudD1q+a+UOuDIKj6V5Ek/7j4CeIqB7V0+DaMrfCQM2
77vmaMst5ZQcXtzH16Y2HLEmNWnKUWXqw9IcdDHnjkkv7B7T15zOYB1ALjDScjGw
ldjd0fEF/MUQY3l+V0nacqSNF46kLxqLYNmshjsh1ShD8gHQs+gX/IW7Y1eJNzHz
fprpqPPhClX64v5/XCx9vQ/mDXUw5eHyW12Jhj+jDBx0Q37kZ2IbYFeqcmfr1Py5
cFEQvCWfZGLfbMlamEpsyTbqUkNdV6V2xzI10ffiI9sRkZqSnip30L6X0V1N1me6
AVQqp0zIBNQnLbT9qTy4qaNs6lZ8pLHkqZGdBGSkhCvgj1eqbsTsJE7VK9CcKt5G
u9jl+ZENwFIzb2yeult5lroOTQi21cLeYwtWq6kjSNF8zw8w0EbSZ27pCo/bF/xN
4eTWIl0nx+rxbSGJm54ZYWn1n8vFaLX5z59NlcH6chUDN8okBUzP1KqCaOn43B1p
8XMa9q1ykRQDPLlyZWqpF+EBKisEy0bLhDHAMESXEG6I/3eukrBraDwFEn2vdREt
4Kgv5Yw5+aJ0wumL0lPv1F+qCRyTyfBW3dFQhzg/nsX+vj9HT3P9zMKORTqM69Ui
//pragma protect end_data_block
//pragma protect digest_block
Ri+Doz6n1XaCuMehRH2Qu1sDlMo=
//pragma protect end_digest_block
//pragma protect end_protected
