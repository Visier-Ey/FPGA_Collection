-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
oQi+4hoqFzLj+FCVA4sVClj6g9WnITwV2bjf4Msrofs9n1o2Av4N0UFLX9Uk1mO4IDH/DmnMK7dk
4JaeJqMBY/xtC2mdElOuhbn3sEXm8EXut5LAkt4QThteSDJNTqje5xb+ljyl6uD7o3uOS56nS8h7
FvFetKnpaqxs6hTPOSx9aILCV6u2Z37i9GJc2SnX+eQ3iKl6Kj9vbPYYeGq14O1zfBB2/poNpoIY
m7xp1QKIG3sVBL5XImGX1/kAKQ+pto4QfThC42RQ+9cZKkBT8X8XoXBvCOUGool4upwe2UXZYyhz
zCx023JOT94G7184SRWncpHiAbWlb47wiG+wiA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10048)
`protect data_block
trRrRIRDLCe8PR2fh1oHKUrN8kG76G1jm+Q6HClT+zzlKgPx1gv34XYJe9neX+p6ePGV8K6xaUnX
yv4/HNsk2qHDx1N3g/m+JFI3RXtrcas1BqOmzS13tCjpv/WR1+xA40Kvdsu9bN3lkj2jKaBIHZVm
9rv1ECGlQ6wHlVRVHCXA8FBsLo1Ie+idd7+RwfPTSrAGasZ1O8Tez/xKgmC9hrumYUQlxqpOVdUw
p4GhbPS2IctZ/kll7flIuSBsClT45A7HHr2OkkA73tmTBY8Me2+GorYX9tAGxmt3YhCF2dzdr+b2
n85cfMk6KyV4CcPSjCMthyTYhc4Zu8MliEfukj1wLo8hYSssBURKGpftfGkYPeE94ko13t80hH+1
cLhHRiKjoh+x+lcLsMnWpna0VMNGIY2ALrnBAc6Rp+HDlGGwAgUaCguygmwMEKPhaPpCHchjGYwa
DDXtOorVEczae0TOyBFMowwWTyjDe9mdWFDLwUWU3g4ZaBTjaNFduyeZwLXFAvrCKsYSz3pE80Kn
e2Qz+5ikVTashuZMqADB3CVmyjgoZ5j7fUsYgkkbGnlIzLHnkJ7V5ntHQpQXz2rgD/AJnVFgK0vz
IK224ScOrTI8pMeOi59A7z+Ry89YMlhc3EH0C4FBbpo70SlgBYx9rlyBd1xo/vvC3iKocllHs3S/
NOvACVm/AV1UxSpctXHNj+MtXmxC64Zm2gPtr9djQnvZDaTRTQzGVUehDKuQXQh5XAfDO9UstkiD
4eDWBbw4Id1FNi4cUYcRPDfSevVH5Tb++Oktc0cljOaGUgVdetOLbJTkL5/1d1yPOEe14Pnht9sA
J6N3UyIzQ+KTSBZu7T/LLwPHHnoC0kTsz6gYrdJjuRJzJA4HY2Gj+GJfxAJlZRTK7lzJHSfHh8AI
1kDWx+vVSAxr7eIkAcInGBqspyM/MM9B+QLLl3f4RTu4cdDq9B0RX9yC2wM0Csl02H+pS+/VUUhB
/l8MByK0WTwDFj08SMwrzfJbpMONBL1/GOwlutIQmK+ZKLiKfA63ViPEzRLoV7gYzBclmcPEpX8S
dGJ7QteKNWDlLhQfxLlSQ5bWXZqtY4PFUPoP9QhDgu5g4f96eSv8Tiiu9MfpJDKjmtpGrgZM56o9
lAGzdmIIIDMMRq5+LcpS7Q4WubaBljO/29RfyrbPo7Nn2vgHiUlQs3i2jopSQLzosQKvvP1UeuzY
F5tEwOUcJjNS8MJ59YJuO2tYvtWyPytUhUNQS0FeN3yxv8PzoSQzR04L+DPlE60prtE2K4F2yGAC
22jkVsAZne7aaFfxrfpSS4S14J72RpU2yZSqab6n2YBoVydAkJQH7cb8U8pCjepqEL/n8mfRnZcG
78yui8AlYEX1xoKzesqIkHHoQHNP9iZAm4qAK+ivCIdCs1JUyQGrOFkMkgoUsw/x6ABLb33SijfG
il/z3l2VwJfhON2bnBi75GpTqG4caZmTaET4D7rh2fWTLxK0NUv51ubGNf53ITrQzqD+wcrSUdF+
wB48ViVK2xZMXe0ZNfOUSNiruFrfGzJEeshoJdHIY+5+JDuwjPGBNdlsEddik8UoC9WxATc/v0xN
Vh49a0A3VWk/iIvDAxfX96ZpePZgjhYvO4/WZkO6uuKFlfApQaRTBa4+rMvcde001h9+lvM/gTgb
91s+DLxlp1CK4UuJbhipo+X48yXlUNcC37CftL9amaIxm2Qe6vlC6FD5fgfZci628xWLTnyJQHpL
VbJi3UMERcoteBwytGsnK5PEXqQa98GCO1Bh/CK4xZ2pX28JgdCnndjOmBacI6WWRlT11bp4PwtH
Pxkyrd+TrfubEBl07U4jtP9Nfe4eH1kjs4jrwqddYaP5667bn3faB09pLrbvBDd1IcfHUSI6+5TE
ItNHV8EbWodpE0sqmGrIB+SVghAcY1ORF1ZHzCcrclWIHuXCcJMwisrGytQvDx/sqN2hdnW/H1q5
R+6WPBkNw7A5CIGl61puPlH+m30XQtgPPWRJYQHeLwbd3rn7o9zQLJYoi4Xri4OjQzvS0T+oS8Xd
9L9r87G4ysE+LudO9q9LHrNSF/FUQHqTmTyVu3W5nIvGJmEOPTYU0sm0LBxErC0WAd1IbRwM3KZM
Z/VHP7LlpRFqTp56qh0x/eB/oJ0ZdwUZ/bPm8nGioT91Fkuo2zew8faeK0COyoHLLnOC/ulYT+iS
1Lz0F8BUV5SqhIEWG0RkH3QcVKb0cGcvY6dzXqwcY4dZPnXWg24dq8/Ed/nCz8rVlRgG0rxsZWV0
rBpKoIFwapILILZao7Zf8ySXRSGFGeM8+bLgl7VywbzzdsIhLz7deZBHNJAH+RZsmVjFtzYbH947
T4cGplncQCKGci58Wzz2pZTQLkki35dbblL/fhD4vG1RPSyST1ltJxN6kGeeXsvUneyGjW6IYMSf
eEH3uQ48ARWcxF90oWISl27WYj0JxyrdeJxinhJA7WF/nqTG4NlfUpP5l67MbdWmSy/rQuvRVJXW
OJIZ7s1in9zrfwa6bwOHf2CrzBIQy2pSSNEVkkRGhz+K8OvO7ff9j+DoIrP4qttcJ00AqvGpShNG
t/bgMwOuuqZk5S3TaEx0MLkmpFjIREQwfiht1hRoD+ijIUAiPPamIC7lhHdbahui54DCeF32OcDb
ArOS6h0kcAAShnFB+ZipM8SAQPDo5pmVb+O3gDKdKaEDujcuIeecf06Gry2dgFU4H+QyttumdKGE
H3tFrYvaaYYp6jhnjZMdiYj9xYozvvz7+icWqeeH5xjm9keaQem/TfnUf5pZ82UegTyzHTzCaQzx
/t6c9cNQpQ4gkPLCCgQS8mfhB5Z1ej9GxjbZ9NQxITVQ4bB6EJhkdk48fb+N4zBzcuy/M9D+LTzp
sW0vwm5blUM2Jcotkx+hGooQbtOjrbIbN40vRKb08cPdlTggmsb8jFoULHYm/y5jZWeGW4mlHCen
NAn2rCfgQIaIKwGc56cZ1EnBTfpF+LqaBOICRP+xNJ0NYo9aEY4kyiWS7XEl/srA9ZCI2Z1mBaEl
zo/CzMEypMGIYciom+zZ7pMhFcv76n3MzBexQUt5r/K2KtppnMwHf4ekUcBIoJhFs/2iBo+8xOKF
tn1ggoCpSmqfdTTBxTbe2nZhRmw9olQ9aE7/OKabU3XrWxhkkL4gOQHGVtZTK1GJ/3sKE9hzQPil
s2AECh4aECuGfNq3sAD+P/UOlObk72DPi4Tsw91x6wAntVbCKaHJr3jckMnUmZHlB1J2HucSlZNY
28nwG67oJmBrLqUHkbackhdWJUevLk4/s2IgpVXUla9tFRCtvkpusJw/Fz1lK4NzVrpYKroPpF6/
FVVKXcYpHfUfmQ57ekHSSaXaahGtx+WMykbIjrgDjqQ/zpX/4bTYLHGBWjB2vdW9vNqCaBvwDNim
ixCoidydehRPWOdEkXuepvxV+UrBlz9+7iIDDthv3zVUWj3UAoMF28XPZPGl7NDYKGXi7sqytz+4
glamKIVdY6JDnwK2FIWL9HeVc4/s8JVfMv4EVXqTIiaUX7D3hCKo0r0Zknlg9ajTPyyKITaUDIU4
opRQeSKegJIDGHvpALxCV3uWoYQ7EEHi08P6PmL2bDKJhWLkQeTOtZ0cxOcX692Cvu2uRVyjWSxj
aJ5HkSID013DgrFV8vS4RqeKGeo20tQFq6dThLRehOKXPuf69CKFLckFMoz1MF61po+RDUHQXkKS
NgoMOvQR1SgFpgwyNJVYAExQXd4Ku5Cu8/g2AFPF1McV95bm+qojdtX9j2w+qzJcaNINuhy1aeyK
LK94bm4QL4cGhzz3VHEBbBv0RWiM/KlE9OeiPPuVh5i5+R3fEekpHgBbKMZjCqTIKXNPtLP8N/gj
6WAKwCMkzbsG8/5Wy+XFckFRroX5rnx1AndSKvsTZ+0vmT6jSJd0Nt32NLB/4clinLmAApWFePdr
9Ht7gbg6bxZoqojHZyPVSZngfB4eUmgABv9hGxi6uFDRc+TK/EJqQBa+YczpAQU3jJpbHU33Wxo4
AijHHTGlmU7P3ov+dS+q6+7IA/ZGIC7+mYJF6wriwQdYWPNNnQLe57GcMR4P8v9LYyt0aG6wor0v
9N8wtCskzkzE3vKKgI1+G4ilfOV80lpbLp7oWUwINXIiXLYGdnTi6WWwrM8WWCf9hPpedq0hOVK2
FabxF3nqyi3LQf/mga7ywf5m8tnggnrk6kJj6ybYTArFTsaSZKCUPnrr0mvx/+X8svPNNxldDPOk
Z+XTbbuiavKrkk16KkVmvydeSFThH8NoQlvdUgW+CTMDwxpHQb6mXmk8rU3lNMTNcYmzIdCLzwsH
+ldEb7PPjv9YJ4DJFG24hpKgT6vjH/V0gQyOEcMIOzNKG/yT15ssVE2JsbFY/QAmurK/p97qELBS
GMpJnyYR7NNYQXq6vtpKwed+p6qyMBpiq/HdJrktuN6cPCg240BUnchzTiSNv0PIYy1xOlNVJQcI
D36Rpqr1KPLRH/Uv3TmslRKFuRMj/pu/6ECJdm1sCc0t82Atd1Srcos+Xuqee3mAxDTb9S/1whm7
+UuRaVYlME3k4321jerv1gH0cc/KNfd8aPF+d4KuxPJN19rqcrYu822jHbSQeMJVg9gugQ37NMoV
9c7MGrfbBAW5GxDuJVur31uTTN6dqGBHFglghqEL2WLUzx61W6+yw4ygCoKI4NwE9GJEXahkV/mI
LlULTACSEEQiCcoWoOKCNkO8BsoY5i9MoNhc3bUhNCvMbtpLR0pi45gtZwK18b3UpDW9wKBeLxJP
ddwqDqw/bDZwFDxuIvxRGW/v6cw2OYDXI8xTt4NiJPDeMNnXvLZ6Ebt4gL6hH6ZYcOBB8FK6Sz/6
2bEZT0OfYtufO/WO0ddop/8Z2ENXtIJSCTv7QVsxwLbd9Yh2n4VRv4sAKli2XM1flrXjkvhfsshW
oydHN3m0twww45AXdxcMCIH2L3bZd/JDyFvIWJ59udr14p1f4PtE8+YQ9PCdwNoKdtwQQ5kqnZ7X
ze8TbV8BnJY+/ZZhUVdriG5+5sIXQh/ggxG9bFxoWlKBIcUlt0LT5dwIb2Hll7KJ+UA0qV4wy6PF
S81c/Y1AzSNop1bB1MGkW9Xl72DM6VuT1E4miKdAMved/ZjittAQ0AepDeXrRnw5ekVuWuBrX5sX
X/j39EGgdjbnuJMV9qpJCIJ+SFtPrvR5CWP4ZFLw0xLBRrKNXL644V7gLKBD//5bLcuvPSnv1T+C
Zyl6UjrFq2jHP4RJcQaDAqDmphdzAmNaRDnJtDuIfUzFuZdiL8NCLlHtm9XNEK13hZPrJQIkSOIs
fc1yFo84du7fl6ZpeVq8a8PTo3cdMTxLFREqEtJRtSl6zsrLbJIUvKhSOP5fe0eE3vQbn04wGKr5
tUB7c73n+tBssOcYrUCGL8bGw3t0JMRZSTzcJBB7yHGYf3vfbSJLM04n1AZzvyUWNIZWRgBuDEcG
OotfXnIc3DKIQ3wXXRbFjSQslUScebvu9rXO4PtUScCbgyBp8DsyJisJRi86nbLdoy6enfNCoZAX
5t4yCbTtu8/HaSRHCy6m1pMK6oqqgtqRdczYd6HW0TbNzQFKOeerjHrnP8NQ28pDSWZZm3SFeYUA
cQStjX9chUbtLc0BIUyYXkyb5TB7sL1mGVhBfGgLmC40O23CVCQc0+UNGscJeyb9o8S/DTt93XRJ
OzzzPhqTZcZAk7e1B/V8SQidLDjg6bBKsSF0HdN5ok/E9RV8TbNLXOaP17xrisdBuFPqZ2dqsbrt
m9l8fPYllzJR5CPy3/ulH0JFJFjznNzzXDf0X7wgABc8gNkTRdAE8aVopYkAWbI0POqYoR/yVLCI
Zgh1Zjq2VoNCs2rPtPr3d3XYs+ZHlGUL/QxmIHKjHouIHuHKklAuQWP/kJBcHH5i6SfcRzZXYd2N
vYj6jYNz89NLTlhHMym2rCAJ/ed4pzYv6VYL2FWuVpItL8A8YxuQthtVwhJZEoSyxjqk575SKBuC
MzYK4z0ehGSUjJ63y9cIzVv22S8wJDQ5vz81g5Pcj1b5vNbeO/S2hEzFOmJMePTAdKo3eZ/feIVM
W4mBkX8dHmICS8iIT6x6OSviYnyrX2nsJtEKjbch4f/i6TBfGMqOuNuqFT5RcR8fiLpl8yDsu7q+
9y0doifJmGk5sXxDpgy3q+JGW6glXY5bsTN7pAwuoseSHtfcs2eEiRAGlOxJveTSsq19yJzRd1kS
RG02Pzko0tIZxKg7XmQRTC6uO6dFW6XrGMnBAsGcumMLt5/yAwjxhNeZY7IlYgTx147tAyAOQqbf
2U8LfhhKdtF8NgICmt+l2t/bP4yY29hlTOGKpWwNOd3T+prnPmRtWnOvSjNWM1Bwx+pb+CXOAcGH
mKbGevtZiIVzMtwLw0en39EmyiUOPkhB5xKegnc9eCo9dci++0HgQsdPg0o9avhIllvXZzbq+TYz
n72Orw+0R7xp4+Mccj2Ipov8WZUo6CwOQsj929dWip41VXwR3l0vzKbUqzRJ0v94bAElaH/zuVEU
CBCeRNLxgZ6dCc6i3oZC1uLL0FOarYuiWf9HsF/o2IAoeCGSM/ASsIu+ZCWq8pPc7A6oTw43IKP1
flBF9tswBxn3axDbbmKFZYlAqUo244T5rYq7LV1N8a25VYzki0yhO8hfNghx3I6IlDNBl/B/7Mq3
TDysSTxACROapatoeUtuF1h7lo5ERy+lV8WM35ns9P/jAP4JKA1FAph5NpsktTZd3BIKVekkmglf
H3RqMERnIN5xUbCwrapUjoJz1yRwrtg4+cuCiMZ4Z/w3QFdZ23No7NjGv44P9a08YffE/b6rkCmE
1VseYJLx9cTjGW9L3+67/2MttBitsJLOxBh429OxuKPeiMk3kmsa3ZPC3dw7TxopWuDHDwaWfZdU
xYmmYQQqL83/Y6QhrYxGvEG13r3/oyzWeC2nXJmf4ozsC+5eZNPaFGvsaL3nnTm3cwJ268nOEvYx
tzPLaI36mtqFbEM8T/jWB3rAIfR76rldBQ+LxQuVdsDGp6Qt5ctXmOS92OVih5tElQ1BViGY8EUc
60ZwmjIFkBFdlUqbyQC69qUmi0VLtPNWC/yz5XjT72wMxbZGJKsrKL6okBk0SBWdigYI1L0buixY
qbFlJnFhreRn9zWh4UoLgY13hVVbCuYqqmBVPf050qRekXZ426ngUDCEjzQDlp264YNp49tpBeid
yJHWrlxaPuu0VIghj2wLTTRbx08re8/AwwBT8fP1VkVdiVWYf0b3Lyo0NvAos9UwWMrR15gqkIEm
U2yCnjCKfU5r3t4mZNtVvhHFo1fShI5v2pmNt7GtqMc45+Y13XU93tKOF5AjbUKkjlFUnjghJ2V0
ud0QIeiZTfwo3n6/+MMrpI4N682N359JRZmebBElQXMfLhK4z9LDRZLAcSngBI36n821QiPsOUEt
+9N3D5WEbDUPNUvyXFHk3IHiZiKJ0Mf18nLPjV2B3f+AjKGpN1oOi9tjdmjIcGJX4cjOodXYFl18
dyvZZmNAGgHkDplE5f94PpnO8ewnbuibX1qchzuV3SYAIy7VfGhB55Vp26HFSWnD+ShW3Ft3Atp1
ocoqLSgnlw2kLu7yfvBraFATk1bFgTtSuyK9CBMrAiC6vZ7Q1Y2izwAFf/MiGH79or8Liih90c6n
JKAa2c5lj0S7m5pZgsPUI+t7WVMmlFazHX1not095J3Xq5fm5w820RWkhouP8dHg0FEVETNeFURf
UoScuJQMOLYyGv/m8ZhNja+jrzBLrbFe7ujydOLztAu0UxbQoGz7gjteB1fVakCLduqJrrkicS8L
9btbm1J5NFJNdQuPLRYurFwTaDETSYV1JzR10yuqhhyoQeAzFIT7zmQWORbNbhfdY7RB1aqs9Pla
YSR3H0915bQhUuhtdocwqAXy6Q7ZP3WSrYjyJiM16eozMw2JlzZHcDbTLDWpoqS0/s4JJuY5IhN/
sydRq5gS+nDI2LLOtotFiD/0mYlkVYMQqMT9jbdla5XWs5p6DaZv1cQxP2bPM6JiatdU2LJMK+Yb
h22YiGvhKuqxLycIBJHOAE1NagxYn0BWOcVZT2tJq25CY82PVA2wcNd1ubUB6zEdGPYDn0mzVE2r
uw909M3EN2jmIuL3K18jbxg+Bcj7ZQ7vhMZ0JD4/RnnYUdxTvm3ztIYVSf4t0hErhHS9Fy2ZHG3G
LY5iQ124nR6nLG97/ii/3xiexHAvR8jqO/ZxEhDue4d22iMCpx/NYI2xAMZR2Bf0rOPNM/p1XWmk
3Pcb71XkRzyPg5Qccp6YVzS2AIV2+ImVMc3xmzXqHpRszodY1Fuzllcx2ODaZMN1NEBeyNOxuM7+
ZnASm07zN9rLbB9muyT0ErIovHjXpXyXrII1Jo1Qr5Wa6gwskdRYMHEmFLKikGYvtieArCj3AjHz
Hvxj7ZiFqSryTNFod+wSCnsMt6pTAlBJj81xhUTnDzDYGZIqtObmN1T3Sd5YQ5r445rn888d32ua
TkmeC6nAzO2I2zM+HSTIqf3YEZKHxiBec4YkQ9e05SveXZrvwMcEePCoiTbo5hYleGkBNOIv/oaK
gA9ixThrzs7nnwPVi7EFRSvvxQR4TUnv0m98J5uX6R/f9Nv94lyaCM7lkcgjIYYEnvsKqqdTr7xg
0TEQcVO5s+WgGID5TnrD5fq7VQ+ueN9oIGEplAWsn/UEKLQfMPX3Rnk3zXr3M9OwrnQv3gPx9HLy
r4lCNDFBN8sfzByztFFH8h/4araZ1lq1PDlblyZ0fO/piGRORJpRc0pihck+BT2gVbBMrdwE7xwg
Yr//ZWS0/IKxodEPmg+yW12yI5rejsGc2xV+eYNWOluI54jP+tPdEmFfwd+KInQ8XW/YFXAr/wlk
sdY7a5Y+Pa5K7WRzri3ts9rthFoN0huoZR/IhACJ6pHgbAmpy4Ug0+xsEliVj6ZFliPJLOiNqOpI
NBYBY+i+VLRpHjVLi9PtSvGdIm5XMAEie6063pZMTX+o54RyIsRnMcE9uT76pRwp842ppqNX/UdY
Oz+iaR64M98QKYV1G0wVfsB5o/L3tLAmI3UY/Px12rmWZOP8gh24IvBqPCqag8uiOV7WWUTvKCjN
kLkSI0Vm8QhVejj1wrlarIA1zPW9jT+coqfJKaIo4R6i0h94LYzcDMuB3ZJcwZO2Flkf/gKcAEn6
z4YV0U2LxOt+P2WGnGB+JnlZm8WdSRCkRZtehoIBD8sq//9BvuhJD4dj9fmPp7e5YfBgcQX7kdXv
cmnPwLfLafhFQb6dwoX3QSGV+mjTiqXzFXfTzkoYwx3e1hQ3cyFNTsla1HS3BFUCO2vuTN5+gxM1
Qvp9uaoses8q1Za5vewSvVjQuIUT7XG6u6CuIlmQbbfN2zUOoLRx770HsQP7yHs5QzdNm2kGDiJ1
vwVoCTGy3D45vCwTrkjXBJy4DPBJCCECgpjPAokjdiu0EhT7qKdQr9xv09F6pbqsw5plZGJm/Fxd
q+2Z9ClwGvNM6hGhGdCZAfNvmyEclFkg74Ptx9JU1viCifQDZItm5uR+k2K2KKzuWkVkubrLEMCn
wcn/AE6QnX6Ae1bj4x5eF9RpW/pJxjoSbrSo4YOuAQGQwJgEKnK86BUjIjrvm081FYKwsrkSPWTg
AsMVF24cED7MDqCDM423RucjXUKQdj4qyignLFfyJEcsgFmU8jWCVHO2YXMY3pbWcq3+lOXUjpQo
5GMqSZw1S918UenWic94YCtW4XegRTJNLc0eu4M4Q3j+3RGo+MIasyQLfmlKpTpM2OB3heEjJU5l
BB6rCo1y8WduzVWuGzvj1OoXtXyK0nWop40rVKMKk4gXmYNv5xAH9jzcvFcWrBC1QKUgD8Zo2y1j
6Ylp5zVJbEgKW0hVi5tXOSXjxjNnfjqC/n6ysbfxzGLj8cqOkqYlb/SQi+qxR4diYEBUa2tauF49
oDvNed01GMmBqSv+O6FcyR32YznJZN18xlGiycbbYhhleFkTCkH6XC4xThKsickciqvGkj0VITO6
uXCagI5HeO7PGA+0LOi5nQmeSG5RYkM/bsSaWD9jUL9fYRZ8lzo39QcrxJ9EOLUYW9qoX4jNxSzD
Eed1RzXVSF1fvHxmlpmogkH8la3h8A+HzpOhPoA5BPT7dksp065d7h24uS/3N+LwyPiG5TKaQBVU
+diVaTzaKZhic2mQN8poovdXAqu8nbek17pT4qEvM9rJCSRHXvWQIkioIyw/23xa6eyhrbYeY4yV
sLo0tnTkIpHNM3ZwL0s0mdVCPDM/HBvqcCQOJ8qwihT56F3FNjmhJ12U46Fwkk5jO9kpAMjmLnKo
OAg2otf3UjyIM6XpxW0zTRzc2aMbHZu5B150Z7S49Gp9ky+Jkr6IC0uRmstNcj/nQTbCh/Zo7JRZ
/c2cBPWOUyuTUMhE/Saiq6LKu4AdwvQotgivXKxMY/TuaqVPpgrpz/54L/sMmRMqn29VPcgWW11p
znm2DegF/2IeJMyNEMlTtLsyHEc3IXiXeNCFsmUoPSx92O0pQ3QPjYKad6z1odoXwXjh+OnTCxW0
SZVfoXzk1XkffODeWKKRA5n+nLKoH6XLIGeAJcJupJZJ/IrNtyCth+PkH+tDqiH+J47CvyWsDt1o
98vyImEWnBVjmHSotbmpB2Gwi6b+0RA8gBxT6ik9jtxEnARHLelggmfhZ4e5AJYxdhYbfW7yUooK
PZs1/l7xnq3kwHGA3BDReYzXtJvuzssB/Nh/e3efkofZ1CVXs7YB8ZB1tb8bgNU0MuDac3/pHCvn
rPJWRlrnlj39d+0xm1PctKIFx9TlnmY+2jktT7qrnyLo/hG5WHof6wjDtolFbSYnymXr7S8dOYhD
dZC9IXp01ZzWXkJUbxNaeKmIGrr+v9olOTSX6X6cUlW5pndPxLkp86mOCq8nvD6YGemqC57J1zcL
4gO8nA0hZ88zaYJzdiNm8Gxp2GBhvUis2DoM+xOXBFShRx8k8mqJR75qLL8jljch/OAE2iRbeoyQ
bgDVFwHCjYfJp8IQQC/++5l8pIJ9PPdGkkoKfSW6etGkORItIuadKWqcFzpDauARzjC/lEUtasLj
kTKo1bMD2hV8yYG0RUtBkgsCPOBbwT53Hn3eyuXjxoEm4bBJMmXKdUaQHM6jNYRpKeHxbPw3E9Wy
FAwKCwvQnX1hDXOi/hM1ZAw9f6mPllIE2cysHw7eFb9rARxuh+PvJXIVrzL051vQsEnMbwsrI95Z
l5TR1mzxNlhvJ8WR8i79NTrK0FHqthUXsbg21jv12blmCU95dIE3rvVR/IRusC2NC6mmCqoFoG2K
//D1psSpJrwrRvqbW6o2QAJ/vt8GkMufzdy/oWWHuu6bydp9Moa7IGHVUX2JFtGjtJlj6OdBWk8t
Eoap1864Kr51IoGzvYq4+LPUTWtUqdYH1MswV33hgjhKmqlG498cTXkipBXwrTU8QLsZpgA3zPqO
5xU+hHCwMHyZIGNTrayuRr85eiQqt640Q7A0smwKvSQ3MG7v4y7/vLBYGpkNr8nVHN4wYoYYVazE
ySgdk5qUZ/FE1r5C2+jXfndQg0RH1YKI8xLuIjbeAz4z1H9I1lya93/HfFVsdHXy/LUncDqzbzJB
MkGmeQ94xtu6VeFegYWAuUaVmtVmZYPBfXJxMxNDtyaeli7VoQV053k5E4FefSCDwVtdPDxP5qr6
K8Slx5xr3hCwTTQwkPeVxa73AzcrT+bsHnChrrVFGjwOIb0gzAfSJcKyTfCzyX1m08q6aHGqiJEY
0rS25c69EAKauGjBqc5zslSAUWYQv9SaX2i3ppIEqR9W4mBmGu9UYvIj3KqiiT4G6KP7FFxyPX42
CTf/1OKzSpuflRCYhzfhI9O6udAxTq+Ip+iSZj4nBJBjyB4Bp7eyK7t/I9vT6nIkytdRL11RLuzq
4oZYlezrF9pDYGgGX3MyiKR14S6cOqKE2rb2J5fo9fm3r/Z0SGXShYfsbWBJ/IeT7mrkmF41bSCd
O7g44fSeJOYA1E/pZYLMrXfW8svD6Gywbp7dFm1pBCQjxTBSXf/Ur7ddM8cSYb/eLL48R7NmTOHW
Zrn7P5scujQelG33U+0iM/vwU2gCkZ+PaPViK8s1V1e/iEDSoOeXyrgoBxGg23ZYbRQpW5Oy29Fg
SPcVtX+gLM49KEH3N+P70qFHnOYxhi2wrDaPmbxxn4VIP/8mkE+rPWuAg4eKc3TO96+SwQFQbSjJ
6026G9X+Vrt1Sl/jcjNUBqGGw4ltFaiUN0DzORUQDy76kI4KvTBP4S4+OMb3XnGeBnVkbEQDVG6k
iZmcJqRT2SVzj9tHvYAS9/srgRRgSLCXooPf7pkYIGjUMws00ZFz+UrJDy86l0lZ4dUfl/H5bEQC
gMuLMcuY9OGc6JcO9Q1e7QrlrloaCGuKXbBxFYMHR/Vjb9piyN8ulqxLyRml9cP/e01LYYkEapiB
DHwRjfkAlCEuK7RG8bsix6sDYssNLKzHlmtJe+95ladRIi81NWcAazzFZemSjs92EeroTB3QOj/W
GqcDMkxfifkivh3tMYUgU+Cq95z2I7S7V0ndmkB5z0wF4vonSjvbwV8zCRMEHctr1eh46OUVsFjp
2g2RjooD9oclZAhrP6d1poEo65qoQe8h3FMLtGPKN5R20YtGvxc3tJp1DYbnf+zFXe9xvnjLW2PI
5UB2M8uHdfK+W1vaYUVJH93pfybOJW69qHmiTltx18T3RSl1rlV/MYh1qRC5kajbDQKiDc9U6Qbx
LTOTJy47ALOASlLnKF7lxCGO8uyjA9bwQfUSLbVjP+A7mbYmAUEI4Dm5l8wllMYjl2Gdup6xucWZ
9tknOaYgbm4X2yZejFTGiKz97bDX2jfaPklM3QwQEQB3wRpEgn4CQtfeLSotBq4fiYnCiZMz77sC
RPXJ/ovBTNhQyvse5a4FDul77qSvgHkZVAqwmROcP8skB5TGo08cAehoUgG5U4KK7/URj97kluRj
A0XMFAEXQNv28L7CuUd42e84Ot3xDUTSmmJ7q6ymqppx6YbwAqnoxi6Qh5PPzB8vPlIskOwATg6K
kCaBpgQ7/L/7MaEn3bUMS8AHshaV9xQ1iAACv2oixmggHmMXyVs4JhVMib7tgpdmol7s3vU8kBHL
DfT69pT7FsDxuJG0vaS7DF/QoDCwykKgw+p0f7/mUO0v29LP/zvlPalWs/qGyqwK2BV6PvDix3OF
vwf0Zhb/NCsMquGchkfl9DvJw3hY3dd/DGYedc24nLb+tpdcGycGqfESIJqDy6IzI8pj+jD3j1GD
Tb0GZC50tWAlLAAQvelK9lhumgfP0Q9nEl4MaFY6LlQ1F/Wn7oPVoJiCnlJ3B74gqunmmVrT3e8H
Vu37E7k7VdaUP2KwVJyo9Q==
`protect end_protected
