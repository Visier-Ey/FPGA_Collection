-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "N-2017.12-SP2-4 -- Oct 23, 2018"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
pB/8ajgU1gjHgxZuT1eEMHKM8YPNb/Z4+UxbLPTDvJtGhux2imZHnhlxSIptmp4p
4d1MOpMiVcK3QoZzEl1E5jvMU6Wc6g6R6wRI4fCPKXyCZnIbq5k0hw0vs4bTsnCI
43Kn12JpEPiEm4wMNIU+axSU2JRuCNWxIMB8uC1v1d0=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 6336)
`protect data_block
/B30z6q9rquZetl58IB6GfHyCvqmHar7cyL7oPHjn41auHOvqTp3KfQajCONnxIp
U/CX+RSuIjKJ/6obls9L/ZEqCCfRpCaBN7qEb5VzOAZNtXig+aBj4Gs2ONkD0Pas
aVNxKcPucLDO6KBWs68YhqNgoSoHa+dXDOxMmS94lODGJgwLZkNW6Diq61VWwKf/
b3vVK6WUfKznaHpFCH46XNHu1LfJJolT9B1s887yJYNHWpsfpO+vafjEeEi4cmlS
T16cC+Ta6Kg2FjkxRv/2bTAeQmATlXdSuRA6BPNh+BKUrWDl9IX2ocrZvQmheyLD
MzzPunnO4HbgrVY0zCjnTbIz9RJVb66dybp/80fcSEzYpx8yTW2/Hrnqe254j4rp
YhhFeRMS+b4d4JaZis6fkJkg52EeVZwB8rgdxveKzEtUoDLbjy1ENp/cqg/wSCps
o2I4ET/y7He2yqN3B9ky7r2eiMXk/G4P01sRILr43Dd3U7ZXEGyyliFTOV4ryr2K
JqCNhGChOgs7dANObAmt4DnRhK513iE8GQVOhhPVOoV6VbKctS0ZrzsKMEw9wLK1
8kq8AAxCcgxX3nCOJX4ojNyqhCcB6xa63DziLaeYMwKEFeSPlC2GS42ScsmmhZig
z1/+VzSZpmGw2ZZqEW1ZGGRIizRd3XIpK07DuMW4f63YYnn+Rb/D19C/S7AWB0eq
vQjDKtxQip/omHu3xSro+rWqRovgsY3lR0BCfCrW/WVmBGnYaWCgilVY6yD1VEx7
1dunSE8CPdPwTqcuFfuq5TDXfTvU0+Z5WfJLWOQkdayGLU3J66z44vo7qy63/dLo
JfTCk2CO4Lq012vjZ0QLWwpE9eZ80UmSbTsisoJBYvBW//Up6DlF+yIcUaDWM4J3
8SKQm4+NTiEBUYG0PhwOVP18zSzcQLiTEdOMQ1lwFGUC6mUOciNyJfS7NlRXa26e
0YU9FksrkGXetDHhrKihAWn2/qqvdezFEzzm2Q1IcMQ6GCrOYPk8MjPaiadgiqf2
WrTmDdP03D+3X+qtKTkbzwzC/egtRczDBn2lCiBg1mrXnYf/Ty4wXFwnTPHI7mDN
bA8fmG3haRz3kvFwSzwO1jNzoNA8dXcByOCHlAA6laha+kPD66PcojryQBZN7npl
cCIGb4nfKakIhVK65nXq4leiJlEIomDsj6d73GAaZdq2qUbCuI84b/hbXGpuNpAf
He1ziPyvbFugOuSEnv6eAao7Yb7/k4ab0VzdQeRO0EO4jvC956jhO1H7mYeQIO5v
25QGYRtDpd68Sg98u6CeBx0drO+bDtKoIO6Vr29TrqG5MWOxWNTUcZER88lH04be
qLpdSwM4feayCFfG04mGiqWXjDRWTVu1zSDwjYOcrKyR/FHr8oYCeoMbZoYIkU8x
uzNuQ6ZNhI5+xcMcW8vxWWdz3Iofxctl3Q7XEgM5JBxTGljCO7XXVBB8IImK5oav
ziSfQiuNG1TuTOgkMju/SfY1ULvbE5vzLmcTDdl0v+1W9lTaM64FX7vh4wbrTtVx
1naVc+nitQDN0qc1bZVtvPqql033bvSHP4czSzioD4WcwlJQrZIQUkY8JafDcJtz
7p0wfrh4zzVO5eDXIrExxvxQnwc0QARzQ1PnmwjzFoaZnFPqGph5CYxaConaMa0/
1TVZRSjrunjz4pEFVJ0lT8YwvAv+2YxqnQARS6+cSx/LTMbGIgufoz0QvjpN0dSs
Dv81F2UwtkT3OKvNz0cqDfmDtWbQNRvPrw+MWqFMoXMY8XpCE6q36oFBTvXrHYak
B9uXb+iTSfdtmV+sAGcxXhbdse7lr1JxcyKlbVJRL2B+S+XkcPQvBR4EzXJegETF
YuZCLzz5a9RxTYe6/Z7uV5+CJI4VKMBqcvyUjjDwjVFr3qGFY3m8+TxeDqt8uGCD
ajEnFNnDgfxF4SWtA0bazhhmUDJNDmoPnq3VA991XegKW+f/kGGMHNu2Q3kLwZNH
BJFkGA3o6YQVK4DWMfOfknHnVEshwWlp6LyJeS0kKbq5fUmpVP1590RANi5p9iuW
OUeBGUbilbcsIMMgeqapI+hd95RhMDb5QLwYaWwmZSkyG9i37Yq93YTWg0FIwl7U
zqYm7qT8pSV1CXNmIbkl/KgcL5ZRUOjUeDc2w0hH2upyvzd/N1K+qKVfX4tUSKYi
9yufdYl6V75UQqaqWuqZeqGLlvtNt5WnqqmvPuKfpcrQXPFZZFZ9ptluf+lWy3/G
cFiFaqmPH7D8sIoSR5vBmFn74JYW6gtl/7LBIzKAOF0enGgxIjOM4bKPlWVytcxr
dvQVvlvKzx4WYxKJ7QDOOrbQ0fZ1juREpY1U6QjMlOs7O09LQINxDoKwIfvq9vwV
fX9/4XPmfAXQYvymf6BolPztHer2vU5v/bRYJcGFhg3HAtKIq8XP3ed3lsIZ5v4G
XgTXDr7/IRlSN4UBN0Kj0l/AR+EUBCXCkma+cj5poIwTHclYdKy/V/alV/hGtvvU
F1WLkgOvdiGO0U+G+Mq7vLj+CFpVG7saSb6C21egPmiDWl5e/7IW9Hhlb5XleJpE
x0uRf3D2ptASZhWxIO8kIvv+BM+H8YoMqW8KVbzrx+xFfSdNUF3qEc+jAy6xpjN7
dglg/yNqmNasfFHVV39Cg6iZqErYTZBgcfxRw131+VDXL6aMuSHHFH5z1nhKZH/v
KkqVBstymZ1YBM+sgZCOls74WMr2EqHzNMjAh60Nx9E1DwY85BeffzzTn5GchyQD
0ddfwGdHvj7lYo2D6eViKPmx4qk5UEOx3Z2966ir8zHbZMMR6ATDk9FEg0UbmJPR
HoUQG5oUx/ngjemXGV7y1Nxqbi9uk2k74EylADRXY1uAmEE+xQjYIxXurwy5Z0IF
GWtVAM9hweHF/9vXouZQEHUpuPh9pOqP6OInNvo8Mbi76QGR0hBaXHAm9tFY6NQA
qZuzinnlL6j0QscxHZeN15F/twfAcH1MMoCw4BeNOnChlSmtNCl0Hetn7NT+H7i5
Mu9MEG23tiNsaUDG+3sT2ePpjoVFD8+dLvBp6nLO7BjjDJLgqETkypH1RRc/9gfs
e4heJIKdAnpxWJt76WPI/WZPuwZVFbEQvyIaZHLjN+YZk86J7dYARxb0c9JOz0v4
VLqPDAF8bGfoVvu2TGLYFcmQ08a3abZKD/jB0PBYSnrYipc4HomdzEv/X9DzACcs
jAkeWbgeDqG2ynJZSxaFIG+Wg9sIKrw4O1qHStNVFWVwad+0yeb9SDc9LH6aLf2p
3ge55b9jw8gjbe5HO+ZnwRBONWr7r7cPUTyfEUNR0A/DA2sipTlaiJWwhDgc5A0v
hkpKoBF0E5TGikctYshWMgMbP20fTvDMWnqqWmLBzuDRc2wGzBodwRvyL/IjpaH0
RKev6CkSo7MXbneCqYjMV+HCqqLZec5d132V/Y30oYSxoUOqoJb4lDX3IPV7JyId
nI9/fUWLPxypUjgzFTSubZBwsqwD1e6PX2ev37FSGJHxeR0jj83acDBSVn53r83U
wv4wKB/3Zfumw/HKbWrs5/GBJVO1/9mbU2DPr+cggbyj4bUminxY9foHnY820FMz
a/QNec2b+a1X/K3cOIrcxYcOarERDDZkMlGAfJjJgsGsaKUBDNUUW8l0uEP6HP6c
6MRRlU65svWLWsJr7LxFzB1VOkMQjgg5+i7jzzU+lqo5WRxvDKeyH75dkMCs0RF1
tdN1Wz4O4OM2dHK41vfauYGauXFqDg1a/c7r4vCSBM4pRiTZ3YzJ6tPwXQT+K4xv
8rHFdCLkDb8cnIFj+tdsF13wwcukABb0qvpRHWyfoA9HaASvT0XZysK3QCIS3OJH
bHdZb7BRWNla0isUzDwV0TGbpS6pIYFAB5EMo0lgjPmUYAQWCdgVzOzwPKabdXGR
j3/xgOenz8QRUoyqjkSgVNg/WIHhGWhAVgVIlVJssuMg7irVHwkI7f4tiHt8v8h7
5VCWdDKfiO12Okkw5WtjPguv4W1lKf5K5tbKpiOz+N0RdGUUEaH0EH6QhHK0O/Md
lkWtVvvEfIVD+ywLFlTwxMKS2o6cEDh3f4QF3FguMcM49IsWKTdc2kar1J8x3kaP
S2VsGSuAhXQbfu/kLu+oomgzdb/kZc/Czh8ReQx8pO6r/H0sDwCGULE4hg3HC+kS
YoCwfW0VO603IWAZhXOWBfzKS/vD7/8QmlHFny+PugaOCN+Q4Pg6Bx/r5wfaFW2D
qnFuvWUixCquIaEYo+jGbOLGNScUXHa4CK3UBhaR1BYE2IGqQP9+2eOfU11Ap+Ax
Ag59J/ikqNxXIoDkaD5VY7vnvmXKKAM1zRkDfDIBobve49t3yN1Sk/6y0IbK1YIO
GSDjzZlF3+PhKvhxaAYd4pZU25BVMw2Ed6uPXMD0kdDq94fl2uStApTqICptGO8n
n9hq+Q0uEdYyHYX8Jyw5OEUul1uTCfJB87g9XjfnTCWMelNziP+zjieH/QV55aU1
VNbalU2e/9GKueQHx3scM7Dy0IZ1GFc7pWDjsHVUx1apyPlz9IrGzhuvldUeisb+
S9Q4kEcWmILaw2swuEansYBOWtfMXLoryDTzTlBosPSlnK63HlxmxM0d0VFGhEsk
YS2UjVLwfFrUf9I6yNXNBAB6+FqLkAfVIZTECmKttwHBofHaFyyw+uUnKgDvqtaZ
13FUkL1bq0NuK7T/81dcxM4ixMLY8CtmqCIDLr0eA8vMkHX52y6N5KSIKA/QKOfw
7WAPwmTLomJAqOkrW1kxuQfpWnKbl7vKrGFdRspS22s5cNAFfZBkzqE/U+GYYxR4
sUMoVXbhp0+K3d7mEqumfj/N0QNkuGxsHury1Kdw8i4Ij0GXYIOlE8/KdVi3YvDw
Mhzf5TzEaPVtuRF55weWsUgRctqoxK61DWgMHkzoog3eZJyHpnyqGiKhgwbfFbiK
maQ7SAN/wqYWKa2PJFy0H/YqvKlxjI7waJxv8EvwZF9+Si5s9k4M79DdNEqIzRnX
d+MAq6yvFQ37kohSNyDod7PIRdQ809f0gmOfjS9SV2yRi539Tn7G6FJ5ZTwbtCr4
2/Xim1f2jqgdmy/PqmnxxGBDAW9CWa9NmE10eo2FfQbgrjzT4O7GGrWSY1Sqv1ye
tuY9R8/+iuR5qlsz4tPZkYLptBEEu9M9FrYzx1AYvcdYrNuyJx879QMcTjNVslsK
BFhBI035RpShdZ+rBaJmp8nYUgnSbwq03IEyCOMODMi1IFGQFaxHs6jz3t8c119w
507XwfenX7vqBm52JZOKAKlQbVWnVwkqO1P71mfEJAcXBXsLx33LdjAgK8CNQ1nz
5FKmzokBXzjyETBFVxWXG4+cLdq7KkoFfqIMOT4nxwal6Ba5Z0jKht+qcDRq48xk
KTJy8Y/8jWcLHVRTAVkEpwQksccM5F7HZ6k7wHI5Ob5dzLD5oJL2FPryoVFNb5kv
hpeW8D6DelAA67FIDaU1JvG+YD8oDnPT0aNN/7p6+VH1CU7HZN6E/4ixq2DQ8YpK
TBH9CdQksaLTItWOzFYw8Evtur9OFohBA4+s6c6c382Aw6d0RrYQNomwCttqAtCz
+icUWcRpvSFApski1/kwlxfYNDKTWbz9lI8Xc6dWQRyeW+YdbACtC5x5WWJuynWA
OT8/dbqmOzNGqIXI0+dsvs4FRYhV+0EA00vwJLxXNllPkSMGA2t4Qlt+zEnyawkS
oynK0h/eU2DF/VVrGz7gYki28+5ZrKE0QeXFqsuOVRjtCK6mSduY7TSihIc7ix0d
Z2273ISpaDQR/jhSQSC727LKkzAxETgIQN61C/T3qJEBuXBxFosp9mPOLQ0oYmQc
xGNXa89qIE22J0dX4hpHlPtL2FexrPmGbhakgX8U1QzgsQm7Cpbhpp+yq4fLBXyl
Qz1PNitogDu6sPtOYzgFAllAGqC5ABwD/rlj4hxMBuzcWWNfKfSD8r8TEs2CuI6T
9Bz4SOfPwQXb6REyHWyZQ9ZT9SehyGh++sNu451PXNY2FGF4LntKsL9CMN/vdROH
vyx7gdocXwdtBZeHpwOiG/nc+m1JRt/Azjl3yx5P3dsRd2gMkpuJWwilW8dJ4Isy
5LCnNJtLbUE0yTh0jCqZPcprbR/m+G99+04ys/lxK3tiz10oooIdAYnMiEQT1a2y
maoHHRiLDw8qK6EE7XHFq/OdpIOOZ7ytPOig5wHaqarWjv1dY8dvPX2+AeMJO6GX
cYnCF9yaD0ATk4AxmomEoSFmOVsxdGFHBiBHbxfCNS0khokadSGgq2nP3Yn8yJSm
dYwj5DYn5QXkoZR5oYoBcG0aROnm2Il84qoq5ois4U0LYRGLEnnHqocG90e73yYx
sJP2P0LmmPG4LDQ9SQeQTnn/AuXynH45Wcwuz4aPttvs6kfFoZxchyJOIEie4i92
QJM0NvfJR4PJmZEGrv3coxOqRsTFjcw2klEMHHIDHKbGDQWNnGQb8IgLt+3uQguN
/OeEyHXXlahzQtz2MAQg3Jp+nTDxJMigFaiMputaH0jNNvWByLdg9kljhJSmbIa+
YUNRFn/Vn38Cik7EW31FFjkKBVlpQBCf3tRDhT+wVy/Cb1xf6BZH4M2nMcZBB2/5
mllQ98tF7uZQTuUrd3rJtBEZ3s9l3qsIjxTxFk4THvZVuwM0l/RuKV+lYHs+5Wnc
eUybRpLO46HURYvKEqSXRF+YYm/zlIM8Qd3GJjXnT2gtS/qBA/+DQEQCdp7lPcCn
UwlT1Lnd0m6bRlMq06gWFe5mr18VqCb7oGV1jnwoPp6L4uGZ3I8sH94NWUsvxwi0
iOplnaiEgUi5ePPWNdWicRkaP+8h7pxlv9q227ogCURn/qZKFQfQUITmzhjT2BiV
RHdUFwft6fWDAJ+PH1rEIpcl3T4aytptbB8rcn14+gsAAsmKlf5HlAmvjTBugCxg
Ug1KdSeBziFVS3ckZ3fsG9PEI/8XsclPVWzUSlwclPqDCo1TJMzBuB/KyOfWrlUA
E7QNPxCrIIa83o3/4vnxdUL8aluvVpn7LTAuKmmqjzf2WVrGl1nXCm36s1AgoVcn
K3357HncdMF1k9e6xh2mL4IibpHLz21buuoEoRarwtU9Ca5NUDTevfAV6gdranUE
HPhswjYeGuBehvysu0J/6f0XVCzIgE1YbywtPR4F6w5seqPp6YivD7jYfns40miV
wIGHZZ2rFey50VmQI0fhlXLuFhPlT8l/FglQkXtg7Shs2Megdg+Unum8au+FKLFJ
dIV1irXIAynVdpYe9BmWAEE8uqZMk21zOelY5CGzYeJ+ZMBTH4gA79cuxOx2ASos
xsh56DTcQGfxGK/lCELXnV0u/vKfbyNJO+AMxrtsUigSua1/hN2GImfNbNMswWUC
gmfuciDc0GA6jvRegnqHpQPQYx8fJJ+X6dNfT3DBycjZ1vXvjsO22TaYgpx0CNpb
CrxB+O4m6fUhwjdKPKfRB67hdkHXO3Fcdt3NCuzKBImfcv5YId6krA8erR+YHjr+
OQc7eeex7N3n2rvZ6x1WNvDUyJjtIwyyVgX4chucaRy7ApYtI8SXPwYU4j7YAVDn
nk2sE09zBc2cogrKGgwvAYJ+3UERS1xPmyGw+cgCcP8zS4/ZD3MnRGHbz+d1grdW
T7Z5oVtCl2TnZopo5BYfNPAx9FwV5t+a8MYI6er2M7/oy8i+vM0i0CCFWjMTqiwA
ERC/QkohGZ/EYRZfbYqs5w/Zw9XwrBx6GhUMRODcHDbt1i/FIbRDAbJUWvhtmlzL
G2eWmrjyyeUdQacWZFZfjgj+l7mIVSfd7TcxEiEpcL9CSILMCMifBmIphCDM1GbJ
0gB3RkNPXG4E7n9jRzb3at6Vpdl0bzGjpfbgy1LfDqDzgvInUMb9JmpPQvPjDemc
O5hkmYULMQpCERBcsXxrq/vIaxqVMyuE9dm9UtaU6/vsc772AsPYkeMteMhmuK8t
Ca2XHRBqw4E8A3A94uGfjQbi9zT0elzZUeKkL2nxrEfwQDiY33l2Q5J2zVrXIBOW
OHe0LpWfDobCyQNLBVsL7xIvnwDaWDp1wuZC+3rGuIHi/DF9nUs32Fzre6jiopgU
/rfh+6zoEPwWMFfHKsNkw+/9u1zgumnnDAdAA46uplzXE+EbjoRGdMNBROcTZpkg
LVPL2Bpb5LYc7fjg9dK74ZcXVNsA7/AEap9dFFLBVk/UkLQGo8PuLtWD4V6zzbuG
7n7za86ta2EUhmoMi2lL2G/Mf5CGVYdqHegrQa6S7DQrqlazkhfU/BGJmED8UxRY
atxRwTs9JMVqlB3lw6bF8FyN8AfK+esla+pmp5FVEbN45uQdfasu61sw7AUA0/VR
rw6vog3YFeThRenW1plOKqJJJ1rs44K5e0FzJWsQpQBHsl8kay4vu5YJW7pemc1/
iQoFrl64yL8FFhjLs9vHmPUIQ6H1eYZrL/M5YEmHsxq/O1IUpeMmxI50ftKBEl3S
`protect end_protected
