��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F��������n�BJ�F���U�FW9d����T�+�wt3��^��r�q;\��af�י,��9NL���ٴ�[�Z��^��Jy���0�T����l|�x�5#B�o* ��J/�CO������|�)6b,P;����t��ew�u��5�v�u�E�8����R�oIk�����Wb�A1���5��r�5Hڜ �r�n+��MS5��n��þ�|R1��������E�%��0E���;%�6�׸ۈ�6��:�!�#��L�jT�a�S�N�LS�[�&Ϫ���]/��nm� 8K� 7�H�be��
@��1>��?���X�U��&��P4
��J��tz�6�^�O�A��S�������EjS�V�6�$�g)�H!�uA�����.����c:k���:J�G�y�*aio������6M�pʫ��QZkw5~��ΰ <�z���i����Y�T�w-�q$��k�d�V�5i��[�r6t�`?�.�^�v�
��l�;�y/��y6�]*T�۔"N��d�V۬����/S[�B�U��7 a��p~q������~�5�LPؐ�V�T��?*�ؓ�C�r�����	�].o������߽o8+\i+�`K��+darwEi�JI��4?�}͍�<<�,�j��'��u��K�C���=a�X̉��37�Z?�(ȣ�$��Yl\e���=~�Xa��s	 -~����w�N���,v-�xa��$a2��hA$]��g���[\�7�x���{�MO|���1Wc���C��e,m�"��<�{����LkQ��O��\�ȉu �U!}�=ã�:}e'uz;~4�����K����F6�=[�P���I�v�%���/�?��yְ2(ݡ��I�^�0Y�)��wg9�.���9A�Ld�Wa�ɤ!8�>�B/(�z lE�d�V|.S�Q�q��b��'t��"���iy6c�%g�X��K.�,��������C����{���#������9O�
�ϔթ�4/1Y��pt���F+y��{N�ǣ�|1��.[wZ�
�_� ����CM�^�$��(%t�c�z������8��&��M����ؕC(f���kKD�~2~��\~`1l�f���o&T6�е��V���]*�A��I�꣡�g�����" �Կ������g���׿u�ط�	�l�}���]���!�o�o���E��'A���|B޼R��Goa��W��Ԇ��:z�ĭ��F(��z,����`��B4�O�`�()��8���&A��M��;8Bo�Irbیo��N��Z�IdX3�ډ��jI���ۡ7�i���7�	 m�#"���L=���o�?��
��&Q�򊤍���DD�w��=����t�DJQq�����äR뎏�#7����	E#t����0�<߿P��-:�7��p�������[Ad�X$��5�)AɴP�g�;^z1�i V���5ƍ�	P�ru��8�]? �a]n>[���~w[�$لٰ���ry���
f�:?}��h�h�ܠ�UݹA���|�1�!n�>�l��[ͪ���7�9Q�@�w��n&�s�s�{�H%�5;�5���^o.��yc��^�>Z�w�з��2���.�ZR�C��9�>[��1�-aI`w��v�e���8��v�w"$O<Q����\��|�o��g�N>��_�:�y�9Y�@���\���pEǇh�3��DjFya�$\���*��U�g^G{��#&[�N�2��;X�5L��7��(z��'H�v�)M ���3O,��.٬���gc��E/���6	��� ��Ԃ0��������@2iz/kN�A�t�NPd���~��.��]�����e��g"�w�[�]��޽�v��= E���*o]F�/8zsN�>0:��T٦�J���
;O����N<:��$��d��5�5Ņ&m��X?�c8�\��;(,�"�<��"kg�K6�3GC��u��"���@:�d�٥<p��}*>6+�Ipw���w�Â�f(d\:��5�5�P������p��#(%3�2�L|�l���;���'�OS��ѻ9H��+�Y^V�q̄]�g����F�`��D�;� Y�J�֤�* �����7�L�I(�#�pNj�
>�;�H�H��T�QX_3�����-P#:]~O�������r��z�Z�;x�k	ÌY;�p|l�"��(�fN�w��'��\`~��I;<�%�^��	�xjb��JauxTѼ@>Ҍ�����T{v��R׭ٟ|�Nm�������nȑ7��Չ����� ��4��rM�W$+��9�2yM{e���G�;̲,�ʻ�u\R�#�8
��öb�5ٗ��7��`$��>�˫q���LL��\0�	hW�r=����:���<d�PG��'%����������}A}�L�S��^��+TG2.8��݂}����UGݚo�th��c)�����M5��{U�F�=����س��?9�#�h~"�/�l/�\ia����i���=���n�5I�)�p��xr�8&/�n�s/�}��Zo�U;T]R?���}h=��m�	�q�)�&�n����8�6��b��Ѹ�O{ZW�W�>����wx����$^�pφ(��_�K�N�O������t�,�w��1U��y"�����m��cz��p��}@���l�OWG�'OJ(��,��K����@�3�����,��u	���1�����sot֓vb$h��7�M)��iK���uk{6A�������5HN�I~�b��2�k���ih�1`��g3ò��@
�x»��~ho��������%1�]p����#{	�.W JW�=�� �NK����Z~j�`{{�=6�L��~p�8�T
{&�{]�ܧI�-�Ѯ8V�k"�����@�D]l_4��E�Jq�,�Nv��V̟v"�:�\�k5��f7Q)�����om�����5�G�E'�o�1��� $
\���4�r��a�i��2Ў�x����j�\�b<7ֻ`��n����J�5�Y�*:K�֏��-��+/��0��	O�/�N�o� �'h�����œV�e�vp�O@�� �F���7w�)eSuB�����䵈�>�x9�5c�c�k�m�bN:�Nn����8#,��٨o)N}�i����Gy�f<�)VwG�DA	� lc �}fzh?d��b߫��b�,�Fǈ��Z���AṔ�0�V��u�^�f�.������\�z�� $��ތa���$��M�I~��W|��v�9@����)�%G ����k)6��y�0�N��k�e%Z�c�^������.�ͻB7:���Y��y��V~Ԃ���AW�wP��HI� 5O+4��2�k�#�����&-箚B �N��
9�2?,rb��=O������8P�:�YoRC�B�4�C �_~.�ҲI:P;Y����X�dM�ό~��0���f욳�U���+w���5e�$~������P�qfe�
�Q�\���W���p��X���~�߶O��2�2 ,r��jMxK���m�(����sm�SN��:�k�����1O����#l��J��c�����3�s1/;4�(
���H�`��~��47�������(#n��<���=���L�t�>�h�Ғ����f��j�?������p�0�w���� �� jQ$2�]󿏛�|&�{-*��dp��p�V8<����d��(,hJ���0H߅RW�|e!.g|:*�=Q��ǲ��Q���4��'06<�l�1$S�d�S+<�Tq�t<�t�wp�ly��8$S'4�L[���zT�x�Wd��yϼؠo����5�?��0<<�r�TOS  ��(o��TC`��h�h�k���9G\]���1��7��y���{��zk�̙ 5����uob2��]����x����U��U�Q���[���6$�O}r�@ь6���מ�:�Nk�7�V�+S0��9��4ٗ��}H�lNOƈ�,)'����#�@�N�:��mB0:�/$]g�ǰV�=2�Y@��U�ΖY#>����C�{��c�����2�C����~�`x��?3b�
ǟ�#+Zo�4F��c��s��/l���_/}���\�FB���K`�[�鼙��b�~��;*��T�_ڞA�H�^�u��iҡ����[��<�u���Ã�r��
b�U̩�6�ͭ$,��&��L���s#�����kѱ��E�24NA�u�-��P��#lo�l{}�Y=N�I�U�����:�mɆ�vGfZf14�d��cjA���Z���.fpq:<���(�"'�'�Ma�f�+V���l9�f|���W�7��P�'�f�}C���?���sy:�O����a�Բ���<�������n� ��5טG�J#�eP���o�	m�����-K�ҫI�l2m�/?�#�8�S[y���-X�"|wι(��{�3G.��v1+����}�ҹ����'J96�dQ�xe��� ��w�-�FC�w5?M�J�a�iBOe�H�5�=�άjw{*�bG|&�7��6�CV�k���sG���h?�)��Wt���f��,
K;�%4!e��kD�L�S5�,b�#�:�9D�8�A�<V��)�>˗������[X{:������pcl��s2�N��N	�g��iH����Ã�,�یU�Y��#���f�X�ԡ�+L�>"���G�q4��|N�fvq�u�Jx��K	�%��pŒt��e��)t�>Ȝȧ[H<��+31��O!pP�(���y��Fɼ�0���;le��b�~P��7��[��G0��5�N���{G�En����(�S�<�[�6��9���\m-�\C2�'j�첊zw����C�y���\%���H�}�R�FbH4�^�f���~�����Y�y��G��GhJ�}CC�=+/���1�lv%D���XW��' %Lޠ9�b�Ţ�/=WlM �G

z��n)��*.�I�/��(`�WJaT�/x���n���hD�;�^�$j)���g�[(
�U�ر��yF7x�R��])V�����T���F�=:�N�R+.��܃�t���9�h��YuXA�t�E�i��h��O�[,���<�U�K�A�4��$-8?|��i���d�!?H���J	�[V���_<�AG�"�T�酟���++3%��T}�@Ƣ�*j�aIt2W�1�DX'�D9�.���ۥ$��8ְ/�3���V���]M�K��J^a
�ם��\����ړ<�'z�9�I�q�ψ�Q������^u_ک\~��ɺ�K<�a�`w�[(��OĐ��3@v�%s��$��p�췶��2P�*�g5�Xx�=�X���%$^�Bn���x�5��Έ���B��mSѸ-�����*H�\zǳ��(�ɒ6�ʁ�c��H����\ޕi]$y#G�kV��LC3���h����V���')��
��K6"�O+`Hd͸�
�d�� �]x����=0��~�@V�Ҏ��~W���Z)�]��A�8�n�=�$qBO��r���QS� )R�`��r�Ϩ��8\�s<�;��*m��P
z�^�~cl��L{���ڑ$����⡮//�4�x���;�y(o�H��^���Iޕ0e!ᒖSp>�޴h�އP��l!�O�����ix�-hI�I#D�]��<GR=��<+K�s�t\�g	�Ze�C��)�
_xT~�W/�<��ioӆQ�x	�$���˽��ƞ��M��B�ɍf8�ݞ���!I¾�[~���ݿ9�@-*u(���Jd��D.UqR̅.e��A����� ����A��vwf֋��ct38��ִ�f�W��wL!h}c}}�9�	���&�)�3#�H)�����f�c��r��՜qv�MZ^%��[bJ+_��1�Jޔ~:S$����
s.�rFJ���`s`�K�.�{�*� DỊ�[޵�~��Xj��XܽU���!	�CO��.f���Z�[���,��eL���ܷ�"|�����\��q�U ��&D��4��u�:�VnI	N�A�7kB}{�6��bI�s��jd$*�2���@�I>>-xu`.R(���ƴ�8� ���t�yN���(�w(��l�!ݵ�����@�?�"�Ƈ����}3D��TH���+�L�o�{�`9̪�%��XU8?��Lq�k}nOxP�%���@om6C�u�w�& ǟ׷��/cj+��5���0S+,��סP�G���/.�Se*K�'����.a�-�8�����Q�0I�]�5Mg��ku�0�!I���	Eh������~^H�Т���R-bJ�@�2U�{�d?��i�?�� �VGi4^+;�]+i1�~�����
��E�,i�95����ã���	Z�M���`���E��x��9����͒�S`s��b��M+&���������ڡ��%{��tp�>缒�^欻�w>0�f��ӻ��[^F�ӑC?mn)uq���<:���9�)��Łۯ���hN��;�I����z:���p�|,��~d���2�B:�N^̚��}=0s����u�`�E���|G���~�������l���� �,��^f��.>�_4[\vq}�R���c�4�Lq�tT����R�����^ώ�_�����Rr�W���G�4ܝa���zNd46���>�� ;�?�B�vDǞ>�Kc"�@~z+��j�or�&rꁆ@�M���|�n����^a�>w�v$N@࢓��e"A4�`���4�k��gy�N��G�P�΅@�M��x6Z5�c�_�?]:R��?3Z�@}Sf"�>kw<e����jc�p/m��K��	��Jh�]�����	P�G+���?x.73���ȩ:�i��؅��=a���]�����s�L$��4��fr��s�����K��]�l 
)�y���m3�*|�6r�K��HYs̈��!�ɾ��n<0�'Y����h��·�I����%��65��7�]��
5@T��q�{���#j��d@=tQ��*?.��&R����.o�5��E4�;��L��4���0��t�����X�����T����?I���F8�L�#R�ϵ�v�G|����Ox2���0�-�a�HI*�j�P�J����4����m�=E>�%sw=����Fst��}�l�v��,�Y7��� -%��c���WȐOZ��q`�\�����0\����-�F��+����k��V�5�oG�Nx�%�Ys��gx�;>�M�U��.���\E��Ώ�Rl'=e�%�PW����J���i2�s��7E�1�i&�P��p�Y{�:�կ�3��zo�3V�!��e�]��rPJF=�N(��aaU!YZ����y��j��>T�#*Fо�*�=��Mm.=��O2+NӣQ���M_���U	,TY���LQ �G���C��x���S׼pZ�J��҅���([�8P'��+\inn�o�fN�n��a�V��Se�S�|_��iXQ{Q�D�0�F�)f'@`�Vo�� ntp��l�kb����8d�A��#�狺M��=^�q):�ٳ���$	d������� � ��~N,����eE��US>��F��H�ݒ�})Ν��4�����M���c�$*��ϠM8w#��uם��`�M��0݋H:g5����v����3z3�� WIk���EWE��}�gF��9��b��ߐ��� ��N�u�\�z�H��Uo��'���{�f'�T�ec]1,.��v�����#� >�Jg[�{�!d�/h��9��H po�K����N�Pbc��zqAB��|�Y���\<���EB�v˕g�ը�6�0(�{������9�j�p�*r��P�Y�� ʎ��^����9	�/��O*0#o-η�Cֲ�Ѝ��2�����d#$����f����-��}�b�ʬ�dF�n4�m���忔{�&� ��2�v�����f�#]}�8[q��G5�wyǤ�<�h�-AF�0{I:�~�1n��\.��䑝�W�S�!?���k�u\���)���P+!%����y�I?�����X�Ry���[=[ݨq�4��H�g���rЊE����H���=�O��O�ي�mg�8^���܂����[*��R��ptӼ����aX?=)���R6R@sL��t�--J&����/�FL?�kt�����0vء��mb�Mwdgj/��`�[$�[f������O��S����k_�t�|�� ������Qr|:��*]4���"P�/�T���^4dk0f�A
�c����F�I��b0R�SI��hk~��]���������޻�<��T]��������E�$,���aq�?�S�Q�ą)⌍~ܿC�b��W��@�-��:��7œ,(��7��ā�*��p@9�^bASz|���O�;�i�e����+�^�{���/:J5af�=g��X��O�Ur����m}�FO�s06G ?��}�3$��'c�B���9�b��}����dk�W�1(U18�v	�*�]TF!����Н �/P��V׀|�/B�f�r���z�1Y����1^!g$��IA@�e>b�[��:�.Sk�]�G��E:�F�$	�M�d�F2K�
d�H���'8݇�	�g��[;Bu�+q����������.o`ΰ�YԠ���)i�Ap��*Z��V����?���?%-ܾr��j݉�,?���=�"�C�ME��n�������f�0��,���L��9�D�[D�k�f����H����~C�U;�[T����G۾��,JB�GBE�)R���$G��(*�A�Dˤ�GU��w�!(u@oY�֠^�$D�܎�K�V��2J�GBsZ�՗`��E>�Ѷ|6ez�p��	XlM�?L�v8�n�f��������gxp�Eq��]�I͠�,���jt"^ć<��~aH����" ��qg
%��ꤟ���$�Ol�a�b�� �M�fs��`��%�-ɠ_ʛb?�|	}UZ#������#؋�PA%���n�8(���+��[��֬n��K�S�f��w�Ѯ�jc�n���%�G�i<�Jc_�%Co���9V��e��Ęs�RZ׮�l	���'��i�!I�\��*����3"<z �cw�%�Q�e�:9N$Onַ�Ҁ�a�6x�h��X#�=���ґ׀���,ADA���U��F-=� �f�-��]��U|23���IF�
�*��)���n��/�u�lY��߃�n%V�rc#Զ"nVG�i��r���Q��&ptp�w<S�'�9v��TP@���Ȁ,���u�a��J
M�
�Y����%����v+��9XD^ IQ�D�Cf�_lE��cTб��ŧ�=���b�)�����qOQ���<s���ߟ�=K�SP��o����,����?7;��@0�mp����ύ;>;�Mݗm��w�i�̌�bj
��w�G���:�*D	�Ӽ@k��#@�/Q'�|ו��	2��S���N��� $v=EYh��$��:=ĝ��-��(��^�Tx,<x�Ao[C=������b^�r	�#w��&�/+�v�N~�����ɦ�9�u� �>	��P�?�W#����A�w.���S� �N��0gưW�s�ŉk��w��'#� �h���2Q�OK ��wbd�9Da��MfSϩ�/�c�`&[�o!��l���"$ !��k������z�χd�N�O�LH����O@���!FzOq����g���{E%����$9e����� �`d�K���w�D�������b��w��àˊ�8�`����=���f�R��8��Q҄WV��7�(�{��^�79O"��>�qz��L�[?��7ͭ)��}�*�C�i�+�{�M������^�5k]mu�gz��}�
���t�h_��F�i��#�����W�]&�^�-���x�F�$>��n�� �k8e l����؈�-�F���<ms.��x������яS�~���K9��-��ÓNU��>�w�u\���>�:�u�����:V���DD�:�)�eٽ��N�d2�Q��Ș͕]�gї:#���=�����ͳF�Y*���о��68o~���%ECf9l����
e�Ek�T<5��mys���E�#`��m�6\%׺�B�iU<ƍ��_��� �f�M��N�'?�qA�8�Y���a�ģM��ۗ�k��1"����J�4�0�e" �`�;�D]��~)	p�]����hht��x���l���� �Vd�������6�A�;E�OBc՛�W�Ãଋ�o^i�#��kBi�����9,.q oM���<�8R�ȸp�2��7�����a��N-+��E����K��X��OuE3O�,�h�`ڙπ�6���#wL�L����]$�{?�`�C�s{q�$+aȕ�KLo��#� ���������첫���zo�6��,�+|��ӓ��{���8���,+�i��R//��PiQ�Y�� �%aG��Qi����¡o�Z~3	��'�� ���R�+R�eD�!����q+��=�Z[B� 09��
 ��� o��w�����H��KxŃ�+֡���TFE�� �cj1(����qN�ĜF�����'"?�07*k�F��������[� �~��J����f����$&�b���Vx/8��bH�H�����~Aߐ���?qU��u.���U���'l�f����N�#�q�-oT�-���*z�-�_�#��?����9{8��������-C�-�@�O��qLY�0�"@�v��4�H	>�%iey���$�bT�#W C��#@�T��u�h�O������58���8�_��Ág�!EeM�-���Ҿ���8xp��eu(��"�����^{���zQk����1_�T�jnRN����rV�N�4�a������$
]xG�m��-�t�РƯ������(6�fc�4V���ԯ6Gآ�s�~�
?�z��)^�tK�T�N���e�9���1��m�ਏ�\a��4���)�:�.��A�x�fW��sc~�G\�}���3󛷓߸���pZ��'�ȹ<<�~��tF�d�A{i�)/O��>�ʍ�P!�j���f� śQ+��6e���n/+���)�G\�hK՟I��JK>����WԱ��<b)#g�Pޝ�2js�H���D4�y���l��$O�c}|7Fa֗2���D��{�o�^"+�~E�̥l��AC5)z|A��8�x!h��]�
�wo���1�<�{1<�k(��Rfc��Ҕ|�Kg<
��"4��߆%��//�i�ysn���\/���@'��N)��Q\$^�j�u��J�;g5��?���9*���$=u��uC�n����B������ѡ�݋��UZ`ȹфo�/�O�/|oX��f$"@Ὸ(dʋ�\u{�ﭪHQ��c�˧��4f1�A��1=�pAF��w�v��s��l��f���g��Q�A��I�M>�{�9<�����$-ވ�
vl:c_�Z���=p#��� 5Gu�����(�%(�fl;	K#k����wz�MB
R��!��X�$Z�K�n��s�Q��nP�̩�N��@�ɠ�����|��p<�T�Ӑ@���ܱ;*�I8����Ox�M��TMȂ�y�	(<p Fn�s����e*��u�9Zl	�z���"���I����xh�0�p�6�x��m���r\�u�ݟ g|��<ӣ����oW���'�,��P��qx��ښ���	r��yku�v�u/��湵�?�*�_]�"ӽM�������[t�t�x2fn�yeO�F�$��5[a�Y���'��C9�f%��8���ǥ�;��y�y�j2����H�X�	9��E2A�Jr��b ��/Bi4�̭������B+^��q�k���e���_=PG�����-�J0l� d]�˄�T�?��\���3�3���Al��^��k��u(���ʸ�H��R�[`_�E:<��Ȫ>�&R���(C?�S�V��Ԇ�:��)����������n}���S�G�l��!��[�Mn�h2�[�
l^'�k�� Љlt1b�4�����s��>���0-Jvn����NV­����[P�}�P%���jj ����3��n���_#���ڜb���#?�]��Lu�(��c��l�t
���S��挶A��4��_o�䏜��Ջ&✕�G�Rɦ	 86ڬ�ye��p�Y�x-g��e�x��I��cXf;4�>� 4���.&F����+� S�D,cy�?�5֒��>_q	kF[A�h	ضB��F�j��q��$�1�I�tx�u^���O���4���:��s���,L8]�k+-[��Vs�$�N�02ۅw�^�F � sd a��P���F�e�o@kAʞ�
���(I���Ҏy4�W���	F닓B/ӎSh7������t�Vs����(�w���@��*�j����ւ�XA!b��+D0����r��1����-5d���qJv\�N\��ҹF^�?������
 f]�U�]}�;���uuZ�
G�iB�t�܎�3�gwtz{�]�<.c֢]���Y�;�t8�6���=��=ΆN��D�)�c͹bdP����(8N#WSQe!U��[D#$'�{��O���g.O, mX��u�B��~���k�_dTk�lg6�YɊ��O�>@�u��Gz�O6��f+����A�5�O�������J�sC�^�t�|�4H\�����DҸ�$��'�Q3����%�w?��>sr�A�h:�?	h��wб�j4�

|/��Z� B3Eug(Y8 #Y��!ͽq�����N�`��eE�?��R�p~���#�?�����c_���
��jxi�)6��� d��eӇG��T�;b×��PB9B��e��L�8Ü���}.n>n�BB�.�F�t��*�Qq��+ؐg[�FPD����q��Zo���r��krM�n+bIT�7
�71Zt��L~Ҭd�W�E�����K�6�TF��?� 妴	9��V ^�8O����,��W��|.rϒ����{�S= ҫ��ajV"��>I��d>���H���}Js�&~ �����a|��H��c #�H�Xq.fy�6��ی��K =��m�3���7�_8�3$��d̒�0A��+��(�~�%�w8Yü��E.{8���d���Q1����oID��G������|��X�ժ��!�Tt���#Hz�W^���WM{�Kl\����얤k@�ZO1����[3R��ey"k)Qt�Vȶ���L^;����jV|��YK�����h��9�8��3��Ee�R��j\<X|��=�D�t�
(��̇PO7 >�{�����ڗ�z�6}-ձ-�ԬV����k)!^`:h��'O��o���D��r��h/y܀61aT�y�;o�|������iCp@�u��,&�P(:�pT�υ4����JU�㹄��K#��F�&���i���������,!ދ�����qτ��S�`�LIqYf7�D��a���i�\�mUdӢ�ï9j���+��Z��-��ϝ��%�hѓ�؜���-�^b�[�44�$�;@gjŞ�:3�i̭U�ҵ���;ڴG݄b�=��'�Y�@����rY n^	;$ˊy�L��؄VVoۃ��%�=@<�k�+�ѩ��M���P���of����w�>��˲0-eFY������,8�e�`C�@磼^�3uF����d�Y�����y��n싽9��7a����,�/�'� l���;�J.��<'DX}m���|�Wr%r��3e��S�9��=J����[��!� ��En|��ud���֭Ca�S�o�]�Ť^x}��4���J����H`)��V
͊�[��yX�㜉������*R�DΏ�&zY�+��xw���3�v���r�ȗ��@{��-��{9{|���L���3�U/;Z�}���֖�*=�x��-_�$.n���^g�'e�������ӫt��)�$ǖHLL�	>�q�Z�f��낺��p&�x��V���%}�!�~��Rw��ؠVؙ�-!޳��sTOR��$V}��ġq���X4f^�e5��H�����7^��?�!� S���_�����%lL�%���L[�J�KÔK��^0�\��E�/�E�����2W�"�\Gk�Ts�o��x,?�;B�N]�>nS�
�o�͑2/�y�gz��+Vz�w��qOh�*��J�/ǏX52<�C��`{v����oc���~/E(���;\[z� c�f�V�2��OR��
�e	rV\d�2Zi>������r�%>�_�a|p|�Q��}�Kα|�	&'�&���)��;���V���n����POJ�(��3pP(Ym7�~%����Q��#�T��>��4Ȕ��i�>���S��f�Sp/s����a*��宵]"k2���Cw^PF�}
��P��#��/�Zk5䅊���H��֟�v4��⣸yu����q�v�o���+\̪�e�;���_�$�D�5*e�[��d����*^�d��J$�Ce:���R�2]Ț~�U]J�}�$ 3����s��ߌ^ߋ������p.�H���77�y�h�� X�qc/3���V���u<�&�v'�=�2#$�]�M����?��Lc��$l�2�X`,�P�lL����S��9 7*����Pv���� �Z��ɣ�3��ntn��>a˼���n+�0m:SM^>��:k�z��^bn�zu�(����$)�8B�d�P�-,�^MݘNq����R�~>���Hi����Ҁ�/P	��)11qe�§XZj��':�)y�<�uG6���9[�}��Ǡ"8ΰe &O�kL}U�������.�8t�ۡ��	U ڽ���$駅�3���#�&�
.gE�т;�Ü�8�%`9���^!ˮr�ڽW��H��`z�)Y/�����ꚿ6��1bL���A����_�}�]���v���+���n}����b*B]��s���kʵ�բ��Ou�ܩ�@���-���+�2�rDh�X�?�5��n��B�nH�j�T�?��ӄy��0n��ꆨ�U��]{,t���Em�K��@~�|"��⥦{j�f� )o�T���m
C�n~k�-��h�mx��tbE��$	����|��z.��"�i�+�7�/3��x�"�޻�݊*�G�/�Ʈ/���%E(eOO�W,n�[+�b�Ξ8g�$=�muN8��BڔuΆ�1ք%}���M�ts9gc��;ns�|QE����P��Q��=�F)Ol�	6r6��􀅜Ɲ�6��V uM�����쌁o�D�WD��̯����Uev��)@h����`R�m��W�ܗo��*k�a.�E2f�`�`V�����TߢRs��3h?��l((��c��g�^L�j����o�o��4=l��By��"wyq��h��>it���� n�"��'����]`]�'Q!!a�z�����6�~�7o� �w4�"�Q y)�#��
����i9�D���r0mw
4&�K���R������{�g�鄹ݷ�Cmg
�P�צ}5zi��g0?(Ө�<ԅ�VvRq��ٱ|r���H��I]�������7�.�7�?�Rr����i6jE��њ��^hr/N�x. +�p,xі�Ƿw,_�Wծ�ӱ�ʌ�@AȽ�A�D�Wf���y϶�wdjg/=�L!6�c+�Wc�2g����(	������]�п�;z�[�Cu�K�L|i.]x S��2�}U�K+��k���Wj�5K�PQR ��E��R\�����$�L�C�������:[y�C@!��?��=WmF ���}kA��|�9+��y1u�Fjm�܎�%H�7��-r�Ca�贰gM푢#��	A��]�3�H67�B��R`$ͷJ�eI������sd�3UK�}e�
)/Bfq1d���W����z�/����������P�f)n�U۵�\gj�B>�0�JkΓ�T����2n?��,o�����!����x�^���.Ϳ��q)���E�X�3/�]k|(��#ip�#y�`w�:>���$����t�Ԭn ���W4�j�*O��B��k�0�,�2�ق� �W�I�i^}�a�q�
���`���e���}��帛{�[rfg���胊!��T����Y���+�_�P3O�'���:�渶��5�X|B>�����q4����/mf��I_)���M�,2e;kٔϖ�`w�Ȝ����*'�֘v+<l�.5�'����h�$`yu�|ӡ�*���zIz����'��D�{��� &mO�or�P3�t�D��Sy���$�1r�|�
��AK��tL�h��Ɔì�סԠ�ѯ~�D�@kgJf����!)��	��b1w��L��5�mIP6�5.�PzuZ{N�ixcD������{�\��m�UR��l�?�"�'a�TX�����.{�\Im|��d��
����k��)(`��9�3��%�K���81��c�մ�''Q8j~��P 6ܕ��Vg�qk�O��&�S����Z+o
]������o�T�+j�BS��K��@��uN4������:)p��{Q�a�Q�=��� �v*рד��Tq �b�}��AR��Gf��S��(RW_���{������ƿۉ_uֈxDb�Ti��.�uP�^�)jR�y�$yzU�}j~�Ʉ��'Hn���Y��r"�W�=ꗭ�T��M��a���#F��̴ ��4 ��#�N������?�iB�eVw��iG�"�F��{�y����
-�.#v�n4�)�|�D�>@�^�;��PU�|������3;�\&p"�C�fKbY�	�&���:GFLO��\OW��\Dj�w� ߚ�-��K �Rr�OX�8�<`^ʸ+����N�]�ާo�Y�L���O����,��*���*�R��`Vc�.�X���C��������Y�E��5���kj6Z�J8�"��Z��4C]����S�Z�s�k(Ϣ� Ϛ$��Y�����vg�p�0�.�k<�ȴoT��D?˗�ڏo~��z"��v��`�aT��]V%.�T�B~�2��b$�V^Y��{�vxf�Q�7fpQ/�̠��(��Q��-��^��؟�ֻg6<�\�]��{��%r���! �(���){�E���j`X�TQ}Wx��(��jl�0����R����{� �o�|'ܷRdVH���+[jh!��U�]Ej<��H7��X��q�(.�`:�&�����Y�zQ^ĕ�pgY>\]�koɳ��ȈnYb�I���rk��$څ��N��B����1���I��[�
)/�vgr�&�J ڛG��v6�6rūVߡY���gc9�u�S�d)��O�P̪��k����a_|�7%Y���P,S=Ln�9�?]�k�s��Ȍ�����5/zSd��X���H)Ƽ�2�΋n2�,L�q�F���SJg3>����M���� ���T� 57��F��bW>��4f�a�QC�htz�����$P.��'f���$W�@�*ľ�=n�{��Y�k�ꯏ��H��gIa��S� ��������=R�@�s7p~�N*��˘�)7L&`iGWíJ�b�s�<����c���o�W]:C�3zP��Ȍ��v�t��{�.�9Vu��좷�2�p��×���E5�h����V������ �����g�=��AEU� R$;rI�}4�9�7�˞����J;�գ{$��K603��s���{7�;Jal�-t�S�d����+V@�q&�ܹ6���[+��:K�]k�98�lu�?lpI<u,�X7��7��s�����B?"�D���2��e�,��N6v�$r?�nd럕�o�=�)G��at�Do�@�ƫb�����nTj����j]1g���m{No�j!:C�H���з��<�!�9#ow] ���W�Gl��[ɟ:M�K�sDjp^$C���� (PXz�8�N����<p͔,��B���t�~bm��6�]j3��R{z;�*lƮ�A�D/��/9��8������\ix�uh>d��(��3���ɉ,��X�Y�4l��_rv��G�~��&v�>�
t7���Y�_�%\�b����@�dtI�~���Wb�OdD����!7����>�}O�.�|g.^B.9�>���'G�ύ���%4����	�r�E�N�|�����׌�i�]�.��F�ڗ�q�QXu �a
1���X?�>��(��3H�+֕�_��P���!
EM=yHz�ކ�ϔ�r^����+݅J����im�'��p���w��Q@S�ׯ��tĵ8N%�-d�+`�#���Qw�Zo8��}WV�}ؽv��������r��n�F{�C����8b�[��9s�������Ϳ�ᆤ�ҹGo�P:'=�����:�H7c�����=D`Z�t��H����ym�_ ��À �0�#u�+��R�&b� u��փ��䶅�QCǽ��{��W���qp_������T+�i
��3�@��'4u�`�$k��y��$������l�V����0F��-�(�I�;�������/�l�%�����#�l�uo��y��1˦*����| ̗%�f{���`�o�dR�`v`(����o��"F�����!ݡ�&�L���׿���,Yğ�^�|~���3x;q��Z���~�j>��AC �����b��q��Q�U����0�;�&]���v����*��߿��0�'��vAZ7��H��FmXϷ�)�H_�%�����W$H>��X�^��j��p���r�k� veڷ���2�����^tLA�+�W �B�iz��x,l�{�':���	���(%���~��z��Xy�解wN����O����4pTӞ4jy�|_|w��6U���w�+��.&A�!�M?�.'��z+,�d��݂ԥF�E�+zVp����n�p����4ҕ�.
���yM�F�i��H���L�!KtB3'�`'P�^;Ǉ8�>��s<��"ɗ=5���#(�μ��d蠙<p3�-Ga�)��=T@�{� ��q���b����bS�N�f�|��1t����S4��>Y��	��0a�,��d�ͬ��P/�QC��
� u6-�k�<��b5�3Bo�4�y�¬,�e������MHZ0=֟�Z'�y��A���JI���V;�2"X��×�>��x����>��c{ߔml�:m�T���|�mڀ@�^�
���^\�3y����NPɬ��owH�ϷI~�ÊB]�К^8��*'������:ѡ�P����'b<;��Рէע�J4�������v��3�ޓ��ֶ��}�M��hp|G����i-���h�{=Ğ�Ƌ�+a1o�R)�+�Y�jF8e0�Mu5�(�	|��؛[��B�N��Y���_��<+�FI>Eڬ]6��m�����a�������m�ne
�z���E	�H����I�W(WO(�2Ç$X�p��[�no1\�pi9�i�,V<��ݗ����q�7o�B�[�P��G�=ޚ�P �S<�Tk�
��;ѥ���^I:؇�r+V���4��&u�B�K{ݤ$EWi�m�r��z��n�S3̇��yPC��A�(�N:}Alْ�����|E[��:m�!�L:����m�QMsg��Jɂ�x��l�r��_��Q5`:�ؐ��Z S7V��}�/=X�����_�t >�e+wB��׼K�iXԆ�W-/N�����H���QJ���<���J3���N����� X��Xxj��i�}�0XvQ��8+VSN��g���'�2\�L��h��pC4�`[���LI��y�@�*G��K�E2�c(�	S~?�#�\R�Y�N ��6�O��iJ��������C�?Y9rr�C�ZH�E30��3��c���?XS\��S�`�����>m��(��w7��׍�~g;o@��A0,���:Z�m�`S��3�	j,�8aX$��}�z� y��o�gz�?g����o�eg��W�������um�sɠL���n���ûa���A�>���AD��&vu�� �Wl�w���ˢ���0瀇{�/q�~� ����O��W3�iH��J�� Yf����wf�#t���`^�ٟ*�p��Y}YL����f1��x���^|_�5�$L>�}r4��&�;���%}}�q�đ���@)��׈*/��
Ƴ��ϦY_u����)h>�}^��px_��۾Ll��~�y��G{c�T��@����p�� ���0^��@_�8V��N��H��)g�ֱV>\^��Ƅ�ʹ��r"�[;T�{V�~I;���[�C�^'Ӵ$��yk���\�6+�Y�7�f���57�΍� m�HP=l���t(��,�H pW�%P�І��ve���B���ȝ���_[�0:�0�WI#)I�<�:�0�&��O������|�V�x�Z��2���O����� 7���k�(\Z� ,���Gg�������|�%�܏�1@#r��{�n��擗��&�=m�Zde�܌�\e�Ȍ}�9�&��"���``v��e�^a�y���F``t�~�.�r^����9���k�wq78�~#�~������Y�H1F��oIW4{Z���?��D`��a���odg	|9F|2�$c�9@Nj�x	�݊R��w�=2�(��7D04�_L���}u1[������Q+/zHnHn&�l|����K�f�L�d�+ܛ0pH��ia/ܸ�4���pd�]ʍw��� �[�2�s�`W�W1w��p�'�М.���<2d�:X!����3g��N��%:oۤ�� $��=��Fc��x�D�������;D�X�t"�[�K:��Gx�Ү룦4��Y�uO<��0Z)j�o��'@ڭ?:�X2��y����^hWi�<���cڙS,9�V$���T�n�qn�c1�f	)��HWߖ�yS�Բ��O�ڵۥ!�^���T�H"�o.=��7l`GW�&uň�V	�����0�#]�~�[��'��޴;9�$IK���d4�u�a�����K+�b�,L�k	�c��ޕD�����H������ΐ��n�!����=��;��S+]����t�~EBL̼I����N����]�U��(nitm�Y�>�GJ��;�<�C:\���K���������
-5�K��t�m�y�n9�q�d�E�\ae����Oi{��D�6�>F� `��KF\�5��;uaE��_��z�kn/�=XY~��J�]9Iۨ��Q�鰕���SUP�&��Z4�q�����Oʹ�]�Dh]a�$���$�H�%4�%	.����2��1t/��X��r]��0�(��r2��'����B��H,̡�;���a�r����!��c�(F Q?�Z!>3�C�]�_�Ԯ,%��B9�9�Ȧe$'G�QC�f &p�Q��J{}
W�IzZ���"4��;7_�\���d[fWl��e��Q �oR`�̖7`F���l���䄶gѝ�i2�I:�E9���i� B�[�faHuZZi.)0�U��Yd�_ul6[9v��J_/��?�V��\-E[�B���&����$PP��ק��CON�\�V�լ���8��Ԭ�4
�ׁ�;�:尵=���V>q#��]��}M>��3��o+!��/m(]/����M�S6�◑mH�|����W�KX��V	g�K�.M��2���ʳW���y8�$"��\c&a9�=�y�*��9��s���zS]�xR���K�����@�8#C�^(��y
Y�P���{�Qp��\�Sփ�Pq^��z�[T2��BnZ�}nz��~뚹��,\&+�f/p�;6I�c��qq"h$���<W��FdcD��H>����z�<��i���+us}kY��=�c�&wL�],���m4�N�^9�:�I���t�W����[�*�v���1"�
}�h~U9J��F��P�s��=�����a�I�j=D$&_~rIz,z�x�&";ǣ6�2PVvB���+Im֫P�!(�$��H�3��ֽ�A��T��~0.>Hi�������2�Bå]!ʹnP.�����2(=g������|^}Y#���I�&�\�&�nLe	i{�}E�SptԹ/ik܍��A����ᐴĎ�}H������%��@io�ru��]���f���nMW���;Zt���	�k�̳�ee��޻�0d�B_i��;����'��ƛ���;@����Z�E��*�q`
2�#4mB�}p�z�F7+v4E��H.�o�� ��b�W���M�S�,��20%{Y!�Q.blK�xV���0l�����S0��h�#�!��.��������Z�i7�K��[�EeG�tR=����j�&�5~|���N���"O��r�,r��o���`2��Yڠ{�ts5�0S��ߊ�;�$���a�b}\��=���(�ڛ�0�0�T߀��IVk�O��$+	�
^Z�U���U$F���eRF���f�4_�D�6ז���0�C�1\�<+�<�V+
��p��x�X���|�S�=^ĘEr�nӄ%`
6-�#8�P:b�7���f~I�ǒ �Tw\3C�P�~�q]�
�v��׭|�(u��I(9���{;[5�;���	q�̷Lh8�i�j�ʅ��=�aiy�-n����z��ｿ���g�PO�5N�p��)�ػ5r@�_�;R�&��|Q���u(e�`��#��%�Tn��	�l���bz�p<za�>ArG!�+�}=+�4za�`%+[��(���s/T�5F��T��O���X�V�ȉl3\���<��qb�����+~�����%*GRW/m��P�J���ʤkHP��p�`��9/=��/!GL�պ��M:.���m���v�G����d�C���oj�8�S?e�XW�o�a!D`�lL0���H!ѡ7���u�a��Ǝ�Qu�k�W��0���d�`�k-��S����3�DX���E���0L�EA����2��2�+xax��l���h�4T��d۾ 0�� �(�۰h`���$�@TIav��W��	6���1�?�b�Q�2�c��>:&�`t�Z�������#��)߽�6��>��M����K�/ۣ�5�U(؄�ؿe#*Uģ��3󚞛{����+��8��q���
�6P2H���)0����d�ܛ@�����}�<��$P�����5�Ά�%��p�0틜jc�Ó�+��SX��-��D��
=n�lяu��y�S0��y%��p٘V���,"#�Uy�Kk������!(6��ߴ�s��P����u����s�6|7�uT1�$�u	a��6$~�5t[6��k�w08��R��Q��\څF�x�p�,�E~�T�YiD"ދ<��q�����ft��!�ࢧ���94��pK��������^�5&�O$:E��c�`x���`'�u�^��ojw�� vM�4���2&�B!xÏ��9�Xy6&M��#k-9O�� ����.(#�fQ�@㐁�@�>���Q�)��S=��
�|�붌@S�3CUc����C��D/�d��&���ߛ�#��{Z�4$=�҃K8ǵQ4�n�k��yq.�5㛹���W]}�2��������<#BAB���ȍNmE�!���q���R��aev�uh�<SE��(nL���ID��9���![�����/H���K[�N��Ftв���ko��"�`�K� �]��>�CP�n�˛��x��zI8��kʬ�[<��M��ay���M�]4=���(�^�H6�Y![��n&Yt+�Yi�S���"/ü��\��oJ��r����=�1�X��-��^�U�&P+�s"�O.�(:J�O�a����\]�,X�Al�Eɟm��3E��xۀ�>b,@���a��7�|.�0�{�"V]��Ӧ���e��꘦=k�`��Drתz��Bkq�n�.J�N#]��v�hCMǅ	��
!$�\�3��M5_���o�&�ԃ����9��;���P|���6�ǥ�����x�[�	��h�\t\���Z'f��ɭ>��wB�M�µ���)��GC�v�澠9�r��r��-n.��ؼ#�E�g5����uav)�~��&|k������xC�-߀kbM�f��r�,�R/ �d�����H��=�m4�����֬�/�y���-k�鵦\�{<^>N�pIzO�pc�tg����Ӣ�vSj�*X�Q�غ���栞���u����7�\�;=M�Y���ȏ������>�vy��I ����΀^V%���F�+�&�E��"m[�X8��[���E�����V�b|N\n̟�$�;�+�G�y�j쪶�#�8�+�D�� ]p���4+3��U|�yk���Uふ��d �k⡭i����Z��(�s�4�*#�- Oa�����U�a��s��J�Y����`�}j͋��Y��.��ki��͌4�k��.�5r+Va0sҞ���p�OKC��R�N/hx�6\[��f�C]�t�e�r��O�$�?t���:���]��G�W���^�=)
�2�{�YZ=��z�j^vJ"-���Ѝ�t^nF^T�'���C2�DC�zs'!G12~X�g���N  /����5 �	Tp�%�;��&"���� �(�-��nhk�?趾X�Z�ꯛ�C*�4#��i���v2�rh���#�k��[��F�-��9H�x��z�E9g����2FwJ0Qb�ٸ�Q�D��?fߋ,Q7��ra*�_B!,���ЄȓK�W6��V��˯�����E���"ϑ#~ы��N�O?���|�jy���Z����h^�c,j��L�{3 �|O���egɊ|���a�R�s^��6��\��&��v��Oy*8���~���T�]��RNV�}��[�f�r����d�o��|4�O�p�����NxV[�=q���42ݛƨ���������]�ꈖ���<w��I��o�Nf|�wV�,fk��'?|�
�/}�rD%0t�VQuJj-��SOi@��򝯳�q/�vz�C5�va���"v��.�i-��u��h���C O�"ц�Rw{0��6y�5�}�9��w~Z��C?����f��r�&�,_���1���9�����^������H.5���)]���K �e'Zʽ�4o�u0"6$��В�2!=K*c�!w�/��ͻW;O�����ß���(���t�ʨ�:��,|� 󄧖){�ԣ�(�7�o�3�*%�?��ԑ5qNn��Q/RH�ʏ�zҒ�l�ii�{ŧ�+�����+���y�M���h��N(K~�vt���:(#��#�0W!�����G���S��&�����l'2�i�.�#��<���BAL���랰�Q��v����$�cc=�֊Q��>Ŗu��e0	%<&I�9aӶW8���+�*�C09,Kc��s.��c1��Qn�nc�۾N�X�y�'�T�4?k���u�wn���9M��|�g{°}��V��ْ�9�f崧T���un��B<_�ų)8j�1�?�-�^oo�����B0�ǥ��(�ݝ�į��w��UC���u��쨱1����Q�^�S�0�Y��~e�-��4�,�t��O@m����2�M4�qj�l{���ЁNݮ^�M&|XX���d��ǲ���L!9Z%�݊��@/�'�n��fB���zq���O����>`M��Z'.��1EI4�t�$S
�HA�Sg�{�C��;[c�]�F��"�j�W��L��u����w}��*�CT/0��bz��V;�A��Yl�%��cTӅ�Q̻h&�1U�g�y�e�E:%�[_vN�{�N������J��Yn�Ԛ����F������+�F��:��ȭ������0<�n(òO��<E���,r!;0u"U���,��>{!v8��fH��
�D.�ۈ����y��M��ǒ��;|�����"w#td4��SCh��	���T/s4�����N��g�����B����6P��<��@�l��w�a+$��Ϡ�A�)��h�֥mfꝌ��a���6T��T����BKf�e{r}�5��ۜ����B�S=5�(kB�	�3�k�H��j���8(���D$�g�u3�@5"�ЭU0>�X�\��Q�9�%�����I�4�F�m��|o�+�\�>͙3
;�K�i#d�^�RBn�}��o";����o���h�@a�~|�;Gix���kCVXd�l)'�q��gs�J�U�j9�
���L!)]��O�V�����zn�A�{�b��q��`p���.�7������͸�4׋_�\��vĈ�TT�ż|#��1v��1��S>E7���7[[�& �xRd) ��KfˢK�umk<.�I��4�p��9�Wv����CJ$��BHg�,F�W�t��p�����<�<��\-��=��-	���H�@�!�m�/et�x2��oq�m�\��C�G.]\p���G_B8��7fZu���}諠��}�]e�vn8������q���\�|ؐ�#ȭM��my��~vzg�RxB�wfx�}<{�i�j�5���U�ko�D���Ĺ��חbѡ��A�X��,>��|(b��,Zh���Ճ��p�6E
��;�ֺ�b�R��˫��_����;So���<�bǌ|��b�����k�g)���t��f���P�%}�k�O�͆D�F�؈6��Z)DD�h>�}��4�T3KH'7*�_焋�M���dL�	1�6O4�P/~����L��.�L�^EX)Y���Q	6۲��(r��ε�!���;�Z��/��	E��<�/M�g�M����EŔ汛��!��`1��̏�4���G�v=�a���8d\�i�n�,�kyxFP��@�H�U�Q�'��a'}7�a�z��3�&f!��֌@�n��է�i�*%�<p�2J�u�t�}���x���yC�����M��<��+�OL�y[soL�B���O^#�̳�6�t�[�Ǧ�2<���o'�)��l��>��@����ɟ�����
�� X���1���0�(k��M7��$����K�Ar��8���[�DX�ƚ<g�L�8��!�lxe��T	e,i�#��N+`��检�-]��y��>6���[��(�B�Z� �2��K��@d�gԁ�gh�O#��!7���i���b��\ M�8��9�ȑݯ�4Ae�D��o������!�>v_Ha�.N��l�;�%�!_:D;vM�C5�(��H��p�����Ef��w��`�0֐��R4�e��"҃��&�qV_`TN��5�9��_�qt<�L��rDL\)�n� ��\7�2B�l��Jp8�sqi�݁�f���4�f�-6�����үJ�s���L-� ܒ��u�Ӹ���r�d�qJM��=�s@��q}�4��Gj��@u��^�&8�5aj��Q���B'��=ս�V�éd�"��_��x������\�ӆ��G:�i���w�a �a�d�z�$z�j�`��h���K輿~��[l�O4�s���˕��TPQ� �4�Q�~�q�B��i���[�3�x�3R���o���:}Nk��n �W�ȥ�fF��j��tMv"j'���ț�����TN�|�b'��s�9_G�G�lV���ta�G7X?���ZL�����=�>����9U!�a+�E���BZ��h�i}��S~��p6��Ƣm��k]�ziGr4��4y'2�R�G�Fma�H������~b�}��u	#@�! .�+�y#���D��b���˼��yCz�#�Ll��1�Bo��%��e��v=,=MD����rb ! tP'�[�W��\��yD�_��8�tS9
������1�Y�S�.%LG���_��u�u27v��*� ?~�Ol�N]\�� ~fӇ���ٓ/S?E���Dm���4 ]Ƈ�����-S�Z���P$�����'p\�/.��D0��� ���]�ƞP��w|W^��"� {Ou�����:�tɡC�����k�X�X�8}�ő]��"aQ�B~�ߋ��;ݘ&DøY����A���9�-��O��,�*�A�������j�A�o�T�{������x������|���`�NPx�!�p�&Z:I��_�c3h5�9�$)1#�;�Q�5��f6��p#��6k�#^�v�&JeT^6������!�����(]�'�ƾ�|���1�]k��U��eڑ&����G�(���S��L�=�#z������O���뭘�1��	Uǧ��cn�Gw �oE��fBNa�q]��e�EpYo�<�Ï�Cyֈk�O��e�1VH�݌DM4�W�;3�Z0g�Wo}6ہ#�%�A��,!�l$�Q8O�A�>�p��&T��P�셚m�?8�o�#	�^;P%�s
�^��D߬�,g�]$�EX���FOE�e7�Y+=�~ЁZę^��E�10�4v����>��0�A�f���V`aS-�,��u>�Tȗ�2���`� �l��!ِ�fG����N�#[~�(ǇP��Uat'����a'�{����xe�qYDo��̦xB:v��O{Š�v�h7ax�7#�y�疵��J��������e~%�h]W���A黾D��d�h_y'��oTH�Wy�}`����E3�F�i޷)R�
d3x�G��3���V���
Q-/Sb?Od���(mh�0����6M@�Y�Q'��M�wq[9�<'%�E����(�����O�J�Y1���'�̜h�s9��m��.��p�ȼ���4�f��Di�f��x�w`I��犤q	D|��I�]ŋq��JY�T]��qRߠ��k�G����7�����-NL(�~ҹ�)�w(k�����ޔ#���ޕ����M�h��,+ D>GP�V)R[9�w_�*Q櫺�]u�R���\���0|$���Pxf벫`����U5#1?(���� �-��Òtm���M|Y\��X��l��ޔcf5)E����8�����?��Y�e�t4�aW����ض�F�0�Y�5�{*g���ii�/�D���kELD��v�(�?j4�P�8H��p��]������m��-h�7��uX(����1X����_#�;�s�[��/n#N`t�"�%�Q<!d?�����?��rx�yA=�h����+ci]N��=���EËŮ�Rm��w22��T_���,�������LÈ^(|[/J�4B�^�h(ReyZ�4�� :�u�e�U�ґ�Q���S���$AI��t�y�ǆ���w���c�6�f�P�[��6�j.�^I�$�9J�MV�{ܮ"���yG�oɘ��(|��2LT��6�V.�]|o�Y�29YS^�yg�� Q�MT����w�����\��������gDh��&�q%z��~y��K۰ R|�	1��Pi�q���Z�?9$���%FHk��H&��-]��M� ^�8��#����ʦ�K��`s8�!c:Ơ��;��B
�m��� ��4���kr�w2�m���<W�]�כ�`{�(��U�X�������{����C1-n�x֣r�'w<�d9�${��qn8����h'��~{�A;/�%U����6���^;"�~W�����"^H�73�*�Q����2��= ���=�_J�?�1�$�yd��?,�����ڀ���"l;��y�m�1>+?E酫Ur-y0I۳�̬�CIq���4؃ ��1�������y1Z��m��/�5��Qy?��鰬��X��x�V��[�ږ$�O(ʛ�ZPq��b�)�9�U����TLGG��I��Ѱ��}��V��h@���X�>=w6��b:*��-*ŏԕ�ߣ]��3�����?���cq\��D�˼��vF:�Z/y +�.�PK.����yE���;�v��d�"��~ 1���0�{�]C��ad�9����t�y�b��.��-ȳkX����Tb|ShD7B@%�/F&�I�1�Ԋ��˺(�U3���?	B��MCqSK�0&�}�ףRS��i�`.ƴ-S���d�����[�x�U���(:�-�@����]���9�"�T��!�2�^���+������Rw^���V"�
#6���l�"5-�&�I{ef�wX;+���;6>1��-6����L���jڃV[����}^��y�$;���Xz��*6&?b pU\b�,b�YODZ5B�{�^a��D�JZ2�X�t���+�l�ǚ�X$�����]���H�g$��5��U�c�'
�ad�?�H�:���Ǜ�>t7Fᓐ��Z�9����֯_�~t`��,k���e�ڭ|���n�cI���u��'����:��Q�LJZ{�׏�@Q��՘���r�Ѐ��1cd)��0=��R�������A�ң��b^�ӆ<jcB��V�=���ξ��/���rwǤGO(�~�ށnI�`㮝MC
L;'���ѭ�!��n�%�sU���#�=2+N��"%�6d��-���A�Xڲ�Ʋ�Ȟ��[fi(�F0T�C(�H��'ld}�_�}�9�,?���g��w��6�?������^��sռTEk�~|�ܵטG��Cyn��N��S5!|m���õJ�1EA�>�ހ������Ut;.����T��xFu%s����^1p(#�Gɮ�^�x��h�@xwA���W�۫B���b��"��5[���-��ܗ�A��	/����9j���y�m�6�g�����ɥ�: ��i�5)��h4*+(�( ލ�yhC���-�X9�j��@sZ4jVKAY6�nP����5O�rfl������ʁX	?��3�3��,s��L�Z}��X���Q�ք�����Ў�r�W��*�S/�:fv�a&zqah�Vb�Eڼ����"��9�Ez��:�2��B��.r����_�_q��AgӒ�o�� [�FPD;Ѽ���<�y5:�m�jK~*��E!�E��������~
�o�����p��i�y�m.q�Q�s9�S"����X6:�����4p��<e�����?��ɬM�	R���g�![����������b'^��~:흠@N�հ2���h�	 �̧5�I���w|��ˮ���nJׂ|�f~���X\nt��vx����6�H��(�z�1�':����\S	�Z�>1z٢�=Q��Ϟt/:�η$jȉ|�;Ls̖>'���<ɣ<�*�V*N��CP,�F?�<���6�����,�&|�g�*�_5u	�O�d�	��fBƽ7�0!�c@���޾�����D�����j	�|�.������@��jC�%�Ά٠��C�c�5��X��ӝK@f��uF(�V�M�Tx�4ລFZ5��h}�3�M2�$�0�O������|(�$?�|�;X�4ޔ�Y]�@��M��k*覈zOL���'����F��W̬�}�?Z�91�Ė���W�#�@�~��=jr�Ͽ#��Z�q��ܫ��rj.Ŝ.�j�B�m53����t�*{���Z��0��Y�S=+�&�R/~�ƍ�k��!D�*U�hų��o�i_^���*.��l�mK1�n��a��� 9!��7�?ey���'0>��tt��/���o�e��&����a :���[D�.c+r�_C��f(��s�$������ּ�OΎ-<��;�ɟ�G�E��6w�٣�f7>42)�~dJ@?7
��:�:^�����HǞ
�q�� 5w�F�x�3�e$ �t�h��a����Y�f�����綼-7�,���	�D�jsQ��A�`�H�L �m;���Ŵ��r0!������|��m�l�#`�r��r����9��W�vl���B�������b�3 �C2�q9`�������' QD��0�ȵŅЉ�pe��"v+|ѱku1K`a 1J�SA�3eGk�,�1�O1y�ψ��M�*L%7����u��`
��|�`���4Rn����U''����@�P
��"%W+�]��{RtFX!���`�nmc��eR�
aU�GzΆ>�AX-� @���\�mG�Pԙ�����2zV�m���j�<�o�x��Ń�y�m=���Xo����/�ߧ����V�>z�g X����5�V��_<��(8M/��m�y��t��LF�����?iЩ��+���%=p���r���Jܫ�� �]��}g� ''�Q��c1�3qI�����g8�y֢�&�l "_��u+)o4��z�����P�C�&�I�z��U��Gc��
@����9��$Y�@ɾ��Z?����j�%)vx>������u���t��Ă'�s��&%���_��z�% �zh`5�ȻK�4�iw��PN��Ս�!����1����9˝���-T]�5��Ez��*�L	)�������ϑ�i�1�K���\����4q@�-������A����h�2��I:֢)�h�b\U�w���C�5Gb!������e� 3����ၓq�'��Ӿ���.7;?Ǯ��^Z��H��Se<~>�����[��uhfŞ�l�kR��!��m��XE2 >�^��̀ݛ	�M��c�O����< ��;<2�xS]#���N���?���bg�0�5�-d���{��>0 ��I�V}��?ٕ"�(`��]F1H�WжD��b^w�r���DUY��J�^v4���6XT��[��bˇF�+�"b�}��J`��06�yl�ŊA+n��Ed'�OsvА޷ۅ�w(ո�K����
�
(;H19�T���S��ۗ����(�,D(��c�
v��4�G��f�w�$�"A�RD�$���j��0�y邮l��W��@�75����t��tVg%��S�!���&��y:�t��:~�v���
Q�4���y��ibv��EQ�r�fӽ7R�Yk������/�����+��W侥R/��N�SP�g����>��&�N_x��_	g�����D�S�-��#Z,ՖD=|�z��%0�d����7�w���;CN�d���T��~���Ľsʃ/�L���k�Њ| e��i��("X��AlE��-� ���A��j6�Y��P�8��h;tE���In�.�<&��ꖝHv��*��hƾLE�����2=�fR��g��n�qU��5���:�
붉����K��3ٗ�o��X����1ݧ�邳�3n��$Y|:db��gûa��p�}��a
l��N �é���qD4�܄f�g�I���i6��N��U���#�_����|m~"�� 9�F�C��g��6L�Tڧ�#j%I]��g.�=�k�X���-��0��W���h�X�4�7��
���ha
�&�O\�H�C���0/����Z�����-