-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
--pragma protect begin_protected
--pragma protect encrypt_agent="NCPROTECT"
--pragma protect encrypt_agent_info="Encrypted using API"
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
--pragma protect key_method=RSA
--pragma protect key_block
TycRVtzYeYz+CO7JZg5uEv90e8udUgJ1LDe4WFrPpJe2o62ubD36f36LEXYpGUn6
ifwPUu0Rt1wa9d5OZV16uuNgXD7UmZXDtfBLqHj4ovFE7sQFWohXDQccqDtHsHDk
Nqt+G75FMf2r0K0UCtbO0EDE8Wj59OVRjX1pZvwYQ//VabZu2qgJ6rqN/utMjiai
CKOnfHpKkzeBhIM8kAkByy2YH7FQgC8+duwhwVDPH+Mlkj3+BiCInrJbpIm/uQyf
9AKoKuDQg8RuGnpodzz7ChUpJrn9rSXQV71YwRi7F9HZVAg3dKziHqSAJYMDllgR
OIJfAZEqH1D6EqiWcKDSxg==
--pragma protect end_key_block
--pragma protect digest_block
erTIssKPJXOHUzTYoNWfJ8w+hy0=
--pragma protect end_digest_block
--pragma protect data_block
Mxe6nMt0c7BwTlsM2JqOxpIHAatD406G2DIu436/XQbFk8WGuCkfZ2+TTBkH2UpD
7EoZBCfshUh2I6DUk0OkI8zo99ioG494cxZpRlkzDxopH+p8e66GXVaBkmIhzZlk
hb1Nsslvc61gbTwgSJAiFbtn65aZ1JsC7Ln7YKjmDSJHGNy35oD+rM2Cotk8+Xq6
qvrS1zOl5QkBxCN4giTl4wj0oIEB2k8+40/WYENV5zIp/mlKatltdOJfuU2ONs7H
GGkgmDqHOGXcKa2W4J2w0l9DqqbO08VwDWRAblYHwFKy1XnHVcKm6qZn7n9vcBPT
nCmiW0gKvI2XsqH3mEHIfYk6lvCnXyx1cU8e5cm24m7zcNhdTfGSN561pWytkIJ8
eRbeAkuBW2jUvkKaFfEQ7JD2LkkrifYCJ3XR23k4JcBfMfD583iWloSWDiLhXvHa
cUDTOLNxXmzWQ1+QKbCN+31dBFruoJGxPtLJBFrn1i8X4G0WaGQuVWHJ9bdG/+Jh
7RW7BkkJ6HRSuttLXYqaVCFXNo1aCsGFcGqiqwccKpwftPqYL2a8u3tKLe3h1xrP
Nbz8/8uW1CM/J5JNt2Zex5zHEuWw7NCxNJmXrxRgMxa294gHxROtDZLvJUf21lkm
90SqRlEWFDg9w/gSvnKup/2hseej0VJTTNY3ZPc4wwGuLY0n97EPrvOhLV+Uzz0F
89lGrpC7Ke1VntEE1CzGRPidKh7Hw+RrZ4W+SXfCKsUlkcrqYWIM9EaSfz9LO4Vk
BFzOYm0wY/haN3F/PF0INminmsV8kmnET2SrAXzDIPp2kSUVmTJHMWpxW0/Wylgg
hOm44qSFW0rLpdmsuk4aHQIDz2wc3AsIHvIoRyENEQuG4xYzqn4lkfJ1VepeJOB2
2Mpsa0/tgcFi+oykkdxvQ1IHnwnojFYPUYFhxnNQhdb1JkjqAvSvfxJHv+uEH5IG
M2WpH21qNIGy2BWpIa7pbJDB7XPFjtuR9eNwhWRlqfAeL8MDljUS0Y/0T3NljmSv
y9ngfjhPiZPUm5KZPcAuzUg3E7my8oHE9P64K+yBjqxsO+UbDnZZvuqNLEJU2x4w
M9bz3j2XX2lZGDFGEF4Jj6gAAsx/uA+Yx4EuLIlmQoIkj+ZLdQcsYrEOZyeVYqpO
narWg4XsIKwwpC2ZNpHzC/dUSjRpjzSsm5euQlXoaY62Ayq0QK0cI2g3FGatSGKe
vrjV7F568N8w5MezXrMIW4c+4U5TkyD0v2WMqV3l/LqgaUDmomDotqdOnY7aZwIL
XL1M9b7dpc+thlA0OsFR7YT8aaM1/Ib4RTn5L/MiOTCTJOwvbUloGMDwlYSfOLtf
y6WraGnzMth8U2q2u2Ed3mJgRisfXVKpwCaVfD7034+po/DtNiq8rjLQoXl+tppv
SF0gMDlO99iQA6aRIdEckBIvrRzzs6Oq6SgLjiwFMrUacXskZnhtjciHUNj5fvvP
+pvBQsRR1QmC+cp102uUJDIBNbKsxDteDdzrYUFag+JZX6Ok+9rX5HddgLhUgGVd
Gi66odpf/BzC512hEF5Nw88+sekK/PbrvS61dTZ7OA6sv8d0cDiVjs3kB/AP9OGg
bLbHc/pDAyczWeEbi5AqrdHwNitn5k/l+Io1i3fwQ8c/LgCS1wf3oMiiv0RQItKL
0LYjBWNG0XB4kzNHyXQs0o/kmO7jLXlt5RqemXnwUcXUbc3XTq3LE/XFEsE/Dq2s
ary1WypfQ2fUjOvyA3x3XmPu/RrWf7J3K5yNK+Q7VVzqG2PuYUybjmpEHjgQnWVp
2cVB0FGZMBu7g0Jc81f/c1uGjqhokJFqxgpcMAGIGmz41VywhlvS+ZFkY/ZB5REU
LN70hK5s0angN7Lmf0V2F3jpt5IAyATJRjd4R8OywyciUIx/DWQTdxA2U7fNSK0P
nqoWXmbtJ2LdT4VzcogaZJ4+74re20aa6l6zxGH9fiWQt4Cra4EZLeV1Swfk66Tc
3HyQKZFWpygjssQ2pfWPLO98Mlj2+80qrXeyU+rFQyFaKG0tZ5/tFVdlkRd5v0NY
IO/Q2djJHECGiOvNHu4x8vNhabBgaMDmBc5jAw2QpTR25LyF3QswWh6N8RHX2RxF
VB2dH3vDl0Z9ZxEFipv/vEJQHVOhLaboFGUw81O7Ou8zTjqyFBxhMKps00HwS0rR
I3Q3lLr5CT8Z0ym8gV7XLaNuphGQ+7t2zI2H6QU1sZuATeX9/ebIQP+JbJeyDn0U
q+9KZsBcsRIKKa2LVu+NFu0aKUFql7SsmBxponjR5egQ864hKy9vs9wAwHDcK4yu
wDlKWsxlfH22nAZ8dphm6H22J3XFopkMxewqeKvMSqIvHPVhjl7Y/fxzOkjA88di
lzinB6Mn+2ehGQlhuA/5pdPWhM6zqGHRcgC96OsSz3QLwMfJ7Ns+XJI6iXdgKgZY
fnAn4ADTTyorQVZ80hKBeYqjlY8Fn1JPY4AUzW1v0u0f8oT+TbJPy3Il659LMTZ6
R3ush8edZdsldbC0PS0k1IaacsXfoXazfmsY53gRA7R/FHUKV/FqJ4xoXGqPhVXC
xrTo3wSr4bgH1rW5yL4cBCHNzglL5KxuOafj31g6bDl5h+Zwhr/Z+5jnRwSz3ZTR
HdgexxxSpNtzmYV1W2apuyW/lqN/xgKlZiWG33FJqHf+6eDR87QzQlKr3gy8bds+
zGvgWygxDO2dZxv8m4zFTDBd1lz3tnmvB7pNIhxMKaNaVxPJTmo/4twqpzP8FK84
WNA6DxDN2p1ma8d0ZogzyeT5pD2WMSyucy5ckLoeGSwcl8NMSIW2KqGpGZzouzKs
Z4YYhx6I3zqJ/OniKvY2uyatO+d3NlZT13Ilxg6o6D4HfJg7uwrE0N2+yaQcDqWJ
lvt/BM3wUPsfC9iZT8lLNrAPLdRZmsMZ8GM81E4H8phPXAkrkveHAXB4DuewVWvr
ruYJux098T2P9o4aSFqg7HlrY+l1C+RqDeq0nO1guaqbrlS0H5bd06XCXOvhLP/i
ZhB8PLrrq42cEAl6tQUvZPHeNUGITPO70Xc8UIonCNUC4NgPp/bbL9R8j6oKkGXC
1R970EkpHUHZ+74bn1badRWBEeNaxDZR8tiD+gNKZSjM3RZDw6ghJQCyLfwLuktL
p4WI0Iy8CQ7OiGgSyxsK5i5hwDuQKAskTgv2K1QtprKeXMrEWAlfM6hDP21IY65f
G38GNlzT5VuRUwLlDq96RE9hTz8PK1J7/0A7ui9EYc3GWCt1OzKjYaUyVB6dhxd/
ige6S8DaNyd3QBwWvb6KfmGbhYECn5bGDNYavCh+OXuTYFqE61bI94J6/SVdJsKh
OX1i6UojFEITcPLGtV5brt4NhMb2QIAM41UrMgm3RL/6kO3sGAc8auJFbuXNBhHC
bjNmi69QUQ1g5sIn25PlNs7r8CsTkA/PVqWi5PWQ0KN5SLsj32mybW6/TiLplRQs
nesLawHn2gvo8WcQPQGhbsF44r23tOsBuUSImCfAPOdTPdk4FBWVIdpGoii/SoVE
afP3K2VUFi54LAhLp72O3v9a4x3Ia6J7HlSCq8SYXNe0BuiGOKfriEPZn/4bFXyw
lWU+4xmndOSE6r/oL+yoMxqx2VvXuFeNITXK+lfajrrs3DA4qRYhvwqvfNyi8f8V
phHbxtMlIIXRgei2GGianG0g6ceIaOmbpy22SdixyKL8bGmaZLYxgP1GdAdMZq+t
U04qYKIpIXVyl+twlGS8+n7zivxIO1MIEOnTr3QEfctrGyvVT2MhZ6UMPmm7LC4B
ZSIFepstmI9V/4hoERu/JihiB0dlL2RzDxqZCeJeLU5rvjcEqHdhqtVds05/hjKp
jV+Axt3ed/PXnScv51KtHubnmrrBetQ4Pl1ocRJf/zPIYGs1Eww/TxeKWnEHy25D
zvO9oq18HY4gnu+v+tmDSKg1S1rBUbtenJkpSz1CG0dCMb3tGOfcRjE5l/rcfF9U
dO8bIiAMja1K7rs7LXNBDONnVdl37deMlAynkcHNBQn0Ozm1XdLybF9/W8h8q9ks
SCR2Ro4r0h/+ye8laFqpJeEYbkjl83ovopnG5B2IatDgUrdxRicSuni7QlvrgD0n
zbJRTpL1YEUU7UhxeRiGVaFIrmBpfRLT8wgojFqunE6PINOVCFEUh0wTjlvuc7c8
X6JrnUM7Ypi21NibF+BG3RIb6dh5kV5Dv7Pzml7UlhitYY70AhupumNrPVVT7sEh
F2c0bzBlx0sMjBdSBgydTMSSqxEOBUHmyHDwjL8R6fJq0YjFQeOcbi6xgPoA5qfn
e5pTKM/VMVICFrcu//mhBnlADs94ENfaRhT9GKoo+TYJ634OgFjnwKTnsIuLsb8m
qywDJ60ioKEjlXenA/71IajuyeojClkM01WzluI7uagbOZoHFaWLEqL+Po/Yygmu
JTKLBCauhsfjB7r+EOMwODxEuHC801FXV2gTWzeOnJJ8TvKWZw9AYMqpsFoqVi4y
Ch0g5uVdG8Xp06ymv89dzHAyjsBXFFhbe6K/pMlRiYIAD4KQdI/TVwtDO+hXUOGA
Xc5i40FAO4fzv7taxnuAqVRYL84eKNB8g4kRSUZGjvjGdgz75bXAXP7FUypn9yxd
Hwq/yWlp+lmCJdB0s8Vfc9eZYTS3gAObUpMTxL16d+Y84izAUvKoKNxLXLIsL4xG
t832CAwlUqEWFhCQwUPC6qL22JZNH0p97Fob/mZcd6tqlg1QxS9qKaxW1WMqHVsI
6FmgGikQyX+boXxTvDcXZbxPaTSaoUPdNqQSzcUJI2MAnBT9ZqtSP1PbHN9i8NGS
sBiSalqT7ipDjOySG+sHKOpqEIB1T27FXHxYaHSCP5TI728ZLtAMk3Bw8/dk7yBT
+D54K312f3xrkFO6ov+9z+abqxD2yrNLKZa0P1TnSvG/+mtTMrPmk1/z9nbKjx5f
cQaaTPPe/CI8d5FGaNaHPDdj35LTSw8hJd3j8IKQUqSsbwyBDuC0/Pb1oFvKq6Rq
PPy5jnRmxQ+8kxZlVVjxt5f0r8LmMJtZpwpPK3lcMAN+B98uvywCGt5IuFEuT7Zg
SkNPOsV2uMsqJ9uXLYzG7MmdCcOavbLn0/H8IrbO9z+woFB8xqXXg0zo6ikALUAZ
aUFpBgkagzS+fSjN9dJQj/oRzskek9y5xCyKhVu8p8iIDo1rv6PDyZ876neQ33jG
WOSyR6CBaQ+6MsKtGGoagPICUtjhw0fmaRs6oqMj9qmVSbP65MUVp9Mz9PdMcneL
XXjXJmloQ+S0nIXvv5qOPrkEaE+6NNZhn9/92K2DQVIZMnNbkRcczD+AH9ttI63U
vftYVGF0JOBTBpDcJ1HBX4qBn1NPJpd5WrO3aroYzdC/0CtZt9e1FTO4pAOkCagT
7CcqYXmwc2SosX6gaxjRQA6bh/DjTRlmKhAJ/Kei+hFCigjq1wjm5rtHYWLv7wtw
ks9XDssr71D5eEkPopQKJEbplTSiLFn4xC2HdQV8eBLcuPBC5qWyQDmWwsHkhblG
UTULqD2lWoBrE/gA3wAl9jXs3r64/1nGJfwiuzyP4Cc8nbtxCzXZYa+Us95ne67+
BhnA1IF5EKySpXHTvW+OrZB/P5leMjtwfmBCw1fREnWY4TO2wA1HCVWPrxAhXWQG
9qGiV53KglEOqkN+J2PkGV4monLUl0IjxSzNBKsQCsIunKQO7PLSxd9ziS+F4OfK
iwbVnubLa0JBTZ8XyiCzPG71/2NwW9xYGshmTPqJcoO/T1mkyURaWBTcCkOGw65N
oG4jQVfPs+hkag8ezvpDVC8SaM8L4XU3MnZcv5Yko2pTfQz/V47+AB7Ld0ugXyJP
VDKE8hnzEAAEvh8CeYua7d0dfL+ypgq8tiHMXB8KlQhljI2+ymq+HwGqTYObwBUL
K+bvQAMa16CKn/fm3uU85eRYS98lbp4kXba4BIbHchq+TDTp9OsPM5OHIf6z4sFz
SWH3wED++XvohzS8X17BEyl9JnPH6FO7nVe1r/k2mB/7kEP75fSX10KtZK16jSuy
au2ChJJexLmUnG4AUn12Otd3xSSz+CTBBAt4NoFXe02Hox/JArx2jIgl8ps7+Hl7
doe7oD0VzGlEaqvKMh+i/hfAIRBOZDwRqrJ3HC8dvFhaOVo0ttR6MoJPPMIGfPhO
EWGJTeE1xDYv4IjjHrqtETBmOhBTkax8mcFjFNZhVDv1TVEizZ+yffr9UWSIKksC
GTDLUAw5oR5VRmhpBWb1lpXBpfuXjPBpL2wWZDcMqOtzUfbsWiaYmiftZOexZ3pj
0kvV3zV5TljrNQfCPBEnHqMQ3J8gPXZ2ebQQmU+yrwXxe4MT7RGlM76ilJ0EsJ0r
n/kwq3Xbu2Qn7o2SW4wwd/gZKvg2KntmxEQCaGRwYZQ8m7Bctuzm5tVCuBfhQAdl
iV3qEzWQ6h+dTIUpjUiwOHgzvVZhkHElC4//3cq6k7SDEjiyEopvUtvKBxsehdJR
oXFLVwnydVYX4nOTjg/EpNpYoLiqNOssFVlNb2QpFTe5q3EY5WL6ScFhn8oRezLJ
hK0bhF2DPF0G+yDLaPNtSL9+CjbNIEWM+2zfRZhOni/fVlWvy/oGMlc8K1kx4+/E
UA4f588IX6LWpuGK1HZ+RjKtHMmza22dTUgszAE5zTeX0tthhYzJH2DHlCBnFUhW
/3bcINibfghPtAyFPmJp9EJ2V9I+1wwpAzb0PZjiqUTDeByn+/VekPSQkyX562Xa
4HcxBTOfG7bnjW4rSPqvV6QkWQgjGpk6z0eBS3H5FKQcLHvR2fladc2YOs9PoRzg
EsB2p1D52/CGrYwlzJSj/UUK6wAAI9L4+dpJmrPvnJs83cm2+GCQCTrl/PFsHB3Y
hg832iZoKXy7CPcVeYA8zSkho5l+uXRuXSZzL26QamxpUH5H7ZquyQEYQ7f+Vq6L
Ewy+VEpVkPYlMmQDPQD+99786mNsIVBemfwYvPU6vBReaRaPIXctT/tdlaE4Hs37
5/rIzjEjdsCoSEkYv2250pIqwaJqdxkdL+kZ837gqLPts8f16mUp30FQ3/CWr47r
dW204BC/YNPACK1ostMgkWNOffq04I4442MrwAFs/GdEig+L4UCs223ZWCDrmfz1
cmvhKsXGT9IrkSbQbAWq1dOxV+46aMNyoeU7IPd8W3MeCIFyabjuUDQJ50uUhmTP
brz3mj5DjmHnYzokZg+W/ZbUhvNPTFLC5KjqDh8UM8ambMqNJrVAsUtRVCr+SzGS
057Liv1zojf1Xgq7SkrFvpIyneHTp0c0W5Je4b+mD1NLIgZXmkKgdEOERKmEInz1
XQSQRt+9fWc3N2ySt+ajWQDYS5bZU+hAvmEvh3a4dy9P91MDDnPMHN/1PuBgt+DW
EBYBD5SbQjoZlWGlXp2DABgvuaOH+Xqfz8ffaYIbLeoki6MYSW2NsH9ZrBOePN6v
8MiWfMFKwILfstDgeAR4c8G+0GUoWh3v1DX1a6mH/rVjIv+8s/QC8gOkI0oUvCw4
R9VvkiQJpZHoa7iJOPMB4Jv9smxdq6ahA8xxH69f1kQzzWvk1hppb8fi9DY+nAXB
lwfijLI3KD+Ickc5clfvVyEVqz9EgZ12Rbl1coeKSv0f8Fb5pvq6qo0DpKpXCa15
cmXNckgCJ41OJ5vCrv5+XtRZ6s+Nu7LN1tjJ2GjT8apAnheqorJ9z8+BA6kV0/Od
TE17xVvbOiUXgW/ETXQ65gF3OyDBTUvgjKdqJ/r8tQBU4dbDnWjGI7A65JZaoTiy
SdtJi5bUX+o+gaQ4/JupzM847bfcUS3PfzXjLY4RDePX4NkdeFxmVDXBhHi4IZOl
3QZCri9BjKnNHpLWYIWipI1DUTfkqA9PgGl849yL/0s5WKU0CZXVnPfmYwtI8aXI
5mvkaeiWGhLhuWmO+DUTvKtR5PfZgzKjWMes0vyiL4LHRLI/BvD4UgDUZeqb30c9
N5IWeeD0M1djsSMDS9wRVRul08ao7Ug2cUnQGFtKdlo5TE48GYXz4k9TceP5ez9F
vjNE3fjB/pzO4ShkEe/4LRoU4u+2nc71JEe4x02Lm0bJZzwgTTJ3CSvn4D8ES3yj
b2lCX+YWDfQFpUIjZl6LpH3bwzmtwpIZpnznhx4+s7v1A2UsBHwnTdR63+7M4Gye
gYDTBNItTjDFEq3KRqsS9eGGusQjiyIheRTuRSmgn5MFQ1k/UcRX05EbBvmrQK56
Ds3JFOSm5F4wpEmRs49cZUi1nifOD7618/gW/hYvtyoH/qb4W+leHiCSKgxw6Lyk
T+QKQJaODsPjEUedVaO3tKG1pieqnlfUVERjqJwXADwKJqQBRSvUip5RyNblR1Rm
1YH8oKF8RgH6Hf5WbQFaz5QmGKhPB1oWg7lwiTSZs1mnmasGegGw8mUa/Q4G48eN
pKVkyyFf4wjpAruanok5PaiEq3u0KWRVMjVuLoMpSI8=
--pragma protect end_data_block
--pragma protect digest_block
B58DmZ0PDGIEnt9gpGKRRPbwEN0=
--pragma protect end_digest_block
--pragma protect end_protected
