��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F��������n�BJ�F���U�FW9d����T�+�wt3��^��r�q;\��af�י,��9NL���ٴ�[�Z��^��Jy���0�T����l|�x�5#B�o* ��J/�CO������|�)6b,P;����t��ew�u��5�v�u�E�8����R�oIk�����Wb�A1���5��r�5Hڜ �r�n+��MS5��n��þ�|R1��������E�%��0E���;%�6�׸ۈ�6��:�!�#��L�jT�a�S�N�LS�[�&Ϫ���]/��nm� 8K� 7�H�be��
@��1>��?���X�U��&��P4
��J��tz�6�^�O�A��S�������EjS�V�6�$�g)�H!�uA�����.����c:k���:J�G�y�*aio������6M�pʫ��QZkw5~��ΰ <�z���i����Y�T�w-�q$��k�d�V�5i��[�r6t�`?�.�^�v�
��l�;�y/��y6�]*T�۔"N��d�V۬����/S[�B�U��7 a��p~q������~�5�LPؐ�V�T��?*�ؓ�C�r�����	�].o������߽o8+\i+�`K��+darwEi�JI��4?�}͍�<<�,�j��'��u��K�C���=a�X̉��37�Z?�(ȣ�$��Yl\e���=~�Xa��s	 -~����w�N���,v-�xa��$a2��hA$]��g���[\�7�x���{�MO|���1Wc���C��e,m�"��$�O��
	��M_O�~���jCL�"����V��P�h�Jm�_E��HaT0CS��&�L1<LJ�ګg 9Tp���N�Hm�}r�NBa<��9����-L��s�/�ap6@^߇T��!�3��`�[�� [ݭ��O�>F��� ���&�	��A�A��.V�Sk^�%�M������P ���v׮���w���>��!S��'ho)���9�D�oit��Or�/;W֋{�_��}�
l�pl�ƃ(�Z>�(+���Kd�W'�s�@~NT�>��x�T�QhaKtO8�F��e�q=Mn��Ɋ��0��*g e���<StQ�w��ʇ��p�q��˨/����pV� �s;l-T�{I�G��`��2M���WW`А�9(b�Pt44{]A��蝨�W01J ��	d�����,K��/�����Y��z�sI�;%���#��ftǼ�����X2f]���� q`+�b�]��Vt�1�!�+ %��O#9�M��O���P���п'{MQx�͐�q]>��4*����\\�O�O������;(e�����P�H��c+�|a.�0�"[����F!��^wLo5����rI��&
���}Z��
:�m�{}�'Qn�J	'1��.IX&�z�N+!��Pd����Q
�H��M��T���q%���S��]�\R��N�|Ǟ�Җ�]�$7�I��6��@����X+�EYٔ.�O?��sX����g*$V� |�|�H�@�h#y	�p�Ǹ4<ٍ�`(�+����:F��j���#M�9O�2��A�ȍ�v��Tw=e�ڼ���2��~A��Y�UUV`�Nc�G��y�6�K�*U����� �'��$�����LǴ���uW���~S�E�7��ȾͫR�h��������\�y�SH�0_AW0�[MP�!���ȫRp����*�|/����Yr�&��ϙa��е����ق��ɞs(�X_��ɪ�p����K��8�|�ν�F���t����b��O]$:T�\j��"i���l-L���-��]O���>x��H�+�!�L�mŒNj�NDep�M`=ER.�4rh��͉E�؟�@q`�;j16ׅ5�������?�Y��,��Q8�-�B:7�����4Fp�ӥ ]R����0Fks�`�ql<PI)C�6ee��e�Z�[��+���`ߋ�k�$Jh�]�����.<��ef�y�9h�p/�/� z��w5�<7Nٸ�<e�R$��s�楤�d��>0�Ϊ˓�e���ZR��N*�� ��[ȱb�<tp�A���ő9v����^��&�����f�6��A��I����1i(��0R�}��^�	��g�XƗ� ��?�jNg��.���J�7��g������/X�ĺ����dg��9p."�8励�[���~R�a)��[�ȯN���v��K�n��ba�z�V%��%6���E8�g[:��:�1��85��ێ�oJ�b{�;ugTe�҂��K�d5H����R\�8�A���0�����a6w#�q׻��	슌!�p6��3b��E[e!
����=���!h��>���봁=�������$�i�=/����n夲����H�F�򧷛�cs{Ú�/�$zfJ�}O}�:7,dʬˏ�d%�y0^n������u� �[P_,![:ԶJס[���ڇ�%n���S�)S�X���է3���9'a�G��g�w��z��?��}��ȘL!ޱ�6O�;�^L�[�I�EP����� �"%h;�M3�ׅ��/�������	�z�MTa㹛� DJJP��FT����73T<��z�q J�MG��m���v���az�#�>����{��H����[h`@�-E�D���d�,6�/�GMQ��R���|P�����o�<��Q(dg��lXI��WA��Q�x ���t1���������^�G~���꼻9!�ؤ�/*��j�z9�^�6D�rg4�#�Z�U�ĚzÂ��馛�%Mm/�0L���/ϩ��棬�QF|>���{�;$�Gñ���!��������}p�ı���gm�1P��`ݵ̯B��"��X!�(ҽ�Q4���R��֥x,�=X��m��zv/�3Y�,7�xT��Pe��֒d̗����(�Զ �*�ye�/�l7B�<�
���Ç�XE��e�a�牢���ΛӾp����j�����¤$c��Y,V�76�jЬ�$dX���f�Kx��b��G��S�O����䁀�RV��2 ��"Ԗ�lՅ�W�!v�4*�%�#*�1 |z�G�hߜ��Y�|�����U����ۻv;����W�m[ʬ4�@�ι�7�?{��HI6'm�s������o�T!i����@j�J��=�������F[�� S6�~��+`{l~�\�k6� �B���[23&gyl����'P`B�s=��lI3��f�U}fV@��l|\�3*32�	�ƺ�\o"��:Y1�Џ��Zv�k	ÅlM"y���d��g��փx{��J���9��	�D�,�Ίp����C���� h�J%�	+�m�B� o���5i}C�'~����Յ|T�� X�K��-W�fL���<����}��=eX6�gaFkc��o})���y~�����n{���te���~�th��X��+��o��a��:��mL^��ɏ��!�3�l7���e�ݞ� GX۳��j�ď��7�q�^]�<�/q�� � x�[B+���]�)ȍf��A V���]G0����h˵��_<1����T �z�Z�V��-0�[�h���v_��%z��kފB��3�l!��-�^k@p�/-@�(��_�����5+�:ʨ��[�\��� L�R��%R�ܝ5��>D'
#�n�T3H)H�բi_������%�D253���E"���\C�8t��b�����Dq��-�(�y��&�8�-��w4��1��� �s��9"1�@��d������Ll��ƣ}��ɲihǯ�q>5����z��Qu����em;���`�����Q��F���l�^wFA�e,o���L�YD@��0_6�޸zC���<�����m�peh�Dv�������V�Z�	J��/��*@K�9���2P�*)������K�Aj=�J�8�U��Ldy�Ә�?���O蚝O~�t�l��c��S������b�?��Ͱ(�s.i���u�N�M�ϻ4��l�D����\Bm�r/��>W����WO�R���d n�w$�1h�O��� W? HB/#3_����jŽ	�K�8<�+�cl�2҂댊p;���`�̛���+�7�q� 	�������9�[��ݒu2�i����0,c9i����gf }������k��OxX~ϓt�����'���9o��8Zc���7���ݮ�V!��K���:$�N�)\��Ϲ�.ש��v�xK��'}jJs��"��V����a~-`��Z
�gQ�Ԁ����r�IbK����z6�C��+{��]\��S}Rq�}�=���܉Z�wGR��ƹ�¹(C��2�ZMn+���1?��s�l3T�v �wUQ�p5R�G#Wr�Hp����{=��	���������
�%���OJ]$(�:�oװhGڂ�����uo'�qd?���}J���ր�(#�$gdw��n�Eٮ�d�C���L C���B�؆���G�vW�En&9*��zYB�L����n��|��pg�g	v�о斞Q&�Tu;�'V���U�l�5+8}5G�E���0X�s@4�1�f�ۄ����ۧ*H�-*E�ޥ��6!|-~	�gA.��I�m۩YPe-�RU��������#d��Q�l��x雽X�b���.������I�֩�����k�U�[��'����d3���L�{�?�YٸVV�L��+�]�J��E�&w:��*���g��Ʃ��g&��ƹz��q03`n��v�����;�bx�\����ڙ����3d�37ܨ�D�|u^���k�(���*|!��b!�o�pYq��?���kzڊ�!h��ҒB������4�^a��S�le䀢����򌠴���(�����"���'��J�Z�i�^%���dd��v���pS��-���A�[q�qk�1�?&\���HF���N�i��,|}Pi�,M ��2e�żZL�R�e�Jok��#ϕ3"�r�E=7W�:̂�-QeX�4���p�fR@}�`ѩ�`�1���[O��^+�5OW@A�6K뮛?ثT��֔��8G��K��C��<@�A��U��{������f��r#���4Ȩ�����W_�n��g�J�5%�3�X0���|���J?q,4���[x���G<��t��\w��/���g�ϣ>�i�iԝ?���Ӥ%p��c��(k%t�]�b/�&�ॽ�]�Kvh��z�b)v=գ��C�ȅ;n�����b�Ov���V߸3���ز��xG_�L�#5Cc�'���f��������+�#x.�ͩc�l�szC��~."��VdI�o�Q�a�W;ې�Ji�N�1��e������:�A��v%���H_��wﰶD�Y�^�� 3��k���6� @]d&$�v	����$�� �"�&�(l�-�r�X�$���8ANi�[�>te]P�U�		y҇�A�����s(6��KB��g��}���ˌjSԢ�C�H᲼c�V��}�idTK;�Nz�Uø;���\�+������,,<(����=,E�Iu���8	i~	��NX�5�PP��hLѵv5�[8��<���X�]�����UFh���{m��h��f�Af���v�,s��1�0Nu�u¾����x5L�K>d�L�lW�X�_�)�Ŝ��}٫	՗h�����U�KE�O��@}�?6�YW�Tx�㯸�䝢��G����N������&�S��8N�	C|
M��A�p�����ԫ]���v4�r.6�����)>�*f~�Hj� 2��&�/#sE1�Z���o4��Ǯ0z��]�vq�i!Y�ޮuߣY#�=6�9;�>��ʷ��o�5�R�mF]�� �������>W`ސe4}��o�+��7'_Q��dy�n�'��P�\f�n����4L+�� ڊ�e�r�N��H�NI�Qw�鶈�ʇ��q�ӛ�eB�i�2jie��u�N8�yI[�v��B]��}�N^�m�q4�ޯZق&��E���B���7�Ү	�����=���0��M�%j��>�9}����v�������K�UFc�D~��<� �xM�7�.�4��:+�]G��)#�D*L�Sy��Z��j�,kQ����4��DZ+�̄>�BH:��<_�]Tt �͚He5��&�"���6f���ia������ǿS��\��]�x:OӶ!y�n����6u7�� V١�.��#�tc�C5ZÙ8ᔫ�2����) �[�I��X�<J�Z���|P�S��C��N]�P2�3y8��;M��4��ڴ �\ߏ{Nnet�g�_���z.4zZ�!veg���7�'P p%i�v����Ʀ1� ���`��b=�V̴s-�Yl�{�U�c�<�,]�P~U�~���]��;ٌ�f�[]u� ��5��.'����ڒ�z�rk�J�r��a���Zd� 0ֹC@:��=��:�A=�����tHBG���Y�4���1J����)�zdK�Mr��R���}��v:�4c���J�;�$�3	C�1W�����o?{^+�����	)pM:ߴp����IXNN �d�Z͐��ٽ,^�Z=�N=ҙ��R]����k�+YsA��-�8S�w�و�o�����lT�4�^;�uKe롗��ۆ��a}L�Ʀ�:O�y���n�H���.�ڼ^�;�Q�M-��n��a�v�	I�� ��h����pm�ιc�`}&׫(�U'�tQ���D�w���������K�`cq����W �9���/'^��/��^��SDA�H�Z����Z�����'mBMi�:���5���S����P�f����?��Mv����)�e6��*Ύm&���u�y[�K5�Hޏ���v���sݫ��rDO�Kǆ���$�Cg :r���{'���)q���AMH��N�U��F��Y$�`�\�+�܌��z�~yڬ�w.q.!UVY'_l�41�O�%#��F��濰ꨩG�p��_�t�g�`T9#0������+Pi�̾���tG��AcX���p�h��g�+"��Z�S%��y�XD�j�8�a&�3��5���w���r�3�PW�Y+U��W���^#F�,�'N��*6JmI��A�)�3���7�V�L��f+'����h9�#�y�6���Au��������W�Ar�N����8�_�w7�⎁J[,���� vN]�㓽�G@��@�?�v���l�Y_rtg�_bS�#؞���)���l�����	<i�3��Y��fz�~;of�x~3��N��mU�� ��C��ߣגȘG�����������GS�r<����Sv�\Ԡ�k�t�r�����K�A��;�9TFw?-��5�� 9�[# ������HZJo*0hZ����.�Vh��H��2r��6��y�0�2/���������g�����l�(��%�*C�x� tF�oD����l�[t G���2۰u��>9N�/�s��Å�_`�W�W��~���H��ZV���+�\).L]T<��.d���E l����8$D!���Ϡ�f3a�&�Է6A(#��1��\�女������;�Jsz�����)	.Ƭ�J�Yx����NӁ�x:�&9�7���Q�R�^�#p�����!�"��\`��s>Pw7K%*��-�M9�)�7�ؖG]ث(�+�Jdw�
r�w�J����8��7�q������֏ȏ�I@����r�b%��*ϸԦ�V�u�zp�����eH�b�>8�]���($$�ank��~ ��1Zߚ��	X5kyo���p��buz�����{��ƴ���>���k��� (��֖�(<Q&�4p6Y��\-�#����i�[��K�s3�:d�$�Q��G��7�-��_0���1�}ga >�5a7%��+��>yBs��ੱ���\��VwU#�>Z�Zu��f�5o(v$��>E"]vR)u�C��@/KD��o���#��ū6"��5 |����×��Ն�z�La��}K��lP8�[���n�Z�27��l+�R�N_�ғ=0�R���
���qc&ֿ�[b6Os�TLk�j�X}IN���� M�c�f{,^��u����LKUz=놑XT(�Q]�S�z���c�1�G�"�ؿ� [
5�� H�뵄�QJ{�:�W���	�F���A,ϥ�q<ܴ5_D^�Yd���v>:z��\�Cɴ_��f�����pT�����  �+�j��=4��Y7����"O�Oz�欩~S���͹$�d�J�(^� �o�4�p����]���M-�,LHDhy�	
��
�_}�V������}o�m���DO���$x���_��G(ѻ�/U�O^Ñ�v�Q;nȱ��w�
1��@���;\F3�)a�8�z%�
Xzȁ��Jm� �Cz��7Q����3oHCY��#��v|�q�qgEG��vNԫp�8}W���B�P�˒J��2��F��Kh�m���JifE0����߄�,*C �����Z��Җ�[4s[��u�k�Z'_�1�?��
L�������Z��ܓ�}m�������x�I�wu��n��Z��;�7��Bu�m�^-���D%k�!R��I	QF=@�Tg���Q���|9���}����㬙ү�>)U�
v�)i�Ee�P%�h�8���N=�s
�k�v^�\U�N�������m����`?��9{��+��~\3�g��c�D���0[��w���� u���cLϵq-��#�3�3���W��R[O�sKcX���^�(BZ����~J���]�NZ��3+�3�����PB��(zU�� �t�ոE�L~8�5�e$a���n��ӑ$�.����̲$�j��C,1���Lj#B�=k gxބ#��h�d�ՖzzMA	�S�6�V��Ś�`i�ȵ��)F�>ܵw)�W���,!����AP�Q?gK��E��	v0�D�hq)�Cpȹ
�晼(ߦ`�B��]�6����2���Y�t������ 7!��V��q��H��[	�d���[���<Yb�~�n{�p��TsT�]��n5���B�LS�On�jq	�,���2�.\�\��}N��^S��j�t����ayN'y�?���Dr�P�Bcco�a��<�-�y��?�٬���$6Q����!ю,d����tw���oB�R�R�˖��i�Fͱ��P�u�:��_ViЍ��c�і���at��a��)�jw����ky���V�W�}f���i�i1�~I����(��|�X9�lه%4(_6�Q�ۣ�ARp#AX����/�0FG�j��W��]��A�k��*�9��'{�J��NgPc�{��
kd L�bZH�Q���n8�.�n� ҈�?��)�KAZR��j��yƥ��P�zu,�I�l��zT���m��Բ7NwbۛA�'�ß{�([�L��j�Gt� 8� +�'��+��%/Fpni�o� ���ns��������g9��WX�'S�uՀ�}��/y��,�A?S��V�K��V�!-f4?��g3ܸ��oߗ#H�"$f؃�G�}��X�۳��Uw��hl��1�|3(�J <�l�FF������	9җ�٨���g�Y��ۦ�.nNsMY���n�%�� �(�� ^2m��'�v	�$S,/��~͗U=D܀VI��TZ`|q��j�	������s�	�U8�FN]V?�K�r<�$�1I삥��>�i��ku;!%*��~r��FY��
K�ݧ�0�v2C�҃�ޙ1(�J�B�z+9u�!����33�,�s�V.�p�X�S����m ��ј`Z��b\���@���zVr�O�+d
��yF4���A$��3���<Y����D���U���l2��,4	s�u�f1z�ܹPʡ/��!ml�-�E�B.�b�́���r^&rE����C�G`��A�kvx䖛Y�E���G:�h�"��H̧§T��;�u��F�0(NH�_�3׾"�'�L��w�gd@���Q>x%�j�B^LC�U�j�1aIz��ohmm:gm
���+t��-xܽ�R��2�R��P
����P�� �IN�x�i�DpȤm��&@�]C
�O�)�ۯ򿽍�9"����9I�<����{��E�x�w�a��[���/�G�̿~�\�� �c�q����׭����BZg�l���uGy~����=���;=��ϒӥ�A����N?����n?��hJ�]�՚�X�˅�5��*�4g�)�?��Rc�؂px��N��+k]����Ձ⃘ ��_�y<�R������5�[����L�ֽx���`�m��Jqj1�V�]�!3���P�w�bS
�*��`�pKq��[��ڏ%f�������;�:������w㑓�Z�	ee��)�FN�6>�9��� ��D(7��f+b�Pe�����[5��wp���bƠp��T��gM)�T���omNҜW�ϴ2Z ���z�)%L�$�<���Ȩݺ�#^-=�R�n��X�Mn�����'�֚zd&MHg+*-,ô��"u���&=�q�9�6�����61LKfxg���e�{�Ù�<�;Q�tD r�!W�䳽|�����2ky�����գ%��d��9�e�T����dh�B|�/�nw�&�
�-1�q��^����׊E�=��8٨�ȷе���r���zB�C�O�<�� �f�wK������L3$?"Q��Ԑ3`���Eݽ\@�W�Z�d歈�_N��_1�6޺ I#��Z��I�Y�����vE���7K��a�h��3�n�|��{���1��#ڸ��[��izV��E�R�b!W
�EԇzA]���k�޾��v�O�(Ģϊ�/p��ʹp:׵5L"�X��G	�G�?W�ov`=k.0LX?�j�z���l��p�,�t��+���ˇ�S|���8�7�*w+v�|��idmnf�J�K�w�r>F�-����]t$���p��e]t( @������.�ʢ�y�	����Z���E��SJ1#��ǳcQ�,���ҰhySMx��Z��"�hl��]� t�׆,ؤ���rE���c�{�Ήr��N��.�Yjt��2�`�����&Oy�E��P������:ұt}X��|� ��4O�S�T.F�+{?	�<g��ײ�mTҼ#�D�9�CEM,�7���w�qL1�<�X�:���ۤ��#q��7FIWy$�ra'l�A�k�/g��5��R�{%Q�v���|�~#'yY�zKK�E1>��YOml�Pb핸~k���F�+6����6c�qT�(T|�i�����G	��R�Z&6�W�B�Os��&��m��"X�
���34$�o�:��n�0�G�=f���o�O�9��j�D�al�^t��N�c�{C=2��V�%���$��o��9��4��n�\�+֖�d�D�a�<�KU�)��2$#*!��@w�p�ǃ	��>����x���~�#҂��V	C���y�*�^��E�Bf�]���#���"�/��o���=4�v���y4y�$A��)����P�[A���r5�aу�i'oԣ�n�E&�9i�gdHk���A�"^ϰ��W5����lƿ���t���)1�ӂX������l�k���y]�ѡچ�����oV� �b�'3�e�I��w�q5^�{�g'Oz~v搣�w�D/����J��p>�։�J�����Qo������܁u-R�D�c!�a%�uA��F��#�W⣍�Y��1�&z����* �m��4�q�b�N_ч|%{�--vdh�U��*N���Dvu�W貆춵D��0�z�����\��|Z�$��4w�ԥ�O��Gj̯�s�����-�5�����<�o�*��E��t���<B�q�i>��`%"1Z����)socK8r���Tk5M�G^��u�8�=��\�>�����swUo$^ܞ�p�o"�;(�^�E��sߌw��N�}�g���"�^넆@�����p���I�H*IV��[���l]TZ�4���~��i<�F�G��C�O�q��4@nC�X�(̽��P|����^�Xa��r*��yOG-��VW���}|���[\��	;��������-Zj�o7��'P4cJ<��H����@��v����,������H���1�$�IP �mƮ�x�o�mf;,�gP���]�{!f����I���kA�������C�l����6���E֗+e�K��§���������������lbU�
x:��k��Xށy� �oCŹ���FjNF���vAl�:~���y�Mˆ�(�m� !S]=�rڤhjp}9�<C��Q�~/,�
�I}��p²��#G _��7E5t�]3�B�"����LĊg��i͟
�K�5e�(�0W�y +����|�_��y;73���vvm��#��$��3(��6z�/�;��s�`d3gأ��h�C�))G)Z.���O©�w"P@�<���ݒ��� �s��kT�Dg�u=O &�$��|<1��e�_ո͵�f��Ix�+��ڠ&��z��R��9���G�����hx�����aU�i�q&Nߺ�x�.\���\>t��ښuiz���(�ͧp!�_���br��¿��"���ϱ!>���+6��n��FL�.z�$�m���;�I|�%el<��I�_�d�
$�z�2���z3L�TT�$.�u���>Q��8����C=���!x�X&��Q�j�z���0Zc��hy\ǏE2�B9�k��ko��윐��CpFI�CjӼ���[T�J¨�J%Av`b>��(��y%�m���>0�Ⱦ�@D5+��Q�����jKu4�L(g��z}��K����PQ�r��C#�U��� X�����;��R��^��� �z}T�ID1k�@V������VO��1͵�zwE��F�4��+\����	^lٕ�)�=rۄZͪVVN;yN�a��>�-!���%O
���U�N���#^v�Eb+��v�+�)ͱ�N?eV��gKu ��З�r*��E�O���L3��`	I}��LR�A��h��Y�ֹ,2��R�bU�����k����[\S�WY�( ���Aβ��Uc�?S˄���74.7ޓ�${��'�����2�3��p�~�S��1����]��I��_J�s�l�fM�����X�D���h�ȗ��9��M�k?��*��^5	69�Nl6��Ã,M�_	����Xa;�,�(����!ݬ���
M#Ā*�v�Up�b���z��Lݔ?I\��q���1�;<�b��s�Z�Fx��3vj���j�6�r8.F�r�:�⦨R���~��S�Bc�fq�X�{-D�~��"�|�n�}�m3l��<��2��`sT_���P���D ���a���f$�7ZFB���ʫ�eFαʡ�vc.��9~�FD�;^�
@��
Dj��#xm����ҵ���U��#�P��U�?0Z��\*-���4�dΌ�F��Rv�xV�3���iG�\��ou{z
!n i�f��m����X��(�{9
�p��f�(�G���^�sp��n{��7�@[��s[2J`��a��f�H�z���8�D��r5�h�.4`��k��#�@�;��t�k�ґ��k��KR�������W�v)����!���sXW��#�CC���Rdv�~z@��`K;��l܏׆=�E�G��O�f0���V�0�o��I�#0��{���[��
��A����&}�����K*�*�`{�F�6��羑y����g*Jq�tصh���-�m�Õ>e�4}<�$gכ����42hk�u��B�����[��a8Ki�
ВK�L9_�ߜ��ݪ}��6���̡>��1�/a�1\�2]�4}�	0|c-(^�7�ͩ0��!^u�bs�ыk�F&���v�Y�8�����:�F4@�����h�'K<�%]E�k��~����2pdFZ��l�q>Lы���=���Y��n|����0��rf�&��ѕۀ*��;hFuJ3]�R�	KD$��+�o�"�Yƺ�=�P�����pU+jH1(���Z5���S
2��gQ�И�H~JAO03r�ڋA���V3�*��~��G��|?�<8'k*�>Qa{o��;�ci<�%k!�a\���J�qw��3ێ�گ��h]�Ϻ��I+��G��������rHk���SY�@ӍO,[]�O�#�)Җ���e1WU��(J4��r��S��X��"�����ԫ�V��d,1�+д���à�}�q�u�6[m.���w^ճ,A�V�Tώg/����0���S_iFR�&�j�,I����Ӝ��͚%�:A:ar�b�Ft[�c��W��6}nz; ~Q= 8q�L��j��qЗ����R�QV^Z��_�}���^$�p+�%��'���C,Pca�9�0ڂ�����e!PQw���ɕh�w{��]D	�r	h��r�[������H���R[�=4��5�OF��r�4wnƦ��b~�'���?�:�\�ӛ�AujɹU�w_�b�^4��'HngC��C��������@"B�R6{SNn��_�G���G��(z=���P|����lʉ]n�juށ<z�DG�Խ�fw�~@�}D�^|&�p/8�0�l���
S�e��.(�(8N�����b�`��~���7	���rq��A������������,��L�2S��:y�-��Zs�����+���A���bu�4ұ1y��Bq�7�)���K��d9teS"��Y�Ұ�F�B��.�#"N�Z��By�X��g|�HRet	"ʟ�N�/��ڵ�6�������E��|�4d�x�N)�)��-��1_0���D3�<;�'h�C�4X%!�i��i]la��Ӌ%\��7�#X�R��15��ܱ�YnX������Uh����_���dK���:@�����`M�s���ѲmV��L4�e���%���r/N$xR_��#�2�m���<	���+��o�M�`e���ݥ�W����V���q��^��J\�M�`l;F�g���t�0�g��D������5󾾯�YˣU�9���̻۾V8���h�/ې�^��l0:�I�?��N�/�ڮ�8�؇�-��C��6C��S�Oj(�uՉn.��ȗ!����hk��n��[�f	ӘD����o4طR�Oc�{ ��H=�~7�޷���.�ft+�ŞM��"%���R��pQ}2����-���ݜo�qԤW�hk�9��Vْ�SCB���]���f�v��H���C��e�a�Ċ5[��x��v������
R�� �s�����7����&�er�Dh���^��M!�8``K�^TMa黸x�*ع���,qB]�W?F�V�V҃@�������g��8���Vw���D���;X�	*V$���y9멞EjП����������Q]?o����:˜��5Z��R_���,bUѢ} ��ٰ-[�O�����>|��	�]��!q�ce��f��R�%����nH�
C�=¿n:4Fp�))���cE'=��;��C]"t���?h�C�}���,ԙn��)q�GFj�ژ�ꔲc6�L�Ec3���w.�4� �	W=���~���\{_�y)5�FQ�}���OK��%_0�.:w(��vE�A�2�`%I-��d��[�d�y�~'��H��Ҙ9�����U� ����V�ٹ�Tz��B}H�ĮRu>3a}���?k�I����a����TR/�Q��2���ܚ��L�m����E���y�/5����Dw?�5�IU����E)7��,g���L��IE����ּæ��d�95�q�dxps5�&��Ȁ2��ߎ≆IN��)o�A��舷."޵�V".������β�����yjpo�%J���!��(V�o$��hlN=a�0��"Vb�a�}d�$N0ȇ�lc�z�,��ׂBih��+��5o!���T�.�w�Y����Ν��\Wy������b>�%3x��d��\r����o�����k|F����9��9��ә�J�n@�mG9���̾'��O/�)Qd��<�VGg.��y!�*����&\F�(�ޙ����/��?D���E�|J=�c�;�)����a�}����/�J{�d]b�����X�!;���ʅ���%Z��>L�K�g�t:��_�n�}7�N䦴��W���ZX�q��_P���g[�-5�ȭ.��N���o
S�I���uA0C�/(`�d�(��=����U��E���'M�/rT(��o@/5�1�`�A�t��$�<�/ �۶�#��Z�1·�m�������:$���Ȗ�*�AS؃��g^z=v�������g����`�]Br�cO�������v8�Xx��@�R]�2;uw��W4�د�Mjҩ�s嵖�s_&��,�͊�mHW�x;t�L1�9%�'���w����J�ګ��|��v��YD�5�Fcvj�hQ�B}t�4��y�D,+P�`~�rM�"��������+�C�L�����׺X]F`��tV:y��*�lg�a��A�h��v� ��5�I���^2g��|�{�ז���F��^����4Ԫ�>-i�����L�4`s��wv�iH'���@�t�B}���1�۱�.�[]{�M��pG����m�VҤ� ���nd�A��<��U$���a��"K>o5i�H�9}����RO����~t�{s�P�u�F9�fTS1-�v�GC��:w�|��c<�2kN���a���d�cHE��v7����Y\"g״�3Qh�e]���tvإ��.�b=cM�Xt]{��*����)Q��B��N�fK�������ݞ��E8B<�Gȧ!_-X�E�82۸��G�5lU��T%�����X?J�ѡ5��2 Qپ����P�'t���$��u\��.x� B����K�7�Ńa��0�AP6�q@c�o�����Tf��fkM��t�����N.��$�4<֎�x ���"��V��\e̥���S~B��%���vKZ��i �����ſ��Dط���'`�h]�������������9T�S���r��9D(�4ы��.#��3����20���������#�`%����R�����L�����qI��l�:ʏ���+K@P��oqHY׍D�����Rj"�B]^����P(���l?�If�[S|�4�j���UQ���W��ɔE���}73Ҿ�����
�����T9��#�gK�X3�(q���̎�2n���~]i-M���󰝛��$�\�g���svjy���cz:#L���X�ף_"V~��9�bf��~T��{%�0�;(^��T /)�ʈ�?3�m�z��1ç�2��ݺ� 3V��ر���y��B�1��oR��T�gGz���Qr1G�_|IR4{��$]A�2BgaX��[�w)B��&����[DV"��)^�cf����8,�fGQff�Z�~���2����#&��6|�(2�Q�Ta��վ�QP��Ѵ��<����s�ɖxqd���*0G8����7ߺ>eOv�-aJ"���U̲��6i;d���L�0�a۴k*�=F+�BT�2X�H����j_��^�'�N��؀}�F08�чQ'���@����U��j�w��׃��.����E�a��3"
�+��ݹ<��b�35.1cM��z��&X��Pdo�U��]���z��0�C�ZQo���kP�^���=�~��c�+v�s�9F����i@��7�"��g��bt�v��R-'lOL?�>��`��R���u�Et%���g��X���}.�@�R��R�+���/�.�@�<����ټ赻N���/�g&�t�_��B�c�<��чI�ɜ�r@?��kc:�\yVɮ�/H��-�I�?1��|(2&x�p�TdE ��ci�@���Y؊(Qoȟ��!2'HM�X�P�Ξ�AM�Ȑ�I�\!V?�\��� �*GN&�p�㨅�o����f˨�AX|�!��]Z���(��LJ�C��j��?+V�S?D8�AT���7Ӎ"���g1
Q�:��J�m�������7��p�c0��Q�|�;zLD`��%��N�z��:��1]]�6�� v�>@��w���h��~������R�7�y��L�XY>��-=]�MVK.�� �Ҍ:yDu�R:1r*���'�^kg�5���J��S[�������H:����U�鸌#�����Q'3k�{-_km�����u%~�RQ�D�|�>b dhEt��������'a�6(9֬�鼣s�[���-�cѷt�jD][ݿa�C�C�C�W�d�f�9�	���Sԩ��8������n�H�А���驞U8z6&�M�Π��lf���	���O��b^�=�Q���Y$y�Tx?�l�'iҧ4�)���(HD�es��kZ�l����C�j[/�l�h�I��Zh*���&[xp�5�-��$�?�H����7�C7���Ȼ��ޛ�1�@����
�Ϧ����=Y�JE_�l�+Ϭ#U4R��8\�s��ψ)c����&��*��a�[�,WL��y�a�U� ��5Ŕ��+�k�������b��VV�A�j���l�sWF{�p�[������5~A�l� h��TLۊ���|��olZ�g��f���J{ ��V8��#���`Y�
��&�������Sa�%T���Q��V�#{8x�j`�͜X�.o�sɤn��g�g�>�jH`�@��޹�D���%1:N��n�X	�P_k>r��L�C*��NLF�Ϭ���R�`�b��A�-Q�o	wcy�нN������[x{���=�/����B�4z)F��|pW����۰/�`M�
����%��K�e������cr5!���A�EsT�7p��B�)��/�*rK��mj�L��Ԅ��A���ǌbSMf�fU��y	s�D1�����c�.���	M�s�o�ގ�d���*�@�9����P���E��^~���$�}��sw+��t��?ԗ2��Z����P]5����P�}'}{�j�����\�R�޲�@<���b�.^N*iD�&�F��	�����v������a�`m$�!�@sW!m�CY�j���绖��:Ӊ��b�u���D!B�"����G+m1[e^o�WD�p{��eq��ȳ��[O�|�3����1��kR���ת��i6�������sʛ����u�w�������B9!x�W|s��
�~��y*+�J�㒣չ:t��[|�C�.$������{H�W���gͮ�E��ѧEA"�M=#������Q��ҙU�S��"\������N�Dg�Fa�jU�����ӓ@Ũ����7<����P��>���䦛4�ªO��
�)AS���vB%��2�-]�!(� �M�ٯXkc�:vJ��z�veJ����p�+��R4�	*)���dJ��'~;N<����P��~"P@j����	|����ۗ�[p���eąݲ����ؕ����9M���/%�"M!2p����m@<�+������0�],�.v@W�9;�K�+G�䈧����&o,����n@��]�&Y�v���ͫ�DW��x�V�_��J5/B5MK�Kqm+l�t�!��LBB�H���6i�b͒M=+b�W�%=���0Ft��o��A+a��g^t�f�5�q�`��pT��k�nɖŒm�_5����(��v1��9ֺ��0��
�����"�q`U�H�+w�FsF��F-��@6H�������_�P\�.�h�&��������%g�|tVK��T�+�u4_��L2�ECT�wgJ����;��Y]�u��{I
�RD���,���l�8w�3�*ښi��?	�7N"��$�=���n9Ed"�h�K��A=�U"C�b�����Nn/�����,���P����4.�d��ʛrd�� [�t����#A!���_�WM���N��e:U���;9"j5o�r�Q��|��ʱ��W�H�MZ<��[�d� W�YadZ]�Y���'�匣���%�Z�)ieH�Mȭ�^#�a�4n��آ��i6��M���@K��V�!ɧ�~f5{�5У&hKg��=?K���:g����`�<��U2*3�0eMC��[Y�f��L�6���?6(����)�[�LM����P[j%bqc1郭NY�ނ[27Efؘ��zX�o��FvP�.���c��.5r��	k�]��x|8Λ�� iFw8�
���P�w:�>3���6�\u�����Q��ळAhYӋa����(��S\!����|�����t߯P���%���$}���"�&�@���9e]�F��i��%5�d�6�b��1C���]��8�����^9 U�zEkd�כ�(���\#���1-y�,�����k�ɣ����5,{�d���WD�ʟh~�]
�A���>ٴ߰����8I�IE!%i��� �;q��a5�_#������L�&Q��h������W��2���D�B�l:�*Z��)��`5��xk�M����#���a@��&��n$����aoy2����S�%����T'��p��7S��_�pr0�'��=�����~<=KމD�������|�u�V`G
�e���A�\����,Jso�de�w2��4:˹6��Q_0 r��qL�;'�^#��{6�.�Zq��8GIDRX����,��ە�/d<�TG.��`m�=`S�C��c��tq��)z�G\@#A'�z������Ugn��ѥ�,�E��}��.ƾS �%[�궀:�U��O�Qo�,�s����Y�O�A�@��7��8�� |{��O��)���%�_[�^�j���6d����/�oj���9~���3����L�GE��������eN6�<����k<Z�}�X��j�����m�v��$�{=U�iCpq�4m��6<#}G�1_#�aW=��$��g��o�z��M式8��t��Z^6>�j�c�E��r:���ّ(Z.Bù�Ih\�s��GūL��e�:_($�,=������`~�(d8F�OMow���m�����rW�fB+1ۣ��Qߵ5=��W&H(�i =urk^�@9&m�\����Y�J?O���xKl�k_ gW�ʹa�JԷʗ�R/���8o��toe���l>/��E���(�db��c%&������r��^L����*ůmr� ���s[��xDHf[Fj�d9(s0���x�9��ߒ��$5/o[0��ij��1���|�*���c�¢����n�ZrK�Ҝ���Cr'���7k�q(Ğ�$ʨ�R���\�q%:_7I��t�T��n�����?�4�Wy����!!�gb����b�<�-�r�*�6����]��(�-7��F+~���8��+��U�� ��� ��`���J���$�Eu �22N�Ӱ���`S2�.�i���U�D�.۲���+��Ũgun�\"	��j�C��K�����2��}�|�1��{���+��3�DW	3+�+��c��_t�����������峸X����F���J. �r�K20����7ڽ:5�{V5a� �c�F�RVl��O�6����6��=^�Sp׼(���Eq��L8+��RI��PTD/�e��>S\ս���t�J?��`9�Ra:��4������f��p�o��/G qʟ� �p#71��!����>��znR<�\_�-(��Qw,9�3�zU7`����� ��pc�>��Q�p� Lf��R�����N��|��Q�s���h��!����ݎ br��m��+'��hp~�@a��zm�?Q�F5�Aɮ�_A��U��0���0�Js�S@j�E)�0�r*2��N+��49H&{.�vK;~�K�Γn]&k�X����fB&,B׫�m�������*մX_"x�Ow�"?ӏ�a�d]dF�I�B�g�O�0:�7������U-%�˼��E��t`�t��X!��,�9������2%����2�W�bj�Q��Ik{%�`E%����|���y�k���k?~C�+%��9j�*�d�<�MR��)_dX?_:��WV��L4�1�'�.�NY��ӅCm�+\̺�.�"��C��Ɓ��IpGN�����GN+VUH���X'0��)�^FD_iDMm�&��*'��4G��4�=Mw?n��azpA_\���!˺�j5�Ȅ�d�'DU�*���
L����U��~�rԐֽ�J|�>���T�[���ԟ���'��_�r���)�)�M��n��JE�KB���~��X8���cn��}oJY7�=�sC�}�T��x�1ŕ��?b3�k��l�m��H�5uP���ԳӍW��ո��߽f� O}.9S���a�F5�x.�v ��բ��3�.p����*�k��U	�=o����g����z$�RN9):������dgꪮ)���K�����=ޓ���m�{�|H��i�l��U��e��tհp�_�%�cֽY<@�N��l%�/T�U�������`��jX9,|�e��[��F{��~��(=��9�X���AS߶���y>.��$|�e�KDp�ti��c�_
�,,kJ!���G4�1��0Ar*�6�Q�#9z(]�Tߥܛầ��k���}A'm�#��{� �[��4%b��ώ���[��z)L?�p�7V���gk�X��1���"*�e,	�V�ਥ|�!^��kK|ެT�v�=wi�e��L�W��4jSE�g�Q�Z��X'��"����I�a.���C�^u