��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F����Z4��#����m�ǵp��}��a��1��qh8��ɞq�t�m$��?�Y�¤.��i̓X�☾�}ד�^
*4FFx��:�o�""�k@�n�H�����s����F #ʨ���~\��-X�����[��Mm-;>�B0U�s�Z|;�N��I)4�][8x;�Ȇ]�i�?�@%+�"q���#޼��oǎ��L���y˙����rcdFNf���������`M"햎p%��=�Y�����,�8#����7�����,�=ң�q��8h��H(�[ҭ��M��B�E9��Ê>F$�p��<y1�G^Zp	kk��������y2������%GP���a�;M��0���n�a_3� ��J�u!�9�������r�i���@�X�^Cj�q������j��))���ϐ��\S��k�4#R�`ʭ1����j�Y5.�<-��
AҌ����i������J� ON��*��.(9\�5����K�N�ŮeЕ)�;���s&Z���<v�l��h�cܬ��@�3{p{�
��������A���cT�2�I��k��y��Ա�m��`�ݬ��h��8�E\m
u���(��}�a
�j�'^>ٸ3�t{��ӯь3kc'ɡ/��c�@A���8,��n���<��=|\�S�����浽k�g��㉙C]\�Gk���+���*�@{fЫ�%�h�gBf!z���|�_8zX.���J�Y��
�Â�L�t�-b.1��u�� eS!��X�x����t��5`�mp��CgS� ޘ�o]$|b����e�\J(^�FF�U�f;��8���@�Q�aD;ض�5���@��AADEȀ~V��%��JEB�i���sY>0'�\�V��ӫ���\V��yY	�-��ԱTp�&6dϚ�hVNk0�# \�u����P_�K��`������y���,j�������q'���=��g����W��u�8������F�4�!�|u��. ��tXNɥ�"��:���Ca�(P!ae~DW̗MǷ/�+2%Ꞙ%��9L�$��p�v[�iR"�;��d��n�ϑ<>r�"�{�ik1 �#<-�$��h�B�T�)K�5z�)K���k�W�l;��5�%)gn �M��)�	=�����t�����E��>(�2?��nk��1���W����q��S	���rB�cP �*�nw�*
����h�xi.Q�F�I.�#�<�
�I���<������w�oYT�ȨYM�;?H��(��VN�تD��2�U����fu�e={M��O���?�o�!%K��_nQ2합�ߒ��h�+o?��=������(�"\sT�����6�.}62lR�,�f��bId��H%�:޲����q����')�J
"^y���`�V�l&/c7�Bd�o�2�?�v����Kn����2j��wx/Ŝ�S�+�	�F|�k�Es�K{�R~G�Z���4E!�Y�~����xЊ�������V�MU9zB�ţ��j&�+"Li����ʄÂ=�e�麣R��J�T��=��-�G�#Λ�г���JK�=o*ð$PYu��΂�^�n�M��j`B�An#�J�9�J�]�2]��
߼�M��DT��q�Tat�R�}�7W�	P�7.���>�w	�hsv<9�E�ǁ�A.�xg�"������$��(XiQȱ�65��d��C�ۖ_��a�࿒B���b��I�~�
��ʳh�f�%�y�H���s�ʋ�D̞F���K�d$�R��S��J�ר�z{��&�(�L�s?�AᏂ'"uf�w�S�O�Y���U>[�D�T��+�E�o����6}Q�݉��n�
`o���3�v�ڦgsb.'k_������fE~�|�r��gb�18�Ck���l�2s
)�?ԕ���c�%R��L�?�� psy�y�%���:�X���Y�a/W�!�-T`�%����8-W�d;&2Õ=��0I2�=�odh
�A�����mW��#Ιd��,s��ۈ��x��{��3|��T�m�3�?����1D�s��$y	z�Nо��\ Üa���C�)(�a6S?L���������$��nAYF�������$�<����!+�C�� b��:��ql=pg�6�"9�pe�,�1��H����*X�%���V�o�/���+
j,���zZ7��U{Z"u.S��Uz�`F����0�Ad�=�����  ���U����� b?�vx-bܼ�9+����{g:]�)��M�@=���9Y���z���L`y�R�3,�Rٹ0M_��ص����>�˗��g���zw�,�z��������0,l��iq�@�F���X��4���z*O�N,r�;�	��3�7	dΪb��.��X ps���p�Z�(�{��Җ��7/��/��&D�K#�|<�Z:����Yu=�Ǯ���] 	�mZ#F��v�v�2 �T!�^qD�o��?�c�
o�+���S��%��w��U�P���DME�*^A�������AM��O�Z�������)��;�
X�Y��[��i/��
f���:�iDR��.��Z���dC��X4a�>��?`|ܳ7r���ᬚGI�S���R�nрҭvW�ưF�L"�ߔ��jOXQ9���H�k��(MZ�wWPVlm{`�1q%��J�P�l�g����,y���Zr��Yhj`�]�x���E�g��j7ܾ�v�>�hϟ�5��R�"��Y��ڒ�!�{\7���-(d�������3��Ҏ'R�<�]�3M'��x�J�ʿd�H\��b)�j��g9�7�^#�y��N�c�z��#׬rbV���·�����J�,}.��V(�u����B�î| �#��'����6���{l
���]u�Q-��q͠����أ2_�動"@�Lq�=�"j�$�ֶU��vNeI�s%���5"����<3'/���AH^������E_�|��9"I��1�s�5֙-8?ю=���	z_�%����-�
�&��"�:�T��w/�)�̠�Q�����`�.�9$j':ו��g+S�\b�8ӹ�O�N���J��)S�����'�ռK�E~�П2���wa!e3{�³1I�S����[L�.~�WX��H���th)G�`�t2*`���1�� ���mM)u-��2`��ؙ��츚���i�����-k�F�=�N��8P9Ɓ�y�<���e$*c��C�!ǈ��i��%��q��S18�U8���������n5Z�F�k_m��4��s������sv5��fm�Ńn���4��b�{(ܕ7�&�lW��%	�}�m:w�����ah