-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
kCj6EF1EvrxeXwWZ/FMhY4dM9BFecp02fEiS1PsfbAiETKnTc8MB5793jPpQqHByfwESlAinJN/L
CCXXZZsZ2owjpZLOc2Ql6mqWEysqW3l+xUq+1ilEEA7uoGcq4exnXTAX7PT9Eak/0OjeFZxZq/55
2FVjGHZmDrmQwtScify9p5QUxhP0wlYChfKOTTva3yUWYQy4uC0VB4wuqpP2hYvwRs+/17ouSWCj
CE4wG/Nii60ydBQWpGk0LDKYQZTaX6aAbU0W7RJqZ4Kjk8UUBZANecIriXEyzVpgeI02zpkyp0MZ
Jam7okEwpdee/IIeYEgvKhzmp27O3B6mL7dpPA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 27776)
`protect data_block
0OLq0AunJDIoWtVYrAVqJUBxu+fq0Nbskx43eMS07EG55ytwekW6bjT6IFzddWAK099wZdNXMzEb
Xg7Q4aCDygnndmGiNWhLehNpYJRb7yHO2JhYe2h+2k0aW/f3glP6rvsizZGUzEaB2IeUcdLeKyJa
M1j7Cfly6kNbtAJKap7p6Nw1Lt5W6nIPXO+sRq1c3af6raxIcoeTSzued6H+BWM1I7EH/wazuOFq
XrDkNNm2qed5Fz3Ubvt9DpQEc2rdHgNp+bSsz0WB24njjWFSAVExUBUY3Zkr57JoOrBbykQujbaF
2nautAplRdTgsK8wg2vnnG313CDdZSaMlum2kxrN3HNsQW5Mv1OccAfsejRnS+jj1A3pUV63ybM6
hnxhXcLPPiG5PeP2r0gdsprKRhpKKkAPKVzAogJRgQ+Jll51FTLtZX23v4T86bKpKDX+FsqfCUpJ
/F9cSJVG/z9IDER+q/ljzt0sqxkSY44cHlEyKUjulqUE+Fwg8eVbcVaft71J6gnGx3CxPuftsMdr
ufGTGAg0BxuPkXVbHgdtLu/SRHSvmG26jib7jYyX8fHisknboiiI7t92Du/N2Yovs193lmEwkRnW
1VnENe7fCzwt9q2lgppOz3z2MuEaSikF3NTK6jFAqfZ1pVjd3CA1BBusbBOctsCud3Wz0D4Sx9kk
fqtXL+4XiC7BWGAXqF91aVYoGtTA4RAe3/l++468w4zLzlwcU5ZWYVJvk+K58eaPj5z2d83NtF4D
GJisz8rAywun0IAZlKVFCsP443KdLRMW58/IdWl1XjPm8V/rqgvJ3nriws/XNpQ5qiFRTDDTm2z4
7EXAyamRwR7zMqPo1nGaqzx3VHU1ejODPvqS2cnuopuDuVTlySLgXgeBS4aeAaHrYRSrOV3HsSX9
v/WTmAGPGYbVzx6KWcNG4u2Pomn2vprhwV+AWAJWel1SWGtVbpwPbkw1UYno58uPUCFGyaJr9/6B
gyUGVpOhwubfW/o3yxDwkuSsJ22dO+H8dhCsYJt1iwCUnrgADnCyfeMY8IJ/AZuX/rY/wPxcMZdY
ji+rHZeUUBwqWpMVJZIZVvLLodhqct5RZMvT7Btun5gEzMoqDY/OjSbJANDPCbfZ0ZRWno/jqii+
RRI5lNsOc8ix2nvDOxzhUgrXz5YpPHUP5CzE0XLhg5NzWvHHQBt1LsH7WLykwH9+i4k0k+pC2wLN
5ZfPQPSWRTEKCZUZhkcQpTMXhBzkL5IbZxGwN5gCvJwwBX0M8vgaId9DKkt8gEaL6xoINNsWjY+S
25L7dSkfRUZuKHphSVozpMAAb2Qlx0GkaPIfazJiS21iQhqVswDUDwH/WrcWV/Zz6gDFwUw3Xgax
gjNuTbPmNTj9ttqfwEJOZFT7Z5u6UyftEonSxiIEgUh+WnG02SlQzRxClvOHLC43P1XPGIsZzmJY
xWLi9En6eLgi6emsQ+t/efDfMXVWH6nmHSs1xrkevOELZJpDo3YO+EplnjiLJ6nc/DK0Tu50WEUl
tbvb9PXH/IKHtlk+NUs4Q919BWpMhHjsD8c0bv5lwXoJqb77e1RuRyutD+iB5K2x29zz41YZfgpq
SAmakrqfHbYpz0A1d+YZbKKkmFm1ypRPXRNNnpLeVMbXQtw+TNqVNC/hY7L5z8N0PYEtrA0tUw+L
HRazYLNvbviPTXPMSbQU3qv+ad+6R233pl5f2MWvq5J2O57DBuewG4uF3HpLVrTyBAmZlup/vPgI
nawD6XdvYBADw2ko4leEKV0S4kYxfY8RGP80axLZmbChPqV3M6qUynEzZkSHDjDBVoVxbG65GP2V
r+xDHJ2iBrRVNYJ8Q9IFY2IylCdTWq6kfz1P9cKYKXiBbXC3JSqg7e9UwGcyusLle6ENU1viGNEV
cSR1fPbAIoiM6nAHxmADJ/GPB/G3TtmkT7i9zyaVq1Qcn+D/QjrRO9668cwW6SWQmRovozuJ6aa3
xMHAeVFPfQX9AcWAdUH4atUBW0wnCfJm8vH640OgCNtoat5Lc2V5lR+8mOJxPxacaGpb36O/312e
MwX2yp2ODN+qqwWEGFsqgPdCa5J2xqiHJcHMf/QHtFgTLtpc3wmL8KSXXZViq2wegP6EPwaw49/t
Kp6gxmX47GFcdfY8WPgISQ7OFIEvIkZ3cgXxTHgDmUYBwuUx8gE9S8doXL9s6aRkGKM48IQw5msH
OsRpSrMKygK48QIngSAuSxEbpthiJw+9N9SQUmoUD6VArFZ++zD/9Dk1JWfe+YJHizD7Mko2TPWQ
U4iayS7MPLjG5O7LejwWQ0TDFDmAwrP7EoVeb1AvKueRUBf/DaCEJTOWKIvjIxaRuEzM6MqiUfAF
ZvDC4oWRCINZjG7ZPnP89Pp3w03/5sXCopZPU2dPJ7l1+vD2GpaXKCzwtlImlqEh05Dk6axoftIL
K7WUCaxE+OFsoF/Wens3qF4I5sVGNcvGucIrrytWcfNpQYLGB6EpU/TvMD8v1LTfOd0Alwjw90k6
VLUpm9V4+qNBFbLkYsj8USHchtHv4LYgHgOxcrZwifnATy0/FdIOpzjxHHJCJS7ZexNu93gYw6dj
lavqmHHpJ22PExaLGxheJTUxgKKeWomnMt2Nz43yf6GvQNt3yAqZZRXK1SlCbuXIZ3J0sRZ3x8et
TsM26fMxMyF742jKDmSDkqnZCSM2y0obmGWdX281D9V1FaF5K2n+Nhn1aP8UmGSmYESmHTe15UYQ
iaMEx03bV2CtI9hRAN/Nq2B6qGrvM8aIPSmjtRuIF7zoslUdQisRecZiV7ngE436yd/0kLO/xwrm
sQYv1Vh3u1Cptd/QnQfmuaS0mXSS/344rBikb+sj1+whtVhecoP4LUclI9uGE4QTDPuXrxRoPPYh
/J+fbbFr1Jwqi2sly4iTcCuX2oHXr2ynekoufy2lh+BOvNU4Z343sH/Mem4DeBhAHS1mPrqXoVV8
xltCmYyyYhD5k6vJKZaNP/clgBEjoY3QLSkCbuNG9KjGNyd8W6/mWhDwsBQz6DdC0OQZucs7HFH/
LbPQfKBcBRCPI3T6xe9jCZE62krBGay1hmDA9SfadUIT0FQwgA6vjMfuIi3+RtDs3Igq4wceHA7a
wCeYK4tSrxvg2nph5hzplBHuM8QO5FEqQdmMaTXnVXtXYw5iucma8Fl+VsrVHaTQyDEaWsGedzZR
3FVGlzCmO5ipPESoI8lwWr0Y7A9CJrtsr+WSqswwKE15AXHiWl3R4kc+JuP2BFGWcpDd9RdegBCW
4vkuNM5VhWfHY0baSm5gbT6ocKRNp9JJORjTRowIYFqnSiiAlWUd/hUgaoqVP/R2HAP/LIEuo/4X
WtPNtwVKDk7BWAASmW6Dw5HElQ6BpVXRZk0XBKLESFto+m/vMdEy2ONv3C9fwZ83iftdCbglHaJk
lD5UQrdHxquLGeYCEP1dR+bMRDdXj5gDPUycy3TokQ33RuPIS3u4L/fl+9ghg43hMBLP4EgFwVqk
exKQff9wSBcichEzroFW9BrywZSVxxupsz7Pq/byihAz0td0RlYRXz3w8qkOWc0bQeU+OS5o2Hrj
3hnka3pDlUCfndqHm/7qrJ327ZXOJMcnxLa2nb9F1UaN7koauEdtkX5ztYpih9Ez/CWOlyAeO7fQ
19s1CBAdQQ5C1LeVltW2a1wXK8Y5TZUvlGyxtJx+2LoxlQnRCJ/Oc/AxCw3Vfzo2dWaM1elpTVJ+
1MVG58K0EqpmT86JU4N+UHyx9M0whqlS8BTObw6j065Z5qJ6wNvsZjXiX1X6gLysUGy2l5JggxFh
6OsWGZv1GCvu02aS/ebg5oI8xgJDtbjvKaTQL+Iq8O8QBTOXUdpCFUCxPFsASc13mBPojihWSfzH
GGfZOfDMspN/GdgsnA4MrNiwQXzcf0YAlqmhLoYLE6/mRYoTfWjjxowK2vVWQM1Gtm0nhiFRxatz
GnK5MfV5Zyh1i2EQxpMTdJlMeNb/Or8IGJ+lnM1raSRqvWwgnWeUwLANTdLNCH8GvosatgjLU/fT
HDknOoXbib5u8uDRCegNUCi/F7LIqQXCsslT1aLtS7j1Y+xdZos613I8DuZhTu5Nik39a23WjZGO
YYg7k4GtkoCuFvaAIyONULHM8ZhCFQ/CKj1hgKK1MkiH5/RpXx0WNtAz3A4+Mu4SXbL4f9GsqBKM
Xz6bztCU0IQtP7S3qugfSecHaj/G/77QNl0cv/n7YpA8TkVBX2H5coYC6uC7rrqCKscpB1Fxmmew
/8EhDJTTSLrHa6xvptPX0SRoaCZpVqkuOkRhFLH3tz3uQJkQd437OVJuQupk3MkjusBHEnjBU3AS
6olM6Enj4AdRSDeGOAy7zbjDByYcWvwkfr+Qs2Z+NWWwLmDRfVqnhDSn0Jt+rVsLLkgSFUfEYnZo
MsZNIMRA82DTl2wwirRZSM/sezBgRRGZZHRBYw7WHO5CVajgQ3y0Byun4F1k6//NNDeg51NisU9V
ckbjydGdQsaQB8kijMXHSgbiUjLCwMfw1zdJBbQANsFECFcHAMUvbw8/0kY0G6UdfmFRa4pla+ZH
T56meGzRSJRDEWp2WAlBQp3mZqjLSMFcVY9CvqEx41OS7QH9807TiJ+U9mGN45QKaPTYmQKMlwvj
hJV4r+nJEAoVXPe+AZFjByKc+hBYZ+b5EBLBgD/svH+dmybfQ9lMOWBd6xcesgkQtIkX0UZ9lZ6i
u9sfFTnSx8cbProT6BhuTronSZEks0bsMzHX+C/75YTvAcltOCOgFy+84eSapcpG7QMqLHezLVgf
E7w6fa2ouQVIpnZ1PBnsvPCd6ZafWK8zAsJs+EDogtfFR35Ii9DA48GYML/57UObTgxFZWocf6z1
kiXc26VJW8YCsWfae7YMZfbBjiJD4GY7l3xXKqA4f3bF4RkPoi22QPNuG88hLcB/2dT0/a5NHJLg
dI3eB30/SjznY1XmHSwCuiT+vacpCaVb2djiumZfyQrrVNXidS3tygntM3HEO7u0aJZAu3v6/mQa
iWcT2fWQ54wSevpVz9ZJaP4H7zg1eAKmSLqUh+DMlI52DOpGhU4GnZ0/JzrEE5RssuIuvGZcxSJP
APKTUQ07dgVgQ7hguUgLHkRCQUeJzRutih6n0oGI2gHhk2+NsFm9Fyf58oq35Wd06BUix5Tn9ucK
OjSh8LRtnKMl54FPidqRqGpoAkyYvVxTOnz/tBkAiAsTGxlxpTpqa23wtERaCNdzdFOkckcGWiDc
lRwbJDLONrnFKjeDBNzJ7uHQNlcKCgynQrU8GXtL6B/b6z7PL7/yyhewjE0COdJLedtTNoPFkNST
WKi7wLeEuE52r9REt/wza62mhzaXgdqhKFk42njlv1Y1AeAq4ceVNJvyNpwCT+VD7Ml71jFt6XKc
WGjkAdJT+J3I0PpvJCIFjh8YNfIOSUvdwy7rlbFgRp4Ut5f4WEPrx+w5+gtpQ3nq+eWwf7ehV9m1
PHnWSM3HbgH2BO2JotZvA+Pe8tuhzXNoJIgCqsqfeIJSs90dnXGEpUNaotD61C180eVvefwYWSzU
xkPPxW7iAmgLZUTwSQJMvnucxxcsVnJtTyFTE3/vLaWCUHWry75yQLStH4bUp6IrlToLzwZiut88
65AlFvXXCe0eHl0VJ0VODhJhZXyKYXXqfbStOPzMcFv1mkZW+OqqOslxIFKmsHGws80MwcUrnPtd
zZ89D4007rr81i6grTLVQqEuCGuRhUm9qN/qt6l3h9udHH2oPaFJZxKhuuApbbmD7vrc3/QqnN6w
aeaqD/statnNUq1fgkAXJWANjvhFMUZcfYjhGH2PBgQJdnje0yUs5xSVeJFtZfrDVxRWJGp3NFvb
NXDEziR81Z3zLZlrbyeqQCg1xW4zDxkmyYJ3ohlx1eCV/W1RyBuk8phgR63RvJ5MEwZiXi5L/lKJ
/z8ZfrHT9oTY90sCR6Nuc8e4gVC8SAPm5hQNIi0amywE1uqEGkMPCgDiqBlLcqF2qih9es8TVcFC
Cm4GTVUY0czAF+BSQqumsipkg7i+a2ifAn9HzjxLFj++fZ6LkpZMDptt5JZEtFcRz8Sxtfmz/ayU
5NkKcCzF1LU0FIHjd+9405tJBJrLYZSAVbehbvK1wEfqcLO34YZnRY3Qq6z06qajPaTTxqk6RETZ
PVGnnRwPWivA3aia6wYNPZ/Z3CrPP/yzT2Po01iiPeuRxFtpq3Ik9R2NW98WWvvTyTpTDmqXqZg5
dGg5vrOZ2DgJZ4PKhzOUc1WcGLf+Mywe5klv8z9KEVty8C8gVuznpZcY1zDzE3RVAPBrEnvgkLmJ
Xua93KrQJndwiZpooeF062qgEVMWe2zFvD9LJZcgOi/77JO2+VpdFqo2vyG+5Gd/VatPbP6yCNxO
N4WYjiJ4b6f1JMU5pdalWNTIlUmRzFfi6zosy/P3dvGvTSZtB+jpzojP1DkgCwxFldackj2p1LiL
WrZSTpRCdAk28fc9uZiaykw0CRBUnerk4M4scZxuszJ30umMUS/Ce1xJQP1VRV4kLO/DdIkAVf3z
fVLLIECqT1Khy3bV85woaz26SH2i43em4v4x5SOr33ZbE3rla7Bruu7XRyQSKE/mlLA2mdb8HYTP
6A0ZcbjhI4dYacuDqmQ0WP8okdAMQwuTPd5oJRRx9ghwG2YV5bBIluMtNH0fV/E0QmW1TC5eQS/c
TM0dCtOx48OccSzBA6/gGAcymH1KBOKt0p2luJZ6Od4N1UiZPnxPug6h/oYZ2hqNe4kRhygol9lH
WLCRwtMbDM+9sukrk/05gfR/igqQxDjlLBCdXcwtwEDOAdq8rkjumP9wzcIIQbZE+FOSTqwDhGYK
7aRtGM8MFhtmPRCEIJJ4auHXo9vYxCkMM63yscz2bX6vZNXdoGBRGtmOrvwDnM1uHc7YjcT/3OS0
3TNz9AAq4Y16f0dNyiZ18BNgMs8jsYRAi5ptcXJe4GgKUb+CemzJ6YdEFoaavebfIG+uz73Iv/n8
4ioeDrqdVL5gUxZVMmET7/yYjtSLSKa8glqSJVkL0f5FJsGaQ1HVgUMZiA2vQO7PzUTT1IOomyQg
gC/K3RwJOoXZclA/TrF4hSWayCO6hfCJL8nOra2omFJKrT1lJ3JVyEBCl4zXhrrjzcYudKjaI+SX
yQMzH/ad1IkES1/NUuHQS42sB9dMeZbcsKZ3cLKw6nDkdeGRLvxRSFd8F5aRijPnuKKnDfbjKrLN
JHtr3q85OIqX5uV+hqvGVOEtKPdEvRYtkNy6HVJXj5iA9/4K7sajDv/++Es1PXLjqzsDkyTs7ZSu
lxD2KMXZGqvHFowZ0i4S7sOWSuB1b5Y0lr/WAQaOf/TmBVELfVLu2JjjUoZ8Q3V3yfgss/cfN9RZ
fiLjBdhtQ+9SGgfVLSXTjbafeoR9STs1r1qm2acSHDazs9PeZo0OtPm6JBIExeGTJKGUTGRGwKm4
dB9kFKrmEhDRTdDLit9gUfHUIGgw3ta42YwDDNrHqMhufcIv9orV1P96VJnAVw6du4PQk7laHu+3
yVrYsj5PY3Tmd0c+fY3XzsIrXePB/xOgAW2X6FrJrLsKObXpCCMGQf2A3HPSZPlnlFJTi5GlU1IC
xpJ1kcuUdRyMq5ANDwD2MIaKEiIAsIGOcm+7x5Vfu4cmOT8UiBf08jozjASulyiLJGdo76XZ43DB
qJhnPpn1Yz2bTi6pqaVElttzDD+azsGuMUK2HsVPN8sfy5/R82xE+To1jaxy05GnNROUTeKtTZHO
dC2dVaFtt0+BG2i3r4rsMv7GN2CC/Vt5rR+i8Kd6WBjEvziVz6WQIfOO9ubHs7ndd26UEJGxnOAw
tzi1Q/Do/8U3WGgViQSSPcByD2oEjJfSVTPT4ISteed/g70xxgmYwwg86IhRA/ypSWm5yDGrxkPc
2ek5zvEgWvZbRNxngU8ON72hDVfWhKh6Zqcb0o83amRZvz/HLIorsfQZP8+oHUMi+ZQRcDFBZNWi
9aG0CT2Z1CvQCUAPO11E0yIQzjscuZS1SqPofXrQOgl5u2WHM/834jstSiRcoH2PEaXUDdVEllI9
VCLXO6lI/gqWUCnt6O64EcP+DfBxipej5bcs9r3GbCwKsix1+ZGfMyOmNdvCFtTNPq9YFyzq7U69
C0NiYbuuGAuNQ03igkzmNB336fgQqi2gluiWUaX5mLaQ+7/Y8TGAepnh2R8iQ3nUaxRnUHGkLYPl
ImYnH19ZwDe3waI6gcOfwaqz8vrIbdrmhnq6aJdSkokQmcJmZpHisaZesZ/kC8FyN240HcpegPyt
SQJb4WBBf90G1cV6TAs4qucphCBI3PXvyISSbLRn7KG4ZE0UaLoP350jO683mFzCkp9rK8wGD2Nh
bD+eXOmzQMoiv0YjCejTmF98I8X5zqfGhr4u2lmyqiQLaRR2+k//ftH+e5U1pRzAezB4pjsCVxSZ
gZbXz24N8u/cmuoP4kLRkkQUPmUI9n+trx3K0LGROVl7+bhZRPYr94Aw1ATueUADcFwCbDsGZ7hc
opdhrPi6Xrd3n2iPJedGEuaJhHUcy1cdzl0e5+9LZHItT4HrOUYNiZQT5wFIr+5wNc4kdp0cEEhJ
ffiRvofOwnolGPBw2ZhZwlZAV3xk1gLub+frBQ+bD2uuwX1yD3tVHXry0jUWtfkPT25BllqSQnyy
YwGN8D+TuvQjtlSQjxTrerqyTU0FonoQlIenpPSWoL7RHX9a4MFaW4aXwDZhnO7bEgbYc3ZNA53E
WElqAOOJAHIxErriiwJBBKOtfv4diwTjkG6ewMyV0dfWbQdYTQZpiqi8y54E28YLfyn0Q/9v/Mi9
T0UMCqj2sTb5g/TjRxwW/Ym6c0AMO/bpjrXNHVQx2zfHEwVQbePaPo3qiVLBDcFhYRXWaBauBDhu
RW1h5boj9sStnbI+1aDrE84iJjEY0jYNCY5vnFqpOaTrIGgHMFGZohN2h6IAmEgVT8LIpCHi69U8
xjE7TxyjW85IHFH0KdNnQdtKk3fjrVmxT5aJhaKMvokHrRNplf1As813UW990RpaqS1artW/hCLC
TGnu21bJHk+Ap5SNVxghHJZeijr0N46wOY6RChQPGdFAUiQOnul0XWwz01y8xw5N46dq3UF6GlAz
dG+vjT0+uEh27ijzl2o5WrpuMEw1bZQJB/VkYMnORrdZI+a1pB0pqKqeAoKQXk5TmN27I3pX0YaP
MUfFXIP+pw98sXgm4IJzlS/I/OOmIKDzhn+Hk6ca0690nIGuRZwW4GdgZEDLl5q9EGCE6osr+z6Z
xHAnNc6NG6T7BofnKoUYRb9PLZMb1Y/PHW/3dXZMeYbrKObVZGAZQtZi2fJVTjpVJjrFzAgLv5ai
eyRlrQm9WCEkIBXPX+1hAQIy/X1XkW9tAqGSrtg+vwWnnVauoseq8WLSuMdKSnRK/v8nANwKXVuj
He1yY0EAvmIItpwPUscYuIxKyllN/h+sO3kDIdWWI6/9Vd8/x9TNUAlrz2bYIiby6j5Ipz/eSYNY
10XQSoKT2c+8GNP+6EsVTOdO8D7KdPyyXcucJhir9khoFIlSwPv7Wn5mNN2wRmvkyr9WX4WVkdw7
LNAjs1nrrNf2071hqLNVjaKiQMXw2wbtVEMruTEroFKlE0qGNSzrjtFCoWQFgd5Z8iJdPchzy6rQ
BJ3GYMMvZGfk87D4poDxMk5eETRCfIbcG87rEsmoi2bvJDXpCLM3sreO/H5sCiF7mHKjVxOvMAM3
zrhL6nGycePazkn2TSVGLTUyq1T3wRkJa59TjhEjG6dMAk1Xt6HxD8/pAUdetcyVdetKBwKzZfPd
lCzCt6PPiM5aIME+N2YChq02ZKMEC39qSDBuiO6hCgL+rn26t9xv3RKpZA6ZGFqgme+PE5GxVj3M
1y3cpxetPdIXOkhRRiiiWvk7UqSB42gPF76818aSgvZhOymonvzCWDdktmtQf3LmkwnWrry/lKdo
FSNQyX3COeQ0saD7MOu7x9A7gPl+sC2913QTVXIkYFQYn3D4kLba16S1phDCwNp7jUXq+X7imrtG
VQdG48ZdqGquHtYZ82n9zgIq+fEVWrYV0US6YiZdPaqgDJSCgXCqlY04P5VZYON/4A4SHCsDBIw3
/lSenNeOcDM6QDdVif+Ru+OxYnx66874La6bC0p87HF6+KJjjtWshI6mp9DzkORX++z+GYmalL3h
ziH3L4iWBJV79FVm8RCaWs4aReQ4d1ixR6eCoT+bo5k3Ui0xqO7H03WI/NtKVP+xT8hM1nFwZXgA
zR3aTM+1cXNqpd0XOVzt5g85hG0uFQW5ZgITEUV3qmLkZ52HQwy5Bu5wsJGLLWI6buaD2AM8Syn1
3dlMP4xJMdBcgBw3xi5y7PyKhToj6/SBUI8NgM/7RnE1PRrlGhPSU2DdoDJmtsAUXibeO39NG2Kk
NCxBbKYK+0eTw2KiBBraGue2refD10IYKDvvEQkREb7vvxUY7SydQwhCZIv1g+m1TpC6IM0UHvoZ
hbM3+zKeE4pspaijrvChMUmWKd4aNT/Klmkm5gX1ZPPLgRyT71cOGDAGWTq9i3FcLoWx0GBPz8Yw
+AgMutmh4Y0uHqIAu7CXtJPmKCRdO0J/vpLUB4d5TFEAfYXguWonAB+G6JbxAn8i9UqDHP48O+h0
pjtztzavuCRBNz+ArUJkIfXcqBicsAUqqTdy9dHD+wwFUENSSI93PBUTxE5EQ5kXU7U7Ock2KWKj
rA1ZDFPSTlMYb9YCjDVvNOeE4a70XRY/KJDJngmNLmhB5S/aG9r5J+LTA/KdOzqU4JXjVEZUZzeG
IlN7fHISyZ+keNFpLqu0XXUw6GPu0oqBWXKjy/1znS64GZNx93xLJws71ZUgX/LNRQPF/mC6FYeJ
3fIfXtDAhi29yrXxP8hLqG8XcFATGECv34a9hdad/Rp9/zAaLyjncYOuZ25MliiJ6y3GoPqVgQ8a
9GVLBlfZtLNCbUZxbB+7IviAPEyvfVFBakTMeg2yC9AUzxYeU8gjSFlCcHfHLOtE9kRYtMbO7v5c
dGV/5BJWvyQV/NMfkiuI7finaqW0cP2ZC+dXdLqUwHb7nyOhL6T7G5hLJFv19N6iaja/PUSxoB64
bY8OcS9lh5kK0UHXCQOq7QTooYEKTNSNxX0Ua9xpX8bhosdJ8oDaJ8KeAQH7saYpi4zrPU0z3FYD
RLcWnfxRpDHMMuWZG7Gt/S4yfJmAHJzXh4Kec90V5VcN8/BaOspP6M1eyX5423QiOAwkP1ILleDU
sdziZaQLU9Lea63TbQ6F1r8+7OEycSFWNETU50zfmwNTx7XEGZgq8bOnVVKR24st+7O7nhDVSXM4
0Fa7nCS7GuLUtTFpMHr3qohWaAmt1OGFLEmi44v8Wd9gzoUCwBwNNT9C0KcqI0DoqigsYCEPQa1N
QskLgbh9bvIE6MROkWv04YDt6D0hIvAonlXxo23bgJpIem0QvyZSWZ6cl4seP+QoL0b8F9mg5HKt
yTjp9+pBo3q3YSWLd4TfKeCcAFMIUifCRg8qR4znVY/GgJi5f9kfRsxWEmaO9t6vXtGJ+9736VI+
hN0X8X9JCkbv6XCN9ZTu1HlvJ5xl9ak5xjgzIEK62YAkGEiMiQLfiEmBVm3CZ0vph09VA8fA9e+g
WgAhHb5b9PWv1Pe/H5gkqCy1p2VchOJR57mVMPc+g6an/Viw53K1BvOCTdTV7Xap+rHRzgPMC2ij
YQQgti4cE9JoJS7+t31RiKF7FlK0QuP+Ib8B97izy4p00aXlyQMWTqQdrzQf5h0MVKUnnTt+7snd
8SehkYHRV5b1szb4jIt0PtCaiAO/sXRlEl8CX9CxuT/pvSYuj/YxBkR6zE9JUlLto7zSqvfk/5b9
8i0eLmbEvHlnbIaMJKMtmR7vnMa5eeGG8HLjgB3yhQoUrjg4q4V/Ujo2oPpPhy6ZIPEwHWsehJb4
yzoTKrE0h6f/cbF/2THuBKbf1bUHXMbGeTK/3yaRbXcpB5sEJD5wwW15aFjCzyPA4dV1xppBpkuk
SptuPAswo3g0TNhjfTH1XgrP/UoTCJJHITTeER06A/K7+D9QgaUQbh3422KyeyhK12nhIwT9dU5+
9bXPzWVv9WqfbEZniG+sA0rCfTbcWqZzbGnHRFKhbyv90jhCexcuWSvWsqpffo+SkElrUTnaukxo
381wazrUQg9XtBbTULpsccR9po06pbgzvENaAvUNcnL2q1CeWwyrhi1KP5B6poCd0WfEJsac4Fr6
b9l5uwz3FrSVT0I2x6uXEELZSYBSLHpfX3VpSdAOc2OLADoRQHI/QvnHfQJbjJ3+uVHGD3rfb2sh
pFxL1S9dS/f57LJqNJbqbqHBgIOL9Lcf04Jy92M51mjrBuzKOa9OgeuAUs16fIpOe7oJYF3PvYj0
dqRNDR0wjvIexC2CFZoqGz0654EmFuxGI6WOsYaom8Yyj/ZiJKFlQLNow1krgH32kykPT5QuVC70
yocFZsl8RbjwkzHcHriQhkyat9e9w2k2KZwnYJ9rQaQUb72UvLv8p0kFlmqhy+K05qPnp54149YJ
dsnTU3y1yBZ1gfXlQzOS3uFhJ3Rg2548ee/3OOsBk96K4lS74ehzW24ZR7IEXnOXqOB4/PYUpbsX
R12ptgxiCj173PlnQS4PVGetodZ3XuTR6juWbi8HwQBpFOP1dN4x/HjMHh1u+2WzN9LEr2YZtV5V
r+yKcakgbCpFGRjALzRMXpM9rw4prrOMPt+VSMA5V/ZTqQX3ahS043ReS0JINtegKcWs5xrBB9eM
CwRTlSOGgjG78GOUs8SykCV0ynnuM5r9Ri6tDtrvl7V9GJxu5Ls8zzNeHu03sgMRPeskzGjtJ96j
mz8OHGZV+sEC7U7i83eYH+vzq672SJ/MPXDdcWRnVVEuZljiqDDEc/7/zndXqwgE7jvUWKTLcN4A
oPP7CebZwds1b6LzfCKt5P2yxd0FXLlv10/PrYeRfTu68TlJEB/v74MuhTQlDaUjVQ86Hz34hcD2
wDQQfA1hU3OaLnfpZEJNscyD7mt24SvLCaNfWoIAvyHD3UbuuAaD9VqIDe3TBbvcvKQY92PQ21Er
6mJ1vYG9zlmdxbm+qmFIiIi2BsYasHxMM2vu25BnC+EG6a9ko7NJp9SYzriIgT9zS/VO/2FT7bTK
Tr2BwJ/oALnXnDoOrwyAY14W6VabY0Pf12n5ArBTQlROZJpMvDUZaQ3O3H7Zmxa8N3mPMyfnmjoT
7uQZ6/94gkbTciC1dgI+WwIQbRg2eAtGcNb2d/0QyPZFvvk5G2rmVwETXdVCUDnH+WOaE/BWYXKD
4uf7y/fFt56rytrEj9l/+IGjuGpNX/87MfBllehyHzyUg0oxl+eEwsJwtqrSccumzLyGgj1kj9W/
Dgjs8snz857wrCYQJlX2TjYB0SP9j7ET5MtRWxWa1WdOo2eriWKWyVp14xs4HHdgqXJyfkSaGEs/
ALB4i1i1OOBP/gorFcQXoXAW5Jh5ACLMEhc41hw+Y+uiGnZL3gUDJKJ4M/LYjLeD3An5H9fADnjj
5sLyf7GdI11cW97DuYICivDV7v8dwNzuUlxOjXrQ7n2llJPLaYlonpT7f6kbYN6O3iWJPlcLEctE
Defr3o/4WJDmbWrA0hezhoPY/i1wVB04Uh4cbQG1SwyYfZfPi5xBOTMMytKUWxzYNl5Ldg05vSuS
Fb263D/5p7wlNVIP2JVIpcPEKDKwZnbXSngMXpElBPFd8PTofapLofKr3lSNb/fXB+yNXYfpl/wo
IsZfAGuI4QagxOqjOK3EbhThUU284Vm652XpToMhUs/5k64td3K4LWN2XxShOX6CP8LFOB5OLAEY
ogD1N1wZUOBV1ebjTylc9gOLZckpF0O5oP1Jjbc1V0BR6XSqjgpwNTY/whLhono26K12i7VbbiPe
/strPtYIMZ/hJ+vzFzgqnZnQ57mgcZrNQVkkTz4t37I4bm33sGpTuZM3l/GhDPW9ZTwggb5RepNY
6UAbklPPbNcyGb7OPUYQFY7kQgHInNzlE+X7zlpzQ3wNVGIA4nrGfliP5czrSDKXFrs8n0FYOxzB
udiNEgF81dnjuE3yWa0165QhBBvHdJhAdqXsitZjWCMRF3U/dXoZX9a73gWoKIYzrTfwuGg8rRl4
KT4QkAHYWfhCNiIsFyLby+6asHYqv+N1hPStE0uzdXVVwW4V75APwCUq1ZFv5YBxrYZ6KhlahZ2m
Dj7yQwWXCYtjqmNGWE2ZLE5WDvfn+OKpuGY5nWxsqzf+AY8Av3KT4Ir49RgKWsZXj6B56/+Nhtop
RcXTKyDVuGTX0Y/GB5iCFl1b0Q1xfqWjW4bH2L3TO0HItqLyiHT0+8t8YqImBaCpCk7KNn7oXDBW
9FRff7uaVZLbW7G9/37jUakRoKdJJMQkF1XZvxkzeBgqpSVE3k4YcNOsn8BXYDQuI3y8fD9h7Ozy
a4ies0RouqrbvCVzqd2bJkxUMsj64KiaJyM60491to0dlkNdk4mp9kirGfH0hgaEKBqpBNSoAgpa
ubif77LzJkAlIkNikTdebEouvTnZJq2+IF+bC5N7USYNUoxtVdEVrHQckxpHjbcBfpq6uDo87I+L
sufFXt0nfa/n2Iyxd7+ntF/UGdSIy8chW/Y5lx8Uis5Zhf5gl/4dbZ6Gw/bU0sV1oafMELmPUHlB
pXf82Ve3i5DXQutrlNE9rYMYpRLlJYeYcmduZmJtjQwVQzASDZpYRsKc9whGz1ltcLo2TmVl1wX9
AXfb+jF0SuCw40/TL273j6MwQ/hfAefJpP2hUjOOpeYGHvAaZ2y4y/45X1SDOLhmo8+lqMLx4JVL
XWrA8RwpuUagkMDXvyr1qfHEAD9Ls1g+IZCp/EQ2GR2yyw2RXZBjOOcw/23JE9Ctjk8Tf/7JcPbb
ylyY4iDZpiTPv6ec6LDB+wqNRPqQ29trOD0PZnmA4gHQzgfI80gUgzS9C8y1mwKYMTpU5J0MnMCE
6yjalUjj1mfcWR/AWqR7JMUHS1xuzUZXav6NFZISpYkLfDZOzAs9jMsSbORMg/AUfZk+3yzWaI57
Ef/QyrWZpo83uau1neMU1R8rIiJjyjavnYe/bnwh/Hr/a31Hx0LUu+N07AC40wnkStLpJ+/B6wM/
ZJp4BOJ87nau7DoBHgGYFAn6X3ySpDUydRSRNr1C+KcKtUokB0O+oL/CIYn83/7sUc2QF2pdkpn9
29FyBWLAxbdsrPN53Rt0kEJujiebyQh/H4Ds6Bo9prwMo8ZOvQEURxJBxzDO8Syg3EEP4w8c4Sqs
sS4SVAPXOiJICR/wXICkbhk7rTN0dHGlXcxPCLdPUYx7blgMTGbcP9jo1EwdB7kO/HHeeH83pm0s
3ReAKUZiSO+pjYl437pJO4UG+4BQCcEm2bU/+Mm1dhxo/m+XJqFUtRE13MdF5QmCqWPJE6KBglUL
OoxK5E3owW005i4OoINQCCWtlHuUPqtUSK5z5tXJqW/WDwKJGlZmHCJKgZMapbn4QRCxOZLjKUGy
W0qnTRBgfbV2t+xCNd0nP+9KsUfr7RRsbi7cH7Rq9WLFuFzW0Qbm9r4RIPjXGJb5pSHHNlF90xSE
UA7izWQ3ykUUGVl6EOEEl1t0DxuxWhIHpm0ZFOKmCv+BzVMqAtHiDpskOsxHRGnfRDaDRwJvWt/w
suIQRTcsLlsaCK6xFDFAN7Fm+6bLqFRY8BRDJdPdQRSFdHKkQHNtcTEAgbWFAnF5iNMlzckcoyKJ
4OaoGVpf9cOKN9GP24RK1ExI0LmLTl6J6eSsv2aR0d9BJj2CAq8Y7SyWOxgJCK7QG8vFnwQC6lJf
aKg9yPAj/+92J8P/vKv96yBotpCEJasnKBkXXKk5ghHputZwZDWeMy6ax5WoeuP8IDoRbqYbfTiB
4ccD8QZos1IcvfvObrIeWARnnxKdSaK64cPxz9SD9GFuFBAnwgtf/YwtxqD3l8No9x70EgPJ0dEt
1HwpOeuNfIsMfc48EMWIvSbC9uSM3tafgCA5IwJA0YdtwTg+ikjEJ9QUTzMrERy4Vy3zIcnO1NWw
fxCJgHD5j01AJnimNKP6hw02rDMa5WXS0IbZRmHRrIUmL/R/Y/yZwpKSH5bdPqaMJVnN/1uvsGrk
Dneu/88ebHWfxZ/Xl+Lbozs+wxHsXgv+kaGx2S/3/hv9kBTq7adaujQsQqWaY6q9hEUyJXq2jTLg
vNtHDByPBojIgrMtOeKF9XmyB+H0Z6k/Vne5sQoS1T3MNlcYOkAZyol9+dVwA07hDYHC6lLV+lfI
Zx09JkTCITEPwG8tGU0Qz7/aBl6FfoPnm8cyKQJ47bae9mkTcGbISiVM3VNTeHpON0L9siwzElce
kI28GbW0oycf/902305UGrmgDNRkIpmdGoc8mrDk4IaaoAiBaPhpjwLMEUBWTbtzulZOcd8nIIEx
UuEoHNoeWuwgdS0cmoktgW81A7Kh3+L4JMg0RpMwojE+MEpbyIzrI1mGH+wVP1hTj7AZ/1igT968
M1SVLSIrWHh97etWYAXFoNOso0xPDzuPcsBSsNom6WeAosNF0+ZZ66UwjXVILdmJOrGpXOmLTH+N
IrZThmwu7bbxdg8cJE2w1VuyiEWYliV6rcfupbXF3M0tppjSYNDYMec4JrT8tQq5zZzHznSwlD6R
e0hO/V60p3nR7mgfhZ1DyP/GrV0wLT5TiA6m1txYvCMsv2HUrvrF/GUf3XQMBzqRobw+mbBSD1CQ
8vsU+PfChnSUTsYZqoGVIIJSP6Fz1zZk1YtN6Q+ofg1t5fIpfVTaTXLIk5TG0+XJTxiH7szRhqSy
h8Gw89evD1fXsKmKeZMmPADPOuPyCyX1LeWJZoxy92s4F9duBXnwe5bWAvwXM1fROY4x/bb/Vy23
ccE39aWyP8LgXhDXV0rVNDH1Ui/7asaDi8oQpx7kcgVtnYVOTgy9dtTWbmCE1KBILdies02yA1OQ
rOYmoZ92+9BP5riPiq8V2TVLtz2grVIzxbcBAKghXjjT2+S0UNYiT5JtkPF7RXhFAuH4bUL2SguI
hrTe2t+0xHXfH7WYunJG27bnLZd+7lM3HKmdw2KC2K7fu7S7RAzSFWxOUL6QhJgafkeKD1f/Hw4u
mNf5o4j35G+vgKKFkS50apoxNdyY9sbR9Jvn5LgRddjKdofTyf6Bwnmml/gpXGQeZN6+F9W772c5
6EBtUTt/EvOtaAxOxfc45CPdA4aIpv6LOILhwnpih5pZ/1rHH5B45A8kSmNl6a27XXhddT2s/xfp
6x4HMJ7qettBsRBCf4+TFoYRVusz/Wlf/vesS/uP24GgY4+/N21zi0bkmnelGE6U4KCnnyscW7Eq
N9GSnAHitUTEA09wkxGbp64PobLxtbDRhUD/iqRUVuamW4Ug2irrcCPmTEuea7kw0BHF+pb1m7hH
DHoYD4Oux/X486WP4Sjos5K6AiJwWDddO1+neDv5Ob1Lws0Z8wWrQSxxtLoOPYTQ5JWYkSpwL/9F
VtBwjGiByWFYnkM4UUMkHa7gsOprHp8h2TtiqJrYEmc9Wqgw1UEsU3SYKga3rtiGsFPPiepASaxU
grQoRHcUCk+igktHxe9bZYsgasc6BpDqpp1q79ICfYB2/jG+7b8MdbAw8CTODtIog0Oh3ENTNttW
Fkh5pVK255O59sNM15NMXWVOws30xjzraevcSJ416SSMqCQFPbjLQWPn5M4wMMxuklzfpGEyAke0
FzecYAgNfV9K0tqHjn81Czigb4yTS6HQGbA/gkvY2v99ct0I4XX2We8m+2sH67XDA9p/cdd1Vrph
L3Rybg3ORd5hSPMaUBZyjwH70QVU6rIuJVvZLYSgiFFi7to0wnu8fjGygMCP6k5j23mzk9rhkCaV
eGO0vAkMnlSBegfQf04/InmH+fAZXXTT+Eg9qC+JVfByuZaXJjewiUHg78EcdNRoVuajRs/54ix/
Jl4nGNATKuI38ysUBFvqfyY6+h5+nxPKQkLXZxuvbE5q2ayzOtKJth6wjXVBr6ISJisVbE3uPpXp
9IxD+gaSYHDOUS1tMihjy9KGGAuu+uWpee1nySrst1hOigEHZbwcnbmbCK8GxOacaquGw7T512Re
DvR1GfvgiCE/Qgwnvp67vS9mxBHONk4EYg0u5588yEg0s7H4zGHocoXCNlE/WU4tGDipMFEx9qDw
GSONY9YMjdmzG0ccie3nVBJm/LIWfq+HMNI2QoHmrff0+uiQ1NkgsQ+Z5qmY1qSO7Mr95y/E3koT
8Z5POFebqVCmbYl+VWD89qZOLLoBsnw1113NiqCVqeSVeBWDqCR0+lDXTCCNw/s03ADbIbKXio0M
dtT+Hkg8jnqMd1Y/2rmUDhl31hdipGceFUrEXJTl66Ky0RzUB2P+MNeOCcw/HDzn7kARI0r5Mt7h
tOGMjAnvkn7bY4CgaLmBlzMXSPunPKgfDmkeyeGxxxjw6wmf1Zge5cVg6mv3F2nmP0zdAdqHyVRZ
6KiE3E4IMllyYnsc2Kcf2LVDNWnxQF9A2BKEeJv3SoPDDJ98sDiCeb5WeOjKBLL1OydnoItq5A1F
86ZByn2iodu0rAAHHK4F8xYH61Y2i8NMhA+yGGb2TDc6WiO/sfe94AQtaP8XVCRDFfE1FeMQceeq
QixpLZ2NVAwogLMZPoOLYMXozRgqdHfdaHCSHUkawb3qaAkTs3JzlrpY8287OE32OoSkLG8HGvAc
k84CbfIGVHu52kGm7C3uBTGVbnYOcMAuvTOYwQf7KY+QH5zHHR6du+JToBODthDm7XOXVgp3nSuc
6xZYJT12fNFmvJcPSERpA6MZb8P2jNA9iOv2dXSEfLHQ0F3+wsw3APBy3kmm7w7VH3uEB8p+KYUo
xpAsknqkTszmh/3UUilgB4YwzOMHSwgHK3gfMTNrESVRnsHZUcovEEJLUQZUyYvr1FOG7SrKlCwf
qIjm6gUjgAdkFfaFHcMeaO31poj67NKw0zZZiehRGxUdmA+GCmI5Ipz2dfdtoW+RZzUpItGgMAvb
+mqunW1ige2wWCsjbFFtuAYhiRrNYAGKZ51xjKNlLkXwuMkXgw/Vavm4Em6d0yf/ENU9UaDF8cSG
fDwn78ZJoXPZth7uTkV44b5oyevBfCh/6TiYsuYsU8Auf/BtkqGp3nCtIC8rKyoEzoLQU4cVzdzV
bOoYw8PIeeoUnMsFHF6Dz3Z3Dj+t++EmLeobOI46PV50C8Dlom/Zr8p6vkQqAno7SCCC1YzZ44jT
qr1UgaL8wr2jMQQ544ZctQHwLSzK21CaoX/vQ6JVSaR/hJgtigWr6454vMPMky93852MYD91lOvU
6Z7Git4q95if4P+RfKZekU8yVh/8wgkeiCOkk0QPcXN1NlzSrYpq1GfhAsoId4YNNZIwa4GWqQuS
HcLBiWJXmfvzl3dUbiE8oK8sGqw/DWF2xXQV4oNSwrYDFs5+Epp/w7sGRL5+hXaXzEUEsgCwiBa4
dzTHaeNhVXPIIDIqCJgqY5vDVS7CHYOpvPSPdUQW9Zqbv39K35JWNAftjxarAuDwevbXS6q26095
/iyyfA3fJ3XGf5OktLK/gFYg+renQK8l4knbw56WejTi436FWGBqNHUki8sII+Eit9J+cXg5GWpx
sdWFz/beL+kolD14fhsBB2fSB/4HW1eRAKOWcp1o8O938lFCkqJaoPGz7XcZnTRAzLMivcZifhPF
vi0Ggtv0NeNIqLcVB2B053dyr/j3HYp7xKWjjl4xx6Kz5x0iX+JTwe0BXlChyFEvtcZeR173/w5X
T3ePrMtG4naCVswSRR2jPiBSBpZKT6kAVaTl7F26T+xU45haRuj5J0t/43KnJ/p5pFxhKgp7ZP7m
GreFDYdYEphEvXLeITpKrPlQcf3gwfnbJIaDGf1wKzPFQZiw4/B1x9I50r3KEhL92cS0BnbF81Do
Fp17KFFHDkIRPVsGQeScnhkTY+wXPW6tawmLfdXB1+/1N+k/e69bw6oAS0MrvB3dc6kFeaF4ud9x
zdnFxoEkpx5xfPHZB/P22MOzt586MGN84UTag3nK6qT3EH1GcmTykxEQ/5PRtkxtQrrPWO9gO4UA
BM29tIZKH6OPydtjNMPMuaDcARewA7HaVuNGL95yZLkcamG5rcKZZtbQyUHBC50nDAo7C54pAqRZ
zzoRTdLbdRPcnrJwOW8B1MibLWr7MH3LDMqgaCaQX48jL9hdrNOKhqSBECe1a9WaqrjbJNz36yEw
ZX+uOk2rUNump/luKSlH70lwH/22Tdy9FfxiMPyisWugXCKUkgrBkQAYCnbR2IT6kbxqa8bm/KME
gkcoss4OR/EL7TQemHIknh93ZYc++n2hfqOtMRn501dws1OxUPVTwINXw3TosTP3fzI3WonGmHm4
ckOYrDIwzc4K2U24QpzpguAfb3wrQ3LgQcy9VOO668NxVUOI8X2vkygSKcvPGcdyop9RPFvgX9GH
R8yvMuNfrgEzYMmyucuUT4J1WmrbNl/+i2m6w9QUGoGLdoQSxGOTZNumTa/LwKgDZLLM51/ee3OF
wtuTGcj38kBxi30oEeDTtmSdulE2HMCWYAlF3lF0HarxlwT6cZ4xSo9vXj//hwkUuBAzDnSu43HK
aXddlkmStz4TjsKWfG9G2yVEe0VgsOpjAEFZH19A8Y8jX3BqZJ6VePeSUHvyB6q9ec5OpO9NCpz1
hfss50tvag7GgWAQr+J8vHd6/GYoy93eKJCHmD7/lX4ZQAW/1FGvahCToo19/+7BLDlyLX06W6mV
aYT9uS274KYjpbmy0SEOKFolhGltIJh3pLKTOvPltaaoHsRVJllaDiI8JmO3cTBLpNxhV8ZDVBrx
rJAOsrsmmC7RgZRpCUYRUCEE3Xb+UhiN1BCVEXnc/ac0rU03QpEWAw66HWdEAQqK8KWjCHMVNO0Y
UmpJgFSH1hdt4UQJpEcofJu1LvnvWVU+jbRDuu0nJPXI0Iv1pgn16HDGhXQ0sQnYad9QFOZWh9Kg
9RbDomOhuAujxxp8UfPdd8V9EjvWJZzH0QYp1NLH/zfdmCFrAbflhUNj6y6oJMQfuZ/GVkKjH1mA
ribbC8NYdqdApn+Nk7gLDiSJIKsXezXwF/9HnYr5VUrNOkKdqsiUJ7CCiV07bPaO3DoWmTEtWgbX
QE3rw8KplKlXQevWm41+xEGGngn4jPt5EJaAkR19BPF7u/WA1HBTR9SwqxMiC/hB4j5mVVrUTKc8
FQfKN3vuaDf8UAVt+TIMNNExb+CBQVviZoAYGch2Eoz3vM3tWlcfrpd4YmX1O44SSDENL9qJL3KW
9vnYh1BVXJKgDOf1D08f1vCa2/Cred2rl+FWdDveHaMhPw/zgytvvZsF9OoiWd/Me+Cve67/npzZ
Yl+ogx3gfDTeBAcOrQKB6n1ZBZDKQI33D1W0xNCvhxc2fKfQnww0nJaPAH+090jgLy+DhE3fMS3L
dE8ItPcqqvznxkOMNsCj9Am1HRjeU3GXXSpM6ur8vlF50XlAEFbwc/M/EOXo+auAhDIGeQRXM6/A
qRglgUeFyezsxeeyat6OHhBw7g/Bi9qnBQJGIxGMbbtvy0Wj3zc0sQf/m1QvZXVpYFN9zpc1U5Lx
Nng8QmKC58kQ7ZcQ6eAYL1ci5COFdw8aJjURfEKcz6VKgUDmFFYe2I4LPe9rUge+kh4E/tEH1D/A
6co1ZFH4Q4gvo2gfGLXgx9urMDbou/hrxRinaRTZ6ZT55zC+6GYM5+1U7bM5iyBr7/F9xx0ofn8w
Iey/F5hM9We3wj/rtBnQ9n9WPvrjTHWxcAIkm6sxnHqKc4XdG0WIj/FFpuPvWBp1MQxwgiGzAnlJ
ryzh2//NRSxHde2WrL8nSYS//Q8bY4EqHBDGBMWJ7n0PAA1Nbsl61PT5n0aIbWRHu5x+jVYlc5hH
j7v7qTNnmNzhgKX0bjWMMBQB/xi0Sug/nOzKpZRExa3+qnU1MEuCdP9H4CDByCZB3TtRmfQHsshl
e3OHG+9pa4rbAEL+H/TSjK/5jwQkKaO4OfUlMDN1tbKw49JO+jGWuLC5VEfGI/qd0fbhiurSYudM
btAUKoTfMzGPod5PNuiyalLetK9L6q5XLX9mhYvB6k4aWR56/pffetXSFHb1NbQB7IGREMBjL43p
NqJ+X7MHcLF5zob1rTt3HioTrw4uTxlvJhBFjAgGTJSu6c988SLOGGh7iKHijbyX9yh/m13JlU3s
9tmNbfaLxIX+l9Z8CCGVBc9dCBRSgYUAbtsxWuJUtPapIeNemN4Ax31UuuH0o5kJADRsc5BcHAjG
cw2+AD6u0x0rvK+o66wvgREHKBtXbZM094fkWYPKFpCWTfgqIVWxktJoThyGClJ4A63l2yM5+4nD
nq2y0aZo+6kCie0kYQSt70NTAzOkPkOCTp5ksGy6zYIdYmno/PGWNfazVbUCx5Z6aLqPUvGgA6aW
VGhLGj+HLPJGgJ7uClzB/xbnqvfzZERq6nW59IuP0tKO0E9ixU+i7yMKRbPYFwDAAkSbCDzbRmNl
9JLXuYaiXvRcJ15bEztRm6uNNixq72LrewvluUGgbAUnSfcKKutwnIuMXm8L8O6t9Au/jIkCqIRB
Z8whx6244lZvZSasWBJJP3GzQmZq/AueC5L4rYjhNSxfTMLWYfWuJoEw0NumesUV+dTeCBxQza/k
2uWDrmY7kDDaaJB9PavcKbEKU5b7b840p+7ZlJwj3sp416Lz9PLGnaynjYNRaaU+vOMz7BqRWfRU
tlloxeDiTPgnSZcmC66zQhAOk9A7CwXpD7tncM5zFWQn4SlHIfWoA47nBlh1HY5Q7H1eMGllFiyT
JUo+xDDiyLPlj71f7CjsTUjzMrO6e5OlNwxIo9ToqjTAy89hCbhDSn1NSVh4MPwPufQH+YKG8/dh
mnWWPIVO9m8P4wcWvUqXpP/CNqrQG7FPjLuj+kiCj/l2hW/V4qXvTXyPl827cLmu05n6PJV4/NIi
LzWglaX3H+xzpZFbM0eOE7y9+P/ps7nXlX6NuEmoW8zuYlgJBvmr7+9nZ/O93jZyDE3sp69CDwwJ
tqposNEa/VEU7JitI50HAdMYlFv+hD13uXvJIQheS7M+iMyy9c/fcAoRIvRf4VtmK7EPtHE6C6GL
gdiBaBpgoioOykbpmrA5RsFbAAIiuVyXOAJcye9PElJaEnoLF9QL2CHU6beantOdgUXYdyzszZEI
IWueqrdhZFyDQnjxc/f8fHky9j5Y8dAAEiGp45BMi5rZNlVlyiL7SNsuNDdF+j5oaMb6+4RgMQLS
7trY+HiIOg20nQHGnE44KsjtgZ7rGkKPsaGl3HZxXDhB/rS4dFsNQc3jiu+aE4anTQyhFQ7v4fI/
SF5oIl2F+K8Hf2N8M91PAemLzVUsqLFntHU5hF5xXYNWlz9LbTleVuWWjKIX+AJ76OvO6HtPzX00
eWC9W8TEW++Xgmmqm91mLT5B38J3Lpr1y7BI8tjOfyASDUB/AWFAYCTqpzPePwy+A+ERuGFsn6LZ
ZOy0HIYTY70FnAe82RGmhozqsZoNruYLJY53RmfprwU7KOp5COQx6mNlGIY0ASAvfIOQKHLU77FF
7KieH1MkUDtJs2gr9jcizIu0IG24k9KaCC7XV0WoBnPV/UMFDxKjSrPkNd9ECfvgi5R4gLgYz2Ml
XOzkWELBdT8EAWyg8PEXy2wN1j25YwHnOIowVx/MO9CjZ5N9dOFdgL6BUO+mAmvqGna/7c05JTMS
InoGXw2UiZk1/0LbpPFRdMKO+EfYJdQYQEzmOSAp4zNMuHgBAQfVIQTB9xfe/6q06VDmwmSPiCGD
gHoFsHZCLx5SIUHYE3II22FERkc9y90W/ClzDUTMi695BnzwjM8agcb0k4cR1SmO2CcQDPrQB0Wt
LOtXgWgXq+ryllb84OuF4QySoLChDWzyUtDNO1SoCd3qJPlRM9g3KT65H63V9zKzQmnzc7GO2S61
LSQ695g9vrv5WlOdAG8axde4nASrftl/2NHuIFcRJrGYVeSm3R1rDAO58hZ8oENC8BqWX2bG3Cxa
Ezogv1G3lz2hW4e+0ZleSRS4L1LXeIB9orq6Ncti9FtLDCW3Yk0i+C9xlBh1gdLGkIfVNq2RHgGP
DmC+6KhLT7y8kuoSD5d+Fg8jxknMZlRYPDSDfIMMS57zqdG4TDL8Wrb86zT060ixzRdUZ63IyIGE
dn3QITVErNkWwlZOtlX2J3+okJObXG42m9rvZsPWu78TEkFFsP+lPo/WFciBiGOzp4p4YiVSC9WN
VCX1rCBJqp0tHeKV1LbVWLg7psmDjFaymYX+gCA03VIqvZQhx89SoUmJoZnydqGRquNeXJqjdTIX
aVDgxXHCvy5Kk3QVY/S0t+wEojv7mzt/SVkmKJbxoDY0j1u8CXCb3GuJbL1SvXSkLvSktgsY/3CI
uxDtGncpcx6PjjdhdvVq20Sdbzn0DuX/C2lqrPSxEskQ9kcNNVeXIg3hTfQqN9492VTxJGmrxggb
aRfOsUugmmF+TJIabVRooQTo18iSVRQlssgQ6458hNf9LlDq24ZJnGi08gfbx9Myx9nFFVjE8yYR
Dl0xr1XnCyXTAzWIt99SltdeZbDdIM0zlY0Q8Y+IdoWtGspd8bZ+jHLf46xVhrUUqJhASBYavjLy
rayzsSOU8hq91MMAiZIiWc8IErxTcIeaX12bLAjYcuEwit+vch4hANlOajRf0DQrFHz8XYXfkjVL
GhC+kwinZDAk5WlbWrmbR3UXmb8cQekR0C73GDwUsvcBIZelpmohA2m5YkIryrRfoYOw9RuTpG/g
lx4iRQMhL8baFgFh95OABydnoKxCZ2PEdRouIbrVHNHC/xZD5yNnazG3wmwJ5MLdGOukm1QyCPa8
dbbBc1g+gmC272HxNrMjQNeIX7jNFhFRGFlRME3367BPCcLGzZ54O3opXeLH2JMjltsVIXp6ryjl
qbApWxAiqHK+6rqUY5oMUt4oi/73MxHypzOyj65pTjTcYDTonBBmAyFZov0ZVcl4nNFAjEqwEY9S
QGYT0FRjVMdp911HQuPV8/0kxKCDJ2cdmcpIrvnK+sbS99Ybln0gIcznZD2R8O4yvA92rIrnM0O5
LhRBbR70VkQg5JiOqBnjVpQTMMs+hPKtIutze0/rH8LqpKnyy9ID5xyb/P2SMD+HJfUYm18gAu6J
0NhBI6x13WtZ+7MF6KPntEp3ZKtcBPArp0tgXnZsYihhhmGqhr8CvOq+jvgucGxmxSKGuiyDK8VO
5AnoBLt8Xp3UVcLcgzQWEIe/xi5MVqGLWClk05PMSRSAfKGtVNb7wIiAw2+mJXR6YKW2/4V4HII9
6+BjwJdPkK6CzqUFGJM1k9kki1B9Jye5CvnPclJ9U09l2S78H5b58u5wfeilmlkRwMnuqKMAx62m
zPCDOkL5N9joLV0o8PAZ9tdCe9eJoc4Sxm97sNSdpVY+lQt/JhyhpOnOWsFbwUbv4Ya1fZFyoCn2
JWRcdoquOGK5sUGjFZKVtAp2jmqicnzYsO4qSYUHcUJC3TGvjUEV5OsPJfYaRJt5N55fOgMfLasl
b30GYnUJarYTJZYCQ9cm7pxDCwXMI/CsTsKd9B4w2dxS5tszA+m8+bH7ekRqjr1cUrRp90aAl9pz
YmbLuCP27Ca9fEXY3+DkqMTRdd0l+QTBGQj5DdaXNXa2jIy8s76xBDj1tk8Mn8mj3zwbB96Hxacu
CeON3LK3z1CtJ+CRTXLwPYKAUyrXn35h+EdTHkypEPKx8w7IlBhld4pQmu2raHoLNHAC0QYJFSx8
dXPU2hPP3ZcJCEktzEC6V735szOGvsgoHW+EPs72KJ1JXC8ynGGzPqB0drlhb2fLo2yuDj7E3IvW
iQja+OB50iyjLtQKCcDfKJziTWY5DFjdtd+3J7pp35wpYzN/KWkwSYyvMI4otRNomi+EWktZ4I3/
mC7Fp2QcLfVmfslflSLvLlrw022mySg59haohUe3HC+ybc4KkbAxI3jRIRO/mtJVVreLG0YbsXOK
wtYB742zoqLbr2eAwOo/qdqG4aWjycjKrsA4aeWQaGP5In2RPseDuwQa/bg9xjgH+0x1f4NS1/ih
g8Z2MLlfPUL7VnZz/1HAvgyY09pEMeZutm5JE06vXixy21hEYMZCpm+8393uvktPRrx2RvxcTax8
p0BgdLBHXeSYJpaNH/fsOlogGt4VpOcGtj8uGQztUAszLZs9KrT7v8zEbSNKcLgZYoa4jEFHWZ/8
xosgCsqmlpIN+A5EXKNVRh0ygksIWdE6ibA/jLe0CvVItwTfwCf5PzuWY+Hq0RFZQtjP9/jKiOMC
HRtaxMy8TrqDvXifG/kZnrJJRvykKdN63G3KhcTQ363PuqHs8TXjgBnAhKyr6UieVVkRABO01duD
SDylNU7/jbTfOHITLEI5kVxp51WSidftg8Tz4vaWER+2m3kR+l61kohYye3kkJ03XE87+yPxgrgg
FAfYoC6oyjM+MAo5ZzoAb8sh45PaRC7jB1jqH71FvNL5QBnxEu+DBwtPN9NisDtpVgd9wYUWvDMk
hP52gMOdViwg4AINeqiW9zrjipakS3+tU32bvpS0G3oKXPGawccoArjAQpF7Qty/y+7y88dahbbE
hWV9obwANgoCNWZA/B4sQNwhGTuwOjhcQAV/GR1oKlpTu/RALhq59h/2qcRLAyLBRXbclR85EgeX
qduxjmxcxScJ90qNMUZ3TReuixnyZ8q1zOcpGpREN4h/EQJfCYZVId78iz+OWW9Hv/dw+74bAKF7
pDj9xMecRDJy/PvUHBJyu8NScrybPg93zeNBP2L3SqoeFc0nNAG00O9z9gVgRuTY8D61VG3asihf
xgmBiwTcg3FC3cK0ZOVi4WK8qUStuePOReeCutuJ8eTiQZrZAtojETzKqMlOhWVGmQfG/5zTH28X
sJUfxMi1Ptie2mVq9BtQXRXntap3HK8HOhsMK5HuCi3rJ9HbG7driU2MHq9uQKW+F95HxrFzX545
fMfYprIChg3PQYHvYMLyoFrnrq2anE18KtZgzgNveS3r1eXDrq5SqomkBDpHlPq5GSu5If6JL0ys
lRHmyVFj4NZBmi7iPY3gDs0O7nGWt3nnAIRMSbKT/yRvnoake3bet6/0rwUNONK+jNuAATn9VPoY
n5SL0qdRCPZ7QvPSSvRuCN+qFPfa0xxTuXrpFuQaOEtFz6HHEAwuUwRpfGuiXYB1rDfE9pToh9BS
/DVK6HnxzpOVhk0NIlmlJaQVhS6OksNcrkmUMvdU1BsPOxHkrlHJ5ibzNWzwNCM0GGpLbwioUUF/
n94gh9TiMXZ56cYAu3L3G+zOPaWA0tjdjXrFpuE+pbhPLq3FbpFuGdvykgnSnwylAbuR5zqsKr7s
QHs8FZ5FmTOm/rOPqjowhsVMVK78D02jG8b4ZXHtz4NvLHPiOTdc+1pVLhHM1lLIg5WINfv18Pto
2TLCSOIVguYSQM+LI8UTGNaMv7nauJf2Neq4Ec20dNrQ+5Ryo+NekRYukRnEdywNHmVDEjEQEAWh
Mdd/j8tbbztjBcwipB6efe7Flpmm+/UUhph4ulzSCRpWoDTZ2whz5THmAsFTKM0YJbjIPRCWqRdF
ar/sehvNTnLR6Ybzf03YjQqrvsgWB3caA5Xt3cQzD8eOEChxiePEuDpZZW19A+2sMKDrRijSG2gT
2/9cAwbmvDGIomqJlDZ3Sjz0jtTTfknmOrJ8XGuWuXqAMM+fzfNA/0PokS2+X2ZaNheSPIzTPkb+
GAO5V+dFbaOB6WBklS7x+UNHAoSi00vIr+9K/X+i2dw6l1lW+fVt9B57duwzy8Fu96trmzjnahWt
kz54xfQ/8zUsZexblYztLDH8stHoTeeCQSZpNK4x98vz8mQ8rCXw4yXCPSixU/QxFESHO3PiXmKk
SjOdFYAwYt7AVRipFW32N1C8i2EPbO/NopLa5rikYaa2mooYzG1DzsD9AsQ9syGFo0nimdRFSKly
1maDWdHpLK+xuT+d/DYk3Qy/QrtVkmWTM3AceAjPv5gvAU3OiP218PVjfJQGeD5oJio5+XHXyUwS
iFGLIy17luQu97/uk4Pj0pVNoWFJlhiCKImTUBPa9SK79tIuGU6HRWTC8Um6VFJW41YKLJGPu4Hw
LfIss2PvRWQ1TVD35jH9ClJ54SjAJkVUsoalCXGo2x5cpg/ofzCoROB1f261KcFvP8thGIc3hpQj
Xjnw0DwAzE75gxYrSbuXC1ZA0arUEjZQFxyeLxF66rPmzJdeV0L3MVXEWa5bioS50QACCb9nvoEP
Cqv5aCVP3HSMGD+VY7nhrlX9ess73YcS/KHl1/4RbWLXoXoChDxI42vsDVbn/BV5uQekvD66crmY
Xey5ydlLaAGAfBqIB0nzpfomRFz9DPDTP8oG1Ll5H5r37lFyagNDTwFyXqqFTkqpznZoz7JXXKp7
h2dmf9RhWTWs/jx5+sOF/F2OrbLRC6R+AmD+rUwheo04kXrvbp0ZrmtPrYdmAAKU4t2gFH3v55hB
/9L2R7nT9ufD5alYoxFKFn8RpFoLpDHUNASKIF8xHozVmExVaEW/dzi/yyv7gWBmC1VNtD/fTXIL
jWEggQCR7c5ecHgYiA3rmjv+eli+1WfbZccqMw3bv1SfVxBzEPKvy5ONmCvL5OjanioLcKdXurWY
uOSHNK2y4/YNoji2rknKhjtX97xSr4BGY24+ycJf9DUh1GCOZ9zB75MPDMA9kU4uZLVZY8a/2t6f
neAm9sfhQntBm9Xs3DDOgJ3+6n51haWdVBOGRcMoTyde7KUyKH3Vgem8q8HKVvif83ovIykIXhIq
c6ygjVhRYG7qg+WeDOqMqS7Jq4zNf0TbkejKl1cvlLKcXglTLswUqkwBiqMMjsPCAcPYVPxhVZBp
zCzBFThqGHXP4tixY2Qf1/CrtP+9U1Ia+LUUnGhbwuRGugVKcXRvslxfEwjVKPjwWitVpmd3/5jV
gVBDf4UPZECIe+NiM/1xcwqo71hKzcbTupy0XhSwFB/IReKNY8Guq9raG2Byt/tJfaS6wQ5KX29o
4ERVAhCrd+WuvbG4RcGXiwHD3ClzrFlkh9NsB/yoTReAQQ4FqB8Pw4ZEpvAoqA4THIPt26/rnTAb
G9Bx0mkFNlHC83lnXZS+JakwSmj4WPS0Hjdvx7kEwdg6weqJdUGgc+VfBczrjMWevb2T3wtjfymb
WGFC3y4CYmFHzjf222bz3ooa5MQuTDVXV3x6UOO5gjbh/yF9cXIMRZpwtk/IoZLF8cMClpbfoIGd
OixkS5YKR0PhviiImWTSpFWousr1c+0TXvo0xt78x5nkEsbaJTWrjHD0bMa+kxM01dO+0PyugNHy
P2nWa4GMRGNeUMuAvCK35sW8It++rvOr1LXLKOk11IVXeq7jXE0L1hAf5Tmuke2iI3Y7R0aAPB6/
kvV00eexa7zzMFcjI9wR1UPX490ajC1L8fGiPivVD5sUy0BZsGfjaxxI/zJKlNaCe3gX0RG2fdlW
Ua/+s6cs+hViadbqd1B/t/sq3rtmt+/r3EanlbiywiWzPO7DYiGhMerhZAcq0o+f61/ZATJTwgsv
avKiFO0oJ77vXcvEKDUBSWJw8joTbNxyu8zFOXkZ/2S9l2uh1q1FhzHCFpy12rOiNYIh++QJWfTn
zeSBkin02U/2bIny+pUwLPZepKJDTiUaPWTBDQ4drLpClkwq5By2SNs785eFpPN2nkBLJxatE1fh
6w67IhXOGOL5BqeldS5+eI1qYi5cC4zN8oBZ4nTApJIX5nFZVCM/FVBVFCtuPYPFEJwCWTU3CFHS
QuiLMd5xi+KuOBKcrkkrDPYWxIbhFgg4Qn1PsTfPq7q4i7RmjTHju5696S6mMocNWZhlqN15sENe
cN7PolAVMCX/i4vKZZBUQPJmgHIwj9DACq94iGJj4B1VQfV3WRdy5Bi0AvZFEKkJO4eh+ewFl2hq
eZvv88IAxq2iRFZcC/C+fNXV7PKc2NbSq0sva6Hnt6aw8TY970yvUTPamUC4TjoMHQXXlLkIU4M+
2V4NxHa0KPtMke+vRjeBiCxssSIl8JRcSyrk4EfIl/aPBPVo4hxf45ihlf8cBM6nqazDL1Ve/PrR
Gy7kkrg9MD1E1PHUQ3g12PBeu2Vgq+e1J3qov7c4cHazs8ZWeVCyijz0Pokxe/AG/46+ttuJkG4v
NyezP7T8Of9E1MYS114ZE3IIyyANiFzbvhCUxOz0ivfyY3vFSB7vVgEQFxQKLUDeU99A7tEfp0P2
hR9SWjb3c2KJrzTE+DTNGXfLX+kBzaLCoBTAu8WkFCPEPRepg110Gg9ro+gKeA10I4zGD2sgrLWT
DtlLER7E4UYkggGqLzE+FeL7QH/HsoOAwZlT/5edu4Mtgqdx8N7boHy46TbXJjnJE++p1CWGmC36
5AnpZSTuWJdo+IAsiDLeeGUry6QneHlg9+/F+Ka5SBak9inLyL3QGH7cPZnDHWL7IMRepMSONrHy
gMw1qysY0+P5Rns97eGRxFudZJvHZMQVL90KQza2Jn9MfkHUseEIwy4x+YBBtHhXILvC0DlA8igu
s6RWhnNoSWzk6Nokp/Yi1//eHKInr5tSM9ljylAiEmWbFZpechmURh2IBjwfubQBxIlxQMixUoR2
UVElwgx9RtrUEksGBSaGBAK+Q8rilWKJiV+D4PHthXxbQyNhGIX3Avv80cdIQafFVpGW3Olb0QXt
uyDJZ6AHizqw4KjYaO5cWfPBX4ZH0y3AeiCgOp7obQd/w3RcwYW+BohIyzdHrl6gtSDunqCl3ekf
eteXWkCEW1yGZDTwQtJgO1hmqFpTzFI9vcYU3o41SMCBFMAfPdx/+1zwKzGXSN9+bjJia8MuPtil
sxbPnoDrb0394cAHpL57Nx/fK0oPnlc8DfmDQljNbmozD9hi/Wki4M3iwLgLS+Gr6DI58XCZ8fR+
Tc5V53xzOTo2UXgaKZLe+FGI5VEO1L2FdOAKbtL22iKOlH3h6iDZ8qiQMuZOQciUbwrnLP87Tq/A
eioiZcVyRrueOiZXgRJclNq/gtnFWH8v0GsXPEpDCaPrv5P54gQw5IlWwOqd2BUB28Ytvj/ltiQm
8JzzZPPlOyvEAn0+BbiJu7Tnx5E8wtJl21A5mV9Rw/fOmPyU5dnjpDf0jWQLLXMRiJBP7u73gNog
zuRc5Gn2ZZ7XMOmDMGLGpfpR340SVbHQdzq9jtIwOFvdN/c7VIU4QoEk82yCG/1L03tVonhM3fa7
kRbG1m0THl1Xq+twoqbgtRV4xkrE4mBg1LU9GTb8RX0VImdJU//UUidJSI7tQTd7ek5hYJwNjSrz
rwSvjruv6czPvhLgBcR2UqA/HTsysVDP5PUC5+ri2w1XlUhwNq/JbcANAcowWLedLbsaEm6A8x4r
/LicXWS9mIqtTAhEIf+JzXpCtN5LOd6f0fHsoSipMxMWGbrSK0G0+BPbdUBEk6F7ZZYW9sv4kvfY
rRRnLa8x7fX2SdKXszmZfzh7mZer/mGkSlfn/1zAfpT5SwjwgdmHuDcfKzETjtytRPSQgSok0Zod
dnDHYyotXXCmZm0hQyMI/zhXILQPhDtjnEX0NPKxdib0PUZHPTR6miZXmlZubEgTV70JHnLTTEjd
c5Pd93GI6DT3wibdenZValSf99gNDRYe/QAl7mNcKiQ9ghPbwIHU6XrLAC6hyCzuDcn5Cgk1j9NG
6fjPRS58eF1IdXZ1MRCfya53ReWXHP0jzUevjWoKXmhRXH1w5nYccv4+OCFlay+dSwvpTy5qDHyT
itCroR54iU195w5zrw0Ftf0wD7mFc0DYAy15bvHVqQizbDrbhyYR4lvHe1ec2P6gESMz/kRs0Hj9
/W9x2tUyJYjV3MovkFz5d/8SUmidVtmmBUAZXyJrJG4VCUBpMptAfa2Jpgckvv+y6LSL9suwVTWR
FxZGjWmaCK63KfZ7jLyPI3lqduAsFqiWCwUwenFhdWUZbSUIjTIiOAvk4mFLRYde0gedxVLHrFNX
OXpNXQjXZ5nFan1qxBfA19C4MwlKDuvrRG634Gmdkcek4LLGDLoO3PqHmqmKZXHDivCs/woo5Go0
nCbrBpAZhRbqK1zbSlsclFLh+mLPm7/qD3ivpNQujduSFcKaTzdRCPkUfDZlInJIlZwYsdY1ljVZ
gHUhkVV6ymaSlQ8836ocm+IMGeFQjg9AReEw/ohO9MZpYsKVjXVXNnhLpmknC/l1Torj+MSsx8mV
Rkko6APrqe+hoONDZya7zSl6gGGqKf+gbw2Qe5GdCrhDobteDNK2dZb5eU9n7cpgiNgE0WTlOpYg
Eb35A1ZcLb4MA4PddwUSkyHaiR4/T0W+PKAEdThozHbls/8hywqtS3V8O3srixKn9HMMopVI9cGk
qPSYrn1+M/ICqp54Su8EexpRpVWKiAD+maQtVnBGLl2Dh74H6anymJSiGjLGLA+6zfufq85xG2c+
Vf61StGHBAyIEb5my5yyN8NY9D/2GXj6R2jKCW0ODZL9DBDiYRpyLrOtDsH/GsUyKG5PzdppIg+g
KJWpm0wiQeCbuTRetzMkzEfpJCtQo8SCsRHw44iBysg9lLtET/aK/pQ8fcK6LYZByxwyemZYQPVv
1MQl6jypmRMD2VJITuQ1rlyLCNW+wUjlR3siXd5n8vZjbKkilCk7w/9yoEI6hq7nBYp+7byZvuQv
HircPuUcVfRgtLAfGVaCILIffCfLiHYGBe5Y5lMdT6FFuEw01SmFNV7TXhm7n2wrVovhd0Q0xwyy
AMLXNkAPtoz1HcP0onbRh74HUzukbR03Yo1lCUxcenjDOAQzF5RPzcE930g8byt7xTHSvBKrMNsz
d/9D/11stbqei8Sw3Jib4gj6BOVoS39RPV0yPLYHaYTdNVmP+mmdv6NOZv1e5q6IBOr8pDymNi5y
HiFBNQe/YE8phKoto757tmYYwNYo/AP35bmKrYMaFts/f83l/qOicVMAJgKKk9H2v95n99TxfusW
hgH3sjQ7qu1P04no48OayDBUmjdvOBQoNAUXJulLpqsdIFnogd2QTHe7F/n6ub1xFg8x7R+bWslU
mbsLzxA85DDhClZrvkr0+E86INzzkmoItly9yDvYJige99GMRkpTfyRRfuvOmJsBVbcNwnOw862A
SkstPf1P/hI5cret038uoIouulfdsOTnBHExbbB0tYAUXLZYr6QInCg2PV0M53SvgL89cwlHPLzQ
T3v1+RQY3XBlpEqBLzxy/QbOB0Tv15JyM4FzEbMwM+PbK1GeksPbTTyhhTh03NA/PLUC4KWWJzuG
S16+SQ6DdftFYQ3yNxjZp6aqqxLTrfMW60SJamowEC9EXaj1V5hvX86kDhC8oKKtZc4+bmE376UE
OctAiXjo2asK5bWb8tgIjoWB64pam9c1UYaN4euSpgjQjWbN++bzkuyj8PBIXJAaWJKeC6BM85Bv
mGmPAE5lArsAo07qj5zd2sRmoA0ZDS2kKPE6LbRxNn+t7hXfuGyvMc+erW4BY2Dpnr8q4zyUCIQD
EomN8VyF0Yf9OmgmsJfntJMXpp37/DzQLZHrkPu/A0oG0bC/QYnaJa76/ZXM3XfqqSbUFGgR0rLA
Hp3y9KlLCj5prH1XQbq8+YopEpGsaIRnNaeuys5x33SQ8YkaRKUoGTBzJNcRtOVksDA5c3ql085Y
zT3YLe99wu1ptQHo6VdAvc1dKkuH0c6pHLCcXk7RevUUcf291dmdbleQFLwbOdJ0QQFePH3S1FHQ
NjaQn1pjAsndtSbT3IBbnIal4OYKkkKZ0sLZqy1Xia73gQN6qelPuE+dBJIvkXSzdm7m7JNJnI0m
YLj9n5ey+MWVkjIivHf0vfCFNcqRYS0wR2Hz0X1VuMP4ji7hTX4vH0eI9nr/7XMfOvql0ruowppI
aoz3yUnWe+4mYrRL0G0Y2TSIHusiiXlAM/kHGtyg1C3RiNnR/Gg940XVGCzDxSLmvxrbStXR+5n7
eyZtXz+ZAPGyxmMsKc7p4K7ZDKjJKYqhvPn6Plnp5ftLR22eZY9fcFlM75P1aoiDh7zFd7/q3g8A
Tr1uXfjK3oOgcqmmLSDhDKHSa0ig7s62lGje0n6syApIfDQwEayUeaiaBUY1kHKMWxV3RGIxLeuo
PGZEzpStpDWe8povVbcguyLN9Ugd3syWF4lcQOmDRMOCYMrtdDQkM8jLKmlfQbqLSfXw6q5sB+dM
rrSzgj022WIMXyQpqdACnCU3nvXqGx6LIPy3FOb6/9WAaiUpCpMKYvnAk82F9rOChj9qt/6mEb6e
XaAQQNdxI/HFw2pPMYatAf52QqInz3F+z74d6q6TvTYJ//kFe24hz+xRati1qIaTdg1yUWAJxFDK
0KSK4mOyCcsQL3uts4DWMmtWt0QoSTnvr86qJorF3jeSbR3aV/STK0lbbTt1aWXIsZzQnX5a82e1
tOXK7e6bMiEC/QcIvJ2MOA9ev1rNZQXE/eeiEDIdIV+iVZpbHn6S1NV39GkAL5ZAVd2jAZIa5ZAi
i0mu8oIf1Qd4DtQxjeGgvMqEMRSKMVmg2OEOSHoAzxrl9IefVQsIK7VNPIvHAyWQfysAKuG2PPlv
JJ+ZgGsUmRbHoHK0i+SlTHk9xrOBud+IBebF5M+wNMN9Bd3bcHKXEUIUa3WgZapARPh3kK8gO4W4
ncNk89kFa4tMZpZX8Y3PcemHho10qrVkdryxfo7wA9XHNadlNtMMDECStE3zwQRaDBwYaQmDexsP
bE3WqMMUKbgiUqKMg8ndPGwRyHgkqlOJlu+67JRqJffSH330dHx3gb1xitooO6uDlXBSigoQ8DG9
sfGck/eySDVOge+buxomeSQ93oHVzkWDJFtoLFGsMRmHAZY0fnw+eJ53f+f3ZQErCDeOnbh9SNXq
hKBB6AutGaGSazD4e5FwSGF2vgIHsoyJZQxuMFqULFjURX7XW8kJ8IKkm0/r1VDMHqCGu44QJo2y
qaIeGLjhHF4bBsdkgR4hwyu7+WzPr46L372jGqT01L+WUFMckxq8vyGCtHbAZKOamerOeeCReUBe
jpAt5FXEA8BDfMozjBc2xtmKWOwbXuaH4IY6g5kCkdEKVbPi+h2/mP49O+EB2oRKVA/yZRt1ACRA
Z6in5VtCm6VMmxqNkQwt0A1NKysDMU/fAjiWmeNkqAVEaLi9RK262nk2HScpl+GpGIub/oRyrNo2
rROOGABA6sX1MGJxVAnPSEQclWR7MoDrhxa7S50iqkYRgNbE8olLHpifXegY+MAOgSFiuxjqYLH8
JNjMxwGGeNp/1JYpkgWe34cptDpnr4QjbbB/9KTpiyQGBek+hG155pMnHkGJ/DlpdRYMrwTx14Gr
92tJ7lHqTdK9HBluCjmF5Invqm8z466wN7QXen9Ce4TO3KXqb3S8K2jYYbTDRCviLE69ns7IMz7W
4PWTkTY0DteipBfX+7/yraVQLjIDczhAbJtI9jMrlasgeopdU+p2fh0+8x1ds1Co7hpkSVWVRdy7
hL4cw5sBmD2/kcXz3fevhY5A6+GAG25uetWckl6H1piWQml7s4tKePw4FGZCx/3U+YXOXG8kayHB
0TVbpPD+g0kiLmaH7VOumMeBp6BtudG1BgU4XV5ahWwFGE1kZVFVcKOG312MnBlcVi/1087cetgF
80r01N27IcgPY4nhY2g6jXrlxgiA/QtU9BDZbvqBGwCVbDINYCC4PJTYCULgsHaNXMoJnDUPrqG6
+0ZD7IdVT2wmvUr/gEgnvQw0JXcktvOsolreQCFJRVMZ0/4lwHrTIcF4+ni1CB6Zawyp4/lMrTtr
t+K/2HlARaACpiN19CdMcIjSrWJuCr2Lr6la8ZsL/tqNg6Ces8jru7LU2D79EO8CAiuEwSSpRjFr
hAu+gciZ7UgVMS0HatXa/qc+vCbEeWoCyGB3KMWYdcFAhOJtP8KX4uk01k7Mhz0pi0QYpcKxjvIr
ENQ4uoJ+X/FU7SwDKXqvOngEzMTyEpyWs8STWG5JhDHTFhinERlbciMlYPUIU47VziDqCO+UtBA/
mU1oT/nWjqplAqS1M5UvKzydaxJH558y2UPgZNwGbXXPZcGy+DlweiLVF96AFoK37/vGijjApPPK
3XCNSjkmh13/H7l2mqf8qWsp1nSBybBrgBOGI+8tIGmFMDhwI557VzDEAeQQSkkCBqSw/03LzwQG
91vShh+v0lDXkbDP3WLGt67fXtjznaB+xhC2EKqH5kcRPsCM1CAZWwor12iUclJn+8vFANxWNHei
wP0uJUlGG5b+qyqQQvRWVCBY95BT3F7A1pZskPfHQuZcd/QpSoxK0LKNtjbmt+P3WlZxyWVaTI33
jovCsknweZY7psyRGWyKyWnMfANHOhsSpPzvnIzZUBtQXr7D/5KNkkqXwXzvWLs15OREUFzStojH
gO9Ul7o+RLN9SyYNRaE7sPDl3elKy//+8FEqyu5rBoZB1F3xBbtZLhWcpZBy/2zuWu905lcBVpSZ
RXfm6DMoGB090MyY1wM6k9y1RFwLO5R7fdQwPlqy7WbDyhWVATkWsXHenuKQA7krFgGcETX5yWeK
tH5+ghjKof3AAqIkk9OxW4xztUKtkRs2/X2ItS/VB92kTm1TN4fzwSDOQ7B0UBoOtKI1WIdtN9CM
Q5+jFO3wbUd8yPF5F+mzxGpQt6PQEGbawGeOFJUty7crOBEjCdUYEc4TZLJF94o4gCGr1w1VAXGi
IpJ6WggjOkESaTL+2oj30jorB249PFGexESOoZ07ToPU3FNeyGMiXkuCLjoUFk0O9pqM2sGNOnLH
vGLUIhCD9EmZ/r4Cux95WKChzBo4UnpY4UPtp0k1QNuC42ym2sz8F86yKt+mBts0ut6gMLjVRnrX
svbL/e8QwzaiayWTRJ+wAiUTJNxm+H4Dg3ZO/mEbBQI52aRD/wONntwEs4GaybuEmi4c77nks1dc
fKOA/qehlEfSF5aqfAqVtuvA4r7L4OevrDZTVrvWZFxgWsBJsD7MUsEtZUIf2oW2QY0LIXvfaICF
0qDUKYAeL+4n3Qfws15ejag=
`protect end_protected
