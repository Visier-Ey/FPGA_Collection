-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "N-2017.12-SP2-4 -- Oct 23, 2018"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
p/Tt47557O4cJu9BFLAhHTj7O0ef3ElixuvWmyrZwyboXijJj4aYStjIEO9dIzkH
VuS+a5l9+GI4oFwu6hmi5X6dyfoAGP1PBRjlKssyLPSc+ORr9iUDQ81PLzE8SSXL
xTptCG7SF+bMognWRoPqmONiIEp0TuhEHhskakWzRVI=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 24112)
`protect data_block
3NN1zrOUrOUUoEcVSNtfPuLF0BN7FCa/55NCsfaszFep+lSfvv30K+4PZwfc/ehd
KFMpfwHHgq7zewUqmqOxsmhuJgVNEiVJIniQe14Jz443Z92kjfErsmelD8UMHNce
IZd5Ds/qTbiIwH+TXc/2h924nVqWy+lG/G8tOmk2ZVJlTvGuWVz/liuTOreXcnt5
AmEUwh0FGJqnYmFzQ38enlzS8DPqBj1iiZFrXA63cuzazDGkiD9ho+bTwqoigIpR
ZCQRanjy3skLxgdxb9BqCk0hYG1+tH/Wd6RHEuTKREqPcmnbpiV7WaiThSI+YYM7
ayN8EcuwG/+eSeYBYE/TPU/aGWT/GufJ+gMBlNLBQ85Gb4JrAa9ZLl70I4Hnh+/f
CrJtSRLSUcY4WnGOBzadvJk8W1dHwXIHbkATHzCbjQl95GEHLZmmErSBC61s8d1J
jl/zjcylL43mC9an+33JVatJx1fphZDAHYKMoenzEXXpL/RhprMvcOyA+iD9PRY5
PqrtuYlnk1P/Kf+W4wMsbsC8piL08cabnDMPDiqnVaJzgj2iO9KuJFC+T1QLlGha
PUVrFKgNLhmUXwLBtxjVuJEPKUlYKuwWE3iVPE080E1+UrHJ7u0GQiNY5Zi4xg8f
Cvey113ixao5v3IRQO7uWxEdvluqMPZsVmx2EhVxUfKS+yex2+HHbgMQNWEHzdOl
mgy0bBF++h292h2MbLCUUVo1eLcZbPMZU6c3q4yZ2f8ZCRIFlhH6TTOt5Mv61QsZ
BaNN0sDlVeL4BQaGsv1je9LGNoM1RpVS90L1BScy+iNVEO/w5oq1S2uHaAY1Xaha
6FnfO9u0UXy2fsPcIWOctKJnJ6yWhkra7jUTUEdr+YROOpkKrh2LAbx1ecOqptl5
KP24o4Ao/eoxcmQ9aC1dsSEqOe+K1ydr/wir7AhJCWuVl2+/d9fMY2z3eXdkk/1C
hDBb3zeDHoVIRGoJOzqj6AAXx3s5phmXokSI+yMyFsawTO4AurvqTiyrQa1DN6eL
HVuxO7SnbqvS1Vbe21pLAF+zF7s6Z4k4hmyeUYgGapFVCJ21IZYNqq55NxM+nBNO
QGnbnezJjBtPHqQCjEIDJttLktBN+5p6miJOtKip8ZcnmIdEpARgzRylk5fVMDhK
82DH5PDf8hEq8h7+MShXjL9yHr5oL/GrPu462ZQGZRVrtYc6dRrZt4kcYgMK0n8Z
45B+GSgxO2xhHQtxRqBpNrqpy8jqD0WvnyiNwMn0eCZjzF0u6tJgG0ITU4/iUNEF
C3Z0PBF2ZEmEf7WPPscLqBYdAWWeBkYzh3azrFtvZuPAVeAeQ5ZwmW9mU2TCMylX
/+6h6Mr7cu5Zy8UN5icN5WqQnK99V+BicFPCGGjlGUHg/puMfNIZFyjh+/Ekv4SB
gSBT8iEUxTHbpljGQWzsAmxE9eO9pTm5x9E28HCtmhRNY6JuBACamLIL8hwVeGcu
04F8PlLRAUS/R5noMAkRIBqURO9DvJz2Jz3GT6NX7kRu7zm4u7+n7K06Jz03nH6N
GGAoMnFzwb+jVTKFu6617HEkWqsYQ6BJ1bqMBFMBJBQjgyPQvgL9o9kFkdWV1IxU
voyiHAuYTdS2kD3Rex9VHueQcn+0cVS1WhPsbVufIFtXdwu5V0ZFAGYA99oXuEn0
RCp9/Ei//reh6gw5KIIhMWeATc9rLzImY7nBvjrBcBnQ3H0BpNB3daWAutG2SC1u
Tocb/Eb9ppM/Uwj179qK2jNh1BnGtYXlBOBuTKjrIxUhPOSKA7UoloIUoGq3wgmB
T4fWih+eVT2sWfkCsFkaa7EHDDsBMOQg5TEujFPkWh403jeHFGKfJml51Ln0nVff
fzoc+6vzPzkhTWFekAjN7531aOEtOGb+0oVuNxNkmTdCg8Y8/4hpp2JY5B/gJqhU
XV3tgs+BGWcf0dFmjNG5pfI52qBc4CkJj5m7zWMsHUvRxqk7PrTEMDv+Li/0YoMy
r2EGJQa1Dc4W8410Ke2h47/SBOM1KmC47UsSaa2M68F3JYvL2bUJgMTnGxlOWb1z
O/Te9bEI1cDz5ihW5Lcymu9hmxSJUhkUx1WrfAf88vUUD9BMohuJA8hVG0XsHRfH
PBSnQrB6EFPPdoEMd8E5xZRm+RBbvt/amujRPZ2FOnHbfMl5ByNe8tl9yI2CssMn
CiI80bjTlFXGh8wGQQb5oMmUkiIzNMoIlH8xRhpnIZo+nyabcQUrc4s1AWW17nFk
4J3evnMy79JkT25v2NxHuNmNR2B7f+tMrZ9M2zPwYbEeR/cdMcZFJuubtu1uz/ND
g4BEDoPCEu5m9CM0ZGyHEQyic3RaiQoTc9cwP0gHQxUTSrPJqgT5lbgEd879v+AK
hDmsxOsqT2ZORpeEarqlncnSTn12P4/wfBaChzP7xr89JWgDYhAeecnPpHcVplxW
dz/8ljRYA14YFwBJ9L7ZXKa9E8/SlMuEAONstAQhDAkbRGW3igokxT1B67SJRyqa
LA9nBAenCRuojt6r2PtIr85fWXXZpisFUPEbuLETi63q7cQL65Ho8kSO+fsE9LCO
ZzdQGW7pfjbgLRZSm5zEFe6QFkOWDbb+IOCvp/OmhkrmeugQF2TN9YdW+LzP9gLQ
5GUTJLAys6tjxj2gA5fCa2hG7eAMnunJhsq74rM/AN/kj0tUW8NBFnFqAnAFTZkO
WggiWxWareCdtTRRfcy8Z9heu+j/2AT12yxUkjr85yLVUnrNLfFzevXOLeV2FExb
W/VHHhYr/aFETC1Zq6Aux8dkuBpZWe7ax3ZzCNh50HmOcx2F06IFPR2k3upm6fSO
ehKtAxtXrDhTGYoJmmuJRj7q2J1SqXd5DSnguqFM5x1Yaf+sFXRr+CnlIIzfW2OO
5pT9bfiJ1KO0/SNOOFmQU/21EthkYXabd28SjAU2lTUShMp2DSh34Yorgvcoqw9B
Hi8hWx8jwqnNBDl1zbX/qtnvVMsI0V2h0vRrZQCp+agHtIAvnd/Fgn4c1IRRD/l4
AN4qXLju1c/EeYa++5QUBjD6/05vJ3XEAEue6CXRmx/BvSsNtfIRcYLEC/+WCU8P
DFC75/At1/09Pou7VjsXUQbeJ4HRh1s7ySK4K6dPtxwmjWiNDwo6co4v3cDj89G/
G5ysVBoPALIt3zBUm9Ol2+6RjaefsMYHbSI0p6p2vVcJAhBoBM5lYehMDyI/H4Q4
6zCExyA0JDRQJx7HVYvJF0wR5uiCF/LJpha1hOASJbf8WmRewWp0MjzFQTYqta/i
q44DxpBfm6Z9INL+N2v+Mak2ihq0LqKaFmYdVnUIa19RE9FNjZBRX+nuJ9ZRxNMm
1Dy9ZKO1okRDmlexPo5gOTyjhxGASzA5wevh/d5qEOfVTzz9deI5tyVhn0/F2ib+
jg53rlDp2iHPPjOWvhq/07ZGUgVmZGPJqEyE9LsulOJzGhzkL0OD/6lhGemTfwMq
OjWx2NpsuawehpfHqUPjrm99wYow40H/dqO1xPC9QWoY6Hl6oUrQuqiMQH0CLag8
fCSDozX8RFpN7Bw+N8WO3R7HTy/X+qYJA+UNv6C7GBdGKSOMruxNXEk5xTJBpVnk
o7lk4l6eL9VQStYFdzp3rrYX+OYM+R2KZ//LSY9P/VTmhwRPC8t70DzJCY1dgCvU
HtelExCYNbQXGWe/5G/uaAjgKqNe0acYgc3rpi51x9rqWa4ZM/VtyYczEwXAFsau
7giRbTMfCmBK9fpefAUQi3rehz2dzUwj7axR8KPeWaqzsYLYqpBLMFQd/Z33823l
Lg8h96Y+LrKxF9bOTxnT2JMZQOyEUVT3oIDb0HWzAHcGVlp246DgsGYmLJEi6hIK
EuLQgcWt0jM+vnt8sXaSGjHp1wLTajVTUykHzx1mBQCcVdqmR1eOZpScGohF5wzu
MtkrmqNYEF8iPsGcZtRkTvvF3/lcd1ZHXZH4WsekHUGF20JpKi5zgPJ/8odiB9/l
kYbIPOo4ZgWjIHS0AkeOVr3oHO8Y0+jQ+nOuP7YBp2LZR5Ektul/pPXA3tKDG+K9
KDpNnKE81LuUNOiw1xwJjWhU4Anjj75wXZ+Kb3/3+kSY0QySdKw83Jj6Bgd2Cy26
kqxHx+W26aOI9vyrAv3cfeaa/TEDLUixCUxU6wGA4axn2ftOxAfHIlbZxZElEGpV
yFZ0I0wvAi9JUMU4+k8blTrLhnDUTqeC7qKsUYduzLjrehX86r6hq0Uvi4dTwIMX
6pmUDLKdx2eiZa/277ZebfPTfgqPwsfOTk/ib49/xQe8xe9r3D26DO4zfUcUaQUc
DMxWf4Hl5mRlSGNlcU+QX1LEIoY5mB2kYyMyn89bU1Nbg/78AJWwfrp7dYFWNew8
8KlKAbpoXLhj++ToRfJOkMl6ER7MqJua32XXLtMbCMdyuJHqhvLapJ1PFWmSNFMB
zXLcfPRUNEDaH83E83FQgGvaY496NThj2D3aBVW86h8BN7SU9zkXmBxsMMkMGKYy
89bVhcpzS4qoCprrdGWI1Ml66/NHOAw1XcoZLbswOgQ0qnaNuBPbzYoLhOSJPDVy
sy1FyZG1lqOeMLh0ocU8Kd3VmMTL0N3f1TZIT74+JazpzmTQhHEuKwWpVWsSt/x1
NQhKoRlvi1Mvph3+kuAY9mjQ4lWPbk7nFBjz0vx7JnSXLrIjjle2UEaWaXE+j4ek
PRpGiM6GtF5A6RZcOEwqUMjKYrEkov5az1CXq4AfdwosGuk09YoHxKQgVzOEM40N
wJ177AXzmgeCCATvrpxmMIGsUg6pLS1uylnNtkPSo7LCMeQH+MhR2IZZVnsnJd5w
mAn4cgbgPfai89D1hT93xCoLC6ScmA6+f0JWsdMvPAWm54lFSGmhLAjTSXc0YecI
/AsSCM3PXPccDHmyFwTznSYV0xrO84RtH1l4ioQ4sMNMJWuP0HPxZRJNdaU3Oca0
5slvx3MootNrZ7KDNjooPfX+oij7OuIkabPdvija9keA6tDrCHiMRlxUEwbrdvqV
K63Cc4ggGd8iBpyzklBMP16aOKXWsTq2Mbx5zlGOKgWFtiHfY1pxw8WMKjJoIWGK
Upc6hl+xan3HIbf4OKY6Aagqi0nGQPLAayGR9lqtioEoZx6g8UgtUAI7FaWofAT+
WC7F18Oj6sXyzZNo4+Du6i6fHQZL4Nz5LR8cvP5I5xoiuvb3bPwfoe0VdscdiBmj
S2cPb4ScC2akbU8Ia+I0hNDy/o5dh7avBbqjuXwyODWW62pag9bgkeijbrTupwed
GxJetWrCj0OGiB+YxauQdIvF0ltsxzvaxeFWvOpW39SuTv/5jvlSrOlH2s79H5dE
whpes+HBlu2VbEIFMLHZmKwBjdJLjB3FovJZUp1sXlkraPTqAssfcZYqIoUXvv2/
1xWFuV4ROfIloPh/HyFImMEFOjU0eGLHxsOEyQ+fheVY8vrR1iPnO8faUZbOFbue
P2xF73Ce9Ce6kNmdqy1Mks1Z5Qjk/hnc2adYUOTxXcq3El7xYMrEQ56Zx7msGzzk
pqFE7eMgh4iHGCs/KdqIXOXni8MUiHLODfASalbuP8Uw1g4LiyfxiYQNAU6hXUqB
DraDAbpc/saUg0NXMVlxZMwhlPItCHxoaT7LYrimUoPaSPpxSlY3V4GncSgpd8Af
QAqf9/OOSRe/E3Tmizgf1OeaxGrQO0Jp/14d+cvsVL5rhOlHSbHP3k/0W2Zdv1Vm
MC+siSumUNqmELFA1CwJ+6n13uPFXLmphQ8bZ7IlTnQwhdCXtW3Md+2coJaQu3nG
kvWaMVoTnbVa6iCuhqx5elSaN2+1webK65XdZqjNUdCIpAo7EMjkwKx+QBF6/8C5
E8ZezgtYtWAlFyJRjEDI2e8HIKCnquohZJGzP8WUkujzCdyniVzpDCt9viq80KfG
MTw+H2YaCMTzeGFEnvzwiITtW14pNP+sTDaFwfuAar+raF9CnmZ+BtGaCvg3t/RR
DUe66fhqCZ0tWl5IH0JTtDtwPoDdsoSobF9SqrjU7oldYY6XiTDINWB6BKmvb/H6
D3D6dLuCA5cGfgymplrIlkATVj08aVPeC/bSRcpNHYbJHm94LOJ5vTjQ+iClLgrZ
0OARN4euLPEL89VjcUxuwr4lcuHgtr4oi9nTw12UMBCair5peSdLH/W8uhhEozZg
caic0XezvXVg/AEo4ENG5uvhUNEiPmnuDFwbaleCqNqsv1yz/5fu58CT2/siTVfS
ttYiPuNvMfHZFwnI53qjjb+0lfHc39DuBwDjdDxHd2topsCZD9I/uzK8iBB2vzWu
y3SQq5I6vvfUfa857snAutgRB2DFLDShGMMh01ayZCetNeRVzCn2BESs0vfgxizr
0wStdZLLr+kE5UzYNrpXc4G/XYD2QB1DiXc2ZKH6KXUQ0j+dHCOzzbBFMZnRnkQb
CXbXdRmXuqz3gRcMdTZdcVWMkXzR1q9UZz0ZNtQscS4Aw9mAQ2hGFnvUfWLjjQcl
ONraunFgPFtAdOZZGBeyVmsdX84vmPUjeB3KPEXOyJiv7pUQAHPgDPLagBOMNy9e
RQXWyGSYj1k6pjRLS8Mgl7ZP5heTfy83wDl9XDChMsBMPKtbe5t4IEh/86QgJADD
IT74op23zCw7ROdbfOJbMH0eyP9atKgV0YvxeQB2ZQxby933I6irN+M9qf6shYXx
YDZIFxvKjI/tKtfRF2eoLXR0F03BXiJRBgWtfisTjtO4c+GI+4rWcm7WQxRx/vhn
1RHX8Lwg2EUml64U4up7ubG2Wd4vT/HLSvBhzN6KknOi+ageITt4uyNsh5qM7bQK
Lc5VbOS6eBjwKagFLi1nIBUxV/4R8ckueVegU4dcwD1u4cXNdbAQqs5ZO+LdwqR/
NYCwb0v835sGJ7gz1rQVrkA6c1GI3IZv9UUQmPaYbLkeHrX8pMbbgWXp8PCVnVbc
fcssrqazJldTI4FnFmDcdEqIXsxi3sY0aLXnBFcrhOjf2HDg1r57msS69yknO6m4
MfM0bmZSeysdRi59wh3mw0+9kMpNwgUUSv+HPEureC5k4RZqQFCdwwiPibJjqV4x
UAlA2iwARInAJhiTwjOFI6EpL+86QW9kblzIIdle4xPfjxarTRT731erqjQYAvbY
8l4zNLn7JYCrrSb63l6Vb4maAtpbuMW+v/t7m5+oTBo9R4QBuRRWq5WQbhMv92aL
bmWVPNR1w5Xdv4N19Rn7TcuYd7WNwk1xvHFChGyokR1Q5bJHlzjNCRRf6hmEpNZV
oe0UE9s9Qdfd1l+upEqTG63SbftD7IKu2gQlLtqVjY5x+wreWCiVblEFProypEda
swHQHB1TDseHMuguZZbh8xXbvyWcJCmHnQhrBrzlSxFuDjrfuECZJT4IdbBbgZc1
Myw+sEUgzyrMO+ioFyuS0doQXpAQGNMYo2jpMba7EMc2fMAn7ehY/NZyFfhxob8J
cFWdipwwhVXXGCRn5rDF3+sFrrkKG/wqbUhXtHmNLEL/bWFSuivgtnff/Hbt4Wxf
Iy3pMq5Dt1YCiukz52jae00K/RCccyCbA4LHpSxmK7iKu5IaeD7Rj7fQV+g6ALOn
DNxqz4U92G7pwCBgi0a3D0EazcLypHgd9aLMWK64v3jn/R8lUeZwYOep0o7JQ7hm
MKzgMdUBVUUkcw1aDiTw0sZxsleWhoOGpTkQnbjCX1x2K4pFD8N6wKP4m5mKpXhd
f0vIIhtQf8dLBgvSlbEVjgJ8oznMqFVg6kW8+fIqnOqzrLOhH0zuWnWVuxV2dFnz
IK5HKf3HBeNFoC7j84Cj8+bvoFGFFBmmvXYRbm0gZexZu/yDHe9EQsSK0I4/gkpo
cZoA23xJ5B38Vga86DaY+hMd6ROBVOIK6nfWnY+X882LQYus/dbJj5ivekSAiJpP
+u/lpa6KpYnEAzBmP6rNgeuSg/PViJQZBPpQ0ys4tVUtkX8G0wuqqQJGAShxzQ4D
vMJuTXY6cbjhIX6ylxnyFyykTtXtPeNcGtY5QpweFMKaVuc7wnQsncExc58j9LTi
tCwb0JcD3Bi5sEXFnI6nCUeaQe6uScfFT2hi6M20v6bul9PeU39DVhYpWKjqrrIz
nOyJ5j8Mfmay8DmWzGATi1Wat86WLq/DOV66OEGzolhZoifE2hlNRXYD8Y2utxXn
VRLUJ0DImksLQ7tx/ndbDCtQAeLPTxdlIBSCYgxyJ8bUzzqJn/ITQ22K37BIngsT
INYBu6ldkNQ9m4bdnQN285illbwZdEx6SUmqLi5GURsixqiLj6QVd/duKmPkUFI0
w9/+KW6zbfsle+yVw2+PYPMEKlR+KYfSF5wdJBGG80k85CcpovkGJh39oVpi42xY
LJ81ovrwoqpFjWsSdIFOHdOYQA23W/yrg9xZJWAPkIjZEE/N/jZIQhBoX5TMOh22
scNhiJRD9xYfTt3LzMhfvwrhZAd8S98LhtvmctU6EQfTFKyev5Aic2ttHyM7xqYM
QE6FPPSwRCUa7XVFDgKIzeGDm9y6ehqt2YSxhf4ofZrI8KVlVzdDrDU/oE0SJhek
hafNYpDh2VSOUokv/Kbl1qY0Q2dZcPUUQd3pTs1V1uJpeixQ5Jc+je9ND/DVjFwY
TVQZof8LYyg3Hxdt3NWrrApXBbiZy7flEmueNKqcwuD++tci0/499zDmZtakeTnk
x/7avCSnM1CqgIpSMG/ys9utwVPDc7TUzVE+EtbjiY/x6f49GfuJM57MToKkvj9R
qyGoNpAKo3+9jDjhY4/dTiUwhlpjuvQmngH583sqcX2OTfVBRLa9FjEc3Ckwm1b3
DXGc42StXZWbhvYQejKbZiIp7rk2S6xkkIlhvm+LNuF7j6X9ylWy+OZqSiCjrtcV
+nVJCd3hor37jPg2zvRdzL7IQjAkLzxF0RS76Hoe8yaahkdJT/zKmWiW30AnzSgt
6ClubHrlcoi8mc5O9K6mwc/x7gAOO93FTOOr9RIw7hGGur5AbQICynlfvRQUtMrS
egcjrb/Awz0kBC079FbCIvmkAvhVD9pwIYgoU+TFrsIJWOoudifjUQ0C41jkNJjH
ubqi7PatmmLSjYrF1rHtNGBogrsLDtlzKDyamTJrOpySzmfeYqOeVBdl0kY5gk+3
SJIcqS9v8MRf4b0p8wxRLin4uqlyRbd5tNXLZ8y5jxnSoEc9eCrLqx+y7/dPCJ+0
Wwc7mhBbNSzBGGq4aFaQNPS0MaD9warK6WzSaPre+hORJcANxKIa52zKJ6NOCZ3P
ifXpJZmHLkygkBRfpl8Bsmw6S+19qais+9qawk+FeosG/AwTv2JwI5aHmQIHBeq5
AJ8jgeAUVJTqrF1YlyAHFPNRAavDcakYgSlWO7SnKda8CoIEuGGgYhtyMMo/9OiR
KUFTi6Mr4h48ESjBQg+FkeZn73Bj9nSPvqRuv8HPRx+86k4tjAnMZ+plaaSgA2Zx
WiKKF3So1UEmsdXPh06lAXjXChYxkWS9mgD5vYT3S9TTaQIwXB6h7KcJDTzJpD9U
iMJecaRDWZqgzZsgktG0OhSy+FpKqSo534034Wp5ljmqMYptRrDeklq+BquCPRsC
Zt9DjkEKR8OhMZ/7fjHevuor6nHKtM6zU0rAQWz7CdlZOLD5G1VecydiQaeaE2CW
rZzZdDouAD/Q7zrVAasU0D6p7ADCaqCOJcXiEOa4y+eRm8+D3CBj/FYhvoQZtzhw
odJ/seuUA0bBfUjOsZoPekZczJKKS1FKcY4Frm9u+aSXH1C+3OqihsPL6ytioT1Y
Rm605Vo9HmfF7LKzDvxeu92oEpnsFAL7Y5vEWdOgwDMlj3dFaHBEkvqPDFacsMnX
Z8TttqxwnwgF8A/XDCp/hAfyQEraaXD5iVPzntdjP0UW1jQ8U2NfEgDd+AOYDTCa
6QZE44mTbaSuAiq+fxEEGKdzeg1CNbyHFzRdVkdm8dYvWwwvMqOzy4GRcUJByAKx
upYW7O5DUKMqiQH7xLgxPlDBS6G/thE/LsZbpmTRP3UQteh3oY+8FGY7lDpo5x5p
/vu/Pf3kaQXUhlYZfyQJ9Sj1veXGcAzITtxUnTdX1IGiFBxc2dIxwVgmoGu+040L
c6oinCWTC+euhYWbRwaPz+bu5c4lYmwS9sMjKd2BjtGwAIr+6XLU3OCX4HRF5tBc
blPqAV8XMSL1xip6U7bwCzMkB33J8tc8uJSmH0/2CfmyBvQ2v8V6lHHQcWniSdOI
i42p41VJegpNBws07hW/EcgcUwIe4HCWBuqINrmYyUVEjD/ow3i+V/fv0JkZZdUC
P+ySVKSTgVOYjY/PfOKHwT8DZspvyaq8p3rBQLZ7MOKi0jhRTk3v6Ju7KaZqE3Rf
/0rKlOEed6uFN/T//CX5XTXcKyb1d3EagtIcEfX3p32R9xFX7FdeWaa6KpyK0BRg
WyC4ZYAlER9Tpd2GwiDALHJCAWdiE6ZLVesZzn5AkwGwx4s/Bw9BsTjxadAMen/K
t8WtRbDg9jzmMcYo3fWqOA9IIkTM1Mpvnc2oI5Us8Ch7HoW+UWFOSWP5EbvwYQsh
XRWHxEDsiiZ/F0xTXFPhaP3n7ZfG7Ir6eBLC0QA9ngH5JxBDG/bIh13BGTqZWw4G
3zG96CGEZYmdciHpJeLhPA3R+uX+fAlfrOTadueLsOb45RyFuzrZM30LeCdq3M/U
/zBZoK2s+9f6K05z8bzJ16DN3HS9aC7bqU2/D3kq/Y2Ukyw0hJiAmqe/yY6E7q5T
6PGiJn20Tp+Ik0KrykiuVnEJe4dqgwWEpBFnk8lSr3cLVVSb9olsQQ448eWTNr/G
jiHiRhDW6csAc40ILNAvNFYjkFBjCeALhlt1LrCz0l35XoLyqPGMpqy96Jf+XuXH
ZmNk30+TFZWC5r9r+zc3Tu20pAv/PLDVzTuP+6y+u0ICuF0ATFEGX03eW2fF8Dbm
5/RcNa1B7CM6kaAKAYx053dPiDX+EBIrTxJlMKNd9cC8dgkPtuwyvlzTzZybzjuH
5/DN5JaJfnj6PZxiUu5mXpylpjIfvhN9t2npPYgliwPZ1jsYLVrSl8s6JIeir9Kx
NKyuVVimFRJBO1sMLqxvQ2rOV8rfiwv6DIfdp+62h5gcRHAB88rRTsAy55ZAv2Jv
bfgkIrzGyxn2KtAbQDrRo2iDli1/V/tCSjWNoBUDpapcUzaPcEVPanJ0RB0vLFja
8nJZFeVTUwRW1s9tELetsiw13XZ/0ZqC4kWnt4jY75H+OQITTN8bono0kK5gpupT
bs6NNCrisv1UvWBMOBkuAFutr/RVg9XDFDxRk4Hj8DNHijZ9XLJjHrwSkO7ih7RY
788YuqeCRFtOqZjSUMowm5uGopwafhXEyui1JsM+JqrAUF/pqEUDYaosSB7SVTTT
UivbZGf6rTxiwRLkbvhZIAqGelU00ISk7I2d5sxUeRjbzriOv8DdHZZZZjqSMeKB
RR2pOw5H99yXC00sQomBJq7Fum6nPmPPpxdTocr8RcCdHYN8QR2JYrPhnOgVPY5m
8DaquIMyzn4NcYqMUSu6+nRy9nmAbeYP4WCWGUxw9ASzaKYLd3QrWRCAbcvR0Qz1
wMxrhT1NI2JH7w23bIVsIaZsSLMSi5XWpQC9u/YmRDoQ7cBY0IG0LhC/HVO5+tMJ
Yk9ThnLL2YYyMn+L32qs448QLxyWovqunqtpAy5GaaT0J1p1KB0YnTOGrZO+SzHj
6+l7GflA9VLc15TTpMvqVrX9cnawS25wUh48+X0dZ4706g2pJeWPW5f2oI84RcFw
swBA54CeJjCbhnzYMW7tjKT6tR8zmoAl7k9+2V7xlxSgxQdFU0NQtErg2B1q4/hS
7IISECJ3nYZs1vnPbgmxFk+006ukH0NlsWEF3BJcfhEBX8yuZFCFHp0YHJRBF3hM
D1oGGq0TcTrdfSj8lXVtb594tXpQ57B++vAz2wreWHbwBCc0jKGJqjqrKb1a+T5+
09g4kTRO6fmwYTTMnhA0BdoY1UdqMG19WdeKCXYKYGw4LRnlMjxJAaBiRCKJjcpX
9U/2y9J5W6hJGUXdBhwVdKomTfAKTEN+1Q+5HsiiIHfTqHT/4MX+t+UFhOdJMysf
XBw2DdHJVEEADknwLRUILMS0GMao0+oBCi7gwwFkYDVHwWzNwMrp2JI6GcTiAy7G
ZgJSYrHW5NLv1KHaXIYWIbZOjDvk3z8G9247wILS0QkYg9IKs5SE/NF5OZBDR7ns
qQZQDEhlEh5yAR4XnHFHgHrddMk6GboJLC9WkHX51NJ4aQ/6X5rb0+rOriekblk9
K1AAcRYnLpUqbHAie1L53L97F6n/y3PQv2MYOYquz6PA4SpgtDHQmrl7kdvbKusL
qAt+N38rVoWt4jDTySkzK2XZPajD1RPyXLBva3gwQujnFcdmGNWCV35oIjeblqtb
KEI6kvKIvv+Hfm4fAQVzBcP/YUTwMtrkwDiNBZiyU4y/MIgqmyj6SLEFY90HRJjE
MSEyhsFH98OhVwgRx6gsCjPKk0uevbQp6ecWkYx1f38VQK5K9coj3ma2ECnuvtC9
okZSoIk8DwMoNuPX+M9a3szDiHnusEWawrX15YCpKFtrWWX/05FVmolOj6eU6gyq
MryEzCXDXtJZM8GoMQlkaA5tRrybCqv8/dbexwQ+ezEacLOwP80hJ+vINJCUkdBF
56IKhUoRUtea6faE0RfGoThPvY/n9QYbkf+e6RMYxSpIbkwNe8x5Xli3gGLV+Dx4
fi7D+lK1Q1FuCFU2lpoNHXpzDc1ENnFDhF2YX3JAMJ/30lrj/hqrOUPkdu1QrIsB
axyfb2Ui/PoJc0F+juQtz9CC3R64xeRiD57N5pS+rz7Cj3PKpyTOLO2fmZuSpxiT
kHSH3iUvQh2Ey/s1dBFwt21cRs4aXEldCjroU0o2PgUEuPVIPzOag8rtmCB7VQdc
maZrMkLkPUS5CR6ffuEQp7KwWQTY8ElgigGiu7e8nUorQu48U1MDB0MZGWsCW+BV
YftoqIWKSP27FteaJqk+bwnIwl96HPYABzHMjJ3AVPxWQEjqe8nWGnZ++u4ZvwqV
kk29yfx1XzaAAFfCv5F7OyBbyUEFFAmB6zbRmkctmDjDnixbuv0HlQmNHJRTrCrr
+mkrRnGFRWPcN6ja7Mme2pitVY7vlveVw/Chp0f8hUCxSmGcp0Du9NkK2tbPyysz
v2jFN5TTXptNRfAkN1ESvizEdbkcbSYG1t68PPKTQMgq+qQn/z/VYHDMXHS9PJ+l
5TTEWcpLz3+VbdSOb1L6b15LwOSJq9BrBZc4pgkaF7+/Wl7ApHOrP7ZzaVZzlFix
l8P1AaW+bMK8HX+9ZaNFgc9Dtt1pBo57rRNLLAG0tFvj9GVFA3tJl+oq6z3/IUhY
LMba9wLPS2O0YzyhIt7V5N7l4ckuIiCSpuzgu5GmT0Qnv9ISQzjhn7UaRkp9q3Qd
oJ8UMigHBPo8W4zruM6/CO6R1EAbs/w8dZN29V89nfA84Vswujjde8sMt0UAOpqH
LvDjczAKHVjo8hOeCfayjhljicSQbJaQS1Owdq8oyskpC5jdqPMh7lzRqfRB32Yo
edvr41ZzMRzfnUJ6/sRFOsNUHnextRHPnOM6MA/4R4lL0pE5uKsx9aW75M43xTjp
KfJ9nPs7EZ7nSEJUer2+33aiPKrIeOuB1A8FGnDHvdW4NhLRv5DR7ZhGuiyHuFiu
tq2t9pYqbyG8BDaq+8QY56MwiVHrpqDx0xuPe1VsQSRLFQhs4eH9P368iYhbD5wu
UgxrYHQymOwb+EgUy8rAlgdvBrDALVQ6i5YEoS3RGkom6Vc5xtbIN6/0M3bdbSA2
zCCaS1/dj/96jACbFMlIQudcp0plbxHWc3peEv6c2hAZ+DIWJlGpJdOUtGczTwy5
XW5x2uOLoRlFcR0lbgYiMHEBuF63nvzdTr4GnQ/4JyLVCeZeCsV35VqjHZhiaUTK
Zj7Yk2VgHUTDG6mUi88MsXN1hUdm5NVKkA0qDDI8jVfDY62hxWVG9hOqEBUCG4sJ
HgdetxLDjGvoS24LfdDDutKfbYwuFUg1ogXafhxkOFhajOdmb4H1/Yv70q1xNGiM
bN4P2gEF/D280qg+cGJvnnuWPo0CRXscRC43fNHJ4cW64acX7ZkvRQHhH/lQ6ZMw
qBci1sJ+HjpsH30CfiLl+7pT61SXmthRtjXQtMPDGY7k4AxTAOkmb8G7zKozZXI3
3K/5xgrAORifJhd0DRGAfpOAeHO8vOkxu1JT6M+brhJLmY6eZyiWiqG7gLEmuNDj
wuZ4AniDUXvdcuUtQMchAKpxkKzB0ABkWJlDkLr9Dp44ezoDlFKJcKUtXe0AULt6
jI/Ld0fV5pz5vqGVnX2HaZoicU7IPgAkIO9De45HQDO9c/2FitpEk6IzbYxxSUYI
QYm76mPHilf93b+QxJ7vRHVUNa9luXx4AIyBP8QC/gvloqmdtPprrUkyLofuZKHU
QYTkflKY48mctSyqgbRCnDKpA+ThWYN6Ka+6enDxosVUSLrLbOPd2pnXnoR3YuKa
YyFS9ex5ovfFS+2nEv925W7A3DmZZY/VwqsP93Sv4WBsX1Z/EkM8R49+Cf9yFSnn
fj3XHxW5DgjjKLdrs6Bad4y1wR3lWWh6pF7COOB8GAHqY8GeTkwYlv64n2auQZMm
vGTXujAPudhVcTvZcIhf9rR5pK4O6d6D+roykn8lo9xDS6Xd5sGVUSJZ3v31605i
Cd0ZLuN/+EyidZ0uLsaGOC4KeLS1/bJ5L28Ufsplymm4681x2CIQa6HQaf1NeVfC
/1JHHMZebIVSVdbsFcd12X+uJ6o/68oKAkqMj3Sn/RzDkqnbSOGvP/sJreA1kUwT
2d8ZF4gYr2fxEKMyNa1fmk6AYKuk65R1rogq8hVVt+VWLzhu2Q3Lx2VyOyT6SuZm
saRZKTFO/v+HAE3FD5saLmoaCUSSVWdG7euapwcUzXEKmMU7ADxx6EhqdGOkmLxj
JPzLEx0Gifs9WbTNqPV8VN4n9/khNPOjFhhnWBVwFAfQEAndgPf9Mf/LcusdtOrU
4Z13ZtcyHxt/gC6EWH+3PfhBKNJeWXvIgszilphQFK2e+JOJdsqo2wJKP6T0DvdX
2JwXh2hNLGKsjwTapnzA9g1uRqeWBF502pSnVVGJpk1UXJBMx4gPP0Dg3zFjgEBZ
q4xOeSWvu+y9FgLbABarphGAcSlbf5oeRaS8eCU9RA0NVVDciqwdPZfiFcr4ny8A
UbCkcNW12M2jLBpzMAnXVGLH6aTB6ylnirMZuD4wGwS3jR5wmK+LGCzgtntvglEi
vaEsicGq72yApuz30gdfMalBclTbpk3Z9T5J3kgL+BUORa6tus9PHIGURl6w+wDS
DJFxTzV85DqK6fAfCy/FLbvBq+xJH9evK/78irb1cdhig5IjX93z98aiFdCsaTa9
RvxSsdgjAGSVnSdGqs9HQ7TFDpzvr2vxLGvNrMc84W+wpTo4hDiuShziA5biYgYl
4y2fNMAqHXYnxP3JT1r3zCT2pKwW0SEdVze0+em+EGolIMzDuab8oTUrSf9D7YIX
9nbvGRX3TmwIOZ8N5dW6d/RIX8cvmcxlwUvtxuUeWpEoot/l9j59sdZiA27B0goi
e5H0xDVapRdes6OF5w2P1SxIXctgESM1V3fcon7C+K8DvUshmT90h5LPzunDxtx9
G0JDS5KjmHRH8ZE9sunpfgXTqtQrO8ocqTXKVJlhu1AHKwA6GcGKeckQpeTvZACa
9utHLxHQ3+i39yBVaE3OE1ahnRs6ms++xHbnnDOswvVydZAUZelOftNsM9t0ayQm
PTLLakj/fshAloWLgkgpuP4VnCslF9NNa6iHFoO615QfzNvdYB6lrZkAO7kWUnVW
EAyqjFWVIDBK0NCnb8SxzaTj070Rk33SrbIDypy8XpxlBD97fMY6IGtXgHmRZQ3R
x603RrsBJQ58P9j5WoSM4mUnGy6iemcRwuMHs1m3Kmv36w7R6lO4UjqPrELXbIUm
/Gw0cH2/c6KE2hmbCCNGNRZgoHCe7MLRQnuAIchdJirS5zLTeHxv0F3sCRGQiqpo
Ng5C7Yp6ylKsJlRprF6QX+66ShSd1SkIBOBMLo8N6eRIQOzm/ife1NWd3tDXKfsU
EKIjP0iwcRlIJmzoBqSe4D1+x4/Mu4sPcuRcQLdyy0MEDY+PJQyyKaV/dKiAyF2O
cdHf2zRk67s0Avqn53qzw2nUSNnyQ/qFNPCZUr6ZGzRFCMbz8tpl5k3NqN9v4anQ
dXBrPcu+mvD105nH9eGD8nivfDURV1l+gtOceAruYXVOE1e8gytldEjK8nnz2fsw
NPy1evWWFXFAmjDJM0U+8XTJG7T1e0yzfQgbdk3Jo5PfXAAN/Z8tbk7oopvIc86y
+MX37n/vtZh0fAeYJ1oI90TxZTJTGrc5gP9bYdXZoZ/mxoOZMxhPFME9y+FmIY22
wmB2ZdWhvF8vzATxOPEHPGDX6vLKceXuEXxot84xqkbDGtz6v4kTBqBlLbCk4FNm
Y+P8CP59n8efxuceFHjJXBJM1V8dmokh4ZkFanKPn1yEAQFsRNDXnmGtIY53A1rU
G0g4x2HfHbO6JezH/751sBlKL/40nVBdE6kSN56rjkdBWpgTlABZ84ElDV5U1uiZ
QemivvElVrmB66Im1tU2p8nDevI13muNjFFVvvS78QUwPlzcNovI1hUwMTpiYGJm
CG5ztVti8CJaecZOmgoRmWvscG+I3mDlBZvr7KsH+JacJL5RruwX2E41lZGp7sho
2hZMW1O7LGPi2+FpPBD36SLV3ALpZqx5F9jsGVCUEFV+vi3Z73cpg2bpbnQDeXee
590n+C+87hoYadBWx++mdIHKbcECJXIZJe3D4eiyeQPpYaklqMRLc30/L2ZdmOtM
geK7j/8D5AEm8RhCfFWhmSAjsD4/ENS0srp4CPgt3mQcFWKM82EljOEzzo88joKg
sc8hZouo6FIGwBAuL4su91clNDfgDjVJSsuxjctdudnpHDK6dZEeo+XkdkzWMjjN
uS3to+AsnmLztL5wTUn0V4NU3gZIDIIaw1HY6pNg230K8XrpaYUN6fgDWZkjKs3j
AZAkk5Zs+VxwhRLKPHWChbSz11KJEaZY6jaGIG7NTxryWCU71AFTJa4DpLplj0Ch
BmexOcQx0Tfdt9DOC4wh+1XNbAcxBbONJSNi5QpNUGtLACelHMStLLJBM3Rad201
qs9w2VPO+NIonAjPP9NdqdzIQgv9pE2WBcEiUPgQyEddI09SjVUUSEbwdeBN+tla
w+xD2NNy8zoIIN0YG+2ecjHA8PCV4tZ9LOUijNVu4MtsI98rFK/S7i+JLTQOvCFk
7CcQNYCEjVe9MwIcWX1H1qDbgutyEahtIYmyCtCzZLfCkkVJzM4VsXl+cYbZoA5b
9XemGuQDCho3uLnl75GnN+517oOp1mN9uShbgCytHE4o6jpfpslIzqBRmBl8CWYU
7MIruUK68cWXGI2QkCOGPA9msYs4+VWYUfpsYc6iYb9beUJ/wMU73b0ryNhmksnG
fuHuJGGILDc8Nb/tGer4n9JRSxsP75osw9ggnv9X9U3Shmp+mXsi8iwZ4YupSyV3
S+Asq+7pwSbug0VcgDhDRBarLiB3pGW1JTpXZ16m9bDCGlahp14n3OUjnRyv6zYz
f+JMtoZ4BpBbNLVzbbanCdN6XAqPfPKYRcJFEVi36JIxOG8yGwxMOfBMjaJTriEZ
mrdej7AJMuYxpJuT0z9iyQl85oXv3gdbkWp8zL8/SHmLHDT2HZI6rhDRP7Mrl0Cf
EU3YP4WgCYPOi9bAsXdqY7ppIs9MKImDe7ijkFD0xtN03p78vysaQIk2AJU6ZhKe
QQ/eflZcjAWR7iyGRcBYAgJ3nK/9BKKxFWarEa8lVR/DqkPuNzytizMG3f99OFTX
y8WHpfTL5vmAz/EaVQo4zZCFSJOCb4r4lN381Cf9asaNrICcnb16l+R+yDvHyPkJ
ZX45x67yHE88JJR3r/sdVW3pKPfvWfcQLSDsPS6NuFmaLt5XU0PRXueCsjqSADnp
SYEvOak885JCOw1hCO9+V8QSQFqXblJsw7WH/mgCniT8j+liynGFXOtOx0/+J/ZG
qRd1JjQ8rP3MPY1i9JP5rBVfFwLE5+lT/S4ddrK0u43pMIPFchjKi9jFEPBwWxH0
/T0mvnzTNF+rJWimHpV3R7L/ADq7kWnHI3NFiuJtAAZPFSKqJ0v785wQGyjfDxhe
Mki+vBe17kFZ2lvl+FRQpzGL8DHWNKJLmycFQ1El084zv+vUk7NAIct8VpBRiTqi
oL8zO2lay92EFBpp3otWKCQwMYU1kA5bJUTF39f4sjyq+Ly2WEz2JyFLfW97lnva
UGBfan1dU9iQCXWmuTYTlB9t3nZjxCw/g4G6XaqPddjiVydrUUjZy86Lwhic1mkQ
eklppj9pMBKxu9KZMC8XxiLQyJHeEYHFmjglmWKWZjT4UspvADfpc+tbUBY7E28D
/meZ9NRcU0GU+v/crSvHApr2/Ibc6E1iSVhYMo9I+NPMeIOziLmRuf7MI+DKgRWE
HNjbDCrK/CojPPePtVQY3cBgx8NkcCb3E1ILXwXt39cMwb0CDbjrz3M3/h0cbWJq
bh2B3Qb24XEhKwbx3Y+FFKYkqX1cJ9uqiLnVOWuTqD9Rht1kpS273u3z1r3qCV25
h6KwXdltke3s4DNcq94t6q6BItUSy0TufC2nzbsV/Ava9lvpCnEwgQd/Xt5yT8ma
vWZM5tkykYZf5CLH0jOGmdOFL/M8B4rMPtuPQPzRdI3ALcS6XNnRNi8pqBKaSiOP
vSKl5/EhXupb7K1bEZ2YOMIEyGYPasUZt+cyYN5Deuan5I3A0RVb7OR+wcaej1+X
rkbg7qMdjucs2wSrK7jYcditr/apRugLTVTDYs+rZIe2+WOIP194eWmiJKsdIEok
xTFDAVajR7Q4hYx9DqL7ZEDuvrprIg/gT2cPklzpEB2mBK31FkUwVh52ei94dgKr
vC7d/jSKBFT9E0pZdgP6DrBVt75zlxnFxvhGcmAFfUCYCg2U6yDdPmSfp3Zox9PS
DWja0wiyoF9XYZreAyk2R7Hoc2N/d0HkRs6FePECioRIMX736AFLZpIL/1IKuR9W
Obo5611nybJyzN0ufbH9QK/qq0aQbAYp8kWPjyM92DQ6l67+sP4Cvnsf4onPCNIz
rpWNxrV7TTvjr2swQUkPWWVcV+tuHel1bGbjDq5AgbLPYiGTzeGLARX3HKl0J8uT
webfpIeU8kgJCT+kRo389TEx0NyfwwNXaEspDqgn8az0S0iJWselKbIZc1Nnm0/O
Sn+2ytdZx/XFhNwT4SY47nbjHpCcPnKnj9Lv/3jY0eFhpJZZ7neWRRV82Z02iQmX
+MunPULzrzZMTii1Pqi6tLzLmuNex6ktUeWELhRWu1EVRua+CPmt827/qnWOjxHF
HVqOniUlgYBC9nHQxamKpvZLJyq0zOLmopcjz3U/opmucveCht2ELaQAklMpYbF8
2Q9tXT/5Qik5U3C4IZxN+yuJWBPoKLNRgs9/GWzSRu5e3tZtZZ27vrvCcrZON2fk
lg4K2YCdb7RYrYy7BTzCBjEerPOOPgYyl6hs1y89WYSLTVYW3ag3q9CcWDvCy4bL
lmNsisR/UK1Am1pW3L6baUmL4wVdAge/gMjeLN2EgvK6Af69N9ePzPK7bFcey+bk
hoeSjiio4vdsEaXLB9Z5QmrbbQmko8xVqigb1cf6h281Kf3RsVVoN+X+bBooM5Hf
YrL+09BP79DuPTwzcN3N19mk939bt+YCpdWWceXI5vDEuJfEfnZJRo5v14234sQg
Xumjn2htPKiiT8SRfIoGhKN0FCCT8T9LpfGd2i2ZqNvLigMsh0wb+Ur0WLb/FfUh
j5hjHiJxU/I2siaBgT93J7zxl3/xvnV/i/CBDngj2lyuKAmyJ2dbIZlPT9HQ5Ovl
Uad4H1kGxTJO5BOpfQgHr1EuxU5agCeFNbWD1rRk4fMEH/vX2jR6sxGv5cvx4FoP
Mic3+bGOQi/fo8W3JNv4NorvmdJDkZ2NeKa761+c6djlHrJp8tyDhKkoGdon4UXE
8gMnvG/8O1JRXp48oqMQyDTB6XEKLbrLuv/lS4hLxFat+EzKkImdQtp9GHJ2YYSX
dsJwuvRh2TMx31WnGXxVEIsZ0Ij5qBhN6MLVMCRIO1Lt4WP/ycVgwW1gIuSGNS8Z
KcpJezqQNgal9/IWuwo2TE0zzS6WUzCOVhW4SlMGYOwTveqCCyctZSHBhpP7/iy9
LAhEs+zMjZlvNt0SKoHVhAfoQG/OTlSI2TDNYVUVsXPWg+GZTnwQ+0YrOi7jH7QH
Hpuv/+OVTTs2LE4jqiQo7d88ditzNww8vdRcKeeNrJxnx7abrXzYbR/FpCPAx3Vh
lbYNV6XOc7EPAsnc5uEHRMV8bpIjHQDqjYNwsf3Tl1UGt6HQWd/3xUms9JrgMC2O
0kA5EdmPZ7DLZDdyPIlRzJzkBrposyKRwS2peYDylGfKN9bQUniY9aIXOGR8CDgt
YzbI/1OHsO1Udc7LhGZPVEK5xSDeWZUJH7rPA58ozgOokf3/WHI4pjwsV/sE9k5M
dBfpFxddsBti+UETiD6wshPAkytIA3cgVUK3Xd4AXQ8+MXiNmigqJhzymZBK/eNc
G12syPcIkdihLAbOe9PQHPNlTrAj6xc33hYtutqGWFIRscUbXcHmNlE5lUEn0WVC
BPoqm7PFyul6AogqPuX1+croiqTkJn7QnQm1ywztWfQ1XjqPAAjId0xzmtyqyQ45
ZEseboZkRGeffLd58jMGp94/dZegXDWBu+DBGDE2KRfdJlruq+3dNjBmfEt+1agy
dzz50df785lCypwFwBXdfNt3XSVZNnDJy86bdIGN4QIqDCLiXP5KUcRT5sBHznFj
tt9n4fykn0M6+x2z9B52WXMkHm7XsDkStEMdo6a7yZvJ4aRegZxiZsVirTbKjq06
H3wSNlRbtvdjHhN13nvpywy/fSoQ5N724gvYKji/AHhgSMTDXuIrqiOZhyYG5CT6
wv6VEUVKLiOtFzH78Fk36xgltDJwKs1JAzOKhacHKz5y+yDqbj00PvrrSSm9b24y
FR0kDEM0YIZa6LYdfuUxxbJibC38rbhfiIWeUcqIaS/xZEboPYlpVgbdedcClnhe
gxwOGnoagYcPLXUWDAC14OV0QZPmrXhYqMMoOTgCPtmifU6CneH0x8MenWBXXgnu
hip3w3nX81OvvPk8+Phl20UWFRxD3rvyZlGhji1APnwDHJapPNZSi9LCPXu2podt
9cCoUO4OsxxIdnpvoE+2ET7PsjX7QWy2pkUE8ZKt3EGyo0ztCGTz3bZLvxOl8Vwl
LXfK2MpJMnPQhM02frAcqsJDLQvWuSO1SLuKldsLJcWO/MZVzdy1oGYlMm82O7MR
4xf6TUEkxITc5+VFKLYXw1V/xGticbfvEJ/CjE5Fpvg/RdOxp6bewlDQmKX6K83a
07hYw7JtT3kf43+eBgvgdT0VX2lCZ3vn1DTDfzkoE+UvMGqamfimsoHmULLkU4XM
xo5JNpQOcLtILmG7jSntjtAd8wxtbzaKexYo8W+FeXICkMj7x0olc41Gag8k8Tqu
1qWXWO2FvPR/hY5ceBZOV+4B6oUOkH3yMR+Hlcm3L6gTOcMsQLE8CVUN0LJNp8Cv
XDVyoBfhHG0M23g/ygOtByFgDX87xmGmdNeIYAD+Z2jGbX6ALpcJUlhxDL0egtg3
ogacIZSrXRphUWvALEfDiZ2GeaggqYxjYkmP4pQDZGE3hDfr80YbjrXMqm2/UG9F
MzJClCkQv5gpGL1y9EYLAwJnf5iQ9cLKoZF/Mfq0pmFFVdxZBbZ2nzL6Zbv8NoKt
SCXaqexEy0SbyWzUZJnNfeDWkIH5VId2ua78EdVj5JO5KVFpGY/xoRET7av91mLK
Gtk1Nd5kmbNqizp8YHahJ6EK8lVNFZIJgQ/UA6wTX9DFRN0wMIcKVMQmtbpstCTl
PQ8YkaJaYu87fQTHzNfT1aSJFk2kKD3R0F6YEHBFifvuvbVZC5IdY//nZ0MCMNxG
C8NW5AjPHUhHgrqzgxSylV0AKMlBmwCkbAjpVdY16LHLtuoyfks4UvFaSdwjWErO
Pg2KcM2OxhyEBLG04gLbbejO2UpBe7wSUHIkiOmbk4XcsoFS5oQbJEBr2EUrkicC
p9dAV9AeyNL7wuvHjQDsRSCeRVAA8GDmw7Ld6uK5gnnZUtSAZ/jDGcAzX5aAik2S
O2u6A0WPLGdqwlPWTMHx3qnu7UXFhMPnqJdvIsXEckHMQbrC1DSUqO/LRboHwi1J
f25YhWluhV6YPTEggX7rhYuEYECi1tPTI1+heKjmuYOn4HXEuy0S8bUYvi+omQmJ
PYL4Z211A0nkBQ2o1nmD3oGmGqFPhqobyJ4OztwF4XAPKWfXOQdSF+z6wkESsxVW
t5nD1fBwSXUgoACPNh3HgVUS2tNnPZs9nkD4MLT+4pwdA4KGqCLjuYMDTV4R52vv
IvCZkapaG3fH3G7LBhnAQQxuesYQoau/Qk5/vrd6UB79V2AohCOZ3Y6NsO6dZdUg
jAQsF2ov1+dov7/SoJCeOHIiStSeyrcyqvCnkFMVR4XxslTFuEgKRyEIeUTJ+j24
nORnsfF6tvHF5SOSnFZzqfXs4ZRhfwuUCaEUnNLoCndndrj4OWSr98ajj3Q+FVOt
2fwTBkgJUgaLcmkx7k1DeIBrBflNA2rc8dz+vlY4I3q5qBxhCuKgZAjkm9cWsTts
OZCuGDCtimm4a7jEIUle6/nm/QlKexSGLEPr3d9DbfL40DAF4xcb+p1QR5um9OtQ
aDVc97Ydxj61lMdx296kVtm5yY8Jcq/cP9JTZG8EcwUB7l4iCEizcH+wrBCOyVLL
sELWkKO27y+84o7MGZDFn5S4ttAkafPO37/Fwvlop/9g/ABBMJUA5w3hvF6I/58E
D+Ghv5UOjQaIvSy/2O4pRphTU2Id/jZ9B661eqfXBIePtIJrM+ABW9vlgNWPPWcK
4rK9f4ym61fwStRfSGNhZ1LLyd7OLnenkI7HqdrME5uMLjl0VmcFxCdP84+bnvVR
4uzPbIjqDwdgcIMheo8JypmxKsxpDldhveSof3OB4OO4xfifJqF+7JiypNLu/Scf
2tVUqErirUlzf9u/bOtPCLf0wBpBUcE/7WgldtS8bE+G0ZbKBd/4XWUJxUgKLMSN
904vVJETFWveENpmy+F5f8nXMSHCWg7I89+Q/yLcVKhr46B/oDdYEZcopAR3zhlK
srV1I/RDOLvFcLVtabs2QpzKdeBB5ChUTgLUCVYjh7DiZatWUGIlVEQ0hAEAq2KV
W2PMjvB40RNscfm82PpjFGBv6k00uTNJkS2qHBnBSD97jnYs9DtY2zOs15c7BGeW
s4np05W9yO2SEIyGjhwkTf6yMdqK/KJM4bFFrvr85StK1LHbTcyHrBbSMp1AdfJa
NVBBxgwEyFy5QdEAvjdUd4u8NooZctR1fNFfujUI39OLZ4gDTjwENLACsVq1av+o
9PeUTFMBN1rPtkTMwSk3xlhHvz8BVHOEdHN9ZX+rSQmr7I0se6pVpRqm5BjMDSsq
XN+p6BZToiBCx4zHQPRWmR8efG2B69FtmrTadW2N65w1ygt4h2arITIJpesJV+Fb
akhhn316am++wV5MRZE9RuPDlCVvQ0RpqkEWgJ23W2bN+toic5nKPLDzFOTk2ETG
X2E7mw8AYZv9Qo1VjZSzXeDe6YaMf3ViegxK/ybJYJZ0UvSgjE4RoW8M0MZEg1+z
ksihOptgrzXjLMfqfabvVMO/EkdVLeShZjIVJV7OLrTDezZaDvKjddsFQsG1KQ6z
8L8hd/Hg7sPhIJT+X7J3mMmaJvnUcqVJPxL7QVLsHLuHzFZeARnsKLUj9k8dnujN
NrE9aY7ie8dM16yL/+4stGcuCkVT5Q79Vj+BXgejBDCfDE+Q3+kdJIuxRBgWEbja
SJqzxXwKn03ZfLQEPxq0QaZiJSIWhhgfd/rpySROlx17SNez58jr9//MJ2D7hVgd
r38eLF9Mq8Bw8NCKC9otmt3E2MaNc8yCLMP7QlEkNfUh3S7K8dhlFr7UAHhsjysP
Y5pAh6cgoiWIpmlqZ73JdIZjYSWQwqMP82pxHPemFzEUyT3v4FbgqIMS7Y+qks2f
SwYANVEOkfXM4ddKMKZH0oWwaI3UcCQXJ8Y7Y8PH9sPLTsk/oqyBhOVqjRgKYOm7
nqROMNRDRvl8N7x1PcVJAHFKkn2KIWzt9dfqo7Vj2BE9+hHfMju6Ti4Il4MLMEUU
hBk8boDnOCPAj2l59gqPDcvsZnpKRJHiwuErfgDZk9k1K9Vd28LLL4+zVLIZq+VM
SnI7w/g2Knkhrf4e79Tx69tGe7KjnRDdtCBg3u7NrOKOHZ88PPPI8j5IpoF8ouGU
Tf/xw+Yz6g8joX20B0TLxnMDJdpR98wEW2GU0IYqpJHWSA+RIl5FECdcGgrq+wtB
tEw1VMKbgFzWVK+JYfIa//p3DZQaZb9t8nnQ/0S1E7a7jSytFDbs5vCdKC2jwbQu
eLJr5vVUOVdY1WwkwrpGaLYJlaDxj+UQukVe+TXarcukmcV5r0N6RuaCgj02d0FS
pdTw17qp43k5IUxbGgWUjztj8z/Eu1zuXMCZOD1ekIQ8nqOPlUxjU/GDaQn7rUGO
dUMLW95GTer9qANWS86uTJHWoMqjCCzdY/3sc3qZ8ac6FLBolwPFGI8fT1CKPaxe
B7XfFz+6vND4CakY1JmyqAloQmG1R9ft8x55oBzLPKESNZBFEBfhd+d8LDBPULrG
FidksLXmue1WdEgTqEaFmf/SfpB9suAyGExfKHZxdTL3vFmR9N8vNInzpu+OCooC
vrxqkYBMRbe1cRanZGnvkmV+Qgy9ch6+9sS1uFkY03r0i04YitOlxbO0aDra0iR3
kAsaudxPfDx9iM+DO5VS8qnF8sr0yoDA9nJ97KCh29fUbDtWcc25zJ5+n0OIPhcp
fuOviI82rY02/BVDBnct8N7Mo7Geq6OKqfpkZJtlYkQnQh6IIILvyvsO1BPDDg+3
3AkImma1vKvAEyMvqaCBru5faxPIKV9aVSNFf8GkyQ9I2sP2ZFkkBabFe9KyrzZM
n1yuo5/XrbJZBERCaENtOFRxk3lm/c+lfXFdwD1MtGGePBdv3WR0h8HIHU0eLSLQ
+doyhKq/8Qtwgaoa0mW+jLHAamktJLXMsQf48xk1UosKS/Lbl58Q/AHTVZrTRR71
gaznooO+Xv64+3n9wjBp51+IiKZkxzCEQfJ03JUvNt+byqzbzLG9Yr2yazw8IcK3
uPPvg56H7j5B7hKoTmc0LtIZHk4fEkoUB2q8vfHPRk8H+otxy6mW5NS71oIwANsT
zi3WfI8U24QL5TjSDWLB9xVmQzp7zh1AIzUnTHe+MiMRY0p/59xGtBjshiQ4ZkxY
bQTR4Ftmwi08bNwTXd6X/M5Wb0TOuoZX1Tn+IOoODyxQAWhmr1yXTn/gtGtMt63p
8xebHH1SG8dWm1r8U9cv9fVoLJQqXmKZ/PkbyqEVoDVZDyBgWuW4PaoAf4pF11VO
JIArq3fCVULXPnnMjZizSm2w20OurowT9/CYkAwRh1IOWsysIQUzcqWWAyuKkjM4
GTEBdoIw4TmWzP5u5wq6C9rrnNZkDFHeCjVJTgf/WhkCEFiyIASTp2ZGhV3VFmeM
Aga+shCq+6gm70nvZEmHsOk+WFK7SpXJGg9DwxDlyW2m4uWgBF2oNGoaYjdp3ou0
WxOD5i/IrURXYbj820oZitfgolAKxNsUcL+Dyuoh/JtAPod6uH2j9jszFtvnrsCN
tdFoQ7F0l8XGy+FlUMuu5swATgGmBM5hr4aQTQZX9hY+M1s3g2jnCaK5uiJR6g1T
dZCczKrwTEHXa5IoWmgfP33WrUmcqF+cYeLdNHc1kZgqhXY/RbyNPzjNv4yvFUEX
s62bnrqeTeEQTzybZyHsLMsMDRPrkHn60MYz3nzK+a30Xye/li+kQuQbYfToedNE
qQPhs1c+47S2ZJPbCw8zGZuSriG91B4gsyOA0JcPX+Age40yahdOlfITi+7sgRdK
GsDROA30gbNrrpFJ6L7pkmnysMDf42Wv5TQuNO5ekmPm9QCq29wwPwlfWKnpTK/7
vNNp79DwZz9CrFZfkxAeMsCcdNhnzGsCJFQWv/JJBLJuqCwY6FoEclg23qACyPkq
5WtxTWQ+brE/YX41NIk0a5W8iCPmVY4Us6SstTjO9CajODsu3KgEYXmicb9AvIZl
loJW1zZldsyrz4tTocySUWPai+OqMd0ScJaf+nc9ASqSPLGFPP4vBvLlDb13EiRT
zQMRPxhYVtMrY6KLNIQg+MNYJmLP1JqoQ+bv2q1wN7S8bYqR8/5/lhsIAAcaRWfA
bB9GgHcgWOreuFZPRtTzEEHQyCtyfuBdZG/Gija0magCgq+lImfBfHdQpTTSTZPS
EQHyA86CFaOf3P1qc530IVpSInH8bRbT6e/9dIDrC+nognyqOayrGy4rcubCxiO3
xVX0/MRxc5eFw3LL+OTuvAq9PakB9jrJI/1T67KVZS8Mgj5CcqKaeZ/7LfAZrlKP
gql6N2sSyT9nKasfRJ0HY226voDN7NSb8e1c1DE57rOZVwNfF1xm0La47/Y8iN17
jz5pw+Ky3g5aXjzjtEkXFRUUMt4d+pZsgH/46O4Ev12D9eBV+Y+QXu6WiHkfCRHv
FwpXqBn+bEPbsEpI8Q6jJxz+KvVmNpxs8ud/Q/XVpYS+WRZZFCrinSQkTBa1HirJ
DcP+7Y2lEWmT7rSLkUWm22b1YMKhfzKTeNPEPYQj4O3T7XPeqci/iloV1vn70hjt
jEFc3nD8XfR9fRqSoOpUOfulorH78sZ8gPTid/ItsxS7qsWK/kA970msq7mIjenJ
UhRMVt12Ipr8PC5RBKNdFk8E89e9LN61wTpVyxivc8D/TnjRAo1/2PBmHsMFUpQr
UiWAfazvA9LDoiiTRVJVMd242BFq8DrVuvk8SyxRYFtSqyRiSiQuyAetYkBcMjzN
SB8oCJejm0MD0QteQNqGnrLO+S1TFJR8LWDTze0UXXUNOAQc3STi6pyd08dlho5L
36q70LAQkNzJslDDqFNqOgYPtzbfib7I45lljtmc3GwfBk/p6n+rXC6T9YtrnI7M
BBkWLSZGASLYq6IuPg2baeWApccslZJSOuaAdNO8FNQ/x/Iic8gl5Lo9Cn2vF0Bv
MwqzEL9WyWRx3x92YIhOUPRu64nkCco6I9rfXbaNf7bsKZL+dacdJ3E063rH0krq
N5Eltxy4tmreqx+efLzk7yG8HAyQcClDPVWDMKbICfuVkA48MXhyluFFIh7//eap
Om1LG9FKBIhcLrmG8//ub3zOIcOJpizJ3tV0jHTcovTw3ceqLg0n8MwDF7MWENTC
//be6QzNI0mDReS53XlDhzXe5WyieiocnGCsG+jsFzyfDxI0sUPIWl0j9DAqO7Pp
j0f56d77oe1/xjyR0eh3Pv+EXUiYShKv2QkSW13jf5TtA669OO57Znb4SbjnsJ5V
gYWt3v19F1hF/iJPzmUTS0xgtBM37sWl1OiE0pgGGfBAcnMMeQZ61Cm4GuBqB38C
s0/y5p2qq8bzVr95C+l1klgFPnLfLxqnVcI9ZilkB52L4UPjZhz3QB7O5eNqiXml
u+R+v+eX1cxJ4Z1apsSJOjohZChDBAUql9VE1Ud0lbHZXTY/IybBbGht+Pkq8RyJ
2Z0khIgqRR59c4ObgK9mEEB59TR+O/55KgsGTtEJ3XBKkphlw194Ty5/OjWLIR98
K93JEqelKow87KrlJ2nh5Emox9HQbGAmZCUnGmGBV2/BqdOsDUxoU1SzVwJB7dv6
kpj95T5Vizd8S0Tuq4Zf1T1x95lSYAX0jPW0H625p13R7JLwjdOvnJte3OMEmlm/
dZtazl9QdfvFOCpQtFhfeF7ZIS6siDXBY+eXmYh4EN8djOxTyn1POY94JPxTXGTE
WPiRVoAu/msttxnpQ3m/O7UlHUQD/UZkDB1NxQaQUGqRSmiap5NfSwtSfiusaAF4
H/NdvLyLaZ5ZMVYZBg/2qw1YG2sCV2V/4vsj/QI9NYnbdOAsKNwr73ee1JOVhlx3
AE+EDt7qoctPjFE0BCYfyIN5mFqVKB1CNUCBKZ0UU8SYpGeht5TNRFrnp1MUEAPI
/ICAzfh+RMkDlVL/VXz8Yl3WZ8lI1wK7P31A3GEzlxA1DtoIMiVYyPomHdufHW7w
HlqpNBLCrmc2hMyNmyCEW9sJsB7bxECysr4lReQtkyFdiXD8TiIBvqB/Wo3BmWYA
yS1y/hj9qB1rh1KSk+fcdKPwDK9CZoaE+RP/LUtr0Buran0JXnJnbC58bQRNiBqQ
QE4j7cou2xWCcMHCWyxp8zMTYsJsZNoIQPwSvu36p+O1Cvf6biQrQhFY7SvCirvi
3kmGKrZJihc7QmUXAjgSmoD0dlmCx83FhcEn13NtGx+5CRpozIplGexXE/4ZHyRZ
iM+TJg/+EFJ17x7FBPsSD9LUPSGHio8wq3jKTH4Qy/lxY29dPLieLfbB7hzAXJwz
S+5+5Rm3JzZdXeXvKiM7HFAlDXeB2ccUji7aaVksLxGYVh4IFfjaNhbw6N+WBdBO
luW6YZ5V7nZxnLqj+YM+ogvcaRC6AgOr1UhtgEnmrLdWb9ZbHWxhJJNjvnI7NyP5
34jNapm1LqZc6c0VRFOCmeNopdRS53bIX5sx67MjZph6n8JdXO+g4pWM/Q6bKBjW
n+g84TiRjZIiDtIb030qd/MyOkHqO/nExibNhHUHXSACWUvLZdjwWEav6pDe9NUv
r9eRt48kKrkLRqvUj/4Mi0letRtNSzYZKFuAun3qp6OW32IApQw+sPSIjm8t0+V6
IJuh744N7fY2kjIBhdCWpW26+yU9pBHM7M1Bt6sL52zZIcW0TOpnZFihuTgHdpGY
i1GeMg4gseyy04aI99vSKgl652cib9jK3D41/iERgy46Auhd9pv9QdiXvDNs5iUp
qDecEi6p2hDTb7mLWdIp8y2lOaaEBWMEaMPUgwwmvp7YtIo2mCpTL8mR7AHeXXz9
BqCQdlxqOM8t/CwT+FKo7uS2YKXaeIjC/WMXVMrvofVqeYtZcsy/fadQ71X84gqQ
OmhivKBu+R5pa+ON22Q27hBRCcfNd19CgUJIGcTH5AsLUyiZtTKfFCOglR/jCj7s
y6r8qyPOPor0CnKhWgT79WguIdOMv47CrzkVQTfLImOCJC+fZUNSYA7hv7HpFpcR
I30Z1ouM8M4Pp1R2RmPspWBb09Ym5N08HgBZ3fPB/Cfm0ytTqeVDO6kIeIVL6R37
CH24knlwAyrDHNAsMaPI7sEZEuldcVDoln9pDza1GIr2PZkbAVnRjbMAOf0qG3Ep
h7ZAmccBKCYpaoAw+S63wKGHaWRcB60fx6ehBAPfFPdG0kLNMg+KCNYEcb82sr+t
UsQbiyKAhqEBeLotZjo6gOWXjFEIz8PqZskFVPGOB3B0K3/p1HQc3piZz6bMN+wt
8r7g2hLPtz1SsmBFeIqNJUN0W+GJzSQABT5YClMNaAGgoJp83vd7dgYqbsFWGR9v
XcFF/mRLWYV8uorgRnbqKiY2lFnm9qauJrwLwXMg/NzqphDpnBinZsCQ6jUM5HJE
eMzN5tSvGNvKK6zs7AdeTUy3p5wUZiN1PTZ3VDEa4gUXrPxJbcV7ANS3XEVdVcUh
TkFU16ujYHBQj5HyTpFNovxOlAV1+Vb/TRzUsz4wPnXOd94Gl6KmFoSULtFM3N+A
H/tmukwohKwruUhn9gD6iFxc8WD9d8CaqcViolZ5+6RePkuomfvyzbIXwMwByxsn
yBzv2Wnp1e44WLrfVux8lroSVjnkXdUfFgoDR1T/29Sds5epEdTA0xbqBGrwHdkj
vSuWMsgO7Fa/Aq+97K1OL1n20m39KENbJ3HMS0QugksNQq6xwRVTAfZ1Pb+Og+FN
Cba8z/bmpp4gS3iOTKSiAu8Rj3lbVwMDbyV5icPL3LsfhTEys7Xj+FEeEkln+vqD
iV+lGR54XuTTQ6UODazl22L6081QOFLSa5GgJ2Adr3Ec2Tn+UuVTnRa1KOLszMgm
RKcQRjILxgjGXPkB4/vsZqeFs0eWAta/JT+zhRzTbCc/UPnhjYQqwvCsm3l2o7dx
fSTBy4lT8SH4TFKEDwjr4jZyjtWLXpTu+LU+7MeQ69niWeh/S0jfk5qNnfNQKHmr
0aF4MiROeMdusVtUTBgjSZh1KWduQFVqOJvrsEj13GHqn/Kg6gv2z7WqRWtYGnUs
kcF+nImfn7K748TCCV9jUQ/HEvHOBNlyLBAyI0bCes10fuaKUuSnSdKQegZrpBLq
Yk+6SsbO7mDWo+nfS6/sINa4qnq3IQYyYPdb5IklDahAmYRqASKz6kUt36CHMc8M
65pXlSUss+U0tgpTy/IyEtfikFipvi0Z5oZnm7XaXJ7YnxKUbJeR6II2ArwJDztW
O3v7mDhKl/qUn90hTyaOsXVeztFj7BybYZMf+0BE8haGE8i/eUgc+RpNB9p8cGey
ZZty4uetTcpJt11qYTMmrW8c+0ne+Ofkcm+Bkr9U9jbgbzLj9ozJ25QjzDjgzVVT
6UnjYWWjq1rPi3sKV9kXgyrGAUohQ0Xw0AfCEzf8hn9mkWeX6fEzBIw4w99nRJJ9
iZyDbfnEncNom2niPsaJ4cAf6R9aUQhxqQnMtUKpbxfOrLx0W6l5XXPXD44LV30p
mmfG3XgJIyQKABbfunVH8zCjkRIiFLhmaR53jPgXhs1P3SpS9nguTeZ7YTOeVXKG
yzOpzrQWiBc+9tlEWhDYuJLgq5FHMCv1rOKROeL2tTmSJkzyMLLgCwPgmw5CNPzy
82RWRWZJkTWmLXoezvmgqEoJkR7xMax7U+xkH3g5rjlcXd0cMdjxhGWiMlvgqknM
59YJbsorNGqrZA1jCuUntolM6g5SYF9RBTgc3pmKXEfhq1XvSblDevyYEsPR1ax2
+xyxGltQfV0IaWD6Pyd361zHZDWiDOfJnhYyoO0ZaFVsBV5pQHTnahIEK43Yhf3U
JE/Y669SVkf7ZFkydeibhFHxscKllx+RkYalZSkLy86aCr/EE9gPYBhz9knowdkc
F9y3x8otFjGpk/YMHVtXKjdr6W0MS4d1I3MwEmLsKcxvfjo1FmekB7r2nA5CyUQJ
Aq3CA8J6MzmtUKLvwMl99cx/DPB20TvPfRgsfqaMh9uMvZCYmywIRuNC6nsqMwqN
D8q09IjivnYBW+RkGsWvCGidVFm5qydMAo6H2NlRA8V6cEuFCDJBq7VRRLjel9sT
YyT8RwxCvc09cu1u+3u3fK7pU7CZfYurck7/n92SLqENz76dwTktTMkjmOlcRk+y
cI6CoWoaWoM7SMUG96BhQx52+8/k0Yc3AOqg+glpKpUyqIIuDVE3OHRFR9rRYd5b
mwJEaLCtDg1L62Znh8okgb9PTrf6+8j6LzhPAbZxLgdO4DF9bk4tiSy/NTm8gIgo
nFxvucaehBLiFjvrWuc+zDoa/dZQoUdPJDIxuqYFnJ6bUiU4ie8C/SoXTGPd02JZ
Mmsd7NRH3TCccgxQYX4Vn9LqijjbXBFBr/FeWuBfM6WUviBC1pf9HgS1z4kWBI16
o2BT97WnWsAvPdAfeYAaClM/vozRDjhU3TtMlcsiTisg93MWfjxLt87R3QCxfhQb
2NPctqPVNCIDtwonNMigN/P5HehsXcZhOuHBXEKJOfMMv1Gwt/m4DJED83xPk+N0
i/cxdx3Iy+bOFuYyWBCiaaXVzFSaZzl2ai7fGbp/lYyKR7jhinu3ZUhSUNujdEnq
nsTx0uOpLZvg40jSDR1ISAnfJUKs1Q4bCVS0H2mZiQvoTtU+v09fTWoL3wdonwE7
zKF6f/xbJ98Bk7OOmWPJl6f6v0Cn1GvQW8jr5F7VazyY3dQTR0lFDSW3NoR2ItVN
ZlWQjLfwBuwAwC0SD1j67n+fTxoV4AbSnKwGe+ZcpxPrjAP85k1KDZl7Uzrv1eQb
/GjLbG98imktOg1GyK5jJqg/YvD2v9hLmqJgB9kDApQpFtjZTkdfz6TUpjPaH2I0
znsy0eDyYr+FjHuNZTe8io3a3Bt6XEX7xndNctgiWMhVOUtes/aTs5QACOVemEST
ojvkjkgG3g7GTyveTcupKQ==
`protect end_protected
