-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ZS/nlDQBZ+uW5WtspfPqCTB0nnvsqMI4zUILKc+fG5ThB0gj/A8FLHBkYgRThFHeNLAWloHwPLQ6
ays8cFHzGAwDldjMdOHN7ij4OES4aZO0sLzO7peaDgzpZO1RTGFoU1Iktkz3SVFT7/937x6wMAnK
kE0QfQ/YJr4zxAN4kTdXh/FOUQewIagwce32TH/L2qSMAlT++5mGlo7L20MWpNxpVy55UFSlpXEc
e2jXihb1P8Oe3NWZdg49XK0mhm7Gtpcn/6/S3FE+btCm5VzYELRbetgX8D4aWIB39BCipPRXYVDy
GuasvF5TMgp0BD+7xTJyKXBH5S1of4+LW+z8MA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12096)
`protect data_block
2EkEbVJn/SzxmWdzJfsJrTIvzIeq7vSWb/j8GbnhXRRMCN6DbcR453VoTLvNdY52HZeml5iUad6U
R8OWhcm7pa3iWPMJWbrN87YpOiJJxkhLjtWwADMNlJPjQM8pyOeTV9fvkJPewP2EtxsBXpG5e/lL
Hq/r+VSReWLWOk8OzS8HC6mJkFuKNI0X99DAwYCpjWwLPbnqay9hgcZ/H/yo2K6pVRHtlJ7DIbB8
GLVfyOOeNQn3UnwtDuSY1GqEQ0lZ5/6/EBEl/1u+zzK6DEGGNXA2fjX3VWuBuvR8dauREy7PEI9d
9aSW3uSdGccnOtacEATFnlqW1ie1SFEAyavTs7wKhCz9z5f60gUKg8oitV0eBo1myYAsAW2BZJQp
WPOzMrMsVBz7OaAIzuci8wixMyhtMLv0s1Z664eRxbQ+tfRzAQ+BFNiy7ivo+ECvu1yhLBNWPvk1
jYofcb68MxYWRz7xQYkYwaQpxuJDMqrSaeUHnXA0FGkLzYiTouij4aFhDubq24KvPNk4TOwH8rtR
5g7ozkhAPyR/RWSUg8t9RIxnjhZx6P7T/RPGBBIbkmFON241Vmh1627kaXYmXoQeBvhel4X94fje
lQAYe+wy0Wzq80wXx5qroXKtV1JE1axhGdb2ETwYz/hSngRHr/HpD1a0cY4FS48hl+ZAdiv6hNKk
WFPb9kueUd3Xpx1d+KllYoghTI4oHcf1RQ9AgxCcl9gtCFxdmMYLk3DVGFRKOo9gCqpdBThekxid
B2CfOo4MAm9w0H2kAxpswK1fB8WXQQPdPcipp2REUFLJTFq/U/WfCl2jReViOfNo6joPG20DU/J1
1BnNRwrNeRtjtRmijC+N3ATMDBIbeW0xymDtVVhmZo2WmCg+RHhbLPIvGSr/GqrZt/CBit1oly1C
05rSu9TXvKBhgtoZUOY70huHQjTmkAhSAvA69BsIv6fVVig4PoUWvu01Nb3rQWD8khass7fuWxBK
rfN431FzZDfDU52tmpAGOr8A8MbktJmWAAuZ5N6MYAvmhev79ECaAUXEoSN3qJgj1QpK9tGjm4W5
3JpTUZc94QfKXC0TK0TUT5VQfAueyeq8qUL+5H4BF4WjBvGUbCiQehME4GMAnPUMDdYCqEfRCiGg
nxtnSM8YwSZjPjVHWAJwdgxCkr71j9m8OpdtvEaCbIR5wfqNPr2vD6soc1oRhVNiKhJghLRLAlzP
OVTWq3WXw4aCMbAGAdeXvMaDNVvRgqTYqSigonvgSC43qVD5Kb3eyDmgASvqJpbvlE/xQdehWihr
5uBUSrVc4n0AHVMHENmNBcyhts+wNJIUY5e0JFsQ8BPQ697bLF0ZRnwwVGH+tL52td2d4qTrdyR6
JuMDKYLn6xhg64/jmrLz/3V8uge4sMlA2mPf+ugW4wrfkdMbSONyjW1ef+HCrQvFQXpfO40EJmid
zax1EP0H6wxRFzD85Tl+rLcDDnTlTdfAXrYB+jdcT9leEX7hCT7JFcrMrl2kePOWX9LKWnEJOgEK
g/lbPgB+KCv985/ekulc9iZ2ae/AlUEN8j12KepzCnD0p1wVVageVTd2mUBtBZSOHRUG2l3k1S6z
eIiSEolJe7l2hrvuju1F6+qj8MvhpKlzz0gp/IdSjKrJVsHARssz2rVKflevFYcmWZ/EgJR0sUO0
1CY4Zy2JL4lgeexzEniRLR4bAr+4d15iKNDLvhZWp8BUTxk9yGX4b4ptUBbQNsjNNj9B426F7dzK
BXrDlSVrXUERyqPerXzjGodiW3OwVevPJc6C5iW1t94i3iOcMpdkI7tbcg4ZoMNUtKwKAEZpiCgL
NG7hvC0U5Nuk9kTRJgPEuixWCWgI86CqJVgHr/6nKHRg4psJ6Cn4wqStQW8ZngVnWC9Ran2FVlgd
CO0v6GuUYiq4Fs9jAsip6CDEQvOetmUKc7pVfjLQH61PRse0R6JpXKAx7/1O+B/Oa7ZwMK6ns1WQ
lg93mf19wLKXB0RqyCej+7o3ycfTj8kz/Szg+D+gsADGLR0qUpVqaEIidm0dRVxSO02INcGKqh3X
TQ1dMD0uoQkcxUzukFK9PaOSR+tstCNnq1HNW0gwEfHu+vZfnySRkb9XfeyK1JimoTXJ9tPQv7jz
D7490XGS+PehZ1ebDpDw3xjmg6WTJYps7Rq61lPar9PwLlet6MHtmpgpKYAhmhVMFkdDH4SttOYh
+AwQ30tREBLDoyz3BKIJnoR+dbVHqBjC364/4tCadIzVh7cnK29n1bziNX1uiOWPJiWdTUbWOwVd
ZHPgoqilLIXD9iVO2ji2eF4xb2shukhtDYwgQaRRW6kxqYRsrBMRpaFA/n2G1R7wF1DmklbULPuG
WCq6vRJj/S4hhwUDu7o2DBcMHpGSsjeJoTJ2GKYNpa7FQ9M8WbVeo+pmdPkVFGeP+b2ndi34wwH9
J67h6bKiLmg3YoqHW/Vw2F3v7H3oNasICO143T8cdxpBOCFmCFXQbERd+eQMgov+oikTN8aR0o2f
T8wz6G6qkeitAkWLk0x9TVC4C6X7k+12GaIbenbKawNH1Y1lhC6ci96RGfCc4EMKvdNaFbEUCBJy
Ruy+XKRzjFYBXAZyrfabohByPJi6BtW2EVFn1t0tn2LWh1ErRV9yi7vYp8jE0m3YtuaH1lFuE4GF
Qc3OvHiWk9WKPmPcD8yp8owLGqz0dN2D+LSQ/lg+6MREXIUHl08VlJvxWUU/Jp9juwRvAS+GWeFs
W9raizRBL7ETRp9j/oivA5ndOsCaEaE3LljYvUxCSW/2ypiTVDIzZXQPnb7daiIIDKjQ0USOZ+sq
/zCqBaw0zJTfEuNj36OY4bxxnvLrsK4cwFli7XxO9U2XEStAGhmtgqZglDSV8GtscM7N4Rgiuxsv
sKbs2lmxOkCncbv2xlP07cbyVBwO1at+OsZ8lRzk4f5u/8Kucj0FeBudxk1SQzTB29YLDaiRjOVe
2XE6hg2apB+tpo3/XoUplBGQTqRVI2g1a2oMEDiLRzlQUe7X2At0GL/cI2k1AgyS5ls+lZBbrMlX
VUf+bAigf4ArFT/foTkr3BNVi3WILv35Drwo0PTNO7SnMJs4UKAlaR+FJ4fb+Hpw/hYHd4EbGodM
XbsiGdknXrSon47dscq9tHn/xmWvMVhM4KlxN7RnRNSJ7ivqVFseA8sCRpoLjTtyFTg6JjFZ39PM
wbtPw4KXAYkrqEkJPWxmZ+phQ7MFpB0x7/sNVwCPQobSoblGv0IoBaXBSzzg9ThJ2ga35j6LNO9q
vS4qrBdXYB+Y8yiGePEO40sUthar4RxEH/XRUPth9uZAzcGv+ALQ/yBpcEWlrrQX1CJnem4ly7a4
fARukwgzSDv9pjTj2pyUHFOoQS1aNRAeqqi/3ob6f63ISCuT8jh6NCtMQ61KDcVzwwrTOsQwnp5x
u5Kzd2ZbIKp7UQS2WbIuH0jMArR4wmlIpmlUQYJc/QlsPPW7RGDii2ez34UTTIAYlS0LAE32L6eK
II4iUFQMGj5KXWTp97vv0tQWgczenxlTWD7dqxriDjsxxZnzBXuZuxQASkBoG1L4mRPecz+O5NAJ
Di59/MoQz9kr8l1Mhm7OvAk5BvnUffOJM8Ab6UDXt3ap1hMWctK/ELCJaKGLCTyOvS9P4nZCfFqC
e3xFRaGgOLO4VJ4pk+edhoLkqHSlFkPZOtKlyNdTt8H+IvDSWgNn2XrOr/kRFsdGPTpf0U17z2rx
UBCJEE1yd7p01AzP79FUiXvR3vzqccAywv7CuwvkvpxYMTX7zBGkSp2ufAjhsqiGX8Zv509yNCwa
HSL0zwef1SfSYUjowtd2FfcQWebDn/vKH7R6qBYvwW40ayTrbCI+PQ+oGjmJunVVhtzJMoD5jAi9
rl/IGqV8JojG8kF2Yl+FbErngDLGq2iISxRO7DA72ROD5JTHrs9KY1WDrvbdhxAENyp2/CwIrGJs
SOqiAShBKopN/sG9iR1luzCdWPF714CJjFzBslAt1d0YSCTMihtGPdEHKKtkHxNoxfL9ObYvufgD
HZDHZQrM69D0LKn6ZOp02G96p/gJw8DLA9jheKp7ZOkfp5kO/kMPITb8IN3Pzh+V6qs6rxcQTAyD
9+2Y2J2T6/RNv4NlyuTrQF2/qsYslY3JvnNQ0BdGlgdLVXOhq/3QkzJ2fXyUIrsJNDETxu7KiclG
cOG4Z7l7dndKVTWoX/BYjAhbMXWat/aIqQf7oHdJluorit3Dibw3XrFblNhQL31PvzoiTj7b3Fso
qZzgTjsM+BnfTHiO923Tj4wXoviGfWtq6q1bjCxiUFrb6QrFPGXd0wcuSPLcJiJMtQaU0b8LNqHK
EXwQW2SIIkos8jkNudVLn/LEAwffs9iC+ys+20dLvn4r/z21iEqKj4lohAVaUDp3+mqAogiS2YV3
yMzzVeOnF4iIfsV/N1RVzBpaMdv0MOJyzWvYQjxOo2AtkSyq3KJ7eKeiVrHkJHu/BA4nkWIHRq31
uPj3aHGgnIYcM8tcETfglPFnQuEgUsE+ebFEu6UpbPPkoJ2hfF708DT2WhpeFBJCiPW7ZqLJ19f3
j/zohM2OQs8dCOdeHvARF778afxIPjAvYhyj6E/SbBYxnGTTW5bKSchcalEk+RNbrYqZQ5qjLLKs
D4tesmWp7mZ7K2JmARgl2824iTF47F+pHimgj3Qas7dy2hRz1GkKUMrbacLAkxL8khaVGgfnbyB4
Yrxq4RbD2VOYIc+SPXsKnoJ1wJguqp7d5WdRi5/FYFiC4Shw6+ikRQKckHGTxiJQ3joGGbnObAAb
9KlR+zh+Mv9MtbwJTuw9HG9l7Ra5v3U99P7iqDu+8BghoasGXa0OLZdxGbcIsGJoHn+1q2RIlZXC
oH+fAxTX+cRBYWYcE5YYxHRUm5Pb4SwRQr856tN7UY20nNMFHRuLBX/dv1xBDyVOIOVvovHPEryh
nQus/mnwLApxuUCapeE+igwLT53DVBIYsijg7C+/36YebTZk1KCAdHJgPcMqcK+CurJuUh4kLvSF
2vn+GN3K6Shxo9QT1omJ/awPk8C+Yt5WNJrEBLQHpTJVIbys9X47m3wiFv9b4mWv7jwkjsx2rk42
t5QrjLgwm9mQ9ZcIhCMDscZJC7bJo4T6C/A4yNQ1pg44HIc0ghx3AqSjzvq4aOXEBZZ1G+8jW0b6
URhgsrvK9dq8cdjI8HMhC4Sli8VIS51xj0sFVZKlGzZ4HL9kGonzBQ8t4mw+rzaNpWEar9tKKR4K
hpfm2DZ4kNN4H7lQon/ga2hmAoJQzMSuWFWMfhqXKyTObZEeRwDDGxSHpnCQfvjT85xsDmX9vGBK
SAEatVObRQdJW1F/gfGosklpdp8PFx4l75kcOuXc7Yj6RZXuI0CWDGTzgcv7ELSVIHPStJePX8wo
Rxc3oCiLR5pZXI7FXdzQ+exzCHLGyjtxp7BVQJAob5D6akaj/9T6qowrBZXovTMxkFhdHgwWFnCx
buFpKlyoRiCGZqfxBP1vXdAxVOA8dHcNg7KOuDrlCu5B9kAIj9CQtKpgRICzKMVYa2pLtL/aJ+DB
2MdEUmxl56ZZ8ykQx4G/nrWuOP9FD9Ajv+EAv8RXxpG0mgFVKtwDk8xtJYw4dd84d0G3IX8woGjQ
PYoXbvDFGrDaJEFjv3prRSkdNzAdXMpyzlOsC+j/79wxzAG+UQvjo19V/DhDp2LT7t9lLni/FoiK
8RUt+6fNFfB8Lj1hLm79YFenPkJjR8UQazw5xlGINsZeQlTNm3GIdMZdfZzaRxcHilIjtIqUrRSo
SKFpoD0TPHjpWiG+3/seZYJ7AB366GMWG02j7rlQiZOEYfowTQxExsDlnKGB8BNqJO3W+Qj/BMYD
wC/VRCuB8FdFErMX+SiQI99oWl8dF0QOB0fWP7/vw6qDIio+eN1KyNsb0bjRa5RXoHCKbpKNK9V9
ae5+4hNxOag1AbO5/UdLVgr5vhxsvqOclcS4CUemeQEzJ6Ef5maIH3OgedOtbkIhAKSv7GKmA9tQ
SnzQnLVyGWxmj9AHzAGWTRoQYQjxfG1/kmfFSRzYs/QNF8awr6GchDqZYMmutr6UyHDzDiyGSbfB
ncOo7LHKzXKU3cRVxlmRds4iSf+4aEtisZh3r8I04w8dI5nsbmzKdX8AQV3sHyEpcnxZyaZiOcVP
aEaoh/dfps6IaykBibP2UdCcNvWyQuwchBQfDvyfdt9izqVUX2G4cfff+sEjmUB+vBqS2Uxxn7mO
BzE2y2A6WbsvjID1T6eUIltOMvwDbaFUaCt082uHWC49AOCaQOip/lZtqhmIId605+wtSdCoZsrg
5S0z3KyG3YFIT0PSYUZExgLObD6VPOvVkPPbRbHAByMLqlhtQ+b+qvsGSWZXr2+HLbMche0mT0Xl
gODgq/uxyUQDRzSIRS6U5G7CZn4B2Ln2goIrAMd4NW5L50e2d52Mei13V7OuC7FMHZ2mclnNauiT
3YY2dEffN+GuxtZsl0j5u/MhPjW/2L++1YhjXUMYO3KMW82t+PzeIpAfC6tAiLOP3ZtaDoyOABHB
YRvkh9IU+0mXeWrbTbIfbQ4sNqNMpSsKyis7L72iS3zpeUBkddDYxoKs3nOQ/xA/M0skF5Fq6OH1
PX4bTiBHHlTWdqTUlS4xElNvU0Dken9zvalEYg6asaDRm/98rEQzBjrIezhRqBGyF80czY2Y2LyI
IIbP3qSt8HBs+eGY/0t6ckslgq/uiN1KUKQajE5H5F+ib/dvFuMyWr6MdGAoXI/Rc4Q36trAzlAr
9S1hbITQmVoHWKvHX9RBzFvS+sYvAee7S1V4ae7qAVZ3YNMGAuGFBppNwf2eLD+UwfqcVTkhphoy
v7QuYkiU/8TCJ2Skk46Gro+MW1kRI7Zz8x3wQ/6z5Nk7oEhOPe4qD7ksm3a88GHDDKFrt+/PukBF
HgHTiSeug/vqRloObkMP33IYtqZeP91afr+7QOgnfDkiJwZrBB+rIxFn0FPwegLMNFGi9tin+9kR
/3eMLCyRRDBODaR8BCaN0/1f12HVCbRdfk0gx6vNmfPvZ9W7K+2uUvrjRED46z5dphLyN6kLdHVg
DMZHEqB/Xs87Tk/tNQ7BzsMBK+tv1FGv2RpMY5XPrwbLBOIPx5cz2t+kzpEbT3eaXVPHXp7S2V2+
90KG5SAzDYTOOIXRTSJXZywXjgJ6ydfcCZThBlmJpJAvb26IcjjeKKhrhSM7KX3LDG9tYu+coyHr
XDP06RdSooK2vcAr27zzj8xKtRqUdrYq/uKs/JYro9dMH1Xi6f7RlOSXy7w5YGH9vqgPMXQ/x7x0
FfaPd9o7U/Ofq+VsSHmmC7faWcxKPohtXyCY4xetSpozQazlE8AKcpUG+d7xPep9wrXOpatHKd7z
G+YxsEojBrzhY7gS5rX9jYK7w0EO8WZlndYBxUtEWtoGulv3ShW+yjscTZXnOLuEkk4lgZvIpM4F
vASLuujrvT4gG5uAmf291cCO6wUrlXhFaKY/sp6gyp78sSIbAREzK3ziVYtJOWC6lsc9KYg9jNm5
lX6yZR76dfRw99nRBvQR09XQXLFxM67rib4mWn618Y+KKnp6S+pGYjHYrXvVSBTHl9zu2F6vVc9D
Q5RRujMJs5SUnMw5JMaZGa5ItdTDbQDJpl1q0g9tNvOcGUioZS8d4ok+cLEy4SKETg5lCbNgqzRG
EyvWW8oGgcGVOaisW/pnw7B914MG+LIsh+OeUNMqnY3370JQVYRUqftjOMXX+mm27yse4iP2iiFe
3Y8Togvff8qzjf8wc0lLkj1zuhzlr1bt36TjSphbirbuhZYLRi055SAT1q396673j5jnM2kduPlS
ciwam3Ox8cjYNFrW7hKGueAsdfJB3HBlJO4iQWlxisar1x5v2CvhD3N7F+1lK8QfP9IOtT332fQj
GqWiQKxnFSEGSyn0ps6vsS0kCwyxW7I5Y2eKtUBMJL2aTBIovAMtEsNTpKTMMEoR2OU3qbqNnNQT
Oqlo8/TR+9zKyGxAw1xVnMw4esSOS6HAofXkm67XEqplOaVwxTlid+/V6j/0lJvOkg2f93wczTfk
fdLP8ggtQlIVIj+/uBdqnckB8/mPD4KzDOB3g4qlFARB7FVgQ5l1IR22bzBZ3XHR5ADfzG95Jk2S
1SmkDldtncZpWj6G5CTbPuI8HM60iJgYOwhTJkHuVGpNzSj4J1LUGoo1HzL1gR23d3Cy0s/LArgh
thUpbcdasAeIIo35h7Hyk4NF8OtU+/UViY5FRKyp0RSrUmbb1PCWoMXRczyFHHrjdeeLjH9+laRA
EurhoZLvDl2p1au78bvITmiDYIhhaKdJRahXbJpLGAjHMrl+RZroFgKCPDLNEqYlMDxDKjEsHhjK
NVmYpzR7Wlb/5E4fvXfh0H5FVWQ9NVQMPVDasx9qfj3TxXmakt8xVC0ckwzMCxvfHrT8UD4E1B1A
zHF9FgWQzIgpWX/2CvF8f7GaSyxcBPR5f0nm3K3fmPJ0Hzy/hgv/K0u3NWBM4uCg/1sYLlerr04+
0xtYaksQmRBSTjDb0M0pBYz7UdKnvIzVhr6xeQN4iNrNW6sfJ+t+Nq0QGE91OUx4ZSowBIK+Wo4K
l4AUxG++E5nlLO4uFaDWAsu/izR68XQRZvINODsZVC+i+HOE8wbjV2T+WMsDWYKYk8YtQ3RxXkwq
sKA3jlYLfLaZbx2FyotRFJV/wZMfVViaG0fWsHYXaE4bTpsS4fb0qbPXz4xHodaT1YX7Toa/lo80
V7NeqfgQt72Ud1tu5lNhbj9rIaX2uDg6BTarBRwAOuQ5TbAK/k/dwieCMEjeOjRALKEvUksGYRVK
QfbxvrFtiSGimgiKUy3SQHHDdN19Kjidr4qqdYbpYZ2pSoDm3tw2DnC42QnnmxM6qEHgsqJKLBba
kpUJNZLKABjxWot6x8Jxgx2TpWhV36nzZ7YKauOR3VN64q1JvgLiin0sPU2T2UHdxG1iFoZ36Rrc
7cYm6MncisrNImOex5jDM0SRSha3eMFvhIbmq64KDVwzGA5tHBvzMNTD70peyqjRGF8MLzR8roiu
zy8hW83UUZNSTyoSBuqiSd/deuh0S5aoNPj1DB4Ab8BO0cBF5OzKW9pya65BCEM8Z7fSDr+spxcf
IVk/h7gtabXW00bpD3X8YN6Rxb4oi7ej8EKn/X+TwmFW3M3pGPBsl9yekC413pVb/n4WhxUEviWZ
JTIVeXPaGAQboNMT/BaAVdeUlD1h8E1i6k6X3ycBZsEqSlTAWgqRGZPfESxvf0SW3ZltajWenU58
TGmr0LvxCmmFCDIGrof4oH8RPuXfdH86fZc6zwLJtPEKSVKgEgVFwVyUkN1liTOcDnUZeyLxrXSP
udz51woFgIk2XYdg7nJeJVWr0cE+uTXbineXM6tlNMTaPaEcGdRd6XK6udD8lII2xqrNOc5VRkcj
W64bhWd312BrxZs1qeqYGeP6dwvm4ezP+Iq9obSTdqX0YZ+3STH8YGMv0Ahm1XAyBYAdctzK06pQ
KLfIealuNaqas2G9XmQ0POU3IF+up02JO3WgZh5nj31KrQycylIs9y6sgOM61pJJY2/V6JwyRiyx
WoBzm9vv4se0e0zvevNqptczutPAQPetd0m+pa8YjNmPX+xuPpwX2DvaKtt19mzWE7EyqXc7qxvU
VV1SMTwtnVd8XhSFHV+EgLyKfhw1sM8BKMM230ecrkHCZapSQRYqIuqyyRqRo01nyciZzlNmTd1b
+SjrW067dEYbPzD+PJRNO2kYgDNi+sHdwG7yYc+AIWWN3IxxUo4YD9WUtU5ntHD6GoBqn6Eh2F0f
CPfRVqqOR9iLGQ9a4Hd0I0VUSehdBs0Uk3J26ullb0puTlJ5ds+gOKGt7uwBrvIh5+Oa6H/e69FG
4/9+ZBpRgiz0vyLBxskrxhZg/f7qEGFeh0AHrrbLSkVQ9s7fn/LoyEqZ4pmCjjYFSkb0kC+ote7F
MGQ07fWo5tfeXvT10aS/0D4XbzvhdZxnl/MEiZosb5FEWsjYOw2mMhx9efqjTMRL8NpZMdU9vJtG
VW9fOI7594ql12thumXc8oMw9pN0aJhatoxl7UJqsVcJ89l0i0C+NHM53dCTbGN2q0nL9tfhbSWq
JZ2AxrDmUE8rVBuoDj23y/itX6qdznTipJF9+oSy4YMWtrtv6pUMxoZDLa2njyqKYrQL69bGBmaI
pmiHycbejaZyOPLbBi1E/9r7bXLSF6zpYu2WxWw4LuIS413u9u4T3XTswZLPn8BJGIsY24k9RVPb
EUTTLJNxW4Ga/iWaCleSvqaTufw+liWkaPBTOAMS0LROJImoTF7rJAe679FyymxWgDcdHtBw9W+N
E+7Y0dGLnffzxj7hGxVRaSqsp7iRWBsYVyCIEudVUC44F5qaBkHiqNwLdQwfObqNKtvZYKSabr2a
G3z330DfvTK4L0cVP+sNvwr6ozM1pEGDYs9dqptrkrTnuoAA0tV44AickK30lR6uYnH1aodBJ6DP
bhh7GFlvP0SFPbyCnCkhbDsM+f5PFuaUiBhVZ/kZZvYy5E1s659HlDWhmRlyLA47yYs8apDiQ5WK
jyO/SEhAogN0ATMbn5QzV4WbWnqSIA2RW6mXeZ7TmiBKwxSj0xCO6fY66q1ULazUDYSmVrYSoc1a
nB9ynnhuVWj43nojZOmd3c8IevH3piTJLEDc5Qf3KKVKOWFJBMTv7GJorDrcbKltlk0ZjYHabFSf
mPVwck6bWXr+M78fwJJHwXENgTMDDUm2PU4uemYP/S25m9xJDVtywvHnwq+CjrIXdbcSsh3l3JH0
1W9dlgqHaS4yzHjjN8mWq/dX8GnpBQrx+hcGRevOb6+VyPuNJSb4wfOCyFn7bUuNCZiEUthz/YE/
BYB2TAKvaTTtpAFt5eOj957YRvF4CN45mlyJrM8pPTcrTzjOnZzuA3PDKavNgvskDFTv4n2ua7FO
FqmhiuLlzTCh0hMw9mrbNFKmEWPAUiQW0k6vlCPbUJAOwb60gEBo/Ejs2nE5IhvzaqELfoQigTkY
CnOz1Ezh6A+jgdaxmnFsB4y3ObcTfhWVzGiyxDtDasiPpKURhiOSu2xedeSpiUcjXKoc1NhdJNET
R50ZsZaMFNmBftKM1g6nSwT3vjMzkMYJG6m8Feikn/ZTzIpD9SHU48Mn1PoTqdMoVHrmydpohTH0
bHuv7Y7SC3Iwp25TvNCsakwqxKiFMfGGSsLPBBSqW6UCe7MxUIMymi4fMKXHJDB4d8QDA9lkqFlE
Mb6VsYN6UH8Wlh587brFvY8P+bohMe/1zGkjAoP4ly3MHq2Zn0YRc4zPt6n9y+y4zRucNXc3NQ6F
ZpjfQF98ulEfWu7p8n60AUgenmeB3/4yCQeO3MN/+kiZPRcC+eshAWeXLmDJwdSnsmiEie5Gar1v
DHT+xczc7RJbedoXbyS5CurkAMh5rUiGUA+c6AsUhcK4px080qRerddxZMv9hnJQAhmOh2r/T8wW
uO+4XOYF89WxB+fv5nFbDoEqo5dFMSEKyHcu3Y0ZxpodQD1YX7ogyan4disjWieZac1uQJbNfjn9
zrGg/2vZwVZb9q6ZLRXPir1aylr4yLU4emktX2mYdSs4oTGPsHIV+GJoDSnRaE73/bqy5LuB5Y9Y
6XkOhBwGaMopM1gwJxSMka+oZLpf53edXYBKouMtq4B2jytJlgGqDGXvC8ZthXo0j24E6V1wu1x5
ak8DxIvFj1Seqv547yvlMaW4uIxqdbAwAwEYuMHAt4fTMSxMh8EiyguGCl4b750ObQhlIi8e/nKq
CGCpp3afQnc9Ltv60h8H+3Yl068HNfQPjbQebTVqiUx9S+q7lHtxcA5pnZa3BRG9AzQGtzhGAXN+
LHpcR1Y2JS7BlMDGmYUNtnGmHEcOQmcvl1iLkatx7AODHOi7eJ9s65nUo0Rdj7y/Uxbkk0w7Iaqj
AkrGGePQqEH2+EkaOGO3FWY4fTFKSDXu+mt5QaOL7AqZG9dvn0Ov4T7eKmpSJ79RXmt5ivLsodMj
P7IGcZCRigqPKkVINiNVKtormrgy8u08qI549KRcfmrez+zNSVC1qHJaFIubDfvdXoUekfpbRulP
Ruh3PkulK3Iq3lcz8nvh1w4a7mTKDKzvrtqXbfomm2s6seVd+KFS9aS+oTaTQ0BPtCO+lHOCwv4P
aQlSBeP5kxLRIhI57rmBunT+e0bQujBvY/2eo1pDmC/lGhp6rWWAoo7sz+i3vUYzgf2ptgG1ovjU
EhKLGN8gu9znrX94RdnGDAh2v4KemNrTV/dOJpevanpk4ebqMuEvNl/7BcZQIkQKhnoLEhvWIBxA
Lao/yKL6TsH5zq9sdH9c2YyXqXKHb+GYIBZxBcxWcUR2wiUlVGnN2QgkXunNzL8qNdZRsTaqqR1L
zJXb1/bq0lJKl1PYEDw9cqeqlWk3ezCBEnAlykSUPcLi8W1bnuEI8gOpNou7jBcgAOwZfbFPlee8
wnph93VjUe1MwHQBb+4Clhi2kH3Irn8wZO3Lw+gkz7PHrEXsckVevRTR6RwdlUincGxi7Z7xO+n4
8wTMtppQL4r+yWzV+CjfN5z/uT8pckuvgJHLKRsCxsb4y4Oyy0kHtA4TAZYQwgE6CjIXOD/wGpkb
/7omf/jc7ckB/e4VhndKYFqVp6KhZmKQMuqP8hRMfW7+czXFf7OznaaZae+gk0vk7ZQwdrqAbe1a
+M1uNvyJCtBqD6Nuc1+rdzk4frKUMFGd2dgMzI99LWpb+xyZwsthGGqnY7X/AFuA+2fzb12Sd2H+
aqsfXBlJRZVE+Yfn15cMinfEcP26LN5Gvp595aZ737bFpwxWwW27OTvklDJLTsVtYUUsrDExkqFv
6+0im8UHiP5dv4bul8H9MowQXQYrVGHT2xoIX/eq9N87T8O8GxBQTHqBzA3+FEVlc90AZsYhMXli
0c3G+DZK1PYklMElm4bSMiSPxOt+Dz6IJ6Tge/6jrVglWIQ5AuMYVrgzso6fG187Mzj1h/KoPTWE
7AVBTEK5V3heqYMrZt1+ECZ85PsFwapBV/AyAxpJOCE6rRPcn/mooNNakuNGjgwawnDAQyUNd+Kt
ga2KVZ8Wl/hBGuIS1+YFfKkEv55mhc5TsuxdrUKDwEXCimPdIk2JXp99g+J0EBpRBPFWrvXVu1/i
H8nrrQGbzlo3SSrO9564CT8x6NiLAW5cHy6sRlA6f5PtkYkdRD8zCrWXQ8gE5tRfYyW7kwgZkkCT
myCUDgQ7h8zrKQHttqConRyZNCKh7i4frsQeruTGS8RMw1OEc0XE2nvqV+T09nv9+N6cfEj07/UI
Ox4HQtKCTJyohyxmkWfFkE+j2bxDKCSgmP9zTR1BDTMDy/9LD5UWqNWGMjXhmh+bUC/du3WnZCGU
X21FWlv3nPkNA4b4RyJSLxs5Xhw2QifqPt2UnIZlQ4AtWdOPIndQud87Hl2HaWOluiu5HJfGjlwc
3PnR8R3HtF8J+fOFl/SMIoVFN32utOEp+iApZ1waQj/pFjhsbNqjdn3hOrw3NlyyXfe723pmr+mq
hA/O1TVrYhhvcRNzmzTOM3cprqPDLRXLgsM/Ehfa2D26rIRK5MG8fRNMHmv56BR3ERPZdNQiS/Up
NzlqYyMIXoYLL0H9cUbgPo8vgraS2Vq7m6Gu6ka+MsGGbhZsgCRU2Go3bM//uSbA18T9SKhXZbG+
rkq5Kq1i6UlsDA7vBaPi2saDfmdiM6y0txVqHNAn2iG7uK3pfU2nLYMHP/llGO21BnQulTTDXPqa
XQjfmHx9/ZrfLkm/iCY7UW7Jthr4+Ma97wV8SIgJR7tBYASBw2F0sycSUu/o5FMjYzwp1JTA4hh3
vtecWLKgbfNKAWQxbBzSO6+2LJXNGn57WA9uBrV7K+5++FJQFflRUfa3ASPWij2zEIuihIZvrOrX
StyE9FE/MPJSjjePny+t3dgOmijgRICnWLCrak0e4A4BGPFytr78MHXCQKyQ4HS4ai2sdif7vwLC
Z3Jc4V34t+4igtuEPRvGIYGhx1aL6I+nOHR7rAB0ibtvwhRj7WFlkkEdO2URbbyze4JaAQOW2RkG
5HE5wQbcMnkQ1CMAzlNPx5zyVc6DYOUqE/sIRTpYandHYilGH37BeL4b+KQVfl82wDI2ctMKwAy3
OygFxLdeCTAIQCOm148ITR6J/xhedRm/zOFCBezoDcCebFsLMktjV0SaO4//8CY2TPodnJoK0Fnt
E+18eATjHtQ0BFf7ldEUBJA9SjJtMis/dikADuUDejqTGz3uU5KZM8juI1r6LBx5saQ1d7Sh8N23
5J/YHFtZjgybjsdkGfexivs2aM5ugWstfVaAy9q688rQn1UchmSeb7jMJZtBLRzNERzwpXxGYV/P
jiFetA6ex4CRXE+wRXgQO1kqrrMyhSxd15w2iw1vs1e/plAEebgZibZOmCQcJJfjt7A86M1A1n7C
xR5279Ss2MWA7GSqrH1yIsrl4ejnveaYN7I94VRPc291V9NzMo38+dXu76IKVMscwMaYcM8QI51I
kmEV/fIzvrs6EcTqdJMriaEI7Vz3p/32bxcSsZEnXcuFwSf0/KuR3UuqPgCNImIieMKGJ3+Z3HpH
zsUN3aRKA/oTYmwEjLc7Vp/LvEUB2FFqHMqeT8Br8H2iJvTRrwzo4Wyu4o2p9GwyurOa+v/a7kNS
SKXCdqSDEEeqGoj1y7gNxiraElJHOufUF1AWdwZeL0fOkR8svRpKe64ZZoBXGIXtSXJJwTMQbsqr
jQ8M5rbT+Xbp53P8m+N1zX5+AZpssmkbrn/0x24vD2nVmHohzSVDSZzyLIvFmEJJTh+DupzGybVi
CTQ4Ajsm5sezKIdZWIC3YRiNpq0ImtGL1ZeqEdMBxIR9dFNyIjVaVyDFgY+NNundQdavZa8jKY65
UHqkwglxRM1iDhk/eayHE4cdcJhw6P6BjdwV66wQ8s2PcBCyWXid27R8FPuBnpqNLCe2qZSqdJmk
X0PqgfS2RP1Gq2ygadaDvaUu+BfyP2oCIADIVJ8f5OmuMkfiI9AP4/hnVfkrkjWBqxj5JAaxsXn5
lJwS6/BJUn9o64luHegsaIQY41jBSp6rlFL6ePc8489L7S4ThbI06hnxhCE2RMLvbm3AjXPztbqU
MApwkKVjNFmtHRoD6U7RyqckQPQYtkR6FpSyzC1mqHdLF4eUwRZ7As4MBOO+T6F/CIQxcSTtw1c9
zcOK9spqB+aK/aiBm+jU5F6cRHgsB5HksvFA7CS7A4kbbs0D2HK8ex8xv4Q4S/RHtoFI3/cJCnJt
tw4zgKzuCyVXIrzhO6HUezoyes97SRB+6rXxYaaEdTFzuLEhN6dm/stx35xlb9hMkiacdrbz9ix2
Hkk7xxjhoC2LCGkZlSB98qDGXDL9YJdE+US8WXDbEhdTg7+Ua1V9OvD4sHfjC5CRpUVYqAVzj1sG
RSFyp9lgTrC0pPNvjcK6kdYticQZDRjP/bW8HrzwG70UaDbcrPFVyJWol4p9BlKms8Y8YRVEoYXR
gWooM+IDkQ9pAEX3HkOUGguCxCaVV17iLhkQ1x0MQIS8YbADumWsuBmphJKcHO3OEwa6zEQXY5Dh
6srXKP+7YeMMf51yIvFa4Q4ME4XgrkBZW50G/lxJdb+407ZMliEaP7QEbJ7Y2XYs4w8o6lcWWGAO
7EP7ekYYqTGvdqPJG48jB6fNwJZJ27zCHfGSKNmFSuyg5suQP+rzaZDivsN+7/XdkS+GXTeg9mE9
jigV/Xth4rl1KoYMA6EqPW9GloJFnc2zMQ+2bZLifnN3I7rWhtdMUg6apE61q5y25ntSrSAOcg5I
AIwMWkYh9Gegcrbk+6aPPrqF72urkNf9cSgKZOoPDImipqSzt2U4Op0EsmYlVoFxZHnstpV+kI2y
QvdkSSM6oea361fNWS2JqjNcfGD7lDHVN3GLBSEPLtoxpzgLW/kKxbcZjAy4dnkvG+Ual2HqbcuY
7tWFIPdU6LHDqckBdCxD8KUrfZYhg55nDD8a3JA+2YxrF26GrgV7UgLHfGy/T9+HeYdv90aJc3io
EfO0ynmL7OSqIrOmjT/ymX204qZrUWRc45s9/0e+AqvdzTsLe0OZBcTiDGF8zSSjCSFo0qDYsuPy
cn5R6V4gJIEjxZiI
`protect end_protected
