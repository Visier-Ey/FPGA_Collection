-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
--pragma protect begin_protected
--pragma protect encrypt_agent="NCPROTECT"
--pragma protect encrypt_agent_info="Encrypted using API"
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
--pragma protect key_method=RSA
--pragma protect key_block
UDzjIGOmNUUSrTEv2nw+WIOD7t4oMrmgpF2yyauj3j09X4+piGOTpeVMDSUBLIn7
6bJz3E4tUrbbQ6UuWUGIzEmVjZUJT5QX91DABPj6pZUsnvXT1WRIGl2GWAIDETg4
KD5hmbq74ngTcGmPTqSWUcCN3tGVSoP1roiLi9vjARQQeybEgRrqgWBR6tRpAtgu
4A/Imic7f5XuoDgx53OYKWUwIR0oBa25H0qQN3vg8XP5L0jI6M8Wg3jg0NOdjlVn
NU3wEsSw9qVqUzUeQ6iPyGTbRluWUPhmsLFE9FtZOGxUpfz92x6m5GapCn+G6sG2
2nddwkogFuIr5DcTvpIAYA==
--pragma protect end_key_block
--pragma protect digest_block
2n4R6P2EpxtlDRQL3GeEEJJru+E=
--pragma protect end_digest_block
--pragma protect data_block
0QDs3wzgPZQkFWSoZRu+53lHutif4jRmtuCAYDDKv3lHZsbppM59+g4qsVkGh+mu
lgZJmDgaNVsvj0dNWDfDivoDy/kJXedycrUeeUmueMKuq/jwB7rIke6r8pPQ05Is
EEgZx5zOoUQzVZgC7CtDrNytZ0Ik/JIELDHkQktGzt2lJOhdh/z4/rpG1qtAzTPP
DQQvI/r2YCPCrn0VXpqL7cPkUZZXGSTGYaVH6LW7aQO3XGR+ofrNPsNdveXoyfr2
9zC+MU4rcQ0NmVoRWjZHI3fpHKIEHbArHsBacGKRaJzuIYrzjIi6/5CRCz5Wbql+
4PKMt1IB64WtCpnaLWVekliYc76o79Ot5PbkcW0ita/TGtuFCbr+8vbkqHAuHaAL
ywcbq7xRuwjiyNf66M/AzebeE8BfbaNZi4s54ZASSk6Sw1TqJ0Q9Z5Booel92m01
y2Mx8bkVX+GGXdchOnK7ooecUAFq0cS6qxBsVpmOvrm8TG3MbnGFZIP42FFTCLHZ
4vF3M6jpq0HRmmfwNSIXCQ1hecWiibu/EWlom9zkO8x5z2jrmUpU1p+wj1+jjWTu
CkzHVE8DBd7iAkZzBUpAmnQJGSDvnKvdwFdpY/5upfklneJ9PMgV6Fx1D1TGiRf2
vS8Py9C/GL2ayspjRbrDm2yDWc3jYKbQYE6ixlZrDaGUNLigJw8/LYDDswh8b3VI
HXZHoVw/TX3DhOMMNCMx0DdehAKtZ2xJpOQi15C2NS8UXMtjWWYYWVjjF96t/w7i
BnC6AVWsQMM/MNFVLzzgHwYob0sMUw5GkTLW193HDcWuamByPGFpe14ziGLc1Q29
Tq5od1Oty0atjgN4p4FwELG4AAAFluIT525atKBhiRMrtbKkf3M8xZXrZz31VGIT
CwIXriBfyIxrJWw1yNN+pnVEryogZSMkTi4jp27NX2uXqtnh97Y2KKUuwAnFPE6d
MpNECFNRFfDRkMzSNFNE1O8gzlilvGwz+RqE29/vsvIJlUsO8l62UkQa7OoGFKHB
SzcXDotzQTtvKp0uyvYI5Zq8l0RLuaNYXQfrm09jp1IlvYnTr9L2rjQLuWRk5Yy+
o4yDFdym9zVHzSUt/OSd9gC07E0+jIGY2pznFi+J8AykO7WhfKmikvOHCoSspsMd
kIadLL3/8B2WwnqYXdHNCAv2baLY+T1UNajChDSWWEfuP351/j8H6cYu6tvBrutn
IKgI8uGdANpRahyXhBVqADu1U6vXSMyfrKDyndI7C+gRzz8/Im3tvN3U/XgRNX4s
h7dGvhgnKNwVS66N2gdmI/70ACatxkI8Fvr2VRkGzbEAP6ykdaI4bTEvg8jrC+hF
3TYE4mcOWKGeYhUwj874Dbe+J0VSVXQBrp6w/zzcHeENgIXhfoBoVUQfCzzuTT7S
4tmBI7P2kv3IjnfFGWH8zbGglK3XCqrwwa942kx5gxjbQxr00+7mYDR3Q+8BoHGQ
eysixVo62DteEZeSo4zEP3xdv6UUpfPOU/cW8vKngjRTmdxm0TB4qRGfEbjBSxCZ
h6qRuplb/uRC2rUHmed2KO34qrhlqxRirhsJjCXbUtSs68TqtxOfIsnKRlSXN7DK
jyG9fe8lpEkSwluvLp56fCRy3w9ewA+Y7sNEPNiNMNOmleRX/NrhmYE3bf7GDX0X
GZcE1MKDZSSWx0b0CN0fEV/wJwkshf9YibmuRNVYCcrSwOP4QU2q3iNZfCr3k27M
oElmtCUD9gTStHPdXMOrxiMjDPlpB76VGWKligJky9A9CEPd53Awq4R+rQ+pz/mi
kkjeOr1ILScxoFQnLp58+mILJd+eFWvZjdyaBpS9zyiHTVqLVKaJdLpyt7I/9TC1
tq2SH8zlhpLWQ41/GlDQQB5g/Z8UOdp2VG1eIKeRgvKQjtH8kltvPmIueGR19u77
haC/b85pVMyHBV2eSDXX33yv+G6sYT1a2tXY4LsL4ZxdPI5CrzyENL8WMyz2vVW6
ZdjJ8eIGlaDMdkp6ACfsNX7vGKHM5yTNgcqb9ZyOcoz3JJK4Ju59lK0JHfoVP7Ug
MBDBxHiGpkJR78kx0UH46fxxd6lVNzDQbjxnPGxm5WCC6R1+J4meAvYNvcKdV84T
TiwxhN7OWMEr/jdwKz9euU1ufGAgm+zl/HZykXAPXk4D+1V8QCmHLhv/3mZMTnWf
dS0bw9onirPYKq+IbdXjHLptv4VBr1GII+ZLNZ8hTQ2TRY1wH89AFq6LwRaqnmnH
Tasw99iW88s52Qbcefj0je/+um9p5R1Vem/Sf/A+buE2XEokmqSVRqz7lCHiqzGc
jwICbzcQvPLTFJ2Xja5hrAUvd3kxusC3qnPGoSKHYcxVz7cliE15iMLnPujcQ+Lp
ZbB2ECqg7Lco0SiTEcR02SSstjgJYrs8U+xf1i4in1EBbvKbyPs7fTfCGs5m8ATG
5v3UCf4ALBc0qnZ0mkCKT80oFCKEM6N2XZXiQ2xnJdzj5lac6Ud1zp6eFri223u5
a947LZTsIANFS7CdwQRiwm8SafZmq3ShxJKf/TfM/fEPMGfS8PKlsnnFYvZ6656J
3xGI8/DKtWe9U+nwvRD3hdP7Hb6U84AfkwmIcjIn0c5ZAMJINp7Gsm9gh0YM6y5E
IRLotwn/joZ3M4NrdmWpWfiVORGItv4Y3qzj4EvZe+tZRcd51bjt9XoXaPvwyyfk
9xRM9Clnr1iuQoNHZsERqnCdS9LCJVun6vukcKATTgadxpdPCrn+BP0NhJOltxiB
dyaq976zlrxAOHMxEEWvvqo4c+/du5Nv/kEazjG94kVGbr8vCux7RA1n5i6+gfC8
opC7GPEBuKsKhv+MfTL7Qzl/r/hTSSYP2GBSZkJ+vMtDw6y7Z6pc7r6zb5QMfPK2
1IhzH6jeH6hjz/xqFtfSnCox/5bfvKCOJ4t+92sfg55uJRoEvEdpJdfhU/f/Mfv6
7f1C8Y+zRiWehIDfTer8bXbU6C83YNI3tmigE+fS7CSjI6oGzFEoeL/H7RlzoC2/
l0x6tlg2KdfOuwokjfgfwK3PMAuxxbaidZMRMyTuifKy6xCWjd+cHC6rdMZD/vyy
t6Tdxpr0ZPyNT2szKg0otvSH4LHwpgJK+vAeVlywnoND+NK58f2oswJAnpllGTVh
Zo/uNZPy95Yj2yWlkN9EqJXq7kl9JI9Lswp7NUAGuRKQzpQAbm5K0XqNyyN/C49k
/gSX9GqJKqvKeInWGcAglhx6yA9491h/poTGpyrJx3m7pqDWTFl5sib88oD0oSMY
pgqhYp96xgZQ6hHQpKsJKC8PeKcaiEcbQfA/BaNY0OWh1Jd8oa/P1k/Dqc2sAcBD
uxNW1+JOPh5Cy2Qx/0O1pwA4EZIgj+4uikKKItP9wvJMKFuCcUBKPk9cKVbh2ZUy
A4sb6nXRFUDr45+Jyt325HsjTFOMD4poTzTHmAzALCz5Hb0QyvureVPGLetJVnAM
3ClDHb3rUTNlRLBtlC+8uDY9oT39ZY/D3VHeWCqOU3WSYNTMACWzCL/1YkHXoe/Y
IABa/L9iyl3w7p9lH6DbP4dNqEwfppMnaaZ4VimhMtuyYm3cb1SXXg+uZZv1vnCa
Z5gN585ovogjNu+sE6g0qdGn5h+ejDqNhnw4RikR3RPgo8SBJsxKEZAAuuZQlT/M
y+dcF/tMI8DPuEhCMafy5qQBACOwn8ZK+pPDaPQhWj6kA/Kcuyv7qJ3sBnmf6xeE
n8lfu7KYVun0mDV04d8fSTTcxofsD3Bom+XVNlJYI2mS0VmDROKX5C1emsRAc8Wn
kooE7Htfg7fFFKsm4li6vuxpRdOffnvCgpo9EQ8NeH0q8OohyGWvsO16n90TRthZ
5OoWXJtJZvmYET3DkQ56zkb37xJ/XWb2JnWXUjdc4obiFBHItG4gGY8yGQc27W19
TaJnmFQATGkXKbLXeNwvOru+N4XRBgS2f82Lbfyy8dzOmT5+5rmJNVJZW4HtguA4
y2jeio4P31oI6iX3t5Nyip6/+33ucyRKuY6FfTnPgvICKmKsHWNGGEV2HScDpOsV
iCY/vXIWetDpJUPZ1E/nu9sqUTlxhnpBpSSPZ+h1fUG9GpJ4Tm9AWT4BtyWeJ320
ERbAZeSXjCQpG61HaUrNdQxkzsdcR4JIM8oQFxjEdoo+vqeh6tT7syczfInf5aVz
LkDOv3mMtIOr1rsXXBJsHw1OLuYnHYto/m3lv1MVdOE5LgXeEi/cFU8jiQdtxEKS
Xnjnau/qF5bIZfQYKzO8VCmcDhQPxm9Ewp+4PUus2nyxBtuVGC1XVGx2ncFfRGnj
jtRuRWwr+FagxvwLe9n4OqthcURRhXLlRgvrbFsYxlFVWN1uMQrJzipNVjQzK+bX
wNY/1JwMBRFVuELvYuyxl3qkiqh30R73JKmNuSGZUxzkPebkbZJ/NegDSqLf661Y
FAfKvmJyXP0WjQzp7kBSYb+FAGQ+sxGYt5toniRbNyC1MDOX1keFZ9JaJcNt40nl
UNl1A/nLDqoex2Jzf90U+sReyIOEaqps4FS5BxWsg8OQU02lMDZ7tLAgFYeDjU2O
5sc6/ynOIfraDFK2ty7AJdDeiOirQdIEmdGjD/5XvbKLBo8Iu+IgXZb8ngid0lw0
GzXQexZKT6u1wLIDi9qHhsPspnLyKgcsy+J7qWp6dSjVUzwbCWTuucN2fqM/oYB9
0R/SbPzintDu1z4Jgx+drjizdnUxTIKudSTTpTWRuibNQIG4h97HcSF0UsfVp86V
sXS2v09BadiF6xwWL7DAobNreGlymrGsiILTTmpA0oannYZOFDDXTTGMvfm4wrRO
5+iuS87BWddEH5BD6VZFRV5nXC7hJCysNT50k9sv2clRrfVs3B1M+ksiJOnyTtHC
GTucwp1M+4F5syejxdt8xMBREdzG3Hm1xD/JD30NOcaXb/Zu3bys18TmSkiObj/b
kZj4an+yC1X+W7Knf7fphc4rUxKfRdl7cR4aBNX5NEkgIARljySK7MtiNjwGOKws
EGnXnBi+mdrLR8JS8o13r7w0WWgpaE0KsW3jsx9i9CZhTtcyzSEldSlsH4VtYB6l
L65ua3bPzv7eoiMswKUh0Jvt9kGSkxwXmTBxSGlub+x3UVp3dNtuK9nITtZQPrce
b0KUq0/+ATb5iaMQ1GlfQf8Mr9rE39n36iEPk5NF2N54Gx87fGqTq726Vz1bKNex
m13dMHecAx9deihTYVTD6vdWxM3DNGniDZ4iVqxEF/onPV3WJvFCI/o0hs1ryefl
YGJ2n/6EIYXWJPB3LrCXdBlnwG1ORMDPmKVdULLTMzwJD9CNIctgfWeeYS1Brd/v
ZU1hoS5g/yat1uIGlPDbIg95+nUenEpSsEK/aHwxUbLRw+JDM9739XVioAnJcvc0
096vbcTX/5xfUDf9RZID8cUHudkHnEJ9ZamRMf4xPog3u9cYi2XGJ1URCkTGJQzb
dFDMvC6pdxvjzQNdWnoG7Gm5K3s1KTaZEMcmLUFY3ZBxVbDOyGyUgKgizir76D3q
us0Lj+mhsWWELQOLr/hHRx1K5z5GI6zJFEfUkFbHIvPEgq2xuzhU8wb7T68k1qNV
2U2HONyEMCroQbDA2LbbFiKFzgO3y7rzy9d/b709IBlJdIMXPnrJN+7+aMiJH7VT
/NZ6lpQWPitSW+BSav5zihV4TzMrSv957gu/GL3X5hptUhSlpxA4m+T8/H1a+iWi
YS8rVGfvzKye9Omu0r1ckr3WCeKIuzCdOnb4xk0kT03yCHwor6cBYsZa38aG4ad7
4DRqjRhE2exDmLZmisLIeGNcE0KhYBXU4atGXkntGoulikIld5LvEXRFaLjMkeS4
pPPdzTlbMox3prMO+Yy2YidyAQmmj+n1E89Iq3Q+3FH9kI25n0oB3ItsqlPylg4V
Efp2+ItfPYsDFLTsrTsGtvtrw3oA7sPaFgeUnR8P9Ci3NHMMQhSxBBuR6kOz4Rs/
t+dSC4/EP5WFJFP88U9lZMYl2T9J/H+O3GY36CCnHyHcLZMiBrEnzKEslahHnPsa
iwfJ5cls7f/Z7UetrBoeu4JSBdqNB7jxCxK6q3F/OVjI5XbQHTW/ub6bGCfXA9SL
0fb760ln655uC2GIpkIvJM9NQ6HmY21eNJ0Ec2Z2dnmFkX9qrGWNAvmGtY7Ef4MK
gjkOlfcK/5rBKhOSkRTWa3GXaoqaApU4tz6bZHeuM76qripKgNOo24H7WD64pbCR
NYFWln4y92GvMBlpqLrC9wwui7nSEkqEcZvW7V5atJoMIFcies1cZgP+fsMTp1nu
6Yrr+bvUe1R9id+RIp3yeEU/nqjBjnA5N/BCMPcacr4GHX1ub0wSFTAkZqK4Syjc
U0a+1WTGb/hFWO5w3i0tkGkMON9SLYMmXivAr7NBAE6yqzh2q+blnwEHGNHx7eul
Dst4kbCpR51cotRQbmNOMaevCVgKG3jtauHAwPG9FthAT4+xWtYwZoWqcXAxpt9e
LMbwh2nYYgOC2BGyihaDjqdHi1J1Vl0WW3OcdsdbLGmqbKjoBaLsi+hBlclyOwOB
cR7H/fm/V6wQj4uAeIoyMVuq40EAaeSdkUaOihubJq72Qxof7uHMYj2NBkLgy6X0
tXCMnaFJ8pAeZtO4VI7M1ccRFjAYyk33VAn6YyxW1SNL7DYM0I8gDCU0eeNASCT8
hTPT0AQVU7khFZHRJCLI3wedlJRc0c+DragfSvmSWbAWRa5QQo549dpRymcUpa/6
wzEKyJFUL6anRkLejczk3qs+WdH+t9ipC+kNl//7WAf3ouSpYNgFH4ihd1LBWqmT
olFpnZYdclR9NIcyqfZQHqCciLJ8sVzN4Z+P3kL8BOugxYZAb4Sxr5nRtOoYZPRu
47qETdm6fJnAyXvtC0FwVcU4wbw70bw1IuuQ/JoEDLrbtuooz6nnLObip8r7vNnK
TrUfojXZ3OjoFN1vAD9hlFird7HfocSuMhpaBwG21SBZvQDtMHxRE+1nf3MKqZFI
r4zUUGaLyvytEvG5zMUyxQbgHx89lNVa9nZBBYDi4iXZ1HVvmT33hemPp6dEoRia
zrnnvBe/+e/6/38mfrsDRlj5CSoyLRl/NtiPlPeLac35ACL2WT8YgIv9X8ZUv5Sq
zgrr3FnIazDpt7H+95bqZmJL9WSjRb+Ncj4JwwTg6vZf1+7/9X/2pZm/dzL0Cf4Q
msEatIk5WToOpo1cy5VHewilPAuZ0Rz01xtbuE6+rT7qsQBZiWs89vhUbDUisupv
huMs8MX11E0/p/Sj+tg6yHN2yhpTkLdIPw7Y6kpbplawquQeupYrcJJZ2ZWMoczU
JpDZj/Jb3DI7lYafxZD3B7wolLNZYvsSdvd1nOJKbPFwy+KXux1npMEQzUjigxD2
HYjyOeuZBKFtKEfBdUqUY8llvzInXI9n+aHwS6hkBFn4llf1RXSlfCbI1XnTlIK9
j9tNRfkeG0QQJ7IuAGFLL7iltcjUYAIuORNp8vOeAyUEzAdMTZSNbuND3BG3iToX
2MeSx1G6lAYx+kdJyrrsXnblklkb9y1hYirWRdSTLmuf0E1ja+K5wILEOFLO4kEF
q3EgTtxIHQN5nHu6ZboeDK0+EKSASQC8ooBOvbU8czGLfRq/PuX0iadbYnEDTdnB
5oH0XZyu92A6QltIBVv+LOetWqE+GkVWW+myNIlFUfpkMCobUH20/Fs5xbRHztl/
g2aYmAzqnZslDRu6MDUJU2dQLsbmxVatkAlkUyPCj8keUHZplKaf4UeQogmbqIXj
KRbzfNdw4LdS4snfdt58R8yDulEAalVWt9pvCI5wBwKDSsUPhRBRN3dh82W1LoMm
ccNO+VpvnefvtXTSROKyE/Hql5cnpLcuruDp2k9HbXgz5pX/gq/kG3QO57ip/HSC
T1Re8ahrBZfSSmSzzxSTEWkUv3+Q7uIH3jQaBpcVX8FlUA8butq/9xbDApvCSyap
K3CUdsAYKgq4r+g2UJQMMk6UuctGWRdOq8DCTKi+ACQlRPwfnRYLbcWHKzfbREi+
tVlvXUWK5/O85KmOGrW2hPuG0YJVAROGWQ1Jrz935RFKKuZ8vmR+YxK7kfk0xdJd
Y++acJHhKXoOsWvdfdXoWXgpNAxQTE2jyMuphVo6kIgGTTbE8sGJH/05xAmAmWVN
2QgrI6zkV3BWpyo0ndstMVXosomIBiPN+rANBlLsobG5y65YvOyXyWV3AgKDDikf
JOwCn8MPbDa0Sc3CGKSaSsLpGSaWsdCdYAVQdPCMxjuwE0+DTTpMnUX2Nwkxji4Y
CfFisBew7XiUlPcLuzvR+6mA+lgsMjwM3tna++qDkDKQAAn0JhBdTb1CN0VgNOII
0w2Wp1W9SlHgQgQAb1DSl0mc0GDqch+uJCDGWcbgkexbWQlaZQ9HixR9X+6haqKM
Lf5o8uPljyhDoRRBCRaD8vUAF209vEDo9Lq0Bm4izKEgW3cQx90R/pfHg98Ntx6r
Lghc52Ct6JGbCrFs+Rx6UjsYPRP8kWMPPOsWZPg9JoH9H6YHSIsVyf4nqoQzd90s
qbq1WBJBOzwHksrKFVBMqpZdmN57ar0PyeddmBjiGd18dzz7c6YQHvHXWEffCpsu
Fe0x0Cl0nliw96wlbduEEA2yMBpv+QC58lbDdV7Oii1IGplwVWBAb3IicrcQ8aQz
pe4U8KIha8XIxYFmiYSisj9X8uHJ84OKuUs5tnz259lIqTEoz4qxonjtJ5hhvMbT
wTMNz6+1Wv6GVr7+JGlz7f/EOZrHwX2lrnybVK39178XYDk1rHG2JWH2fkhYDxc2
t8evDS1Del1GxSjM/zDAqpk4Wvug63h/sman2uo6rR6k3Ekvux5Juk5R3FNFT757
7lVuN7Z+Em4D/Ib/rFky7Uebn9G+h0eNaIzqu3cdtCFvpMJvdzJPMdhmKvpdEL+O
rTfWgbWqEUGC2J63KvCNS/9j1Xvt/XZYjjhD63389Fg2Mgl8PsUtHCAsy5zjkjwt
LHSzzNIaf811d7uHeBs/BOVARIQg12tkdUsa7eP7iVdpXXiLio7swY5zHIUENOOp
ymx3q8Y8GkBts0keL8BYC5XIP59N0uz6zbTX/OUKS5kmumPif3StCTj0M97olfgD
LtNw/YQ7Rz+ltVwhfk1+tDrsTSpZbVfWX0tSu+Feg6EFnA6+OmblbVBLQIJskf2I
swZG3zly4J3vPxOuy+MfCGK6dm3jBw192AB+MyY1SCD+Vsgx4j8Xumw2yuZyqJJT
K1WnMcBhNDDgTTvxePyBzSMPVph2CHGJrKi9uHyLzE5ffN3fxXEn6BVv22ySrSh9
V/dJeMgdBpWKkAPEoQKAHqk/bZlP8ao/Mq7OD4uUQ43S0379jfk7PtzSstnR/SHa
OS67LdJpCT8WjF8Ftkl07VhlGQWD9Rwc0h4qRHV7aYrg7BjT2Ni2Mr9QOdRAtpjd
dqiRkozkAhURoCm8YJiVPKrzkRa+fxT7/WQvEYNWJn/NNKWCBtFJiauQcelQP/G8
wtovmkSWI2lizz/iFFiSpX696z8Azj3QBeteXWcL3VbbgWVsoI0w7oF9kSIIdSzS
TwVw5z1TI3vsOXZ+xHSSuxFwFuKxPlaMJuPrO8tJwOZNkn5PHI7eNS4XtSMw8Xn2
zqrkM/71qaDkjX3Y+fMQi9zauTaux3QZnBuBkW1gKt/NWaZcVSvUBmuXdnGG26Xv
bRLNjhu7re7czenO60o8ZzwDO5KMflwFyNdOQZY0fMzuvnUChvpd3Ky3YHHv3fcf
P1LFjyM6IkRmX4HfZhV1E+6gKpTeuhl2noi+Qi8EXeY7tvEJDUn3COP6aqKMX96F
7CdwPxqLxwakFm+YqjbZZqUhRByDq/hJIJD3lMP3wKnBWPgJijyOKgimzU8JxrDw
ZpyJMVRkkg4rYyyMisqgJB7CD8frX6ZuSW+CIUgatIGl6ILzkjLj9JapyPrEXIMp
sOCAjJoRJ+X2+2/TuJysG42/+vvcTGHmtZtkF9s0NMIzjRwgfl4gwDtrN1pf6SON
AjtnsB7AmMFcnrzKqRBjw/9WRqFHIaZ2eLPWRckkPNpamIE2ve+PUKmU3dBhvfGR
QV9jQdVa8o1LBl3ZE33u8smzz9DV7dJDiF1POhZMZXNgUWKEFoxwCPMTRo8Sdfxh
c3WQMV36hFE0uzoMSJaWe7GG1gm5IG9IVruj6j2yVTWlwWYYUw3rIVV9kwIhqRFm
AU1f3jWz+GZv1WqtrCGM9FlYRRIqmZSa1gBhO1LvBHUlEZpq724uV8KMJQH4YcvG
3h7d3SDf61GJHgY0GQQyhiKl44OLivxEKhvATtYfGPP0fgLLyPH7zrRDDbSEJvMe
Yub6b+ESzxXkk4LhHONAiql3IvC9+THf+dqnvsSOj4aCBPWxZ3aSTRih+aqnK4h8
LrXBmgqMxTPtt9LBvXXUKCp7Q9/gMfvEkWp1e1x7CpbaSba/RcYm72OlL/vAbko2
K66KA0Uw/GlxvqZDyYAZFOQ5ARubTK0uSVChIqgzehJGnczF2DwoYLJHIgF8ivgc
JGEKFgrBtpWY22yDZeRCG2H1ZPUe+D9P2OmS4RCPEw9fkiJnY+sy66uzGp8MEESE
fIUkMRN/7NWOnG0v5UR98+ZC9O07pEjszbE61NOJKVOb4e1VpyX/wknCaq8jkTA4
NcJbPCvK7LqBUcq331aEcdEd/BMOHtJgnv/83Qph36ssGKQHx2UCSaMuYSf9KQkd
/qq6dC4kNWo7Ny5vSNci5m94Gp6cCPRfdnwM988akUfMu/gZNkP+zzHf3aqyYCK/
d3NkgKKExzAJln37NceVlDX0i8WYJY81djPEbh+nkqiINac4vqpOpuw7lyy09/Lt
uPYii37GhYY6dmOgVrfWsyt3tff4/qrtAxNQ5Rkc5QN4VGvicRYEK8nx4tX/7x9H
V6QEQWuAxEPoz3s9oxM9+tDp3JLV7/ug01SHe7FOTWxcNstTnqssyz2+ZNddnpfF
ExYS3d4czlEAPiP+pEfVWqZxss3OVNoSyqTOQoF3YYIhGXhylX/tmvdnxxQEmW57
N8peCbVU+WkektXjn9nkLnGTA2fXdRoXgvdFc9s1ZhAkqgGZ9crMEyyvQDd6/H4E
Sif7ZhwU//pEtoSa/vumMn7fuDuT5Tj7oRzA+f4GCBSPcjK91vTFBvCFyvwKSqSv
SJf2n7qufmulHjswYE1mCyr39/l0204jxuAGVj8EKPs64bppgIW7InecwB4o97d8
cSFRoixMI0n7kIw2rmmdvmAZ7lnwCdtKsU1M6hOTp4alESoPSa7RgJBeViOfDDQB
2e06egF09mOj499TIGOqPgda3xR3bf6WpO99D2XCesdbl6rB+XsRO88RNZ0/tD03
cKFSm/2qYe6PzTRSGR6/TBNkIo5g3HaMxrgH8g3fZqMxoD6Kui34UQurzDu7X9IP
kyuYUOzi3iqXIwNuq68jdd+4Y6JTb2c6I+0ynIKv1mchn1Jmw2ux0O/HwZowRaIC
7iQ1Ky8MfhFEXllxzoxBghRZUc7+iy6tYbSeCC/JdlsdnWyKnFA6dUjGjV1mcvAB
u+sEQUBKgcvp9yJNyTFJwwoRZY81uCLg3DJaVP03kMHFIQi5ce+KeD9TA+lQPNMz
G9k//r4soiy46gTm/orEwSLl1QZ/4csh6hraJ1HDy+GkNBy5MRi9O7tIUfO0gwEI
VEFgp8zj1iXcntDEdjECaZlW4+DgiylGouTFSXnKXeeaMPrnLUUuSZrvxroyAcfb
ZhCgnS7o3S3cNYmpCVSDrsjhlw6IvWy3PjSkeUmYvfhYAO52Zg5Qte/O3olxXVZK
7JEQjxmJY2eZst2Pf08eWAL1FwUSILyKKZy4+xtYO89LBLtQQPB311UDy2d8fEBd
vaMwg5X/EyJM0Le89vOPLXyI0gOLTauE8ZAxfTVQlzcHBSmvL+gsgOPmGZuhNxUc
XN7F7Na6WMm+IHob/rg0cBYMOlQkoLabTQTT9sC07ywYgINvt7NznsyOXJ4o9N+g
jMgCXFsIt7Xh8idSR/ENxj7D7Wpdky9s+DHHQtM3hkdX1v312L4BdezeiUFjayVy
wv0in6pzsIwxZ9tEe5ssIqBu+/bVJQ4JXW8Bf4wvNG515Desgx1YLZso2EzT4q9J
ZVuL9YTIs4XKTVo0M61OoCsLLZ/FZfn/XGk8lWQNwrgeN3aJHI6dqRgnmbrXqLe1
ORzTiegH7BEzBX7ByDqN1zsmzvoVveL2VV9SftOLjRffUsUg//+IjoPT0Ni9a1dN
rzFAAngyArSLUVoJkdi6QmFYOYy8u5PDjFFu1LbuxmwQ9qRRESMVI5o1EmuFGwDk
1hBbAQAg2IRUyFhTGABR2qZ6k2XOkuXXHUKoR4/kiBw0S+onNngQ7O3yaITDjGgE
OpsoHMbFq5HOIWtVTPX6mtCixRDkFDbhWZpL7QZgQSyWJeQ1AaWjRV0FXQZWzii2
6CCtDduOPuALIntx2BlfCc1kgd/8u+oNAN1cG2rYgWtKvDBG1sDBddbQL4XBQ3T2
HjUGIiFA40V2odIzjuUyBvDxJzMQ+e5AX+xX4m4ad5Esk0R/uwwIO2VwHVt1gqSo
N7Nxc8tP8Rqe6wR0ic5UkgwEj/ac+P7fq2DV3zcrmmQVKFxAWnq0b9t3Lwfos7bh
7BAeaRIDka83SuCeGIRBRnYbNMLCMSri+Yr1uP72F/h+Xo4ay6+82vErezsHEKJn
Em2yR0Ma72fHEpuV6/OO+UX4sDaQ6KVsvDmmE/Uas6ZrDM072j22m2sOE5N6I4pA
Q8Avtn4mJgBIkVtsWP6N83jjR5aH25JKjqvhuoOZETjvsBQbzYgsgz6bv8Jnyw9H
H4mYmvmoKLgPcAZYBAPSGcOPo7dsjB/9MHC713TD066ZWHgQviaTaL+HpuZ0ZGEj
o2HIZYHKvMjtQslHQQEPNZf5pe6wgO4l5rynTR+Yu5rGEfn8sXRmUAgoYmeao8ve
jdfjtwSDb5gjILIlaXr6ids2W7YcGXERtPiUlUCIEtFDRAcqVReoQGOpSRiuYwuR
L47fv90K/y4EWjDucwQt3ZUdoSIOhSzufbqlxq+Ybeyikur3SsmNiojRFTme90Ah
OXVRPIGgmAoonggcrVSrwSoa6aFVe3E+6tGpKJq9RdNuaMKZAdoVY/eCPc5p75MP
KrlQ25PARafRp5+4OyqoEwK6bK+yKhOv4WFOWGAcOf8QpObZGeOdbnPzIdGBFqOI
pwMhgBlSJ3XhkA6U7Bi65lzh6zfB3mK10W08vhAq98iOjwp6h8tLdRniEHrvVaX4
ynQgID5C8Iau/4eCyoG8ZEUaxRJkR3htW5qNqbPZDCmph03SgxHFfF7VwewQis1l
17ECh2hwfZ4x/t0QZtSc3Hf9tbyvgT9BsXmi1bdQz755I8s8tXDGhKYvqpe1KyD1
jf6oV5Umu1UVNS3IM0vBpfGwqkYT/r5N4IYf6HfTr1j1iPjg62uVivS2NwJcedjB
qpzy7iDgDeZqRHIIx1+umZDCgFJipmF2RA/8Mr0851iVVuEUITHF7PP/s4p1Ml5h
H9JvlTFZ0ZqFh0qLY/TBI9SLogcFcSMU/ZgOvfs/V7+Pzwq4IIvwWFON+x50miXv
fTqStcRyg4I+E33ge2DFHeydH5p3Gg4QUNGDCHsIS+3F/xoVBgfFk9w5vzX6EOh6
EZeIQ2jfVS4n33UIch5TAY9xlmWX0UTvm3mOFFeODtsCA1yXYVuPBliaVZCRFwUX
rKcZdlc4x5HiJUs3d2fZpBMxZGWnf1CtXFwzLh7q0PxepBoBFEg2yf1ncW0cAU6R
/dhzgpuYiT1Ds1iOmLUylOLEG7NXdGiuvnyIv/gy2feDdFbV7IvwLljiqgiFTMtN
xTES4iUVqdET40Wen6kCyOJ2PPLhGXqoB3lMuDLHZwVqZS9nHelrNtA/cyP4x7OG
jycH6pt8c4+884bXBPBeMqkK2tITcKr0aFY9Iv6p3ZiyhwWeCuvYbcaaIul8G7YD
/p/EwivSc0M+v9ON3Q9iO1Cdexo7E3rQ8yZWHEthZqCLQ7XV+/rmjmDYBrxVmL6V
wPUqTcD620Yxed081O9x51A244QqRw4o3btDcdX0/+rKT2ALSrzwLpegK5RQMyDs
APz+3N0ONFL8qTiaUaJaCDrYw1uJmGB+M8ExJPJY6mtTriT18TQH/upT8HtcObjO
2f/6PdGA23eFLRE1YRbysXKaDcyLAZK4oouDjq6oHmpSSksjC/R0j3+nyYDlpNNR
AdJJaNl6Yk054zwFJKIWma24lHLtx84yiyIkHBMTz5R0jDBh3WB58llOn4zVN0uX
pKTrl9AILkbk7gRFoy/+QY+8wkBUKNX7i9P7gdnr/sQUGszNzANR01V0FV2iDJzU
heV1k8b+YaJwDOYjubBk7a6v7fwcS9zTmDS+5/0U6mgaFWySK1oNG314SRX4M1HQ
tJMhgHGy2vyOirOk8ZnHVzumzq1Ip68XziMMT7VQDj08hG5kXt3Z6Mry3gk1JOA0
YVa9j7Rb5e8PFJxticosV0EC1P+g/UPrEq3mQdCGvJguVqle+bH71vEb3k416t3/
oBbWNllhM9GMi4jR4/XAXNBaUC47Tel2GwqOH7cj7rLy1GIcNilsHncJve+x8k9E
avRptS7+NUKiqnDt0SmMytRTsJ651bBuRlZekWfhj29h65rHMkoV6GzFOfnpxzhg
10rWa7D9j0XdndtzleCjO5j43h8FdFT9IrkTiTClidfoc6t+nYEjnqIwRInGIVpg
DxPqlJc0BLoA/ZkMIKSvyb5c4QQp+ajXvilKM4y8q3vR56JdOz4WHCajkdRPbxE3
RMg4/HC9+S39zeCWRR3GQqDoVNWhsDpoZaimeXzeCx3APzObZ+2onu/I2fD8FYPf
R9RMwqUzmlYrvjHnhpF/EL1gXf7QIdo07RaVBEShHvnSgw+P47vqTMEicF53Yhzc
7PymnrMGV/NdSm8mH1ikyBzxgBwRH2LewmnKQ0xUrAgwALQ350F7ttUGR7q4rNcZ
nrcK/dxmZnIFs2sAt2VM9Hwga2056VMMJObcYLKtsJofzIGTNQq8iUdFcKBpiFKQ
vNKxP9KTHcD/GJFgwObvTOxckSBn3/j8bNjcMXP5jhsITf9bfW0EOxFcoIuho743
8uHesQ5/L6CTZYX4tBG8AAhhOSuz+eUuXMTCy0aX7oXyYjl7Oy59ZPYSu/IQrJSf
9y/dwIE/kgHEnu9vIWeklIlXlC8qxT+xZv7IOkdYfu/Am5wwUY45sUb2bA6gl4OR
EpiXLUi6SToNVSIVirnGXphKQGTMFcGVJN1i+4y9OgeeIbTFifG7l4OYJ9q7lGnh
+B+Ktb3EP5W1PM6IqAph9rHhfHoUt4YD0fKjfaJF2jvzCh7Qken79JEh6xGtT3+h
ASqJz6wq00Y6lfey5Rne+8xxDiyROXvm4x/TK3Odc+WjoosFyVD8OBXGiySzZWdJ
kKr03Fgztr7+EXGeHfbC9dLU13diG8+G7THwRAqb4NOXx55IphzJesoHBuuMNqDM
8IoyJ9l58rKgrHoKolf8mIfUCreMs9UB4P+YmqMn1RTIv9l17vAXNlZHQt5qgzGC
j2la5TbaGLBgoFTKoptemQsXqnDp6fvAitNWm0jVUfccl0SA8ana0iNXs7zwdtKI
veGYge74WfJ7QJNVIC0vKjgbPPtqnTMsaiPvNBc6t3U6ZRhnINtE9B4l0R12mHW+
7yOqbiiq5gYLiymXtwCi+BvtZI06QqmtasN2Mq0iCyQmyGwQi7On9fUsi6yTAA59
bASacXLVvp1drLiys9IUYRqd+pR8OTXYlMolq5jqpMDY/4ZYY8qWMDybIjEPvxj9
UqbOMuY8Ugf/mzrD1VUt9zAnyc9+pamB+1qLspLCCNUTkqmVflmXQIWI8KDzMcmG
0aVbtLkSihl5rN4/b3JIHb/EkpuC0QiotxL8SXorZit9a0uzKVb+6oww45uFDqo0
2V3j4uYaFm1VGUggbnlPQrbDw4Q6w1THVFx0D9B0AEt4iMe5UNZDShpjtS0oybgZ
eMU2oeXn/T3J5y9Hsznd2J74ZmE8CbhBTD2wztvIYBC1Bw7vBV4yV7CLba+DKZZ1
mquZdDig8qbw2oGvSt4PkDNiVP3tE1BFVbcIcbLxJY3sIefEwS/TYIqKrjAZZN6V
dpfNs+NaWottI6FUDaf15O9ND5GAIap8rZWkfIsg1o9ndmCL7mJeuEEhK9lCHTLN
E+tMRpZHxnMsVXUnsOVU18rPjcM2aR6yjdoOudtJdgOkFsJoKw2c+t8Rp1t3oO/t
FsZZvZXJZD0ebac76T1ldMZkjbSZTxHH1HyXddwKuSy2MtpT6c1FngekZHWP2xeT
03JxhNfUOGQx7nJNKfsOkKzyXtljDykszm//9q+3dXk3QmtCyuqVBS5IiUH781sj
d4oa78UKJZVS/HUHV7dfZ0C70isO2PopE5Zl5MIobBXotablYD6ZA/+1x2tVOrou
gbnnZGWu4UkjpkTbrhs3XBxw3IXDQ081FmnMYdqMK271aSXOKwxaQk48PJ5j4M6b
vKddCTjKvsMNNWNE5P6HvPFfQX10GjQ5Y3RxAYZGyUqqVrjAj5gq4mGHto0gsgdF
55LmRkvNvMwE7QcjNTf/brhJlsivDkw7BRHm+XUBOvTzYNnY95Y6Ut2I19Zxbspe
D6aXIIRiJH4cWZLu/2CpocPTb+RxqXyd03UApEhyreysT/fm0vj29ZAbGlOscaRG
mBv99mbTKK5ha8767W5TVTJywxcgl/I++8Az5hS9mtPzhsW5PiE4HlZQu87LhCWY
x0Sq5HsQJCcGCr89MKzv+7pKzfdGAgAFjFoC3BxYVolnv+W+UcNvi814dzrGFvja
DQCpioiJ8MmU33JJXS7YGW5TImNQuobsPUAn2md4wQXGdswyBrHNxpAsUFVEZSnv
Qd3l0CPmX43m6xV9Bc316j+wE0bbEWtr7Wwzgrit4Slt3j4RInKMSwNPbwRf/S/h
Nrxxw9DU3W2IENcUKw36nkbRaMqsPVfqbcHxHmeXLvj+gIq56aQlMqyuKHerfVYD
KihIchdj+A6aybK2PEgJbhdgU31y7eGRPeDl4jxwE3lPrnqAOW+s2WdAMRY2irnD
Z6y47ph0bsLxieky5YdFYE8Rq6ciP8XWPv4lei2eJo9gHD5MIl8NEGkrbH0c8t/n
B4HqNest6UZLlMyay6bsbXSNdHjBT1TwKhEJ5O1r9hoeeYXy+EsRflSYsjugxG/h
woic3HkO3409sCEVLgdUlODrDktFJbvfPfbXd4g53BBETND9uBSFOoxsI/ub5zy4
x1VdK9kP9M4ar8gbce8xV+GKKTtcDvxxTlnvgllVJfoKZuRD+UVcmwKHo7g0raPz
HbsSPHMILKFgCFxCGl6wtu4qZbbjpK+BAa3ESUSSYR6BKj0BqNhc8346oOy8zNYX
Sp5A3uOmXZNpFLg2tIy6n47R7cDS3mgUYdHkm5S6wlWlc1tBS5ANrO/dQmB71QV7
0ay0ifX9pXNjL7+QKbdYr5NGQTAHXzh6keK+RasQipR80iEUN6A/UoxxTY6qKSAU
AMLv3oGrogarByYXsM5zU8LKfdHB/l7iVijda5ZZyE5FccNkta6r6WgBI0aqlD6H
a7bdsMrtXhOX39mf8GCQ88GJl+r+0KdYYDpV3h6kPz4rrbuCJVk0XcOf81I0lSeQ
BorvSI00xQ0I02yfPf8jAFmjFRSndrt+bb7MfpTvXV1Hd6gAPHt/CYLERCgjdrQ9
--pragma protect end_data_block
--pragma protect digest_block
g0VpLahEalgU04k7Azs1/xez/xU=
--pragma protect end_digest_block
--pragma protect end_protected
