-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
A8t3VwyUL+tgSqaFkhlH9Cevj9QgfdelQYzmbQYe+gRc7ua7sWsHw51o4C3jDFdIXUHrBflDBIM3
lq8g0HSi5BPZf0zGfTrTIMiu3eqR/4e2rMhLskxZ1Jdhsi/Navfterp1rH7PVj1kEmimB8QgUZ6y
fTcbJ5AbhgrJLKfCmYrHVnYrjjC3+ApPHUaTv6zyqUOd1KIhykSLy8mQQSVWbrcPULoo+8TOwJHn
LXZOENFrioaskLMX3gHthywEr19jwD6j5Ly/cPZ7BiShtx03dysAjYg8sBVyZZQupBoNo5Tl8v+0
uhvPMOG47eqrkqoc5UwfzxM8Q/U5scoJ21/bVg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 1680)
`protect data_block
HWFPikt7J7XXerlUpFVGH8BN2EgjfY+5/Af7moRpK898c0WHdzPul1qHmd8ug4engELkOjrpjHXK
TMvpxHvJVxqrDG0g23hljaUStnBUvCZqyJcary1GwT2QCZQYQPw2kBjCdvrwR3JGSFroihJMhCch
r9HRnWOouCMHrHOQ6oP0ywFx+Ka4VhF0ov0kEfa8Ye7BbGOboTJKl8z0vu9JlAkQ4o4XexOTER3X
oGvpaKKj88kHO+gr7Gl3HvJUGEPrehYE9+nQErAAAWpu2rDRoCIOcOS9Xa0L3WDHvG2grwFu8rmK
C0N6xUSwo0lPorzqs22acUoGrdWSsHhMNnId5EocK/5ZxhLfrFeiqD2Ho5Of+uXTi5Y09CZaoIn3
bMAikm1fem4QpIB6UBghuqwO3GPI/S5tNIIvNZwgg4q85ns8HrEQOBVgFqAdORFF5u2SxpCa1ibt
ycoeN+ICA499nvKtBq4+9xLTzgx3VppGX6yXAU7ZUJ1724P2+OCyBLnz2Tl1x/PCiV6ugMD1Hpi2
5oqLTGXXJHXSuLXQO4lkVVnErXLbrAJfavMan1layhm0aQjBTfLrschkTD+erpCucTPU8v25sOIV
q0jbdTuDqVD08cr6Dx90mxb4NuxnY00PhXwFZqhAIkJxkmn3ZEkYaI1F26PO/oUPNo9c/TOLjXuh
//sPchzRRz5Vxd9Vlc39Ttp1aNCctsESPZgJ2PDhzNrM36lhVy0056smD+mg4PGNawI2DDC0bE3u
XAZ3nmVbRA2G40OH/w/qrG2xGbRSVCzWygSPofBQ615RctRqV4AKL3b1enmBGfI9dhfQqIo01sOf
JMWF/whXaQ9symMC3uWch9wkKw9ebjK8VwjldfTRdXgz6QsFJ7IwCP/GYwxXTEWo28JSMfeQsCQr
2gzAC1I/koPB45iePUAi1PZTL5fUZZG4dQoWGH0zEQibkRqImH5QFEQIrVdqLXa/dXiX7HzyMUIP
XyBVBrF1fBbPSQZ3iL8xZguoWs4XGPJQyegsHXHR7ZB/UyzwlFKs3LPxBjOEVkoiKaM3zk3C9OPV
bKwI38KQFcREbmLI/Zn+O136IFsYz5CTWFVrroq9u2R0CNvJHsifRznaY3NJx0WOVD+R+OxuBny4
srYIWI33cK9SKo7jLnf1DaSCGRNVKETOahRhisDumCb0GZvW1a1zt/iACOEQgyFfo+LV2F33c0ly
rE3P2Lh20rn48JQZ3vEwwHFE67BNIbcgPSWb/l10NPhmKoipVAgFBTfyNSPCLtSWrE0Q/9cniJdm
rMnWOeOHWLve4VIPkpSHPXXew5s2UuEqVxPc6r794QCApZOVcYvALLq4IJAmQKZvkNwPTA8uCb7s
LI1PmgKJCiXp0SU3wkLRQFOeAI8VoNAbAAjrjYDKbTQHCmmVVu48ht20JtF13JyUTArETaUfmd2R
Mq6cejjx1kLlH4Wg2epTDjxJK42aZb5jMXLdNIkAncPGn97S4GlCpgnkGFD0V2l2y7ZdYd++bBRx
AYUSOhLPdacXVNZTS9I4nABKK2NJG5Kj08qDMHh24rCjpQQfqMXyllZCUHlEl4vOoH6mq1kQoc8p
p9aJNMsR0GYbwkA3aHRSAyCm/xCnK6WoGhsDPcScPSfRiXVZ3QYVm4hVdqamSBT5QVNdwUs7pf3W
dpu7FKMp0EURwqT9RChM3odqlI1rpaiWrnoDd6QRCGsEJc5RqokmYgqo2qMNlqH/lM/4BLlWmQ6o
/TPeYPh6rhzNqKrJVXibgRmGEvpP5ex6Oxs5FSPb+Kt5Ar8slCvrKOicqLuMuWB+UFLcaOla0qhM
nBTXjOYpR1zo+31r2OskXvetp2+iWjr2QMYbihIdujUH17d0C0AkFasQF6msUcbNdR5Y2K6Fza7g
JDbUqUB1aysL9IN3WlpVjEaxMbN0Zgm/ORUwsZJt6ilKvJ+AreZCPISwddemI670y5z0EWvcwKL4
MbEQAcWaZUrbXnVb79xW71mhkcSru6UrBr0g/UePVK12HShG+LGfG0tdS4vPW14G2BuPlHHvuHuc
0Oz72i9L4xKOda78lwdUUGzmubX49uflxua1FbJt1pOQkjCKqirpiSnKxDXPTFuFBrXgWuFUUYMu
mxZgfLFdxZlBs6rKjE6l1W0ReAL1Pz3z+kqqdbEvrf/9FcLNkwacSeVIw6xiskTCx7L/BgCCEisH
uaYiSzvoUdWvEn7ePprWRD2HKSF1CvUJdpT5
`protect end_protected
