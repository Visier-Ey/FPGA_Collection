-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
GFcV4FGdvkz+nMGGXPbDoovqB7ItEZqAT1C73gbAHgcrMB6dRRPcGWls8SuBzKxZ
krKQTYCzPF8Z7azOQYyS2Ocf4FebFlIiR37JY+sZsBBk4z+ClltgNYthBIWIhv7n
QVCCIzYDOYUbv+vd2C4k426Q/PNrchB7sS8LneS5+50=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 7686)

`protect DATA_BLOCK
xNH2TYEDQpToaZ2T3JqWH9uXZYDPOkpHK5okYvO1ECIK9tvDmirO7eBDw4y8OXWK
z2URznhaf4auIJ4WlMIkA5hiwRp7H0/VoPDqCXGK9/Asn0YL+Golverocu2b5g+2
XXeEomfnNVKuZS9LRHcHaH06fVhkebC5ksnqFghxZM/ABtteB1FuzhEwX9Zgupml
KJYV1UbQAMKRnuyurrX4NG07Qvf7WHbgti4PqoBE8MArhNbXErXJLmt6vM+c26DM
xC7kLGqFClJW1YasXO0scYHcMTJ4o5hakt4X7SpZY1nb0UBuA+5nqaJCfcjToVaF
U1WU2J1YXeXsZJajXAKuo3KSVpLOXhsGfS47fGXqtHxPqIHEt5fR+Q0T1dlO1FmU
2u6Ou2nSG3M4UJ7UTVwRUgTFBdotWIQEugrJ9yVR/R1xGsCnLgXZ/wif0MNvypqw
Lo5L0uMWLL9pV8L8mKxZuyQPh7VqvgM12xpXsS6cNZ9oopesyaIwkOueh6Ayxq7r
1gB8f2Uawb9zp+REk0s1vF8SvDr55bLUXYUHLykumSvUeaRaAOG15Ew0sLHlSZIj
qYVxPfiWbS7G4luYCUzxT1lGQf+ksP7ojITJieE4ivsoJzQKqpLepa+hqje1iwKc
VOmBPjb0zHi/sR5f+txqT7JVLOS296UHlRZwQWQkT2Vobqye/7HvYAXtALmE8wxa
je+Ig4FpT6nqguBrCda6Tqle2KccoM+uUF6y/vDPyMFRyxBdp6JksQty3Fe4qnEA
YTdXmuLbPRJ7L+ZaFvqfWa8Eh0cjgmrhb4HK1PeejSAtkZFxLRuVMU+1r42VUXqb
v6j7UOsoC2aHhsC3C0qLWHzfGPRUWniQjispGsZ33rT3WnkWBZHh3xjHlviK/OC+
o4v1QV2hkZWOxGC2H1DK0FaHzwFLuk3DwLAUI7GVRqFtNWlFlzWtY9CjEZETBEJI
j4PRw0CkXON+gb2gjbzdwlNlpS59aom5D4r2D0F/3xPZEbdV5o49tIwBLu0NjVS3
UthAVGTLRykQTNakcIwuIZaEIQFyIG2UyOGF9r1R75vkDC0XD+Ae4QJgetawuCC1
cXFFoNI4TEC532hybDVjlkaVrX7AB9p6wwl/51/QGEOHG5ix5jy1EYaiDUi8Awbq
7p3sQTVorWWnMKzMBVS39W6A1p8OD88H0oTGV3yy/nJ2IgCnxVEuZ7j4mWeLe7Q7
igvClD862Uy0Nh6OG/LsPP4DPo/NMBkTADD6SpveCprUa1Tylnn4/AoFm/5K1nb0
SnYYt5XCarGzmBC42kiwplfgacpolyvXJ332nwhpSClJhmUrV46Zv0EFLVyxSBdt
pvuD1eYRYfUjTgAw3rRa29EvRLCQxSWNRjaXlpp904xr2sIGabarn5mkVAMjYLeX
WQJ+9LBgktXiwTl7iXp+zJ6+oosmNkxC1i6LR0COFlzi8yq2gs1Oc2t9tC2770Z1
qxoKCQ92AQR/2891Iv9tLQjwyth0XS13nFpcltkDhM+cO9voA291lhr7E2dLazDQ
CziskwW5WfSdAmc0sEOUO5uQj/CNky5geTQ0sMCQO+Ud3GOUEZ1L3hubKfzMUhFf
ja83gO9a+IlTULUUx0KrrlGUp1qFykf9ObnZQbCtj9xv6ZUwC7/pYksD8YFuqI19
S5TNIDC5PlVUEPnFcr0aIWdZl66wqNoq4WIniySeymA+PgDeDMH/v3QFH+q3wz64
4xt1Si2Msh2BQxITbDTJ+guMK0QMqPYwH/FCQHrShuPm/VQGyucaqDcnLb+vPh60
be8vlsMsGitOB/v8FBc6pn0rQT1pnxJCor8zFZh+56WKOkcRE24O6hzOJpYqbUkp
iobuk9vx8Q4eL/cn2dF3ndulqjFY1QBsDTyioxILQmL1MpeTTe3zZXRFPpXDcaGj
CyiZPoY+DpmclaXoKdx807LG7H463XVMEQPHDe+GNQ5YPnxbDC/SlQW9Ukvs9n7L
BN4KhGh8aCIpzKCc/8Of4fsUfT91XV5TXQmVO6bxj/8w3cx7BUB3pXnPdEygorzm
CoUKA5DFq3fhWJSo6umCZDWLG2C4ilruRjWTLC9nata/C6/YyAa3KCVBryP+JlK2
SpfzA0/pZd8dIB0DRJMUnDoHH9nQeA71u7h4ZpXv/RKN/7QdaGwCMRePDW7RXTSu
+nELP4JFMyB4jZUb3JGtG3vwgAmeT537SbrFd0AakLZp3rcVaGIl+xudJB1DOHI0
H2FSUmVlJb/v5dwFEKawmfznXklbl0TnNA1GnNb1j+UXBKos9/yGlTrzvRzROlJC
HhWkoPWSWuo4IVXeoDCx+PNhrtigCkHHnPnP/57k5SQfwX1BhURaEfDTlo5GodBX
YNaBwNFjyaMjH+df3S0u2Sujn/LwjUxiNNqv/rRpzxjq3azQ9P43g917PJfelcQ3
GwWPtzIPCEliKU8plbPq5oIvf5Xtq5lOSzOwQhco7Ip0LvzMRKh+d8NTSAM+M8DB
Lsdzn0QCkQnBjgLphbuK4OvxJPv3BTTo6AVN52WRzZF5YC7bcPsh9zplEqk/O+N4
9gvdiAt858hMV5cfS4OwI3i9gt+LTGqs4Vcj7oLa+8VcOgqqWC55XHXDjYjfMkVU
poRjOGtpM/5cObV0v6N7tMrucoFDbc0C2SRfMLuSzA5cT17tBZGW+ln++cKGZhdH
FWKrBrCFNtT3rlECOItx8jzWYlV00LB9XnNNrGJ5f9km87q2VkfB3xclfPQIohI8
8st9Sk3n7vSvWcwOXeqLW8XqvS84kqV/VwUSgkcz4XQzHQGjRfyK4SWYjKuxE/Oh
FX8xGtJUb0g/LFlZHtIA65kwh3xjq74AtVvTn6+XKXsgcg//jkgvHmaWEf5qqpo9
178uAXFaCA1NN783z9PMSKjMDKKXbDrh5wQ3raQYH2yqg/vxjhw8zvvvk5l5+xtR
oj4hSWsbVntpyWNGgxCQYBClCwLUQ2O0sEuvaFI4TeTGy9wJpn/0GVO/wV5OicGm
vuGftkEOdcIVNyOdsk8YqpjHe8QfMTQmE/x10pGhGSjvM7Tld/Gd70cgUyIXVQPA
2NZvIsgL/WrXPmIzvjxBnUDv5OllX5bENXKhNt5JuBVjmV4S+Xs1yNUb9FIIP0n/
/7j5MEWIo6OWpNkFyAg6MMGgeq1e1tq53JbVcR95htpGvmAKkRFyvqGOY40LZhIN
PIHPHkxLdekqZZJMbPxJiyearcTD1b05NSCqFPPdndaDLjWP35kQfQktR7i6xOEX
Il8PzgoHiVFFUz2enk3XFJ5gnY6nJSuvApKAsb+sxo0h1J5kueTmoQmy2uNLLW00
WK9kg10INsSqUH/zRx12aE3MEI3pkfnvQXNc0bx7dRjONQviRbK+TKVZPMYtsVqh
kBX4WW89c6/icnzzIQSbBD9i3lKYhHUtpIlFc1rLZQ9o2X+G2QacJF/xr5ANdNne
ps2vRrbgmJUdA3lZmT4RIINTiNDeb8Kw0oEZei7oOitL5wh+/ZHAhIwUlRga3w3+
49rh50mrtRf7+G5CWeVxA0psebt5t40fD32fHFSkhndf1bIswDhVIkEVFnFYkeJe
WmfFqujbE13ohHKUsakFi3s9/jfqTOCofYGJbvmRv51n/ClojCgSuezaUOMQ9WRB
e8dfGB8lBpebkM3GGGhK06Tk4VP/AeJNpXfp/ZU/GZyRNg4sFy+dtruKH4ajHHYa
Zv1R000tIgAq+O7L07+d/MmADl6+yAZFjHEXKKlx9axU+A9EcHWjztAsqxx9ncWL
1e5vsOjFd4bzfbg0G8jZSTzwEPOifPK9c1o0xoJ6Ep2ActiVhpbyiARuXCpkba6I
5VMZR0VHGIt1w+26g2wdXp7E/wNkSzI//8tCIH2rYEWAFB0XQyUdKPDS1dsdYtK9
+FtlgJemuNRU0HZ+mDuFcFA1S2tdo3p9pkinut6vT12Ey9lW2RIEjH3XqBNu4N2u
mNDhS7sanQzus7tsZ2ZFcU/d0B/TJAHY8Tt1qmasEI2QHDpHQGLp8PcMBEIUcuHu
fqheBl6+pmYMr5RMAL0FnpJihOlhWYUCYiSbTjjb2GtOaJh1Q3D0qU0BVVEFGUa6
kbnQdAcsmoXv+yHBvLwxOPxbhmV+K7/KZhjMWxgfuTqQQJgR+E4qkKQFyOFjTlj0
QAUhyVmhQxxVuRSglcrVYzKStcbEmlHq78muocObUT8X8UbYJTLkmU6nBIY1UHeD
1Pd07s2AldcIgGrEI3fvOsvrprZ8YrqqtopafwA3JBEs6w2jYYbamzYkKQWcqN/q
CFmQCflrcVWccJlS8YmV+lGG/BMnhrLi80xz/iB6ha5W8taSK15walVjK8Cem6He
9sKubHKdz0TvDSK73/eu0uYzlWxwxwlTb0UsFr+2kQMRleNVz4ITAJ3RvMc04cQR
wBSk0oG7jsyLAWO/XFMXToQiv1/C1rB63AGJ067sC90tvSBZacXu4HAYj88o4VT9
qLkPi1eUP7EsuIpTgxUpj/sNBN3uld8LZZ1umSGD8vdmobqA2XFWIGSTmS+OQsCx
byV5kVMbt3vLCWlfmLe/jLhPKY3N2cUDMt7bxosDP5ZI7U/Am3PxQ4UlI/w4im2j
zyws/9UhUu6ESe6LLvRljf9sj5vwRD0zru2JpGtlTe9r+1bOwFO83pBguMF6tFX6
fw3NvkmP9LEHM3dfieAS5mKfUoAzzfChtD1CdHNC9xsLOvr5AXKaGXMJr4LUFfMT
++H75vK4BfKydfQTOPwvGKqctaDhwKvNb6iDWeVrr0wU8pwl2X+mHRLqt51txAj0
fprlcxgWI8ykbBcC5lcQ2mw7Tq4BeBVTGEw9XS9eB2sxt2tg2zKoMtI9rPb3Gctz
YKOnxkYqteYnE7mNbbK5MT5Mz0thE5LlFKPIDmBTefAe98odo6dIvWIBZgY2Cb0P
gR40WD56UHkP6CQtyTmGAP2QewVi4cj8dyVm11cGEKkHmxCIhXJwqt08UKB5fF0Q
fkK7XrPYSDo5ZFi3J7wSID6edWsK2uLt2KzkinXTUGyu0MDPywEvZBXwoTkOW0P4
pDc+h3CENi9H5Jwr9CwmimdnfonkAcCa7znUj65pbnRQlT0lk0RgBwB7UNBpcEq2
oznemBWdhsswLC5uPSjwmQFPgy7DiFvpiVkF7Bxs2oeDcgyiaaF7T0MFrmJEYh/V
0hKUHqrZaz/jrTGueHVMftokzDTz9M0xfcC/rILEnrMUT2Y75Kt8KrBH36jIVXWG
R+PNqvLCD5hQlqAoyY3a4gU5NgiXCzzdLOc8But7QII9ehRKUUbmhu4gRzQkDich
Z9rtQx1ybcA+1aid39bBGy9XGKIxHTEobBYtYRbPxm+J29EW/sDoUD0kMQzm5ica
XvxKcn/JgDBrsHLpw3ezTznjw2U3gKDOK72uo8/cNd4Ic8FPXPQvgIfNy5eBTh1d
45b69NCcLZdJ4fXXQVZ1WemK8UI8owobIQnAM7pppxATI5+AwgwGw8fmMGtIuXU0
ta1wMXYeW4L7Ch5J3sEVGMAEIuVHQhPyiHEoW9fBgvD00w8L92OgzK408qb7pJ/6
XtU0bHgtHc3W8X0LxSf7QZejeJke7aw8smzszEeg1LH7g6D9xzSDDSpnhMANURkn
qOIC6F0cHKi7eqjz7DdVKWajFobXm+aJcJVnigot15NUA7h8zWbUOF4ITp7zRFzI
wPINrPazQvu6PYHKBs8ogT6an525wKVtGjGBx65qdF5g3AjlUHSKGkIJbsI79FFg
3KPazmE2MCSKB1hDVzmBXE9ZJj6KMX1+cPHIUbedM+lFZ69nl2sqDpzJnUDt+c2H
04+3291gq2sJ7q1c2iudbe7tBNH4EiOIY5DVAffYWQs6X9UJ31vlzKPgWHi6kbZZ
nERofe+CRcQIxhwukAYJY78xSGzbsmv1IQIJNW86P738yBpZzPm+Bs8Y4E8ybEsv
6FnOMRtxv0XRNBTQwpcnWiTA2jP8h0YcnNUM50aYP0zYlynaP8L81bepxWH2ZT1S
+DN8WJ2CPnEtXqxi12bvc5EchjrOeTOYgyleSGrEkAHE8qNFIkTsl95KDSkNnrcu
FZHs+cRJMPcwdy8ggqhLoTYI81EyLaDOJzamYb+76mauLTzdS2c8XFIhHn8DL2rH
KBcxMdgYRhpvANi84zuhjuwjL4a9F5nR6cbsRrJkteIdQTk7jT7ONa9LunEYze+Z
dzRwcaURMLtE7RpprcoJHAueaLLNI5Cx3SanGOwo6g8I53lh21d8cFVQloD5zpMl
7KyEViyoikzuUpFgEtOnFXogE2PdHIuAJpTzFOnRMg7i8luPxVA6RVv+oTQnmPZb
N/0LU04nCF+AvUeOjeGfJNui+M2tvmPtMuJ6AT7cf7Ge5wKl2YT7ycI2u7MfRFJ8
sXoA6+wktaI+NjPPojUX9qQ2nmDzJRNMs3d0DHDHhmRZVwddGAWwATqX/yJMFoIs
lu58Nd2J/wKs+XILu9iOYAD9quBColQX9CAebB4VXp6vUrLknSHMWCmaGucmeNJt
B89FhgtLFhbuJ7qzPGVRyKa2BDlBO8SWvkBcjN4lVcDcqctKh0rlbSDtUvfbT7dK
wV9XUXkZs3gQNvL1zIsQTHTTTSrbmoBq0W0vXQksAQEAjlrsBOQ9gTL1+MIDAhxc
ETw/J3QCpGcxru5LlRe/MhZDYNl86mvp4srRWHmQBpiotfLJEMhpysrVGZM384sn
fPjsVlNR7px+/E2RFlENL81NufYAthzk2+ytb11uaDVF8DD+LRSDzBSGclWqn7sc
3gHfBURq6rQIvFmxoQxxIgCDEijRiSUY49wJlTiVokXxK3wLqnQbs03BnYuur8Ee
2wn8lhI/NnH8txZfAZfMkYsfrmP0k0gZ5pRD82+3SWdLSO/GdwAGSyNrM7WfJXXM
NF3k15HfWIBnyw0rpBd4HW/TKUYpH2Zap856ArA9dKCQiYj1rprv8z+qJ55Kkxl6
eY5TizP5nM0XMTdDaX0fCHQqkuyDcfUne/nzEAO5kfvYma3DTPepO9KexOOcSppw
cn8UjlD+Jg0tuXF/5FNbA5sjZ/Ye2VQtJae0AHJvWSZ0LD/C5e6LB26I3Fpl3cFG
rNUnTWN3bbWn+Hlw/WAlKLqqaHcfXZ6q+bEPfQ0ExOB9jcwaGeQzRFN5RUVWbrFW
SesTyiM6rZVikLsFW8zUFxnw0wYhAGXHasa08EThe3LN8LrrAKIWDvHGvgk3a5fh
JA7YwMIl3LqrcFf8B+DEVKF3r0lrdR4UMepkb+Zz5JQcQ4K9IHdEOveGtirrZCRO
jZqUY1GZfV7hASi4Jl1tMDLvpFjt/jc9uN3ZFQOJttXLcDIgFy/rXpBxHjRkopd2
kuSreyjgcKvXXor6b0kLks4U9LkAf+vT4nluxHZLPDT/eRD/U3KmeC432i4sYLlZ
gHJbLYdow4cmulJRy8oMgH9ANyWzmI5qiH85yCw1dBNrvEC543qvrWXuC2tNlND9
4dEc/2drkPxR8+UdVZWjiMAc1jEMmXZjpQRQGxdDYBid63bFROan1XmkOdSc/Buv
9v1qaSlFXGQgLcupVhtOlJAcxIxl67QpXR6j/llt5mn8Zs6H2REHEDlyzkt4LZEo
gdd9guFLBZRUj/RP7o1bKdoKl3YEZ0pjOflGp8mkGw1JCJOIOK54xEqVLIVaHEBS
Yml7c3ujldHIexXZ0LuTfhxGVbDHXlXo1jRvjTiLuiPMc23lFNCAHeYJPUESKvcW
e6oZtecUSK5gEVHdc2wni/ebIZ7a7BhPvokkJkQ0XGCvEfiT8KzXQx7U44hTQhf1
NmxL9d7GRYMG6w36/6zPIDClwcuHw+IeD+TJvrbYE1X70/6gQMR63sfHEq/G+MSi
A0XnSOMEpyEjmU3RlyB01oD80nHLaWv+oXPe0mTJBvUJLWlrXuACkIbWOA44Nety
JxE7K1+33dSRGcWjRotJzaBYHURrlncQDsqCW396G0VMf6WKU3Ac/iYFgUXXyRZp
/TxSpR/9KiybSSxX5peisJMfYKc89YI/uwrBD+aX3cyFxeRudqbBoXdI0FGyyix5
TPuhPUWLp3crZks9iTpkczTi3LNsXfMqU4GBXdcCDS+j+WbHdVj/UamqmHn3syhq
xHdUiFxZ6UXJYr7m0EXxpmSxAfJ8M04bLnUne4Nkr8luZ5IAtZHfCbPAvBY4M7JT
ukOD2g1j9LxbxJp/xq/j+IFEEfCHJr/izuTlxBtW1XkTCX89Kk3rNeAtvqo69ruY
LGnyjb13NFatnmC7qWFHF5O6AGEQfBXnqHEM+Z0xYGiMo2LAhIW//639i++VlYkO
d+5wEpbtXBxckvTAMFWgMmLlL9XP68zN8WaTtgD0FUap5zeAknSQ4t72bKbTX4Ju
VlEXc/MM6bzy3HPsVUouOMDwUJS7hkGprUteZ/n92+0WOd5C9fFcr6eA9qL3BF+v
elQh13zR1nWTUpb11dQVrSZGKI3IiuK7uneAkky/oZwjS9zhlbGAA4SJfkN+XnfT
i9vi9eGibH/4+CSobBUrkG8ZIEM99J7ilSpbpVQE04I3htkPu1QzoSU94fTt9BLk
9ZaJyvT56CCoXzU5Uq8LodTuE94jjP+mOVMRyRHw+FrHVB7PUwvP+P+gYThD5Ezn
19fpTB/R1+hl9Hk4GrVC6AqE/WslYVXdCRC9xVHQXkSD9r9dduhnHZI4Awqq/peL
U+MsKM8aQJ3ompigPOwz+BjLwkqEndwfPyTUGvT8ouappctkTi/sEl2QCf2UbCK7
8Ec+CQNWhqR5S/w/lbE3TRC+EQ722r9aKg6ZL/BhZzw8RRq0grUsCto5SdqGksQl
odw2jyIRWj4Eg7RrqdIxKXu+S/HZJZJyQ46gArylQKTRRKY+hF06EF9gkfBLdR5/
U9XOnLlh83kiOK2zWlrU9OHmvl4jCX/q7MVrZM3ke0sQ2pOP3kvXdw7hWdFIXjBC
uFUPvoyd7xx5sKrhPtJXfEREXuO3ypP0TbLHV8jKyg+ByXMWTObU5c5D0hVFAE9H
Rh3Kel+B6BNwwf3d8G9/YVWo8Om70W90zLo9QDVJdtNcneOv5ibzLTqv/iC496B+
YGE7TahazIquXMAZS7GCU+dHl65malmZ4zWJj7jD92J+hNtkIAp8lOS/2MAFMtM2
q4uwzq3GbVzdvJ+tak6x2C32XQdeIsDFWRmG2p0MY+55o5BIk98mn/KSvAfSldGr
hYfCBnmidLPjIp2cFi/QuAm2FRK0Ue0NUKI2MMwJ6dc9as0BUucKqm0EQwdG5usb
i/n1apedrT8bRuuSblGMLPycnD7re/akgzzXB1LP8lA5l8qarVBlpRcFppSz0bwU
HtRRLOBo6djQoTjLkrXy6jHRRZ2s9DaxgTJuJtQERT5ISBr1N934hkYelVbUX2z7
29lyGsHeX+TLTA7TFKeYlP4teMXJEow7w8gSJK5J/38Yzns5mOcq5BvtDqqO5Z5Y
RzuMfjj5HUzv1xQmO+dqqUVfAPuQblAOSBG9roK66hq9teYPEOGnzAwrocPv05mZ
r5c+G3fJc/pdznN5U81KdlgIkBXPxjcLA8BlV98iUNT/e/dxQKoIPEWymdyDLpjC
3X+J8r6om5uSN6FiOz6wdOW+vlG1PeXllwHvbaB9Ry84HxALeIGLAmY68bjm1BjD
1tB1//as7WQAzw7PoqIVojKqYkk61dVzNtD2ORS5GGaVy/hQ15+Qy22W9xNNTCyY
FGliYfw3t6o5bD6LFLlQyFD0SRQP1UPuope6ltDRojei7aDTS6kYSFIgcv9HWXpX
5oPm/UPMZiBJc0dwoWZtqOFPx46Ic/37tUXbXq/q2hUH2cfSFd/s8wioP7NPo2NL
ePYhooRnTMtgzpcx1P32SWOgYM3F3kUAyOW1Bm5/4PAhveJeCGVLmbOKqWVzSV70
kVuq2VM8ynsx0rtfq24L5ihoT8Qb1Rua5LcGqcT8jqVMDtP1K0cUyUCKqxngtKNO
QO3fTjbHcsUHQL0V0RX3Rzw1SoEosi3JtmhURaMQzJqglTsbYYMyH+oYU6N4wR9z
uBXpJ1GIVMtYXZ7peXx4gLW4pTayt0YGZ4SkyAXDb1udDE1niib6Zzb+PDC/cAIZ
pw1CIjgOc7g4nmY9rJJ47FvNCfkeelHE35E8h3LUwZIOwGWbDgIPF/uF+4WlEFEw
brdxJAjVmUzutZOEOa5ERuR0+sC1HcficvYrU6PE3Xy5UnjdIIVZHpsdBfNiwHJn
jE1fGT2s4Be2H/tTamvdsQJvmnDN1N7OvsMuguxbCzY=
`protect END_PROTECTED