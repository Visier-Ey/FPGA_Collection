-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
zxAPFCSYOfPJsoD1FFubpHkjVVmNCZDIVQePj8Id5P+mC1UlKO3DNn5B0arRIZLjL+SYivT64F32
KUCPZ+1QVW29MCh0svlmhwCmEf9dOmhaWU4axaE2R6yAAZUFSE5PMqygsp3r3tfjE5UlFoIRqyAy
bIXp2oYXiiS31uiM/ExJl8BNeyayQ5FZm23r18RjdIB3/CkVN1n3j2guY2OZY6R9Vdz9AijyFXFX
7mpSmAwJxDbSkyrdpwBVXBDknDn/jXnJKaxb1C7c6H/vaLN1jZViBSkLENZ81bifB8Pkdv9ceVWj
NAP2tv1Nqy0KXeNNYzifBkrp4KIrhFpuHf0DFA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6080)
`protect data_block
Ba+zYZzBzB6wV+YUrvnkoZJG7eRMxeGdehs8VgZry+1IdQZtcb7KzMQ312v9KcsVDSM7+nZnhsLj
zXH1CsGqXekBtR4YBxbVfXGNypJVqGqF5ijIQqN47lOUPwHpDNc7i5obd8Df1yn0MMLnOSb0AQN+
jKVq1zaEQS1gXGaqg/ZJIYbbafAwtIIubZkXFDbwtplA/ej2P04nFB+y+6c0NeU2Si1qWHFX9ps8
unOb1GcypEr/Hb5SkEdS69B/+9fVL9/9xucvBciN04Yr/+x3sSM3+n5Vlbrcocflz9152O/rROOq
c6zKKqOwbCNzL959vQ/Td+LcpPXUJFi3sFx9vfG3fgFRd8jrMWU/riOoWIi3tYpDWwC/cniuApNV
8X8+GcMVPDyyZMTBMx2CPoYw+f/QlCxIfgozV5OBTnUEo4HAfa56030Ly7bv1scP52Ysey/cJs6b
kyfUyOSoazcarnas/VLsZJazc0HuH+1KMl27RDt1BfbJ8k/VWNijsxIumMnn1JecJIjNAzbuw0Ld
hygtuLNncYhsCiDLu/5fcGzXWPk1kyaCwA1omDCCYFPQL4MpOpEUX8e3i/EFA4kYD2b0elrKRwSj
9UT6EopiMzTndTpLylPIn4KpWUnMVO7hX9vNxV1ZHMW1mBRaPs51H2M7pU8r7YRu+67qzEMNri6C
u4cVr/fVWxW7EndIntSqlaYpqIIJJHwSW9x2iMz3qTg10Pc5SFLoA8jZN/S2roUsJHk/UeU2pYtB
Yu4aQIAruA9/lRldWOBvKtihXD1r61kdsPqyvhrOIkJaylZhPW4pJuL1yukTDUeFaQeQr34Q3O6X
xEv/5iXxKzHvJCOfDWN+FWkikP8lcC3KTd8wm8YBe4BjCxrV5FKVPTNQxvWTUYeUiQcjBr1+Fozr
YAztJFhHMVMZ39S2OrPQsdBLAuEl/ycbkd9qdrctcfXWtPlxEohvxKk+XqPupFUrHCa2ssKxNVZb
VTQb3lJR1Wf4mIOcJgysRIpOWwenj5FxJv6XEyqqbdpaFbAIeWddy/TF1F4zPLg3c0ZXta2R4Ekg
44cOSJyzSxwgKsdi6DJeca/UGhOE0v4Kk4mWXq0ng0FHGe1TKmtJXwOaReVTs3sazkERKiLplncI
YDJwkoUxUSAdzb+KWYzXowBAGHqwGK5UU1yf/vBYRmDHsL0IkiPn5biDNL81sT224/53VOzo2IYq
yftAnsXXP579Petqh6CHpmlKVhB+HMKvnIbxUcRzBPb0e3p5VqYuEDbRTuM05D6NEybR1kP3CKSm
m47SEDap0S3JlLTISPOpztvl2w13p30YPDzrWwBbxICltJzTOYxUlqP4HD6VgdeSGhPa1KnqSAOR
R44o9R/lWir0NYFHTUNf8zfxChb4vTMIi12xQyTNBG103Nl//75jCwK9WXfggCMw3hfsu24RKFWB
QR5cog0EwaYR/GZ0/Ej2BCrtLChT2MIbm3n95CCdPYfzafCx1YnbHPyX2eKqtEwsQGq+s7k55c2G
71MV6bBuPn6t3GD5FCh9syhRGD/hCnt6RdkLKL3phB4/pnDp+teqlNcxu4kTZCb+mTKQeDwa7iba
lmdx3dIvafj90/WgwTC1vufHwYXjgULsuis1hgPXWdPEiBWyEVB2yVj3DdMXfBjtjneEzBtQeTKp
heuUdNXQeAXNysjGLumcArbHYKqG7q+HBOJi1oymxwaGOchrFdXyWwq1sdEUlce1NPF40ujwBXeI
lCnPBLPo4qONWvl/GTlGLUE1K4beXI3JOxyfIWHboKqLArdqDHq4dMya34hNFl3HiUcoNC9H3AfK
PLWxQ8E78SMX9dV58sxr0t+JyljH/J3C3RZ62+M/xM7Wc0NUcfDaP5Wh/Hi3SaxRKJJqXu40WbwJ
QiAyEFKeZLbSFkhpGHArf0nQVGZhLPSoaqIo3/DKnB03k5PTGkg+r/uMYSfiG+pgHX+Da0hekJoB
6MORUcBYfbFRa/4NURBnwmqwH3WM7Fg02GUgx8XyFe077lgpYhL+HhwP8Ys8L3IUHPQcFmgt2jFr
t9UXfl6e2ijodAYI5nLuRIwF87DABG7Rmc6QGhQBL+nPhHK0VUwqlhpTTWsFF8bC3RwHgzMwYK74
mZ4Fp/PWydENe4UpPN0Ac9bM8anZaTHDw67zIvwmGItxO4zVoQ/uNzRWVo4bGPS5558nZvzBgP7a
6/E9tl5Ji6w3sqCzUT3TrMci8tc5YQvIRtAoLyGr7kD4WtINGstQLMapW0/YwiQEwnvz7vuFWIHr
ljvUXUIB1wDPLrtCCU9Bmh36AW+MAygBJyiYn2NCXvWeDsswdniHWorams+h+0rYI5CCUMCXXaBE
mNZAufftdhCe6jj2h6vp4dQypw0ITQW2juVHsokMNAM/f94uo+WngHpl743X6LE4h1yEh6pkAogH
V5qMPg7BWpmlzyvVv5BWYxmcmkq3ZU2stivh79X9pin+L0WoVRrfuRulSn3f3gdcHOpc3gZSfbVi
HOKf4PU55rNDRRsNkPY1h/4qD1Durzf7+ayS10YHGyXi6yivwZWVgEIapdXWtCJE4yBqX+iWpaGc
zt7m24PuGkk5WZ3pK1/z6mgyVgo7MuHTR6njIMfqEwS48uu1Inw8B5syLZ+bOktQAMkZ2G86tZ94
BU7xNUEE0xi5h+0suGcVNCJ/oRDlxKVDmMAmUoof6oxCfUFZOn0zwsj4HLm3Az79UKVwBGfbaML/
+VUuQNzttqd7fGbvxetSlLs/0PnVARwjK9x5yA4Z6COHL/I3WZBbNV0XjnuoiYZbllDAiNiI+NNB
0WZYt/M8AwEK4XrZxwd2bYBt8OU363Bl9NpxRl+ut0h47cyH/kFOcU9z1OTqyPhwlfTTjOL8b1It
H4RMzLQN/O7UMRkZjmPMsIrPunJQ0NVfAXoctwzL7y0E6Kw44UBsyPEYEKH6qrjZpuPF8+obNYs9
nfd0R6hNCagr+5QDvirOmUthy+eE1QGoLimrmzUsaBK+mat0MTgqm6MAoENbZEkYf9SGkjbvadPl
s8AqLso1/uzRUP+2xsSIt/O3HpL1Voia/+ek7N3+GId8edNDSXkKpz2hf00sfKZDr4WCqyvzy9z4
DU6rf7y2eo0HXJ7JmXE8UYMFDGLGlfwFYBn2y60oefiOlBr/p5flUR+DE3EhqDNj9+RJn3f4RMey
BK54ekJQZAAnTlXtfCxTIJZECdQiBg6XUt+2svtFGLiOvk2v3hrMdfFH4Bozs3zv0bGugSHUmfnD
eg0gccca9i1RH4IQV3iXf22//Y4D0AlsIeR6vhs8hzPyDcQa0DqwQ3Xki9bgnc/Dsap0gQkKMuAd
bnyyYTzuKN0vDoDtiuPMgiuzVYDiiJEQEIdK5IeAoXW/+6si8+9pRiYquz/EdilMgsZJokypDcnE
lNX8L1DOMu+QpkV4FApgTcM6EySaXj+J9fq90o+Snsvc25pnv1lQvuozoj9ngw5iGSgX0Av4nHK3
agOgzLMADam3jhRlG5+R0CLWkTKEjNDB/g6jAixaur0v+x72W0Vs0O0gR5E7axfWhOFz0jjhvYQK
CJUDH71w9W5i/GhyojdlsozawgJMriAgJeUImB9VLw4+CQgtYESTc+j+B4/n/9y2MCFq2J24kyXj
AWR7CoUiXNnry+PG/SH6C+qtQ4TRDoXhFRxW8ooOrTndJQjR6XPM+W0rdcEYUz7qZCFbSDRsNQwm
Rzw2bUwxuL+130Y7yKN31eYJnPPTnPRGffIh90L46XVr2MFkUmyqS5rGFoDmromZn0YdeoVRgQKr
DUpBCgVL2PF22xyT0HRE/1XWd0ZQ8UnMiCFYUY1YJGfL6PC+DY594QBb9swxPr9ZttvzWGnKpfng
jMmHSrKAJNO4Xz9CTbFb0a0xBfA/P3KNjJSFHfo0TVuLO5N5NFfdViv07Q+6DnVFTsz3soP5E64O
OsQEpjUhwRzqZ0SYs8Wgvsl7E2J788nAoNZ8IGLj5G/7tnSx3hLyqs+eN8xHZJ2UdoevjuKnTqFC
BrBt4I8Bg7TGS/5Yj0r1RKQX6YjgJPGdxcAyedncRQFTxAewaeIzHQpSlUXjZHYEMzJg2skY48V+
LTPQCj8zk4ASrSDxnPjVcjLPT084LlD2WnYzaOmRJ99DahEqoZiSBLKH7c7vT+6aCUfNmI+AiiRB
rPpjqBS8+gsA4BGjOCIo6lRq6M62cf4bd45ayDnAeyrUYUc6ARWGZMNVwJDb2/1mJMTK7TpotBPZ
jadQonDoQpfWZtwmUQwcdAdtST1CEC1WRBT1D3IBi/PShRB8/YcnCjgkYBP4G6URtawNAMtZrWWN
wdU2j0fxCLsg6tKkBHMCVDtCxPhc84LvJt8uL1KhCdigh/5BOeyuhmWhCUL82WFRlxolQJOsW4T+
RVbtMjAXxrVWE+T2oorkU3YP7MZmj6okx6stE5l8H94pojQch9kntsR2yVzrb/ahx6piNqvluiTK
Wbn6P9fGY658CirEs5Vh3iiJbQI6RnxdYraUeqHwrP30AKzLtbFXSxa+86+Wych9+wfY5E53kjfb
k6XiTt/8FeTlxSbUU029QUCkbq8WBWN0ilNWJ0iXt1kk9ra7Ap82Ouy3nKvdF1ZPbgm/kInVJBJR
O1eTMF3PRBm6ecMxZQtYN8WqVP4xbemZqPfuWM6RxVj8CLVyUjazx68psMiQAbRBwi+882WZJoUE
KfWcbH9mgS9l23jCib1C7ePjYOitdXr1wZjjbWY/gZZl6KzJ6bOwYBiKdYhGQwgVPM9MK91JoDtT
cQP8/U0hpzUT1aDtiAZWRGOErIo9uoRDJb/bl4ZtFfH96IdiCJ/oN49IjQ6yINlTnwx1MkJT7xx0
kFH94Pxv/shERzVyUqHq/ecYN+jyjy7D/MpWT7BghNgeIR99tCitsrBX6xp2WcEZNRAl+NScwXtH
ZlDLEpL3HDmHSOnlmcPecUFs9YzuFTThlEnIyUP5CFwRj796mQLjrXQW5fWFH6w/hue9bztc9825
72nGRYlorwBbcgXgG9r2EqCqvZbjB7vN+TdtVf/2rxiNY7/aVk4J+1dDgCmH/5oIikPYw8SS69tP
QFsX2YySFcqcbro25sNf42uf61GpFuXiBRKSTfnuIKlQsWVzdEe3kFr/4uUdrXsbH4K1l9Vy99uQ
hk4wfkHsWZcKz8+IpCYNfnFPNEOXpXm5U/6L2EaHqRnEeJnaczzdGLHPoedZGdVWNB3UoUqFHPkj
WYVb2tMpTrOJDL2GgWNLN/rfBpqzbQtETPCxfQk8rAi/djI7y0hC+Ow65XU8dCF8ehkQCuh2L9tj
Q5NgDjR7KrWHY2ngSwwJ4PHHSq1bQd07x+C3vRXMmgLrEZ24wmeWM2yeNkkJCts26mC+/qVkgI3+
qeBNbX9awI/oqdembE42hHtMkEGpjNOy75IcUEq3bq+O2T61/AUGEzDbJyzwRo3sU0JhMZelGvLK
iks2ZvycPJmyvvQFWLSdmIfv9vnP4WCM2wRZRiK6JVq4gYZxM6T/2p9K9wxEJyKPckhh+YkkKVDh
/v84tCKU+ro+hwhYywI42/MITD/aO9dkHgHtwdTYCAFWmkwZD5J1afLRkMkKC3t2oQ7APoQqzHSq
dGyy37yIyjMg5JCavnBh0DyKA9FovYRFvNkEuKDtHk35J14+x5z7weaZMvB9Zyt5EiAa38XR4YyQ
Kz/PysN1wmVdJVeD3tkdbdF3OpLTWpmbxA8JEInx281a8FEbx7M8w0PaUsApjcWuqkCu6OdWBosq
ps1METgrQYrVKPYnL1P7oi7PBeQE/LlIhD9ikW52J20HR2USGX1Ll29DZoRs/YGA6nRsdiper5bw
ez0VAG7yYhpsuMinPLlS+oJ3kL7aBLvWhJUKHaY0QLQqi4m722gnoV9aib+X6WnwXb/U2Z9H8RyS
PQL3urwkFC2yf6Bi4owQQUhmCEOXWRl5r5c+5I4kLfVqgl0sI+UxGmpgBi7HtzTK2uWcqjC2rGG6
/iP/pJRjFanmWImvIIr8JZwnLfpVX+7QWQtdvjxio/V1Bjpyyox0s79kykNSiVuIS5E/KCiv2nHM
0u2gJqmnvxf8vwulJbynhEkoR+WLizVwaHV7K7T8sRjKbQzjZOPwuHGU4qSDU+yFlambqbKIAcut
MmE/8sDDg3gDdBkuHL70NMhPCkHPQwwAoRm13bcACIVIrnukmndHGNoNUUMjvXHb6VGR5JG9MEIj
F+boxLcW57qTulAnmXubvqY/o47AgUAU0Se4biieHtbCuGWLtvR6UMlrMjduiDmoN4zxqzqd9qVp
gomcAgc4lJCQTX2CnfWZRi3pq8uqSJawBclrgufMU7uGRwqswEDcMKRsc/3jwOGKT7kXnx2BGufC
vU9GiPlsOVGuu4BcSv6vWECcI2oHmNK7CNbND7IgL8GSbZTspzqYWYSyoU28v1+6JIwGjNfR6eu0
9I5EHneFwbHbzeYvcZQIEc9Xf8h02xF0oxgQyfwgvDT4+ePZZPMPjzD2EsSGKUBDXR0znTyIU4/5
MDrWJLcIl0MDBI88IlXc7ACUbz0603KPU95CmHL8VZmJw8CfcrhEskP5bjoDLljRPzHSrEKrmiy/
pznoD4lq1i1pLQ6MnZUKjcI/bf7tTND93jLvd7c5y7/LDbW04cpyoVE+wov2S9/E3P3JxT8p4Zd4
YI3jvoAfiv8ypIg3LXhLO0GoOYBXvHu4ow9iz2mgDH+yXLRQy38KyD5e7X8qeFeOX0u8vsKvyCt8
ZUmE4IY/m7zM3d31qbNzGMUmZsvNt6eT1dd/vy+wm+1FwKX9Iqm5FPIsMu72CVOHynNnXnR0cu/l
OmyZzezzUcA3AGEcIG4fr60X4iRp8eEXZybTcQ4n15Mk5vdNaGj4vHpsP/yipIMR4hHfsSVnBzqt
hjng9MCYTPxxztZc44oxGtt84cg2IUfpIKEyofkpSMzpWWinRpnM0QqODhkcnAAHnx2LhUHvC/0p
JVdCn6H5onnnFOe8swTEpovfL5XWITkuWJyBwkMC487WaKPApx1d6QkBjHNM7pEIVaei3l16+aGQ
IMbRvB4jsN+9mJQbame05Wd9Sr+Pk7qrMXMY5VxVr/8Y/PZUWxkmUm66PEwvt9DzbsdeYOOnCXbB
cfGRIdaWFk1noWc/wVabBV7B1g/D1W/G9+jfOJrQMWkht8p2nKN2AEXOG84j0yH2Phir95lTuvVb
qqnvVhGRQD+scpT1fo9FIjBgmp4482WRxcJvahiI/g4+wKzqZ0kPnBp1xeEN6tafUx7Bt5r0zcAW
xj+x1GF8EI1FTnltVRxld//b4sQu4xqY+fxRAN624ygDWW+FDK+n4WT2D+pVcIoLOUhXuG0Uwqg0
JUTulSymjKW9PsfUcaI9kvHFWzbZVZCCtkoU19Pvkz68GxZ0mMrj5/S/TvTy+KalsxyMqiweUkRv
cal2l0KRHhkghQNmnWVbgyPsFCHD5XorbA/z9Ls03O9G9UknlJhkVyGImyVVLMygXBKkcUJYvKY/
uLwOIrp/P8eRXWs9AdXA7ouW6TMgt58rukfHbJx+WnJr0GHNjqxhg1ehvOXms+mK4YrioIhp87CM
ZZbHMui2cPlDA2kw+FkpLIKcZ8GEm2Gl/EuWr5Wybxl9PLlZF+DxlWM39ZgcOc/DoMtc32paf4vH
vHTKdDQBPUqmXkTR2ifABCM0fZOgmRi5eoG1S7SFA9+nAr+hD8m+lnNOrex9jGNMONTHd1+6FoRP
48K8y+cQLxHGp67S153xpFSZx3P1Vzof2Hy4xhQG1g2n9pm+NuI4pQ6qEE+INIagqdhB0Ogjjt1X
ETIlYuG/ZfUolACIftDBdBPx8bxBkEFzVIO8uO+p/mmTUJN6HDg26GLfDTW8vi0krykKGBBA9Cj0
Afu3MxMZTfpJM8myxZngtsFu8ZKPijt/vi9FbXMlJw43wzSwGEirzrVGVABadZsSz7iyOe7T7Q0u
+p/oaw/Zg0xJgCJzE+VGu7lzWYVE8ESReA3kZB0AbtyIjXcY4MoYu15P5EvBqOA+Iq+Sbe0Ixua6
cAC4ZIUS3cA6eDXbru4GEQQVZs3ud1oeTvA+LYFYyiyp5U1Sc+Y=
`protect end_protected
