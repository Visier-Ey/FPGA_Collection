��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���d�v����0�i�=\��A��?��� (��1_B�f�	�Ѻ+|n��y��Q4�]�aY�����*2�y%����>��������K������ �
�D��z�z��C�y�B����
_�U��hkF<�~x�ܕ�c�[�ק���dI ��Y�l�BY�nyWE��:�0`��}�a��R����1.�_E}�>���ۺ�FI7 D��5�1k�.�@GdQ���(3J��U���6��ɒa���6?Q0�^B���DD��H�����u�Q-�l��ݵC�=������s�մ��<��CANjH]�o�R�?�=��[����g�N��7!��'�E�Ջ��
Lz����RIr(�M/f	�c��4!
���4�$x)0���x,�4�q��D���h?�/iFza� ��+�I��g˵�}�}��_�8�P�V����:a��&�Q�4RtN���ka��қP"ĉ�G]$F�S�@	�Fy�2`�E�J��ām	8�b\v@1��%1T�CY�А��״��t�>׻����K �Rq�q�ꑣ�R�C�L�L�/�y�ޚ������ǎ;�3E�����k���Uݸ�-��F�SwxҴ��uN��sRU�n�Ւ��]�W{
�cR���p��i��� �{T�K��X�nf($[7}����9Q|	9)�`{�q%�f�;��=sTz㉌����94;�����QG��U��7E��\��'��.I#�`���! �4˟O�-iv�1Us���޷�ǰ�f�?>�|�[���U����2J�@�[���0�D:D�n�Q�a�y"d�{hįB�mXݨ���|�BB����?�P�d�崛����i5�;��r�Ѣe�T�C]d�.ױ�K��9)��v��{c��ɠ9��q��I~5|��
�.a��5W�����P0*�0�G:��Q>{�Z7I�Ć���(��AZ�o
4�p+%���A����[6&Y]��f��.�Q��P�8�m喃��)�K@�����^�jO`��l��r����$͊��i
�d��}4�K"g�& *[�}��뚮����S�0F�̝�D]~�y2���/+Y�Fj�O�[ťw;F�[~���e������(�[�مg�fݬ��J^>��s0eF!cڝg�/��a��F�p��Nɡ���D�G<U�nl�z��*ř~Q��q�$���X�����Y#�&�ʥ��%�#n�� ���Ve�4vtv��'��[<����X0�l&��!�dU3�y&}�9�(K�W��k_�*ŽL������U��$�Ǜ5)��^���6�F��i�ժ]�sC�*H�jŗ�  �
0�{j)w�O�ȡw���� ��C�OC:���{���x!(<�mk��w,�U|J���?ɇ]ݼ��U 1u)m�@m1e��A&�:��w7���p�p�G/��QL��uچ�c�7�"_��W��(��\+9�h/C��nɡ�zC�����L�3�P�dSwr>Y�H�/2l��P��%0ȋ9��v��z'!=Lc�� Q��V��o��twU1!���Z�}?�K�E1�
Y`=n-�p9��8�U5�~�|z�|~�0Âm,�ѩ�E��|���hi�M~����2T�t�g֣�ކk��33�%�w1yZ\I�-���A�Ȥo��<��F���O�������=������i�N�mo�I&�A����P
_�>�ne�(e�0��l���ʷ8�/'� �*�2NF�W@�LP��N˙����Y!�K��-�����1*��7�#�&O[��h
Y9=�If��2���1��O�r�<������Ƕ�Y��(v��j5"��e\����$,��\�IL���gI*�I]��w ��{�C�����"�/�-SU@�jt�n=A�aiO*pŮ,���2�鴊�����I����D!|�rPBV�:Aō�v�r�irV�8\_i,�}�+`�3���@��:ʟ7��f�M��ާā9��������ɉ'�f�[�D��$b�ʸÓ �>��!c��OEa�ԇA�`�y���H?n8����������F܄���y�|� �@�J���������Z�܉��i]j�Fz��¬������Ǆ�VW�1��n������	������b���6��:�P'�Tw��ko!��KE��K���6�XF"�.�k�G�jë��:�S�i�= "+kJ�W�`����/��Os�j���'�����n~G+���D�^�_ɇ2W�5���E��/B�O�����	F��ɘ��ޓ����T����
]j�5�1c�V�v2c�����9C,ڑ��ɚKF����e$
��${`��D}��ڰ.�a��f���0`6�ۨ��J�h+,_�&���ڷ��.�d����]�TXs�z)��T`�}�ܒ�l��6t������2����>'�Ɲ�}S�{��8v��U����3�C�e��=��~dt����U���^p_4�|��X�<6N�/`wg�����M��I��Y�-T��7�ӽ W��;�C�~���e���%�|�00����Ud]�`}r8s��4�T�}���Q����/���Q��2%?Z���`J��90=���i^M���C<B��E�J�*��<ۗV��yy�e�Ó�&�Xᬬ"��@>x�@=����]l�awN�£/;ۑϺJg���%�l�X0f�Yc�xM�e�->&�sn�	`՝���u!�rs�H�i��*D�\��� ��'�E�y��ϿO��Kթ���q}�vb��-"��O��	�=ع�1�1�����iA���IxO ��+��!��{-\E4��/o��\,U�䝜-��u��Q��-6+��S?��H=�Y�ur6�����ˡ	Ӣ4 �o�X.�5�T����U�v�4Cʦ	��M3=&:�JW泄�gU����������9�0��4��/�n�W;�bj#bYu�Ӫ$p_4�������P5��S���qmzY���r?-X��w�ƈ,'�T�F��}.}��\s�-L����2H�Ծ�/�rw�-���O[�z�Q�+��k�.��?oG3m�yRJHUz���7�X��CR�ʎ~Ec8�S�1#�K�g�����k�_<b�~�P<�X?_�����`A�3V��-N55����h��휷b�a~�`�A���ՅPr=�B)֞���sϙ���D��A���(������X?P��a�H�Yhu{��%sΆ��*���r/K�Ǭ�ui6�5���׍���X� ~������i�$\��=yQ�*���t���zNZ���n�+�#��k�1�}N�� �s�o�r�l̵��&*�}�hI;�(�~
�҅��N)u��C��*Dx����1�D�N}��v,��~��O�@�I���U�$����`ڲj������uv�~3:�%�ͰQ�X������r��~7����^�/�ARղB�n:��ۺ��Eh��%Q�����!�����2�x{�e��Y/){��aFP�?	KL��h�@	���	m���c��gT(�i�]���ޖj�Xa/7�.���X��FJ����@)�f�&S�+]�5����U#jRQ1ԯ%��w��c�ް�7�fb�����Gn�?jj��"�x�Oa�X�)F�*d�o[-�5l$���^�Xy;
�� ���b>���*;�$�
�k%���o8H�4h%i}��B�}�ˍR����F8?���