��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F����Z4��#����m�ǵp��}��a��1��qh8��ɞqq�Č�܌��ie������c.�2�	�`		_���ӣ�����_؊����=��
v���ձ�������v�T�S�j��0�E+�X�뷙�S�.s��������7��ڳ	.�0�`��k{?t��i��-��F��I��1+�/gn����詳Q�Agm7Zn�!�
��$�Z�+�
=uߡu�z�]-���z���xԨ
���݄�	��چ��C	�����,J�򩕉���;f4 �!^?wql
��	8~�M�`@�����mOp�J��t����,G��E�j�׳=�b�����Ԍ澁��Qѱ�j����~���OK����EF�,zS��!o�.�J�2Oҫ��k@����IB)���V�v�BKӟu������_��?~�^4�.�4PӼ	wIH\��rzi����dH�����Ȏ ����B�a�&T:��'��s6�00�G��=C`����Õ�_��r�~	�1�,�G5x1��'?�w�n�j�F�ۀ��f�q%m	m�O����aЄ������N�-p�	~�b���ͪ�"wt<����{���x��a�M���T�Le\����%�U�x��3��z���Du�EQ�bXK@���V�K1L*9�Փ�:���_|��r��ĥo�wYm�z����"QHՙ�쎱ꙋ�{Z��[�rN�j;E�� �e�w�C����B�="���Ąm� ���=���dč����	�`��h���;�n�՝��s4�h��/�^�7[ɂ�0�/+ڠ�
��I�#�q6����˺�dc>#�������)�
	�����g��1i{�`����Tc(Yf���~fYF�/+ྲ�o�}XӃ�|�$�a}SA�{矛�
�$Y��LQP�ʭ4A;B�A�U4w��iG��P���A�,�h*��:�?���a��om���8�)�V��_tr����j����tʊtj�z�L�5?/�}Q�خ�	��F�)� +ɉRr�ل��[�9��\�+��)M�c Ew��s_1gx*JH#��iK#TcT��omia^UXu�v��{2lvf����fI�ǖc0��X�E��]ՙQ��hxc&�Paǜϳ�F!���p}�e�p�y�\hU`�#��S��i~S�UΦd����XT���k��?�}�)G�/t�?(�>�<V�N`f:ʈ%J���e�y����+Z呟��~�p�~f��K�Y<Y�
�������C�(0'�R�]|�N�K�2�@v,��+;�ґ>��Nr��֟���n�J����8ѵ�D���?uPb1>Yd $�����ʍ�a�t�<w����K�s�y���Sw�+I���h�<�)�UQ����HO��� ǥ�J�"f�xt�CL��3��QT�WF����Q ��+u`���z	�����6�]�a`�d�f�ML��Ԭ�b��Ĥ���m42\O����|�y0�@��9tx#�ŀ���4��Ȃz?�nH�����KB,0��W�(�x^r�I;�D�Z~zUaK�8g�q��֭�Y��͚.�j��k��CАn�~�c�޷:>�j��qb@6��ڿg�ÕG�w�q/K����ۈt,Av���:�96�A�&L�@SX���w%�AI�TxUg�q��1(��[���d[�@�!���	�\�R� �[����i�lD>ve�����`XR�3}�� q��qâ���sQ��GL��F$*���o�r�R�-Q���"9�L⿩B�����3c}�����,��-�kѿ��0�t�������N��JGO�J��/�ӹuSB.bT`��H�M�P"���hZ�0�DGv�5�u�����M�<z
�8�B:4��B;N����y�a���1@�9x�/����p�ý�"#��g1-���Ք�R���Ȃ�{��ҥ�� V`��ӌ�=����w�h	�F� �=� �&o�>����:�5KN�2_�ّZ��z����VDfU$t���L1i�_/v6h��=��U��M��Z�y��Y�F���_OJ�C�!�kb���� x�c��E>R#�h���_�f��A�Ve�aRf�&!6���%���fS0 y�����(�ya�J��SʐV��t�~-Z��F�KJ�+�5����2L�]���5���qٚ�%!!u/G]�4�@`'y=�������`T�K�2qO��T��9�TF�����οPG��#�V��_�9`�i���^ˊ��.g����Ǵə ���Y�w���]N~/�k��	�?���n�oQ9��x���͹��߆6f���+���Ei����I���L���������~\.�[b06r�{pـ�ߎ��[b�K��/9ʹσ}p�亝XĶ��I��p}�)�%��]���^;{li[n�n����{=]�(��|T���}_�F){!UIB;p�n6<z�,u�l������x]��"�������:(E���?Z�h�nd��7�;��5�NZM߭�i$�fBn ͡�㹧�	Eg�����%4��&��&o�Tl�&9[��	ˏI��#�5��:D��f����б����rb�q�yf�E*h߳�<��ljxDu����[يs>����s�~h��p����.Je��iF$���˧a���>=�Mlְ��)��d�J�����x."�ʧh�9�~��[�&��X��.��h>�瑩��zs��а�Pk���؜��"O�j�e���p1Ə��s�u}8�nﳦڴ��"N��sP��넾�PB�Mb[a���:y;�.��B���7��h�2�e,H��7����[�*�Y���w��@|*Y�����<�kV�U�h�}�M��'���E�m^̔�R8�֘f����֕����i܎Y!��� ���C�v�c����\���f�z���(0m�,��`�x/͆,�H�2�[�!�i m�Fa=�|� �w:�7@��N�?k0�.O['�����������+
�fH��������� �E�qZ������|������$Ixk���SA�V�.����R�{@���є��ˋ!��E�b@�v����D��z6D��|��|�\����� ��h�BRI���aݪԱ��>�G�+4��Y(����I�Bc��腭��A��]��W�E�l��\���`�E�r��땆RM�V��.�R�i�B�p�mu��
�>�6�4���i!9��@��������5KZ |w�{q*&+@h�)kDg_^Z=��U:0#�;[���6F�>��WE��K	�(v��%c��<�*_��U��On���Q�Yx��+��K���U�@{���G,��,�(3���)��R6�:�K\vQ��7�q�_L�'\~d0%��BÐd 	;W�bs�i��iڡ< ��Pc��p�	L��(���:;���@s-	�7���A"��v���1Gn�%M�K���q�_�-}>��S��m,�.�;�P�mtʣ�Y|4�p���%�y+s%���j�c��v�K�����K�(�'��KD�抌�Oë�Ï�A�_��{�ߍf�3♉^h� �e7�$uJ5GqvyP�Φnu����gj�P������,��0Jb�O��X@|r����Is�}�%��IwF���o�0�yA&�K��{>��JE\�2���/�DP9]��͍W�*�eĹ�V��h3�_�:1�p�B[�#���%C���c�-jT����`�P�z���WW�7)+���j�߹��&���\����4?�/��x�����;�U0 z���8 �������v��H�g���MH&���]s�emmc�5���c��E+��b��h&�4�1e�|>~P���:c�#�߼C1�͌���!`qO�����x�:/'�G�*,�5e����+�}j~X�d�s=g�B
�;L3�;oz���0�
�f?d���ݚ�o=��&/}έ�:}
OWR4�u:���lZ�1|<�0��hc���/Ke�7�.gM�E\�%2b�6H��L����#(�a`8r�yr�*�/��>(�j?D�'	B�>�'�c�唀ݮ���k�04���zR��I/����`�P0��/��5k[W70Dߴ�uN&�ڃ�;%Y��~S��P2��>"]6t�go�D�r[}��:	T�ч��I������A�SH�l>� .�x���ڀܕ7wis�j@ �y^".#�ʁ���o
�b�K�S�����',/�0�̆%�&o�F���L�gm��I�p@5e�b����2���k����z.� �cQ��-C�p�C�K�ҵ�q���Y?��<ɭDyf��խN�4�v��ږ}�Ȍ���x--e��DNi�u-�?�t���t����)�Pbf�� D���Y��<��R�6��Z���|�F|D0�Ͻ7�(LybFvvXu<$�ɘ��m�\,��L����HԾ���B���-k��ϣ���Fs����X1k]����ξ��8��CD�ܘ��W@��Ѵ��*WA�3�a,���-�cD��HOP^��O�y�:p�<Eq�F��8[�z�X{�`G�9���f�pW!�T���L�@������L�R���i����2�+N�a�.	�4���U��ϩ{�Qrp�/�Y]��~ۻ��+�} ��e�_h���t^EB�2���A$�Z����8�mPۭ��w��wH�(Mu�+�Rj�=��r�8 =B��b(�aU��J�Ϳ�K� og��g�7�G�y*2�(fͅ�w�N�:V�o�N�A���׬-d�]�L�n���æ�e�	�6e��vӰ[��,Twg��);M�ndy��c�<�7��Y@��U���-Ք	�6�����88��񢧑ܓRv��8?�:�:�:�PK�fc���"4�N����y�E$D�*n�ګ�`�ng��sa�^�z��3����o�T�����O�_��eg'����xz�򾌹�V��/z��y�����nU���3K}��D�k����g,=��,�{G@3<&`�]���Ȼ���ID���Y��h��n*#Fp�mo��n�*�S^\�anj����s�KM��,�	 �Y"����ظD�B���y1OFәm�k���+�:���L��*�Ϝ�W����Y���1��������@l�>|��p?}��z�=�d�,Y4d��=?��썘�8H&ch(NW�1��ۦ�N�<���=Uq�A5ϛ�q�Yт�°�X�(o��������+�yk��|5j=�rx��UhI�w�%p���+�ӵ�u=�8�J���v�a������1��q*s��MK�Y[+�;[��4��^L�5l#���&fh�^���.yh+�i�l��Y��E!"�&���/�C�4Vʌ
�d��ƭ]���1=3Ϫ�ӆ��k�VS�\OjZ���+r�!��K��x��LF�����d��i�m8@����*�X)q�GLx��Os��5���8���BN]���7My�=Gq�B�������'<��(@�Ę����ahK��*ק��}���*jjz�oΚ�����.-�b�]1�������&͕g�K�r�4�G٢X��|�Y:��������3(�x%�,Y[��~��hب��g��ڦőN�N�*̸oh��`n���_�Z��d�qR�͈<��~D�ur�!g@?G<�ۜy�,Us>�@v�Z��d�,�!'���	[�*�����tO��#��i���r���E��?Z�{����o� �q�jm/��v�)p��\�n~|?D�r��1
�!�$r��2H6aݶ�"�Hv�ַ����q+$�Fy_�%��t}J4��D*,�h�@��x*.�NZ�,ʻy	*B�>�l9/V#J1m���ꘞ&��Q����ڤ��<3���+�֔X�D���vջ�M�/& �m�bs����.D�ao)Qa�ՠ~'���s�:L��X���[�}3ڛ�����C�Ar$4}� �������爼3��
�`�8 ���JS3*�\2w��
7�A�\F0x�iJ���Pc��;`2����J>E��`"�<���g�b��{�/���&[�u]�D����� 42�v�{$��V��a<
��Юg�h�f��x<T��	#���z�����}Bo���["Jl����lj�q�xcX_��z����]ɰo��/�9�\'� i��A�%��;�j ��Ê@;bZ�z��]g~o���lSQ�
�������X�>Uܿ���h	ao�k�!��75"�j���Ʌc[�o�m��&�\��Å���}�����'�T��!���Q��ZsOƍCݷ;�i�|0/l�۱�-��ڎ�RO����!���6�����\9<�bD֔p�u��B?�r��њT�3�]��2���6O̕��h,t�P����>Pa
@@5�������Ao��6���[�=J�²#��� c�Lm@������,��K&�1l���Z��;0���Ie��̓8^)�3~������5��N��B�~��64J���=��|�H��<t�:Fj!�v����m0sNt|�Ҕ�����"��@��\��P���� �S%�d��!�=o���Ḯ���8.9�.@I�U�a�bD�hY=���z����:������S�\Q0Rk�JS9�@4�����E\�6(v]�fǟ��.�H4%�O����g� ;���yh}�Jm�$Y�2S����	�#h��:m��8�׆�63��(7�|���a��p�� ~��B[ҭ�W,ȁo$u'�n@9�1���	g_9�q	��R�c�W��^����Nd}���9n�Jg���n} �>���a0H)�5HB9D��]�Wv�h�PG9|��u0R�Ʉ��]��Ք�é�/����V���1`L�?���2ZH^W��, %K6We$�Bf�^�i�H�P��j�� W$;���?�ʄ&}�~ȱ"���y��_�����1���\�!�ն՝� �ʾ`J֡���`m�7΁S�ԑ�1[�݃��wp�,�(�]�'���M���S�X:9Yq�b������s�܅�F�?qVn�G7��AB׵�{7��~�ς����1�x�2�;Y⨡���?R����O�Ŭ�H(�؊(���'}XX��^�}��Lة�."��^l�p|���g�Y9��g�f�!*���g!����]���ٳY&�2e��U�n'�Ȳ�{��HAʿ#��	�l��Ө��.��E]f�F�ل����J����bژ)��W�2n�,
r�FZ���k�BՉ��۾*��slR
c؆����r��"һ�xÀo*���>N��y�ø/���t�����˧M>it�B+����Ej��-a1ٸ���" ���q�A��J;�Շ��-'*/]��Zȇ	�d7y��t4��c�8�W\w/B?0!CI(�~̑�6wM�E�yپا�b
��V��M<���g�Zb����C��OdJO~]��)*���Ѝ�G&��k�]���b�}�
&��,��ʬ�e˒,�D��à�ru��5�-ʌ��Z`M��`_���oC�t*QJw�S`�(�1n�At����1��RCp���)�h�k|d;{�u
µ���}lQ��e�����6&�@>�_9Q�x���'���34GIj w����������Ι����q=e0����!���O)��K�X{��ċ1�L���o09c0~/�����q���u4c|���Q�'U:��[�h��N�Jre�_�abޭ	��E��ٷ��y-�"���/�� i��c��h$yl�9�t��O�e�tz�\�qݝD<1�f�ԥ?�/I�ŵ
g�U_��x�ߵT^�/P7����fk��9+�D�Z[��U>���=�b�-��k1��MC��!KX~7���k��?�DfT�q91_��o~�eF��DC�C5Ʀ�����QtK��%ό��y�����Ǯ�"�D�v���D8�z�=�� �E*�/ɽ�@�x[��?��[�R�w���`����+Y-�DMe�<0��ZTB<��v�2v��&���� l�%�8B�w�O��FU�3����'V�m��� &h�_`3��@5D��Gk����_���3���g �$j�JQ|��T�V��\WԤo����~	 tOZ:
=����Vŧ�K	�jn��XtQ�w�����)��p

>��Wq�E���iAl8�?���h�L�5�mQ�tŪǇ_��������_�(��cx5���1<kI$'�����H�9.z1�ک�Q:�E��������<�Еn�)ųiE��gP)X�c�6��b�-0�j 2 �kP�����ܮ94��XZh��.�'�꬧��9�U�(�s5F�t�{C�p�+�t��i����e��)��Ǥ�Z�*-�nz��`�H1YME;q��q��
��O!�𦹅�o�잿
�1�nڞ��8�L��˳�]t�˪D�����$�j����~jF���q_���l�G��0\���K�xg9��S���U�g�����4�I6�X�[צp����@7�����
�����9�}�NQ�g��t�Z�/���cT+�Pk�}C��d��4��"��H�*a�)*�Tox��d�4 ���^*�
�����C��s.����`��N?T��C%6�0,�h�P�m?7
\����o�^��uu_o�˶T����-��� 
N���#� -mQ=�/9�>�M���ь��[�D`���gg R	�~n�+���M�H�7Lx�v�?zD�׸�xě�Ѵd���y;K�w3LN�L�=��_򶭌Ep�;�J��.�Y�v{�4��aʨ漟���'>M�^7_0Ci=�G@�Oφ��/f���#P�I����s"Z���ʱ�����#9�y��R(�P��e�4!��
ɼ��?V�Zd;O�1v���z9~`�_��	�l�{R�O:��A	\�vC*~�
P�%]8/'+�������K4����D0��N�q< &�謀�r��� vA�
���|��Ř	��@l�9016c�"|	!��"�0@�x
���fF�w�nU�jR�wwH ó�w�h�[x{�����5�u����ۄ�#��BQ�_[tv�H�C�"Ŵ�Õ��`4H y9h�jl���A�4k����ʻ�,@O�4г ڙ�Q�x��ƶ=�q�6�3�*��u5Ѻd�Eu�f��{N����%L���?�����!7�j�V
Sjj���Ta�i���n=�y*�٢�g;�K8�4�:0�J�nS���;?5b��v%ޑ�C�"��ho�S>�c�H�)��A� �h�Z���|LKI0���{�#�L�;�քJ����{i�}ސ�*����6�����9�bQ�u�,��+t�T{�~�A�"T�Mq�}	o�>�
.^��K!ݴfv:����WKl��Ó}�����kz=9�ِ��0ިa  ؗ�w=`/��#�!��ob�q���a@�a�Մ���wmw�r"sg_�ThuVyU4h������?�o}݁�ވ�,� N�O�,����X�&�ʭ�΄?�Q�1�7@o̧^�Kҥu�,Q�YU�uà^��֐h'Z���w��?`1����T�Uı鈸��sv-a����j�L��.u��S8��܊x�J����^S�M����^\e���0,�tOFc�n�×��V�Yd�����^��~�2HL��rVцB�!ZR�/����;�c7s��t�!G:�ʛ��dE����֏ZЙb�r� �u�D(jt�|�R�S;	��S��:k@��ښv�8����Pv���)ˆ�d���
��!��=�Z�3�G�|��
wQ��od�����
G�.�јf��a|�\s�c5��ItH���9s�U��w3��EZ���a��h�ߊL
�QW�L��C:�����9���p�
+g�<!;�����CA�º�	#H���5�v?7�<y�5ӽ���,{z2T7T��#8����/�a�j!+ �S!.�TD^/!U(t����|�Y�/\3�$�aT�\��A�I�Ҡ�9��t�=
ZB�`��X��� �{d"g�=�(���a=h6!s`�U��!lΟ� =��^�� ��ؐ�h�� �`R41$Է ^r�/ǽ(��ԈD��?Mpw�cGz�-�)7��,(k�r )�2�!�0��;�����O�T"rj�=�r�y�(�OcU�ޟ�&���O�G{�:]�!��@QV 
�3Q�@Cq�� ���9a_y�\V�S�3���Y旗M�� G��y�
��2���.��|��F)�b���t��������Xϴs�ܺ��6��Y���.�����ZfI���ʲ�T�|�0�}�L��:��4���
�&)c�b%�sS�m]�l�=�9�P�v�j"Ú��H:�~�[���ֳ�ґz�	!N6(�����J�(:/d~��W�:�-I�~	��L[�8���;�'d��T��[�B"n��^��'����Y����[��g��LO��U
�8��Jv��X��Oi��&H��L��n9�k��l�mڴ�:�'�����K�x= ��
)��f�i�NP�rخ~��0��zK"�r3�Xؽj	����L�`X�{]Yĝ	��`�o�� o��u�����wX��#، 8ԫ,��z�v����N�N-�X��e�t�do��ԫ/�t�K[��M���?�U�S<W N�1���L�K�e8�Y���3[|Ⱥ���?�k��%T|��h3�tUY<�	�����n�_/{+������٬�;}�@Z9C�	aJf�}�9Ӎ��sy�Z��.'�4��hN��Y�\< ��3�7�����,'�)�>N����(�Ah��}I��V�!!�"��':BFsg�y��	�oۦ�.g���>]� �v$���_D	��oU��ܰs��P5�ҥm.5��RR�{���B�ф��&��ueKz�'��<�?��T��F/� ���"d�z�!,����5S�.�@��/�=ȹ�1**��!&���n��IS��P�`�!���}W���r�	�Wy��[v�k�v�!���>(:�(	I�_V�S�
��� ��~[��\�g�y?D��OJ���NqP>�˯[�^L�0��Y!G��X��mS�E������y�j�d�!,VO6�~��b��������� msb�`hB��hR�����=�w�w����z��;�VM�?K�?�	,�¢�Ҥ��s��Ă:�u*�nt�p^V5�O�<�5;�U��"V�u5��U�hRK���Աz��/̀L��ߑwlB>F��XCH(�Y�����C
��m)LoW�dIJ	�DIvV/�p[C!�{���i�}�v�Ku�Zr���	۸O�f�S0.��I��O���ɟ����~�I�Iv[�A����@8�+3���ġt�]�	��]WUn8���#��7A�4� )�؏<)�b��]�DKb��"��\a窟���\F����=�٭��Z����_/]��#ͼC��5������V�WK~��w��0�Dn�?KT����ǲ��P����x���z�:;I���X{���=Փz�$������H�(<{hQ� �{��W����������g��a�Qˡa"7m$����O8i*c3}�8���W��H0 �0�[' ���6u�Hݨ����`���Ur.*OJ��O�V�>,�11��匐�����zz���޽�ǂW�T:J(��l�{D��
�X��wa�4zAbxNEqF�v����[�|�d�6Ɏ��*�F�f=�t�i�i���\����Սg7���D�:�/�����R���}^�w�"�g�����ӰZE�7\�������Q��S�7��7�6!�9����@��� �3P��5�&���R�]D��97�9��(5n2!0͟��z�
���*�.�jiK/)��ö2�jd�(�9>Tf�8����[��S�~ �,4g͸��ۓ�����T��p�1�<�����nn�����"��N��r���_ص�{�7�C��jR~��[�6����O���9s�����_��Y#��� ���'��2'Wp F�5*����H�Y�p2sl��GbK�;ɯ2��2+m ��/T���&�qu�b�-l��<��\cG�S��ȊO��r�B�\��x�煓��Q@�R�����РKt)���^!΋Z��\��Cr�MC�6� ���As��G|�7Nsz5?4w�?�ym�Td6��NibuK�0�q�ߩ	 Q��e�D��� Vs�.����W�T�5�zS�%�@Z�	����6�wUQ�9�ժ(��!3�Ѷ�@�[�����r�ܳ��*4��y�by�'�R���+�~<
�`��=E޶N0�
]��KϢe�$�osi{)���Ԕ7�b���l�ׯ8?z������dH"��P�}0y{пn��M�X��05��$�ɯ��sIxzÄ�r�<0�4 {B�dV��X����H��z�ة���b���G�xQ�tƅ���h	�,4�U}��0e�)I���z�v���(���.2����&�4����	������,�H�\��4˸q���cժ�VӇQM�{��sۚ\�d�}���h�8u����P�Y0/�- ��CT^��"/_=�4�`�"_�=!�Fe83ӛA�oq�{���;wts�u`����DJ7��l,��Q]�D`D�-��dD���j�U��Qh0]u�Z�AP$m�7�����&�� �^�����;g:�4�(M������A!M}�_c��
hLYی���О������I�n/@M��i�B��W���VP���<}NC��1�R���p�M>D��\"jAb��b�?���I��}F�H�d�}p���˙a�BZ�o����Vٯגك��5Y�] tK���ܭ>u8m~�B��wS�f#������a��p��5R�<�h�T^�P�#�CI��e}�N��8Ʉt�'�	��*�`W\m���D�����l���T�N#�O��UWw��g����_�~�}i�Px����L~�/��s{ʓn��_$�����`1�����:�m��4X+_Dz08U�f5�����E*Q���[;����t�޵S�[Dak0!Q/I��zqT����Y}�c��HM�q�����o�7�
QO.�R��
�4|�N���~�|���._�s��- VH4�m�և������ �8�>VE*��A���vc��8����joG_n7Լ
QO�+�ְ����i�<� ɦ`�R!P�w�ٶ��?>@6kKo��� �1��å�9�J�VZ�UH���<ʇS��ތ�+F��7 �ݽ^��i��ާrw�wh��qΛt��9��8ABFrc�$içQ�Tlm��!������r�����x�"9�JHxrF���=(��A2��������������^�g�A���'��μ�>�vz^�� @��c�'�KkO	�XV��B�ћ]�����y]{柫 �c��K����Ȩk�5���y�=~�!A%f��H�>�LD�f�F�4s�wnk^c�d���.1�I ᚇ�a�h �MBe��G5���@&y3?��۔3}�a'`O:�G��CIC$K�6�c�W�Z\�
�+�Z6�Q�t��y�(|b:_CPC}4[ c\B��}3����鏕�8P��������\�2s$r������g9���k��v�qe&+"�j	|Ǿ�f!��_K|�7��I������ʜ�x�K,Ǧ4�s�7ж���"�#r�L�,R�w��80"�M�\�b�~�{m�����f;#U���~�U�}0������?t���M8i��۶[`W�,]�Y�R�=j��$m�&�����mXb4)����!���_���0��Tp��M
���b�DnW��}&�j��{���:��8h�M�#7�TKn���[xD�"�Y�J�i�����蔶Z��=�N���.�� �A'�Y��7�܁�^l��7ѹ�K|�Ph)�Q���<�۽bo[�n@�_T���z[*�!&C.�Jp(J�:~�"$A�6�ن�.�}���Q̃+���G��3sGM~�|�d7bZ~�ib��P@�������5��tLqp����+/�K5��_�ā��i���"��ǃ�0ъ�`�I{~���n$Vx��溯��R��lBL��s�b����2s}�$&=�p��ր��,Ea����7?0���B���>�=A5/J���f�ج�{"��bV���wPH��=��[��`��!��z��ei/��&�Ҁ!b"�g�v͡�$�[N����߲o��{�R��!3���?Â��h���w��e�ܭ��r���k+L�z���c<�P����|��4��U6t��c"��B�g]?9�.�~%l��a䴬o�C��<����B��yS���Su�2�X���Ka���!�ΨX6�K�c���Z�n ls_+���C�1�f}V��_ʨ> �ӧ�6o�0Pm>B���,\�\�us��`������r�/�-�Q?�s�v�;!n�Y2�Y2��l	xցY��@�|F䋲V�7���qvd?)��l�h�^IX�}�k�8<�;e��X�_�Āa�A�����k.f�	�5N��޻�������e�O���̥Z��8�XcGN뮙a� ]@O�#u����;�(�V�z�Z���6)�0�+�%+�E������&�0 �R��z�gM�n~eu��7��FZ�b�+0����%�7a� p �6�=��4�Bh�8�'Зvi�u%���\�n�l�|[��]�%�Ed{K�<��o֞H<�#�#P������JDLn%��B*�u�x!����ÿ�������ut��4]*����e=W�[���WR�6��f���9���46�r?�'�n�}d"b.Q�̉�q^��kdZx�ܠÓ�_�̳�W|hU�̴֡*E�A��z��Ħ���I=�N����;`�V��Lrm+����L:��7r����#�w��.�*��zֺwO�Ė�B{^ڲ�J�͈���ª?�C��ErT�ਜ਼�N�Ô�pY�ߥ,b^��r���u{��P�rO+zf�Y`�z�p�������M@P3��XǼ�XqUJj�5�p�v_Mr���;��θ7���E���VK��Q]7�����FG��֔w��uj�� W ��a��4?����c!+�α	D\u`tl��x|�Q^XaN��a�����i�֎@9��6b���@���=�ggNt�N#�w|��v���Z9
{��|Q$�G�/�
�99�A=��}j���cJM9��`:/����Q�DrJ�����}~�,	KCI~{#���
���et74��e�V�E;�kK�Y~G�}G-��|����~7*�8�y��vq.��+���$�gÜ��:^��P��`sl���u�G��³yh\$*o�oN' $���?e��}��׹Ӑ�4����PI*9	}���!�Ƞ�k>�ۚ�tC�}6��m�l3~<��$澷O?���/�N��D�����(8F
�����y��ޫDu�]��[{���3��d�����`��Oi��ZgD��"���E�˨�]�⏍�rvL�b�m��L�������O�������E�q��̌�4$d�5�o��ܔ�L�Z�+�!nR��5���xf�a���TҥE������M�}�=�c������wbHʷo|v;_$0=�����S�
�m�NUϴHσ2dI�]i�XM���qQ1e��cD��VCnTԝ�'�B�N�	6?_ew�$�ۨy�!�j�:���l�J2pF)ب��j�*[?�&�W���A�o��l��iTT疕��*p���K(�G%�C�Z���d�Л�"��h-�N�J��tI����
iR>�1�5/Dӧ�Ġ�A,�p��n ��od���@_���ܯ�P�=d�Ӓ�뼹DZl�Xr���r��_w�~u�d��+'<�m�H~��N V�jR�,����痻	wp�vn�p��c����j�w.��2�MȊ���vU:䃂c��F��O�Я��k����uUC���W�p��j�� ���&-�o0V�虊��#��Pu,��z=����k�v15�,۟2� ��Q�I���_=#�������B�B3�o"SxBe�ә�x�mN�X
g�����=o��Q3��R�g���'�X�2lX	S\+dG����}�.c��*��0�] W D�}m�~*��:�G��ު�TW�䂕C�j��6Ƃ�b�`�x�����Z�@?$����يxgK8�Ƚ���2�`����*H�R�=}���޼T�5+�����t�{)wJ���=��]����/��E@U$i �	Y�g��n��>U��a�G�.{! �F��%��.{u��d��Y�L��%��Y����� ��tq�ߡ��\~\p�?rG��.DhPu��'�uc�H$}�V�?�: �'8�N��%+�D������Ҧ��|`�.�g�/��0�{�f6��B��W��1���ny��3_�˻��T$h ���⻕�T�(���w�e�S6N�`��4Eg���b����OV�Ǻ��k��$g<�����9i�1�#al�����wtX�+�Eᖆ�>��6��}|h�P^ޮ��t�=�Q�UP$��+���gPb�{6<���dk��c:.��&����Rxc�e��<�}g�_�W�\���jo���aU���g/j��ʯ?to�䇵lKs���ln�x�y_�a���m�����N�W8��G�9e�����0��@�Y��]$S_i�H�r\��(gÉ./E���Xp8�dm�t�
��;DYs�"*�|f��3�b><P5�!w�C�-HeW��x���9�3�n��B�I���C������1ꕲ8��:���G���mӵEj
\�����Y���`�V�L�*A/�B
=��M{*�*�̷����:Z�D
��?���2~e�����N"�96��kȱs��7�M"��W��*��W�|o&,�v@��uF1PT���< BU��&>�N���I�C[��N���n���(V�S*�K����5N&�j��\�$�;ɣ�l��߻����k�Kew�?F�rX<ؖ�T�/%r��DC;
���7�0I���g�T&�`t� ղd���8԰���I�M+{;���z�������O���~Zý"��S_�lT@ +?M�|�!l�tT���`tA�,��ܭX�<�O�l�-ϣ��N�S{��	o��ч�WPSc���B�:����)����V!�����u�#��s��VǼ��g�5�e�sgJsOC����E�er�n�{�b�����x���N�Lff����h���͡A�����nY���Y�P�#�:i��4��r6\XT㲶?募))y���-�Ƞ�K�!�^��N�Z���V��ǟUET���zwh��6~��O��}!~Q�n��
9�U�l\��MǑ���Y�pYpzb�]Q�W��
��-(��s��t���щ��M���1��6hJ!��,��DOR�	гe�p��71�3�!-���oq����CFe.�er�Y%���)�uG9C&�*������D�����ˑM��c
��b.�)��ߝo�`����H�运���T��M�D���y�F�.l>m��yHća`4�^�t+v'9�v��o�0[N���`��J0󖘆ψ�]'d�xT�ԃ7 �Wqd7_|�l����Si�)3�߲L7L�P�0�5�N��."�U�n��2�܀V����n�va9(�akU|+6y�738��A�Id6����X��yGg�ϰU>iy�(|8P-Ǳ��a�lv�v�TPW[;��q�*�9NY"՗V�� t�O�4X~�}�^*��Av����i�����"]8�X���E����1����j��Z[u��ݣRc���\�
4���?�e  ]]g�+��t��e�x�+��L�y������.wA�i����>qW��A����y�s�8#Q�O���s�_�%�=�F�,��C!��M����b�J�ԓLfc��)��ĕ�| 'k�ǁ_��RtǦ���n����Z�z)�m�{	'��)E_��f�;��6 ��/�[�A����G5����ͼ�LLM���ǵ�������W2��"=o9e�
�y�f�z����G4�)�]�ꌞ�~�XL��֗\O�r�ظ8w�ಒa�)~�*��2����=�s�x*�V>ʁ��kB�4-�{�" �1yl���+������*q�5�$|���n���|)9�Q�aP'w����~Nr��r��χ�2Q3�Pz�D������<��U���~P���l�ir�0�^�9���A��uΙU�G���[8r�
6�2q��d9����ߨy�p�a���$�*&���oy��k��@���:���+����<��t�e.l�uSl0VN��X=���2��<���f>u��N8���{s���[��>��Nľ9?��[�N������ �p'��?RSE�#�{麟>���p�EN�,�Q�F�^4w-���-��e퐟�;���H���a�-���X[���=����;796T�vb,N�Q��x����3��z-�QX���2}����@"���0��^t��#O�î_�Z�8�;�΁z�P%/�N^�K@-	�]�@ͧ_0�C�:�O�͖��|�A�P�$=���d������EY��.̪���৪ad�[��B'hၠ��S�:�!���������&OT���^�~�J��-[���0�(
w����s4PMo:�3dv�M���y�o�<'�j ��Ԥ�k�������8Ʒ�Q	d���^PO9��P�c��Rf��r5���x��l�NVi�	$��TcsO�����?��jKe��D�]��7�ۋu朙��G���DCh.�L-�P�w!��(��v�:>�\<D��Aǩ�@�<k6z*9i�f3ϰה�2�q�'��g��B=b(�H8�����R~@�M�����8\��\cs���V}�֬'�!s~H�H06�3��3��,�R�p%��Oí��h-$R����\�m��]��-�1�R��M�K]+6�{��u��f���`����x�C��$"���_�q�}^�T`;"�k�NT2�㚁�J,"�ž����
�a)�G�p�w�u
�a�7��%ڋ���< u�?P������.= .��B�� ��aA8�qYU
F�#4z0 �ݐ-��dY*}�UT�A�6��%O�"��Q+8+6�l�j@[0M���I����E��a�̴@�v��y�1��̺�QQ����]krS��C�ʹ�t�E�E/���\�s$cS�n%��0�ķ��ř�YX;����En��u�{w�>	 ���>J�4Cz!;�+n�`�>cy�Z��I(��R��#��X��z�%p��@�d�����}��lTg�HhJ��/n?Y�]�}u�L���Wb�ޕ�����c�g�s�ڍ�5B��1���\w�0�b�b��8�3��4��=���{EBE�~�μ�$Q߁�����B�Fg��V�$F�����3jb��`�c�I�h<��B!�K��\��5��Fʢ8&�>/�z]�mi� �v�Вz^�bm��!�*��%2B��Rzif�>2M;ݯd�7����Q���I۔����+3'!]��Q���ۘ��$��w�Y��AuI�*<y;��c��K�[�'��h �f�������N�([?�}|G�$9nQg� ]�ԾT��L����P�u3�O<���i�"X��� �:�����;���!m� �(��H��f4~�ߝ�R���R�]�����j��$�,]���a��na:�eb�)��D+w� (��{��%p�4m��sdӸ .ņ��֙��Φ�v׌h�6WŁ�*uR&'4}C���)�w���۩2���~�;ث0!���ț��v9��y��mY5��?q��-\�H�L ��
�Gä��XB$K����Á��-9��%� � �m"�}�.�f@3�( �@�?�E�̼׿2��5��HL��m�g�2��*�pWm�~��JB���CX! ��0[b�=�x�z
���9K���1�i))��Ǧ�>�Xx�U��L4���^�ko̞��[���1�Y�`cA�K��~�֔!Z��N�h?m�.��=��?�������:N"Q�࿐?S��n眘IE�^Y�;&R.��ZD�X��.8���,߼c�th�����ͺ��ϷD��i�P���vh��x*Ъ������f�5�wn��*k3E�~"u=��� JIna �>b;���.3:�!��C��0��
�/\*7�(��^�3b�u��I��%�b�1�����H���M	ތ:,���]$�9�B���'3�Zr}y�r���!�
z�	����A�?���PL8�ǆ��6�YS�T_G�G�L�hiU�t��w�]jV$�͙p����=�{r�5��1��?"5��91���$��B�p�6Ić�<��ߛN�dH�f�)��Fei�;�]<u�z�j�i���SR�89��6�9W�P��00k�]��*��W����C������[�&�� .�婤� ƃ"�Bs��Z<�푘���Fq�����D0�Y+�������%h?`NJ�	��-�5�*��|�����G���Y<�3̼Abb����3���#�L�������:�$"RA�uz�_�̱i�1y�����i��7�)�ջ��MOT�fW��m�T��Y1#u�o��?�E�!ʵ�2�h��P�M�������b��m�-��kg�2��K��1�G��Z��!c6@L��M��҂�"I���A�V����{6Ӧ�J�Aؕ�<��(���IacλnGVC:��M|?*,4�:�(�	B���[1p��*	69c(�u����vFR3?O]%���Y�mi�'�>~2����.3[�s�_3�d�2��v���م�3Y�P�7�{i=R;��C�+��빚�(��
�0$�m�5`�n2����>cA�
����8��fGG|�N����V�1���وC�KӆҒ�tc����n�Q��:R:W�"�y�j�^y��ГѠND��f�{`*�����m���y�w�x�p�D��pw`�-{(�%M.��ɴ��)+���̠|�H��|��pny��p���\�4�i�q�9p���]g��H�SYS2��?���8�]�6��a�TiM�h Ayu )Ae��GA�o]s8u�^WDf��Y��PW�W���Cư.Rn�d�hc1��TFu�"!����}���%:�WU`a��54xq�S��dt�f��̗����(�[�M����;�:-Z���g�8m3���!�N�x��s��s�6�,��ҩ�M�F\W\�<f����y�*j����a�6��d0�)�1���h\�
l�!�*PI���^S����d���A���ߏ��K�r��#AW���IEȸ�M����'?j�����9*�;�+i�CxQ �}��a+�'SHDĪ���2g �>�
&7a2��P�4������C ��F������F�=t]-o91�G�����QU5�Ք^��?]���q��ɡW>�h�=WP�ԕ�}	=��?��h��b��MB ]���H��[^T;�ã�V���N�sbI����d���CJ{g��
��[�,��i���Nk
e��Vft����zh~=�vSW���T�腔��~e[�p��\��\���Cw�ooy��W���*k3��7�R(D�� V�>�l"� ��_#�#a+����윲��fe�ˬ\(�w,1{6^G8t���]�½��GC�;5 ,�ޗ�]6���n�9���\�L��B�~�9�x�֕` �6��v���}yZN���e�AfֽK���m�ѿf̂�W�x� 
���`�!��5B���|[|��K~F�� ��^߹��"�q���h�\@9��'i=i�)���|�!ͨ(� �A�$ �TW�X�<�u��ך�׈�U�����T>�� 2u&��C�+�m��s'��۞cZ�C恼R�0
�.�i�)��E�\�ooa���;^�� 9�o�6^�N��|��ԧ���6!$���d^z@�:o
����6���j�p�>�t?�:`�5OIQ�1gKO��GE�J�|��ɃnY��L4
T
j��W��{���;k�D��Õ#����X���	D������4s�4p��<�.��� Xl�KC
ʑyV�N\�Z��<�uQU��帱�e�&�6�;�TS��Z�dK���N�7!R�Dw`�n��2�IS��F$k��M����ҿ�/7�ut����;���