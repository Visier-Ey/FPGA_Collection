-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
a9EX/t+uapLUMNsQAVwfTEHtIBmVYrYkgI/MlmhFiOYSNlDeyHArkeMU0coaE0b1
PECPS23vvHMc+bTPtD+H0t490BrW52oDKy7zkBcBOJamPH8qN4LUGd4QD4eA2TC1
6fFSpYm9gQ+EjOv8v87pvfKwCtztNc2lDVuRVyGudk0=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 22622)

`protect DATA_BLOCK
ZhHDxDNwFUhK3nlCsQs2PXdwOcIf4ZjxO2GI4WjmysVKeFsl9lugi7bEPLbe+hSE
zypq+XQF5KOsHvDLw68ATg1fxmtoKQ5iJ0pDAgQxdQa3SLB5jwtTP0ooz3q4t2e0
QaCl5HRW3FODFb2CrD/BLlAHdO0yaqhASgCMb8GkHa+eOCz7WF6LrFYtywMzHPff
w1UEHS+WfUDq8w1iqcspMOtiLe8zriaecundpNo74Y046jPFoiGPhYHoSozygF6Y
KzldTuSdhVxLff0MjOMqpJj8SNea81C9b/Lrfnr2GovST7JOKDvhZ22HuQgMxUNa
PzXEuePP1UEUiMe8U3JiyUCj3/VELuA0dUc6ZU0OrrqA5aN37T8yM2fikMoBt5cY
bzWR3be2l52R5Uwe9NnQGGT0HDoFaAt8dtKUiywaz1BTCeHibbsMW7KrfMNLmOFk
BlqvePl83vDdSYb7W0Nd4JIDn8Id9FUhBOSFzp0Sb60KNiWIHWi0AeQ0cR9LyZjH
Qw7D8DwTAqPCcyafoBqBA/ZSuuvb+NVV0GQ6yB3zkIrd3Om01CKmfHeKHwwK7405
h6MlrsW532TdE4JKV4GynLe70QuQHbr4Tu59Kcmbuq6lWK1y4QGkjMFTSKF3jZ+R
2M/+JuFtg40kqJ++C/ukCgJCNPeNjVsKMGste48Irw3Zidv0ShXQWskMS5HFJ7tX
bTR4XbXbA8B4fFRe9C+vk/CrW9RnIpQD6CDZTpZAeLXY0M3C7j0t82eZ0Aaa/n4R
HuB9oMcUkiZf+2SC0a0LfYKlPXXFlJpiExXRWJeLxDTDoD7wkrtIAOfOxTN0Mj+j
wPwtMwDm5cTwbCaREoCT1EakWEs9p3DKjNFd4LNlb37vSRMfC2yP1VMKv88KKmdO
RM6YFQ+XPfuUAYDaHmG43tYOsQo7IB8jduRBUJhsLBhvpIzByQzSlBNOm9vfEV8H
Wgmhq3/yogaqa741H8vrw8UHyANug8MTSrZAmfYW2ttByyIvTFYTmyFG+AyFItKw
kLxN5MffwRvKtO8xjNLapf8N/CriEGmVQQZbrHWlVDrZ1ic27Jv53WEZziLuoqs2
KXEFF2FRN/a2tvML0A94MM5efgrQ5MC2tkT7/r8l/8Zvc1a0MW121c/K02GTQIul
ey5JmRQkGAIHVMF9/K2z/+IFE3D1HKLwjUSL9oqGBYpHAyPbjklUmCCMlX1UhO39
gzs/39TPm9mJmDV5bcrDYNDNKHHCss8Wo6RffYTHU2lAhA1cqtRb74F7AiBFNHYb
yQV/5tiM522l5lYl0JmFp2D4Ng6zKtyRz2Y9Uww5s8XzVG4J5PqlVGBU15ySVQCZ
ettrHMrJyRHtklWqHXzpetAnFgykZnk7/MexwZzp3+Kqc/jv3FOfcFzPMJMwTFE1
gomH1Vsl9K+6rASkw9AmTJjALIq35b5I6vVVwiszG/5V/WVmBVJH69sI5wWfTLDj
42gXTdE1LzHkEk81sLje0Uu9NRVr97uzW0EahrMA+tmdF92WY3a3tHHFHcWnX3I8
svUzwq+S6sAzC4oA7NUvlPE8SI5EctjfOiPmIaeNU1i1ULXwSsLbvi5bQ0TAdGtF
PqzFyTHzBlNT7zvZt/a5z7s7DJnjen0J0qiAgtVEfHNIEXoYTycrFE5yq4hb4+N+
UqFy0u/jUHdmlKOovXkUmpULr0ymlbR4AlNWeQ8i4f7PaMSHc3yZX5tHh95pbBZK
QPxemOkjqNBaY9/M/PY/4ojf2gcc41hMf+eQ7SJsxE8Ti1dvM/KRljJzkloqpmFd
cYMB50jjj6lWv71Ez+efjv5PP34ZgfBx23E1FUtQeM1TPjDSPQbJaase1iLbpmSh
jqM5PplUfHRaE7o5tsWCpa2TnuQJ11ySLp7PMSE1+7ZtX7hq9ZejFyBnI91IQmvb
9aihzgNf3zGUfD5l4+vzmFfuA7bI/T15W+Zbb0TsA/1HivVEp4e5F6JeEb8MgGM9
9wIL9BrgG0s4S3LzMqY/LFKY3/TSa3fC/DbQH2zxQ4E41WaUtAdgJC30KEW1iWCN
Fn1MpeAR33z9pIOkI+93dywmJhTnwK0CSLW7U+1jobN18dUWAMQEjXn4w5+qZRMq
qlEbW9yh1i5DHQPINLlljzHmzBrJFf0/jg8fgVclRnXU+Hrz7ADrmBv10WOdgo4R
x38HdhGs0I8o4hdM2XUxnlpkQ57XSPcpf+idXlffOOwquQYPC1P1xY5wLe0KE0FZ
qqi7UOwgTC7ZkvJnZnt4q894GWlmoicLRjKE+oja98Md/GW+X5HfNn5Zx75jrQVR
qwthPTITf22RKgx89oVljt+9zhOhdt9jm8JT62wQvmxa56z5utx9jYU3Z7z70jLa
Kj2qUYsdToj9hN9pO7BH9HR+43hXNM5cSFPS/Qzg1YNZwNWJOqsw6/yVVSRt3vS2
6v6Idiiu/63b78/pKpniaJ85o8vXCMV8GUM+WH22uIFGOna9gwJT1oJWSHf+XdBm
g/oqj6QwRBnZOSbzbAKm2RISNN+pjphvqqb8AJ8WKp7a4rKrqMN2xFALseX1ypRa
0Xn713wedg4IHhluV8MkYIh0TJuWCsIAUyDhOXRwa3tFNqudbB3o2Ez2EixiYoYU
e/qAOLf9wSCw53i5dS1GoQANO7nbFpHCm4s5LEZarKQ7JIQOzksdTRwCs85qcfpa
JQp4pLyejSOUyZBZEXXV0XcgNuHxoIOrJ5PtcC8Jvmp94iEgpKGYJI28IFKYHOKV
L/aA+VwYEsiZGzREX7Ze9Av1yXkL8RWVLmqiQEZPY2jK/NVfFz1hKFejtl1zt0HW
YXWJeDMudRhGMeiol7IZOGmV1FE4Hprt6dSGNl0zv7SRoM4bQ+ydFKJdLyYNHwwz
kVR8Z/ldY3C4RyOsoI3oviFaz0fnPYqcGrUfka3LLmtw2cFDHJVwb9SYme+hdeqp
/QcJbGzi42HCMxnRb5YB4TU7taadZqoKluopS89OZMbj65fnm21nVpsIYYWK6CGd
J3k5bQYnONUQOccfWgcrZDCPIqL/9c+pbZGy7nvjgdnTyq5n7cK/e3/NQNEqCwXb
uJJPHWlIjfIpvh7MfIFoZvIP6LZRu17TpUJZQwcmtPdSllynZ3TpsGhfPEw2VIHj
O4exHhAS/VFDeBze92gtOp3DOvSbiF/FQiKSnuh2lca+lZybPaSF0BIQcHajTXNO
n4Y/T1IomDQ1I/anI9f1IfowxyggmVAlnOWxCjPzju1mlET1TwFXbjqEnz1dk0az
iVFs+q6uU4hyzthctyBO7sqWMGSwha2R3OEnR/mfH3DqVBYIyhAF1O2qOw5iOxVJ
aOjvx/JuGdVHBZ57j3aYx8C+Lrv4Qntvo+dXAPpS/T/TWeVYxNnoasiA1jodDeaN
CmUdHYA8CmrWVLt9fBQRtdx3Yw6kSZmURJ5iiPKOYHU4fKJrCcvU4BP7TTW8sfpu
p2KqA4lSb6d8fDY/peomCTngCEH/SfiT3VmG8oxc/69Gl9pCORmTtawYdWTkAbzz
RUl5HDpzk6+xLO7ZfpVBoahgw3Je3BvW7TICYOeFeN4XAEF+dPBktskT6WbtXwnV
Ep90lZ57C1rYo6z9T27isR1CgVT2d+1lI3nF0PivtKpNTwQjJ7LquJj5P7Uflzck
3Q3YTxcDCxWAyhpv1COhiMnxK9zuzZgQ9Mo3coRMfRcXMU/LKRWQPVVT9cAMC0M5
Cucu8KcCr66/xBb9fyaabbMGaGbu0PKGEuDdhoiwroh/dF3q2uMauml62EdzRKe4
wxNuu6KNSgvU6YixZH5J3X05SIuUce0vFIlmVGRLvdrd4WZtnYA5i5LF/Pxw1ZL2
2T7hdEt4B843D8KcRp0R4OBv0By6KxtxZ8E3WL5HMKmXoyXxlZs/YrLYaNH9JSml
flNibw/I2BDAZ+GRV41ZHT7eq3yIxygERR37wvwdhP3bB3NHx4htaNPhMPftaTFE
gBzdykjaY6YI2xvunrR5ob8kd0ylzcdO1O3Fj441hix4iJar31vS9/HGdHAqTe1i
YOBjL6GdVNmggfV0bytvGzASZlF0Spz5ck+UqJaW11oJLZlSTIVNx9nNfu4xL5/7
BCgCXlkCaJSeFXHSAzP+Rw+GiQfdI+aaiLTcyxi63NLPX/OCWNXQHVif9B0qoOqX
IPgWU7/0CwmysGz8VCV8FeGg9ZBMnHUylRG2ODq3xpkEPCYnoehrjB6wRIaHb3QF
GNCbEw9SAynr7QDUKzORrYsUKpd2/hvoPcqMYHOpLEm3iJ3AxpO8+iCon6M2hZQ2
0PFIvs5ta3esnJtdW78HkwBcQxpe6ODSLQ+EycaT3LKXegOJCkIyKvrajXk68kTo
VttH8xigcbAl3TLYgGxBLt05yloTp6cV/m0nv7Ofl6rHW9oHyEW5U+GIfVpiDrZ9
BXH4lNe2KDovKGsoLNi6YLBLCxMtlMYaiRNUdQEDchbnqcBuAf9nmG3QwABEJ98J
K0ka4AKIUStYjS2nySpTfAyciKuIqEDls8Bzd3kuA84FMgmEwzRRGciq9Mni0Na9
Y4EK8SWb9R1yDFb4v9Q3mNHlwbAeTlb/ceaefiElqTlxwq1uG2XJjhcpA7wJ7nN6
J9RqeUwmW53ClbeQhlRfcDQTitnr7kU2PexHiTdi7IgTGUGZFxEakXP+cDzpwawV
DU/0TWX8RUUJLNG/YpexkhcdibXffLMbqL9cew/UtNW84a3v0tpK1l2Usmm09UCn
2aghWmlYp3lEYK8JLyp9keXNyiLIrbg/SfKyWB5ffaOePCi2szkimjOh0ooYcQnt
BDL6D6kQf+0M2jcjlrmdwk6cIALwKU7yLiegAG6cdzUKiAUNxVwNHkf9EFRl4c6H
dBWueGB8IICT87+4YrYonW/JBk6pHq/RIEJUH1kdtv07B9jJiM97Ny/0LNFHzzJf
dDC0n8G8khoiQdtD+S6nzLWlOfUUz1tQ0fwVksCTyKx17od+/1opH4Q+kt3Vjiup
CJilh0hwKaTL+5AymDig1Mm/oARKJexFwJ2mr3a03XznLFXXWwIrtZvo7ozL22hV
CTax+OR99FtSRjvnqJGfi3tGqrzf/Nh34Wzk/uSWXXpLwDPxKmLuFpfxiesV/kbk
ed3uqnOVg5cbbRJK12BEtyVO4OmC5yIb4RWXfPK7D9XSwLpKJ+D7eAO3EOHa65j1
Bn5bgX56Cc6fkTHmobAruTC+gVeROpN0T+e1sxASa8415pCNfssFONTXhCG3cDiT
DItclGdlkCoHr+67juAb6C7KuduI6uD+hMENxnulPFWduyBySWoeojIZUFymNt8M
cJ57QaX702uIFHs4Cm6k7ZBlmpVrxopAuOx4sFHiTL8PUCmXRbiEy1XM/XlGxqDh
o7oznhz8ux64LNGdIzYzixeJGuCMzt/zG1WIENf2c3LzE/kSpPgrRYd/U0b+Li9W
3yS93g4I5WOpV/LMUVDx63WR/tOmVlanyqvqoyZXHbuHaufPBZ/br11aVJG2dbPn
6XW1X+gdogSR5DQAAgpEnnmbm/PaZM+ovduH4jUVyUUax/gNyM7duNvD0aB5WyFz
sJ+wpEYjtC2JEhUvZnt1xhgkxG0KGqZmUDZS1mbYl1tkji2MHIjek4gdnZY+Gwob
btIRFOXzJpc3E7gf+OarE+m5V3vGySmigm+qIhjQ9cYQDfhVcZ07hfve3V1wkqJC
+kBMY0R0xVDstybA1RzWeEDxe09kEHXGI+H757tDilmQWT50d4uJIY4D91TkMah3
RPjaT9BEgYjhc0j7X/w0eVb/LJun2Zz8MgSSHsmalGwH6uQa09G9twflC96Q49C2
qEBIBYxue76CogXmJqsY6xFQGYlv3PG0CvmgjkEhHr2W3HEeK3WMsZ1gA/mxnX18
58QElTIzoEI+//2pAV7bfv2cz8HYT5SJIeu1nWwv+o+VL/uphuh7CbnSwTBqzYj8
UybShCnzFrcrmHzOIbuUcooKOMaEVU7IhWAclWDUUhtiKS1aVsGrs0pqOjT2ynAn
eltBucRTv5AeK0GjeuOwlsBernGzJMhvkz7CGBBLBTRPKoct48qjj8W+8T/hI1yQ
jYlVUqbYECm6dMhtfzTJjPP9DmCrbPffn/Ty6cKLgNXJugffsTzu2K+ILwNdr3Bf
pEx/MzDQb+RqwJdg0YPd8pPpm++nFPjaDcLvrN0ThFZM32DwCxBY3MlTNbZQi/oQ
Hv29TWw8kV3FZFL16BwTjVllZYictm3RTlvByEmqxFQrT+fDztEgeLtFhPO/7pXP
k8uu6ot0eva1jmENpYDa0TFZ+0vEgTpJXDZbw0vtzNaTMz3cR7nhPK6353hjcoOb
jorIJKQ8gGakVnFNl/WoAk7rmbwezgcaAysbx6KWECiNXHbAGZzPq5enqpmdN8LK
JeUrLLvfcGAQE8x7gexHaXEsXELBi36b9H5BzeimVJTVsEpajmrd2abzPeSx0Nwr
MR3nQuMtpRGQOY71p6S8Y+7MaAYwRBkaWD3rA0Hlmgq14+yecPF08+H5dGLKZUtH
G60AgChokBz8jaseU1TOGZLbI5Nppl3dnAsBUvrtdbWQvCogyh2An3QU+oZwY6fN
aHf4y2t1+l7RQWAio1IsDruAQ8aJXSGm1bPUKDzuVBOQM2T64/jaxjVCA/NFH64f
IHbpRkazibn/Vi8wwu6T4u57a63sGN0HJMEHxgXt5P1/ucWexNNQD5Ejza0z6Y1Q
2INiu+OJwmA03yjgzlAy4PCDb0x+MwiWr5OmzN1gMBbs5hXvCGkg+lxPLC8I6SLd
KCiS/1O5TViTsM499Puia/e00CoSkLHh/YFt9R9Xx9VYajLb+Tx7hYKiB3kYopYb
87n2QVWPVoU92QVoOWswgARZNP+g+B0eBWNyuBcfBQdEiLXkQua3X/X/ubvUEoTZ
/d+Oeod4Z8/9BY8hqPP7VkPunPA8jr+BXmrWoAeyfW9OjZBB4dZwCd180OxmixeE
WOK9SvYTP2Y+QnK69D77t89ohX6O7GHusL8YH3sw4Y/SP1DD68P7tbqBfYq7bsH3
P00g+aTL0V9dNk5V3QDZ8JLIAcU4AFyIudO6DyA1/I6fb2TjV5zEe6otyh7UoY/0
5jDmRTwxJWcH1GxjRoZjCLkDRGsahdLw8LnZP0hJshjKyvLfOAWPPPi5T40+s2WM
TqbOkkp2L6acZm4N7TsTM0ERWD1ZbG5c1zdnwKSVCnT+gsZszje3eYPdQmQ3hckT
P6gwNx1Bnms5Xo7cMKCF284nZ6NxylpxmCcTVFGkY3Yiwi3dYedw9gwtq7x2UBH3
4H5qFENBpIlEW5RKvt5tv9QXe/H85A7hxg4pixMNHh4ciM7gruW6c8uOqVvNoomR
5tjdz+ZbNEwIqhnbhl7Zra04Kxuw5HM+tKw+ZpZWFtf1x6MHq47Lpj8jsfbxue14
Ge5s1yaOcuivQ+OFVNt8D4YKdJKkIIFJaMVn6GoKDwWYcf4xETWTpsIbsNOJ61h8
7NBA9wC4I58OH1zjHW32zUvay63S2xoXNeAHj+jjTRQdKAOhQP20CtKgDk1E40Yy
i+NDP5bpsq+h5ektpGUMRavciYZNvw2sBL5sFoHzHqtKjXknAQruFVuRNwardb1V
sSeV2bNJd0J10XIMjBOp5GCzJ9nJKHR1X2OZIutDd77xSKXfiJUleQlK66wn7xzN
c3T7tuJds4DMuuQS1ZryJKEGfw3QCQGIKOTTHscdv2ZgoUxRCG1dAdLGTyuqSsCB
JKcUBfWUUTRH58OO/ZlnPiTOpLzOOJ0m133qh4aP5ixo+d6NJc8Qg9ZQyWFTq4Uo
NzuYkPOdLEYzqoUH2rUZRKybf+Yfk6nof8++gNcW8tGzNH4mpiHTtlJxhcZqkv1q
C2u+hyQcHBU8IM+fpcEo1ZqSfG360PIuUZFRaF70i8kMwyN+75ApCw8/8LS/d89i
5OGlwvrp9N+IkdR3ybQbV2ERJtBxg+QorExM2UjfudjFGDCM6OheWT+WyvdtC8QQ
MwP0//H/9fyH6Y+u49XTBRKffPiagVyG18gB28WVeuqmqYJF5zNFV48jCkmzsnSL
CA2SNfeS50Hg7tRCl56Rog+JvTsULe3gPX6z460A/8CVb5rh6aOhtahovEaKYNh+
9674Hul4dDWxT7T4SdAHWBQi3vo4+ZxtzWHKd8Y7zrqYfp6iVPg8l6H8l8SuTEXQ
Sj7j+VyvEEOOvQs9STQSdlrkWjlrHa1U1moal62Zwwk69gEPsWVWHR+Y/EiHSCt5
FXjgUeejTje3yt7FVNcDtu3J9GaE+iYt7qYRVZPPfVyOyHHf5Rg2fE/HQN0HSs8Y
wTki4D6UW6saq3lZtVxgbPNlwLWJijGikZzml0x7byUzmr2vil15AHhHJhzM5lBL
r6t1EMGlK0PoW3U++GeKNFcTcwcUqj/Uw5YUdHgVvSUSR7eDxLCPUM7KyN034Iqe
wIty+LTlRw+iJcora1FZPjyMCyYeZNTEhLhY1PYYvf5Xo5QAng1BDQtoMbztxe5F
nl/Wth1SuvafDdYdVhy2XV8QMdcUuqAREEf4QLp3dupkyEJHWr1yh1z6sStsLqla
Ac+xAnK8Z+0ULs2QzZ2dpi4T659doffPMYG4JyeFfMaMu29uY9fkxeK7J+qziNV5
K2MRLwZ3QrLpYWjAg8pl3zkO+BUTl1BO1JdkBz48fFw9TWXv48M75htuFOIDoNUL
Kuy8n9uiAHgMvNL57UsnTCJJ4q1FgpweK02L9z6pPKjVx1vMSxnK9MxnXlfT7QgY
aKRhaBTsrTk6JsOBE3jRD4iJx7RI2U0Tml2xI98swL2SydWKqCMCkvvulQe11W3Z
YRUJ6tq9ot+iAm7kfNH3XaOUd4OUhzjAnMbwQGIl0DjSPeVTdcqZ8S9d7Jgsa3Sb
RQSEqXPL3zw8YEyJ8am2+CcmlmGPzdh9a2mxO+GaWgT4fiSBtf6glkcbg7HxoxoN
M2pI/DBRNfOmBL69pbNlfWAKhzXuXkGDu+ICB6llZqYsmQSniQy3Wj0hLg63D4Lu
O/MkLpKLRvcXFOhkfc+RoX40VnH5QXBRd55DjEofDqWTWxb1wp2nVxkaVVNiO/MU
SZgIdnPFjyA2N9FSP6dN8KPhKyB96K1gny1RU0kc8LJmCEWXhJG/1BAz5jfkhHt0
KW6ctR975vzqQYpaXMaFacZW9AJypXueNKiDz5TaQYeldjlIm/9ghAPShlkU+9NU
za4kyvNWHc0x1jjOX4JUgaClhXm8pwiCJlB8ICEYNSyn6zEWtsvvkgAgB2+JICqy
zh1txuI/76FnKFcWPd+Do32O1eBY346oBfjgcrdj4eo3GsTe1QSoZF8CfRmOxaDH
D4Cy3ZMDWzNi2GdrY8XmtzmA/gdUR8LZw25tDpTeYicoLxrVycQ1BZCfznSFPot4
qCRH9IC8MWpDQ0W5uDsDs1TXP4XZU8/KxIHJTbNbdlWbTHQklAU80ffuRY1pWHBc
NMuUTC/ANnFvz3dKt8DaCi7cjHFE3plnsxuDNYEOluClSR1nNJA7VHBYe0YvklQq
RGwu1RUbDHvwXtSKiutFGWrqgM2N/oK9dL5RL6IJ/mDdukxZDh2Kssu9hn6kN6wG
5FnE2A26JmNqwPbkm1WcYleoMm+E9ubniLGLbegbzTfkxt829cJ5WULssnNR0z1V
W/hqbbNqRerkxUbT+PCU2MkYeRN8F6zCheXpAOTyax3jg109QLD3vXD0H14Ux7II
b5g7UedAc2usN1FGxKIaSD/khN8N8HRl52GzzP54RfsG8gjASdd0FvQtY1X4pUCw
rTljoGmmIH6l0GHSfieiY5dcV8LmS4ci+pWf2cdx2jLkEqF2EPv6VCuwVsOAWTRB
UCdQ3m/dHhRp8Wfi/lPDyCaPoYQEho54EV3Ff6d6xmrBeryZd1INq1Q4vD4HrtqO
1OJPrLc0/tgBalCr6GPm4huEmZZjYfLpXRGLhQqROZeDqFWBwjccgFC/1mX6+8H4
D88KBZ2eNfhgF5evvgSSl5wvc1aA6+iw1W4KUhMEQaX0z09ffBo6McX8b7dtoAEx
JORrY8ohTdtS0LXeeoRcYyvrm5EoKiYuD7OtrqPaIZR0HQ1urJiPzElI2cWqZ7HG
2SY+3Wc5c/RV8uo/0MZdCa5O/WBNJqkqNmRPSqgDJyLj6Y8C3gYWnqtIYxk3BxcQ
YescFmHfljz2xledoiY+tmCBdCzDlTrKwnYeaABnfuezriJSewA05P4S6cVJxeq2
rp5+GYgqY8T5T7agB7D5eFFdjSkt5BiH85YKqEbk8a2eYOpcilopZd/r5TrUtLCb
xTF9DGEvNjAgw7RNPDjVWwrgSFwBJ9W7fJg/yOLG9WWC95MIz4U10EMcHF9UUNMH
xwUNrE1LWAyb5PpXnxPXYm6xwBO7YIkdxwY9uZIkiWueZGuDdQORfFCtPsScmp8M
uxRnA0GGavw6K348nzAU4OLv1mZGeTEZWbY/o6kwTlqXUio06F91rLSQv/lCKfPJ
znNQhpv55fCxm2rR9D5f4zhipw0NvSGycB0DULGi0O0a7oq5XYWK656NRCSV8rhw
ZYcR0NsV6/61a86NdQLWRjyO/5hSAYV0B/S+pHGQmTvyC5KYcMy7osz6dBU1ypRG
cn/izXOJWaLxbVsl9szrgKLXejHg6oJJkYUu7wu5ZZAv0JtVWEE6IaqFHksxl7TU
sf4huuWn/iMeEtM4YUWbfp++cW4QDHvXJu7fOJu6NFaN8+77r0a3EUDT4JQoxPRM
hlcf3clW9GAeATVuCVVYciLRvXC9vtHbqFMxmsksEdJ5Jpw4/kOK1HajWstPZtrJ
dMTEJaacJIh3JorzHuU6RAjH4Rfru3D4u4xvOGVEjEp8KqduseUpgVygPMO2elLp
qkaZlNy/z+tAf43Um57hN57KLZvG74BYnCg+VEkW4U8hhyabVBXCkMWj3msmBOvo
KsmP4rF+o/3pAcg93deao8qrSEmlxv24CsOTjVFbEHvnvLk6Z6XzuyeRzdg95PRA
FeRw3u37O5wRKdl72s0zca5/YNImuF2LierEHZ0XGAxZ2AyLDx/AJZuxxhQLY+Rn
vX+6OmSqmjHJAe4wZW3XNLst5vljES6W+nB9itclGMrehXs+SnT6Tyr5apmhZGkO
Amznldsl8KJMWlonnVtCJdhbKhGZzE6sW8U6LIdlV+pbWGTU5CFk5ut3dTVtrKaJ
ktHTPGq9AQkEDTCl6UhDDvBS3YWicNSKn4XkA5dvqE2VPoaH/r6OrvczdgEZlOWu
VJD6o8Rdg5m5l5B+MMUgEA4Q7VWBP4RMkQni4EuZ6/u4DQOZCM4kh/2lmI7x/O4b
pm0vvSpdxH6D+CDX9vmQrqSkK7/SQ4NGORcfWLHxtcowMa5l32Y/dMG64VyEiMBA
uqtppssJgXJ///dqrBlulQHFCVRyxLDqdHpDeK+rthbTk2Hw0uH9KYVcGVVJturB
XlZJwoed1l8C+UTmrO4dVrkvClsevaSEFdEb9oG7oOrRq+V/+8Dkmnx+LDwOPgon
r1gYkeUuo4/Lx5pMVmqbqvs9/A3VQGE6gONepQFvIIGp8EZWgYdAhXpdn5nl5AWe
Qa4Oc2s7vjXXWbiiz/qFdO0NFJSEOhSrXCiJeUA6APqGPnturn78cpHDIBPzcDdO
KSCgI1v358u6eoPI8hPylS5lqO9y6r6xDDihCS0GpGpIa9PEnsJss63DSPo/Qe48
R4pVkog8y+tX6AFCdL8uSW20m8we+pHdQ6Tx+/DFb/5o8WLEnP2BXPoUaoebebsS
ygpKlmb3Ui2XlgQdWJ11V7MPXD4ZJGpvZ92FJCEbpepbypUnakrEs6xG4vlU6Aft
Kts4hg0YM0NNiaNuNsD4rHjwFKqz3Srouhswlk4Ax9oWEUjtUVU0Tvc16wURhEI+
wBrsOFKIrGP9TSiC85MN6cEYuunEE7k4fg7aU7YtzKXjp8jzzq17fUDf9FoLhnt0
7h9tp7qvYyYraSaZrksp2TBv0bypDTHPCag2Y/j6yvCbdO6YV58IYxwUmGs22oPZ
SOCaannsCOuoTkfA4hPQKUosf71b0qYwtPgYIOl4eJiGw2E9lBP/y+Iak1kVV7KC
ps5LzH7/ulz3L5MH/CIOaYcd0+PjEZN5KN55W49gr0cqwwkhTMRtOZOTPXDozUBx
GOh4k/rWKc21ko5ZXZK9bpN/U0dxVAQsybN9z+6t82wabT+r1Ba2kXWWfPAcs+ZN
SR06JwjOoSTDfqB4+xC9g9tUVMoG4q3+0oUCcvPO6V2kXCKbAhHlpRmOf6Wi92Nl
tcSCIE2cGd34zZwVKfKSFLSe4KoiLDFjnOOpy8pOU40gjfckyIp7G0vRIW1mSk2W
l+h92RUHxs7aInbxVfpbXQNFtbExvPQyaWBlFJrv3UgYtBHt2WGbM/lRrYDAhFW8
v1Njakm9DsTFz/JSheK5e0a1LZyOZTU7IehZXX73WA4R2xhrE55ESIjGaBx33Qy5
YceDtTYCCQ0ejW5hNHd6kKh9LpR4/AM2WemF9hTROwNQLPfVoks7yU8b7fbRaDj0
5MRWOc9FteH2/+3IdLJM3h7bNbECBoSGsvJzE2FN0HE3tNFaX/tkWetoERM7OUEC
bJ+2h9CAQ7qWupl5hFROzPmZLkKpOEhhvwDPyr+w7Oqzp+9oiYKZMJGcXl7QDCQr
C/0vwGwoVM+kP11uemDJ6d1q4cZqOayFzcPmViP1AOST1D6cVAXYpqp5ocglg20N
zavCQYuZjIaaUSkEcZ9te6uMF4vqPLQnG68dLs/RCsQUoNx+Ft8uEbUObXWXaq4i
IvYBKRyFaajgexLtJc9YpcV5ffR75bafzBoAgUG9uCV/7btUyTASVdvgBnIgW8w+
ptdu2hE6QiOtisP14+rZRrd7Q3BlWQG50xsFlTvyDtsCxRFCApY/oXRm9kLF26GS
yhW8v4y+asyndApFzrie0u72LCP4O8LKwraJsssoBQvC3lp6qH5qIi8C65jtgcPf
9MAa43ChCVBiXaeAZtrPK2Sk07021XxVSXB+cbgyi7AsXFYjsPRFaPuSn0CgJ3Vn
MTHytxjtkC6EuDHDKAOIEKgbKG2a9cKd1GBCRNrufLFGDCV+ogPYumqrjQrybATW
xTCMsQdUgJyY4c0MTf85b0uRQtFju/2phftuCsbU6Tlm1Wo4LSaneJ3whyySu5ED
SyN+0Q6XwOp4+0LaxxHJIbLaU4QBfESFGuyLZwPG6pbbtvGsJPDYc4VFz6D4Mz2H
fk/TmEYKfALS4+Bloawp2T7Ctj+mk2a57uh7ZnQh3vC8B6FwwLV96wlE/pFGqlqq
vhnS0gl9yOvvPze0WG1+PD5nCBaD5LiDoqO9hK22FPoCR+MdE+PRPELW6lWKREJe
SzLJSl6I1osGQityT27QMM6ZTYXceUQagZCu++TNUwsnFK2X6YGUkTN2xhyQ+RXC
pU6OMyxx+xsCXp1rgJFKnv2vdVJHHcFb5reGwBR/kqxV9y9M9JpEKiTfFwn5RUam
WwuiJ1e1toijaFUfH4/yxl/r+hFtH+dT6FYduYI+lWgbyyzYmQqqHz8OgaHdBUg7
0wTFcMeqx1cKS4QK6C6FLCymhMNzZCtquC52oUKUbxXK6485LQ717JsbftAO9iRQ
PpZRSLdGfg9+gRxR/okms1Yr/sqQAKzkdK3a8xU9qZL6YXGhDCV/Ad0KiR5j9y/1
l5FLanfsuVbYSkTtb1LUGV/CbXcfpiWWXhEwV11d+5GDaXOX95syUAW3G4TNo7yB
uj7OUvrY7zr7sLketgrqreaotFDW/sru+uPP9U8uV1dWmpCNr+RZ928vchu4BSqU
WHPfYSKCC5ttp3FyqFQk4ygaX8jRq7tcmb/d6vKmIjLNsqC9foWpfOHh5FxfT2kP
7yNklUtO2jSsVONJSrfUDfZV8xczPUEXj5T19A3WYSuSaKRZPw/AWCuIkzlAG2l4
XO3uzfNvys3Jvx+csasGkl5Dpsz52q4KSrlZ0AcM05kOz6iTtE0BKyvDc/Pp8o0S
5MfgF4dPgx3EFgDG+78TilXKYMyUXPW7Hf5ZGNGBwwfaWM/osSZ2w1gnftR8yZz8
XfIUooiCGigiwp01gHrTDwJ9CfARe9hR+6SBtg5qpGc849pnyiq+34ADcCC/ByhJ
S4KugRQclrs5xKx5xTp8FGxmqq23+g4EVKwqYnwkjGnXo9yRlllsWdnQxnuMbndc
hVOXkJZ5y10aFA5FAxtF/vnOha6swaeLtUZQxxo6qBEUzlgihv5ubZtXpNEM+MOE
BVzHE1M/ouHgyfYmh16VjyPp/ZkUv5OKQLFBLtt+bDV/+kiPvmIovrBjU61BU12Q
4jinmvwUPRO6xNMUCP7IKUyAW85VE9xGw9NS7/e1EqzHuik78DjilA20LSVyupxv
ataKt5FUGOZn0rfeFhmN8xp446L/QZLSqKeszREA61fso01u9QgNNUtAqd75LQnL
gV/REEaNDuB8jMXBQkiA4UZwFbI7Pgnrpxx/CN3nyCAEh2PqCEzY+O9moiaIkQTq
2VovkodBSvuRVpZlo4IqpiYOx91AWI8x6h1oDylLUH9g8oVm30vGB9GeECQutmEc
wsiUElRNqN6hD01UmgEb5/I7G9kyzMUOuYj1a639SnOs0ZCso8K/5SB7jt8spF9j
2odiS0nrc1r4bctm/FkQM68V1TVJ0MXj9Hb+Ou6gDsBsoy9/VN4j+GhK1CAHnqpV
gnHV25D/msm20usY9yasrBqzRnEmHagNRJeDSKe/R8rOLv/8dTXnFNXzaGZ5g4Z6
W4ZYeCslmG012PMRd+Np3cegaymsL2IpXcDtIpyApHNLbuploktiNKs9685dvFao
BtOY7xW8/VSESrarAaUMcaM2lr12nJMhpKJERCxRlQu2F3wpROB6wbxeWKktAPFa
fVM3eTA8CmEWhVdKmtAR7JDYyoaGVEushKwiCtVGPwmftUi7YfNhP5SdYumJGxCt
YWp23f1qnMrx4qF/YAB1vbIZTx78j0DJKS1njxUqa2vefWVNH04cZE56M2g5myVK
roqZRd4iM+htwbd1Atm7cV6maJ0ZuTv8LUtDpbIvnW2b0G67kZumxYSok0G219nF
CZFahxtu4P9BsJp9q/jngLM+yaarOVl00DgCKLPzfrEHO8XHXWx6FmGd4gG0ps3c
zH0K+V9D8NkIjf3LEXzhpNjFaYXmtKcf8wM1QMERDsuZTGUrFzF8X/4aXVnxgpXj
9+RLwaW7sGCxyg84PSGLv6dyhKJOoPdxqjkAVqNzQ+ZksA0fbEZU7OsL7eA+47Nj
0iT4zbDKb7mtJfCVErRXVaSrT0w2H+j3LFbzphJqZKEAA6Kuoc7GCOuM1p4ZAxaG
IvzYdzrXXHhSvSR3grgSWVQmJoSIZC3JmQETDkbyx4Uph5gxs7z6wUdXRvZoBHqd
HuTgM+A3dXmE69TwtTZO8gpJY3T1cAVeTiXRbduAzL2HvdczQKBHNXSG3TSkJiAi
x6Ow+9JAOJnJSF1UYQUiz+6ddDz7/b/Gg0TQoRjL4vUgtCSqT5eHKK9U7DuM7V4I
oOebF+nRxLzYrbrjSISVoun4tkGDBhNoZTTEzqwo1BgfVEuMbpOCsva6arhsrBvR
nGIsddhUJl8SiEhmxvIKksZ+sBDuFwBaQpNy2WzhpmyvIihV6Sn68y/CXiNhb7pX
PV92Ve/JZc8OkmhSY0IZOMn1t/MqAsXOF0YsJ/tFjqEZ7fA03A4w45dPCMfww62C
jc5L23TbGSSbrv2lfoMD74StBViEDW8KkXLYISJ88SK/t1GZ+1kbjQojEd9LoPPB
BD57oHyylznXhOTSVcKDIkq4U+1aC1/eBEDkBfuDqkb5ioz7Z+zs1xRpJZ7X552R
4Mrb41B5OqVkudsP49eMJo9t9AWpeHsrl0Ja3sROsw07o6VbIFc6oK67UeFhZ6xF
nMstQWQGoiOikiTLQPdi/nPGPEXqkrCBXWdcqjIGjzTmTGJCUivq4omdAf28WTuP
So1+fJVhQWTVCaliBYmOkCWB2FR8nSxFdIRQHruLC6bIpFaT8wetJJaLqH0loWAq
xaRgqbMHSNN7ykNp/Ncth4inHwDRQ9T8sA3r+UreSuibmszVw1ZRqdMNu9rucBzU
j5c6s0TN47XLzgaIq1ChcHI69rjVBWasmO1jOQnvfbGdS6iwexhlwtWGo6Dn1w2w
EuSEeSLjd0lCGIfR4s6UlnkR19lDrqyBFdzhuIxsz4XzvpK9EvbHVm1kT2NGPKro
kHdY1w4P4cNwhQhXwNyawMm9v82mwQ3WyclG6b+FB03C22/LIRV45dqOyhd11XN0
HL+crciFEyuiTuT+l/vBFk5+hqcWrNdCc6MWtvRBWb+vPQavs/hyeooXBsk30NJx
RIYwQL74r4HMNJyll0PzMHIVfoN5E/63SYegure+9p1j55aA7F6DEq42oJm35oyt
VkSjwGZ8nZPaSCSxNoELca3b8u+30iaRqb6BiOGaIkwMbjMTYO/0o97jn3jHkSHx
4MpjXb+dFORTfTwkb+j6uYHAcEKnwgo+9818NiqSaogs8WWn+p6XNbJo4fxXDhw0
hxwuC2/naYTaOXrW+wX8i8Z2UMXhTwvC3ZexgSt8rigQ5IC6oDNw+5KY0aTDtRAS
ACktW+5rqPlnMnI3qD7ozimWjWnZArBoUlzjOBQ3KxDIRbVfcgBN7fS2pCG7Y2Gb
z/G4HVCXh04Vh955tsqQ1Knky2dFY03LrSuBb9mvHSATnTxeuanoHu7W5Hh6Xt3L
wt+zs9GelC+UlnFkrZ3W6NKiBfeRESSoDfSGzNhX2SOVEfGUHlqqWpA+yYWlyYdF
dbOsywj1p9NKLwVRfC9e3FM+NgJvyHe9iy0SzQIi2ET9tqJTsboNJLqx1rdz9Rec
KsfbR3P7l6wpwYlbtI1jC8oJkIZ3zFCsw78lvTGOwaRxEMmJF6wO3V0BVPcsjAjp
h2c/4fFj8l6+rtJL/mj4yxHdqBhcWr1fUrl+294KQ0Gy/dnNSzuBRwjFS3HXAxS5
bfhYmtudDklWobiP0r/D+wczGh+g1uRuNGZ8Vqv5EKXFE5W1yrRWoO6z7rKN/fmK
hYsjNk23o6xHcHe3WHXiqT2u+AYohNdj6jB5MKGNgWfMbyrnKstw3NcpQb6vpuHK
dyzzN9BF21We6+RTTP8DX3T1Py6cnM9dQSwbmQhsDXrN7ijkzBqVO4uMhxQz46aC
yzK+VIBfL0EPJylUXsejpuno/1Rf4rpJnwP/2LCrhJFYAk0r7z4MLxhB6Ud3v7rK
MoUlAjtBI31ySjm5nQe83jJoLky9zwW/XI9BWV6jbvN47C9f0YR/HBaB7xcNFpCE
0B9CcbscOEtR3TrQC49MTS5kzt2rGCiS15XDAtlH9+6I45m1QiTC9qVy5dhf/2Dn
woXBMaNFP+4VulW/ZMGkk0SoSnVXxBYZ9yZhDITM7fZt7gmF+tO7r4LdRHEO8cVY
jLC4vK9iVk/4O62JV07MFJvQmcJsNWedDspvT98mUXlu7N5SbZkNVrtXikcljs+o
jt2KHBwj+mFAUxknhEIomJXI4TZfMlMLZjIK+EAPSUc1BwtnKEYnbwqbFK4wKLkn
sdO+h/wg93KFeaQRmwPdJiiGQk5COrDTW1FhqEdGXQJdLtFlZgyt7R+Z6Agqylq7
jJGV1HXbA7SxHnGo34BmE0tJMpZfxNLwFdVed386E26KmJwtM9qvO9dMmBmns6h+
1bXvmQWSZc+5bMWLkn08p2m6khK+6buu6KvpBz9/IFqeOfRqNEW29ITPDsBAsmOB
G0YM2jnUg1o5usvFZUzzGRJI6YtVta2KEyoJQxN6kg1b/TuA3UdCEPG0s63mln3/
HX8c7LHmHQdIAONo9wKS8d7jaymFJT/d/dlF7irzFV59EwTk1bEOQ6OvX0aDoUQn
DOkyFWeohCeDoPqDYnxXijdSqPC0G4UTIdqkRdzemADJCnYUJdwwKIX9ZzXRLt+e
KCa9yuWS69drrlAQMkokOLQnMmEGzco+EdyDZoHjmsiCmi5q0DWLBctkIZkqwSV8
G61vOGFtP76VbCZREOuOIK6MwnWnqghYvFb1CwoJ3Wa/MD7JRl2D16SG/FQ2tlkg
823ucXtaKuYBmymVhS0atTS9h6MXx0PXZeCaTAeaBnTfcHjJZiRlNut1ZuSRtaA0
WMCDWrWs+rolYHKCilB7NTLtGnbpjzAlRx2R4uOeakMgCsZbMpB7OOuGBVOXlEne
Rb5SJ2P0UQjUqNu361i+43YQ627897SOUNqyHzIoRoZ8TahMyq4yqVNQNzW3TbX+
aeqogcpgCLvS7E/xx52kWq5xbFLfZwStWwzvj6qXdl0E17tgZclL9TEU4Uu8oPHd
Oy3MdIO0GR3qYzV026HdZC+pshp/+gGoiqLdRVgoXzJa356ACHUEnZ5dFtzvLkZ7
XFCJIFuGWWb7AF0l02ibhG5Ptxt7zfY3xE/Mozd1ArN/Aul7o5QXqNKTOR58eq/W
artSVEL0izqs66Emd1SIyHfKF50NyvNKrl46DnoWmqFKxqVXx10LjIdqaBZSTewl
S1ISO3FjRFuIcB6WeSuVHxXswtMDqJhyrpRmfFS7b4GDgSP9Cw1At74ugC1UnFaK
2cmaQC0gTfr3HVEY16efQHgmUD5Afte3rQOS410FUF0sxwUMK51d7afj/yvnxdGU
y4tDwx5CDB3OyEhrQ8Ef72TwTe4aGlSrSH0W7ZRkOBa0bf0xCjt86DJKwABMtVQw
kAWLHTiix/EgsBkU7ye3EeV+qjaxsteYM5mLMEbnPO6mfaaSh5hnw1uDmjNN6M72
M7JCPoitti3z/56LiJ+EXHe+qZzdjX+UaIABccecqhT1cu4+NvUH0SVNkj4524Pe
/LhEuq+IyPigoL4hTNlAEVy5v92Y6Y2FsNryc080Mod7e72XfFaeTHdnV4hpYzQb
C5j4MZeUTQNo37FWO5r3BaIPqO+TZKrbVtIGeiIwscQCiyYztv9GANn3zdGiiPvC
OO8KnKRRDEjjrpPW85i/so05KebL60v+PH/l3K3GeJRYQjkP0ndRrAh/QdnVIbH7
lZHRr0TXgEEvFa/oAkW3f73p+lPo+i759ruTqVvJeZSEMAaHxpIN1a7ojgpVuWfL
NDgWbCrP3KXQTk1hXuEgVr7R760m+fCHc5HJiYPsQuHNawRsMI2aF0v96XXncw6r
6zFv7JB+H7nq3SY7G6G47Hrvgyzgv+xC7EWFpqJfRdwFTYlq+M2GzIzjTLaJyRFf
pcFLjJ0/2fcaEQP2yw9m4LjGWOO1aNF+uGod5rhVIR/qN3OrOJhFL23Vjkwm0ehK
O8pH3m2rayXjt8m0r/xCaXFFh4gcyyycUADyUV/my2NFcuopVdUCG59sVKTXFPMN
O3VTJmVpIeoBqagSsWsNI36wwJHzvYV3zJ0/i8O1S7W6OZo8cWA5zvk601NgeKNa
tyfMEpOEWeEI+e4MwZMfFew94yg5znztDxaaPis/e6vS+H4zt3keApNN4IO6zKJz
cotEb3v1koxNpd5dxT4yGM0InVXRTSs4BlFvIDw8J1jqXS0v0tVQBvQOEmQ3UBtp
8A8wazNOGcKMz2j6/FD8Yst677k8csb4T35w9MbP/C85k/RYLpWCdp5oIQqselI9
MXFrcUM7zxQRtZGqn7LxnDkAONzMTlrXwDKI6jMOpIPteCQQIKyKelWbG0l47+ht
c9NRZe/+jDJKKM+If3QMzdpejJxkhFAGAGfz/2ZdUdtE8mAGp4CxeuwdUiGvV3vN
VxBOko/E/ReOBiELpOclZmcGTVhN3zoiM1vUoxlmKjVkBMUzBlivHgDiSSDiFz1L
TFZe+b3oKS7MMROxPiYHkHW0r7PZ/yxy42BGhHmf/ual9/DMBKzCxlBxzsrwrfaV
46wwmoJYIZlC1aXdRJvK7Wmnki37uT4E3ebF9kNE+NUjHL2G3wqRw/QLK0TU3sCC
aoVp6GDgJRWDSSVow8usFMeUpzyNL1Jloq2w595raMpvVEa1z7HQEhM0hdwF/Joj
RPfPmt4EaPQ5Ft4pOXtivXcadKPdE1Iv/zBRt6HYESE17oCrP+JKlncZ7g3pEoKw
fNLWmabFf9ZL4HRkVH19+6cEngoNRwb2j7Qst1wgqKvshPCLv6lxdoeeFioXO1/k
cQcpSnnTBcqKTO483h13e5m9ZCSWJjc86T+4t1GBsrhx5pnnLhjfTjpTFA4sXCod
aGxo/yQ40BVzJxDWPucqCTJ3X2B2Nwbk07hnehzjtKXhPvtOqtBggRtWQ+VRDygc
FJnKQJCLO5q3Aa8aRAwSivUhmjlmvi9PTui9c2V4y1gAgHtX1v/JwcQrU9ppIRAM
9JuVa6ugTKSJzaBXty1a1C/jVqzZLP0L/YPL+novGsH+dFueVL7LLNd5w3v06zVo
NlR9CqNhSn4kRU9ttdGmwWPBMhZ+Knavk9tEI8L99xRa4SFeVsU/oLm9FiddZDmG
5esmR0+inavP0aVUdx7wu/Rqm1pp/vns5Z3tw5Mt5YkXXoBVcVSjO0EQMM88QLNI
GrsG2cymZkWtcAal/y/xIWQsBeh4KrzkChEwzHNmbRuGPg3yRH2m+h6AOGP8UC25
uBA+IGZjHZ3/Qk+GG/0FgtmNgCGlRGmRd7gsmdZs126EE1NKqaJrHG+fnmp1ShPK
Xj51w7C8foFKENgtCYu8p3Xe+AZjgGfYfvtlzMOSjK8sEuZmJ1Y/9RLl2adeenN4
1zSCvuOGDV1VFf7jEhyY9ZP3s2zxOz9wwyFEtZ3WYqbjsNwaPwY/Q4uSASxlErnf
xnGxbBFLOgDi5PLPjUsOSd0Qp91weZrlXvn7GQXj0oneCM1+9Ejw0GivRrhdL5tS
QSltN4MkW8cyNL3kQxKOETJuDlkCBNP1P4dbUYLxjxGqspgHTorcpSOfRpz8NPZX
PEn72RcC42lQZlxJwwGyKwd+WIow3tHIkW6en4C12+wd+Qx7tvD5hcsiOOQyukhc
56WYovhAsaDR5JCg75P1o9bJ/10dQT+cjLew3Uxw51ArqWGvSwZHx6rAdb691H4G
5JHB77Mxg3+3Om9FmbLlzpZwluh5xyV+6cncsFTa2hv+y3+k4y9/H+GJnVpLQd8R
Bb/pDBuOHWqfs5br1kZbYI9R/37FEzArPMvm9nFiZL89Tgp8JY/oEoXY2gFN1vyb
fVifvsIFSrAi+f6bXWf1xOpQ2FhZhWYAc3/b3Qzki5//WljFYVPUJVZkNwess8RZ
ptNnemWztjrKp809OYiTKIpI9S7WV2uukSwm7PrlP470l2gTC/Cnr2s07EY4yG7X
gJBC5RRKpuXMuYFPkGHtU48Isl1DCx/EDnWhdpuXSy+iVQONNj2RkoBNuCcI7SRI
XCNnpiBCs3GidizKGRRb3d+/2eplAhfDtGbCQ0aACxJyBkmREzzTvCq+S7cCC4BP
Hz5jXfpLJtWeRPEZVnrQDewEBjNYmjioW9m/ggWT9yVhuiXkmwtIm5yiw/8CapWb
ROHRlnbWYDOljfQQuDCghYXMIiPY6NTVD/XHXzoF3i6hyAU9TocEKcXFJf2hvo8V
17LjbC4X42Q+HjSR5irY0aPKrGDVBLpYi7YDnrCcDG7BsDQkfi6WlYEr1wTUK6ZX
kO4i6cmgvyNcTEvhr/6kRvlo2Tr7vu8KJ7g1Rr5A5cbbxYmRrZtykVvbojCYeCgJ
F7aVf+fu/Lxbezds6sTQB/BHpgGlsJ7lup6oKyiBwQ8n96Xs0LbSWtlQq919qlZ8
BoWceaxk4D8CxG0B/UOwKe7/iIxjKURoCVX9wNUaeiOmM+U7D/pukZ8zaaiFHn97
r/gnzyTBCG0Wd6wZWIBIHQf6t3u5uThCz33dVEqgRA11M20DEICpPAIKGxF/0b49
ccScOWTzOIXtQKYT12giTqU+DTlRRZfdKTcjTq+CerXnYD6QjZEMc7SztoJSmvGF
d3bpEL2vQimXN1tv7O8UAfX1U5cafZanre9RQ+sXMM/wCzReM/GPsgPmD/uN9LR7
6GLrK1Kp5EUsD+Z5MaDNWuvEMTmJGxKTT1aXHo1Ntz5Kduas6rTHoD4+XRAYRnCI
B5kHAToPxBS/2+aavxycrHAUhIYJNRuwaAtDNY4jJM2L2W6dudYEWctS/B4xucrx
nEAJcvyMbtytInL+7mXG6AkRFKewhOUuS07DkYMhMr1GJQzCUOlv3q/t9aPpBvDB
9Dyr3ZLt3TpM3gVl1DxZlD63r8i/BeolUqAmwz4ZslOvhVuce/qZkI1RSdrJOL0y
gFUeUqw3rEzaFxgMlb+hY/HzbvgBjGvis0J5sf3U9mYCNM1SyBHbPmnwp8pQhE+2
L5yjVK9zj2UGOH0Ggh+NkXc85bxy6H1IT6OCaI6J2M/5PzuhidVkr3NzYLNfgkLx
FkyIC403oeH/EhzdH63W1c7GRVo7hR39FvSohnRArOwVv3yyJQdHDd6sNCUcuzuZ
9F4DcLli15/z++kccB8/SsWBYocrQ3RDe5SSMbafyBFdBLVVnFk0SnTSGUquaQSG
CeW9NNjhoSTp3iEf/quYPPuUv3C/XJ1AOkD/CE1XV6EITXOPlchLF/3uPJvltnpC
O5P28tAgTmYrfnF31JR4a0kEHCqXVOD4HD6RHPLiI7PRXmIvy2sVWXx4bjhuD9OU
rxjB7UiFikbUPZZe2CucT8ii8cN6Wn9/6ST9gSPv8HSRK4Xzsg4TcwjzP8yl/O9h
9bULe3g4YjATidJ4FgtprjZc6SQvueUhf+1+oOPKnK0j3ajW9Dktr5hZoRySyZlN
OP6p6f/CcreacZySyf0snwQk1Gsaie5rxBcClnq7oaqWi/g2vnWBjFhqXvf1GttD
G7rEIzm41dOymt/c9ipjUK4yGc6UBlXc1cmhGDiju9HaHb3e2HYcPdioaRZnhh9J
lgYsfwOM2IyWqRSjja4wzHzbzDYrxo8V2DdRhHTBKUFhVoz0QU7lmmf3AzgW0S8O
d/tiqKedu8XVQnKz5swIaTDSg3izWK+WRhzjKurzmZ2IVZDYNm9EFUo1u4Io3X6u
g7Re9AYJZ2WA4lokTuAj10QAKWCcjo33rrGsxLDCPW/dcG7LNBHlNL74FNnBM4ee
Owdg7RhlWps6RPt1Khb6D4BoD0pCjhD411TLwvRPsibKBV6dgAbTXgXQ0ZeG4dZ0
gPgFse8rvHYTaz37MdDcVaYH3cxbvVosOmdgQ+vUq9rufdCGEjGM66c4GyXrtoXw
4g3pS/w4feFuBeeG/xtUUukmVrrtxtrvKSoGdbctW65FevYA6iy5Fk9Lay4tx67B
X4dVEodoMJj8sNYn99vKvbly0FOsH6jcOtjnok45iAH31EGVhX3SCFNPh5RVIRzc
D1nwpMuWo9JL4q7ePr72lPpNwY0/HPaNW98mPQhr0HX67dL8I9KP1FA+hX2Iitg9
VR4DmgUckPvYhjKP5BZFhZtfH7xl17bKatcmcAvLqWJC/56RpCFVUOXeCery4PO5
cg1njljnrA54kuIzffr07f/KrliW5zga3XX3PT+uWOdD1Yb4Bpgp4mjam9UpPs+b
Vt2DM1H1EPozH0Mun0Mb6HJlxyYu95iLuIDNu/FATXueb3GHM2aQqJYiP4gHi2Pd
9nQt+XIajCtVXjNRJe5rNhYMwBOR0EQvwt8C9rOA1aruhyUqkJRgqqis9a/MoIHf
Xx6R+HLc8bwhwwfvv80NmyYr7CqHQyRhyY30YToQzpzlYvynxTBIsNBKuNCaqF8B
IGxeD8s4Z42QMhh/txqm2te/qkcX1fe52NFhOlS2ARhqLNYUwvJuorc2Bw8BPsw6
nJNNkIEJpmpHE1QiiS8ypXh6LG0EmgM1d20vVusi8pr/IpHnqedLofKv/s8cXNQc
nwFeblso7LZ9A8SVkGkp13isSNnQCn7jPb22y9SioQDjMisHkNAL3Y4djLDBI1lG
3s3PT95cgdbSwjNRckx9rdLpa4EftX+qrTqMJbF97rVjgw97d1YIpp6jv5dJn5ze
5+787JRy/EkZWVg0fuQTOD+PCRlBxgw7AIh9LQi0PAvSrSLsBZch33r3qepvpohm
/Tk59WIbrFwBclbeFu6rMauXT1wi0nlWrlfooRfXLNL+Fs0i6nGygGENtOH+o1Dl
KwDSj09tZB/dTAVsuHlyz/B3JxC9g6/9Kpuxqu7gg5aoumdbKiE2E3DroKl9FlVB
iwhVkYcQ/5Z3aSi5x7HvJcoOrCWVEurhoRDU5G9+rv9NtZT3PY0TpgYdoBR/J57Y
QzVrOfz0TMJRqVLYSRBd1jfShxfPc0KhYQwFX42SJ5H0EV65mjnP4CWA4d3PY5y0
HHB0dUmsyJ691Bb2CkTispIw7EUAFAogx0pNBJbKcD9emvmiLExqA535lP02yES8
jn8mnlwhbESTypyYaT5URItP/D9NiDQuzJyo64QWX1+xB0HMeHfHrlGlpKTk6OKt
EA8txpFN0MGnK7phUaIBQSQLAGYNZsb3E9w5V1a3xfFTi1erBSS6qiZjgNJ10bvH
678Ua5RtTYEd8Wa6lek7hDFdE2ly0yWIe4GWFuUdsG9lSVkTRndkWvZbZGaOOj+N
Jq2ldIGVy4ZlD4SUDnv354mRIes8Rq3YekUi1Bpj5mdS7T0vlSQyn+zIsyWJLJox
YTtjEvJYrMzrA7DOrj1jKOLJcxjUQIl6/9z+YN88vX/i+cUGA42NtttEUl1rHek7
WYjGI+XMknloNPLeutAQ7sET5NK+Eanczfg1Tt2qjiKaq06dNJXPomLndzYcQPh8
4cJ1HNoblcu2hsxCm45F4J8zqhBSnFfdNNaNvJTrIPWZB04FvNuHRhmC+QNjWr4b
+3z9qhQR9ELNxxFmjZwK6qY/1Qw4PFrOtplpQqZQznzI0qIlgx++nkAXxkLJZxr0
5ty80gYodRZSRPKAdPmfyu3vLY400vPVuf0cKhXBKLfxG8e9gQOPqleUIhRgGSkU
w87ErbF38urkEwh6/Kr/hURFJJu3sCXPgmTGMUMz8PK4w/q7OU8Iz4RicuNQCucI
5GcNU4rxzaS7d3wAYPx0/JuISvpqaJJLlJEm9NtwwfTjsb5nSJp5jjJ7Ws1W0MqU
qw/MgQWllhIk5TYZoW+v0AZLZbyDvWbHD+7wtUqUMSj2SmUsHNgTK1u/r0IxB+Pi
Z9DBdsSo7gj61h6XhwUq1LVEwLGC0ssAVkEVKCUj+FU7awF7UkNzcGM9q+0ZeVng
HxNHmsLQ1TmeCXcE1ljE3qsvI0438hlH0h/qd3fz4GwjZ/FyPzzOqviJdC3LONFV
E/dZQhSppxqKx+pRzBlq8JdLVPrms9K2fonvqABD66PlcrNQqc5SB0ZoOKmxghXU
F6Z0oS2LpBDoPger2bD0j+zMbr5pnDpGBFPR9JlRp0WAhI30hOQHt6HctqHO7//l
/AKMUMXcaXAtWy61wnw2F8MTy5xx4T1bcR+yXfFwM0ejFZuLRZE8Eq7vu5Hi5izH
6kcylp4Y5UC8yDghPYsuoCTYxXdxeShWCrdy5mPwLKeyoFtyqSUuxfBD64W46aFB
Sre2UROJKtn2OQ/ec+agYt/8uBTuWVsO3KZG5znbes1ISbp1kofOOFD0StyQ6I4Q
VCSn4P2UN2Zk/gMvo2Z7xHcqruELRWpKg2xQowVMQiQEWEMEn0PEZ9cvz1Bjcm4S
mQor8tIbUEShQSCAlffbPrb6gBNGOJ8vfF6lM2UalgkwLvibr73jV2zNpkK4bEIz
HrQoD19/LCr3Hkadpw+6p/1bIrDKZ74T9cRdVUOjFK11RpGO0rD6MqEHgmvlX1/Q
zNe7yIW0aHCqK0zZ3ozHDIhgiHd77b0pcb6pctn9sX6sw1cTGM8C9BgZWZOrSTGG
bnKEYbzJItiZK2zh+SsHkEgjuiAkGY7elfAWT+esWjCGE5RvyWhRUtTOUxZbh3AJ
uCNbZXFjSgJUXwKQ3iBPwPZUCG+Cw8Gz3nsMEPAbcKD9zqXSsxH16yNbcT2IMSr6
tqkFCjEP7ylyPvZT3asM9udrgy6pVk8eMCEX+jvzgmugYxm/Yo5VojMpgBedluG4
IHM+69kfzjJmw8ojk7E9my5LRiMYEUZm6htuCeTlLjUOmW67+Fz7ECSAzTmuYOoN
TjOTSg4P2jQC1PJYNuzghHbEnZnlE3mhnFvZII+h+qlepkuxCTfTEh0dm+hTqXyr
8hRQCRCCBbbc5cOjJtqMNvrfUR2NFXTjt6EbC9LEO1TPHUgittsW806WDiYXAN11
guCDkbfStEHidIAa6vJRJs78DE60GY0O/uC55qFnPwmmmIRjLaZZYfuRmgqGHxpn
z0aV6A72H0l4VoM6GIEjj1GlK4cEkxsH5ScwXsK63+HYo0EYgykn7+l23oqyPeCZ
DZjLnj7JdfsHcoSLHqECGIE3pADyybIdzGQw8+5Ko5Zl4+jyD31RsDksAgopbL03
3XP3RW4EkroLkQHp2IzWHZepvVCOP9nMd4Ph5GZOoJX+Jn/Tb5/xcxxGo3RZ27eC
I0M3NFyRCIKnu6dcL8ODTuPVurFp7O5lk8aHjIGzTxB6gG0vKg7PA84ZuMuYq03U
EtglBP+U8EPWQdskV2SzuNxE1PlH+yJ/xU61Nk2aCcX+pWvUYZXqSzY6+rSS6MRn
GKlt8IsiaMQxo4ez6TltRWy7sLAqENTkq408qHy9pjEwapbwmIRDxbjKLr+A0UlM
BtZuysJ1S4g3gQs/Et7+gvsnnbn37pYhJm1AiUrUpjIFX6Fjqgw5Qd86wOt6Rp6l
bzVeM/4SdO+4YSthepsoY4qDuPYTbsHSR9HvLqMlNvpE18NMOE5gxY9J2sVOksMN
IwarDE6ju2LFQyqOEzhLyt+Ii7+xo8pgjSf6RGOP0voDoFLN1wgIouINyOij3Yya
do3V4eLUd3PzLnB/zpCd/8v3jI8tA9V+ADtZC/tmiKvrlGo7BqCoZ1T3QEVhEMea
e23mS7CEdt5XYTa640xzJ0dQ2dfHVB2WdEvnBs+HnllYNeo5xa6WFlvxu9RFWQ8x
NZ6STl1t9YhYF3NotjwLgzUxv7Af9L30eN9/XAf8R6BK2Jmrvxf/MqMu+IJdH18E
a9VP4XhzNIOoAdRE9Mmjl+GplPMPXvYqwj6o9YrHN9nffidLEr2z3t7eFQeYfOup
Az7qH4ggJpAZu+/ljOA3F91o7Z/vwt+4X9UNRFpiNtJbNSzi9rJTRSD1bX/uPYi1
w3w8TlDHCO6w5TS4XcV7V8MV/Y/jt1rAkOPVvSchDyH9QjUSx91OnXlwenDacyuW
aQ/xY6oLxeQt7ChGx4pFEC1riZdMjDW+ULfR8vBH3ap3SYF1b5zJNLY/YzqdWEzu
w7XNx4VdlcYsL21UO41vzsBgAjHf+DVjRuG9TfZ/zc9IeTqgaOkdV8/mkuB2o41c
zlYyM0groMtz7rvic/uA5y7AIdGelCD4p/LZXDEvl5IVP3ZSubVNt7uvv2OvkpGd
zl4yFw4oeAi5Lm7vsjbscZes1170Q0x1cMAIoQ8GS55gmuraXGRe5BmW7CIVj6OB
3lfN46oGNrsyXHcvpgaW0/hggru/gQ7SjTA3M6xjnoOXDkNLWS20cS6YLL5xO+sO
ibQ6YbdWj0aoC13CF3DB1+d0MpBT7vk+h13ZRrAxWnFEduNYUHqyJaEaO6CUbnkN
2UQ8Takz3Tmnwrf3OmeWJt0rkgaWr7Swvb/LeeME+JhMebIWr0kTZnUfocsQh+yP
Hxi+0y5SYtD4NOZtMZzB4yS8t4llGoOV7pmwi4RUweBYtT2IOB73Aq5D4nonEV/9
Yxd5bSXImoa1zE5aB/MKudCEUzuB2F+TaY9bvCm+JhYFh2o0ZRAxVo0Xmy+RZLue
Byb7vBAJBnHNCajyTb+KFLp78H7OzH8dtehVSTg3SkCZQzn9hlnUBBK/aSS2+2gv
eapFS2LZghQEA1QehpT/WHGlzW4qbwdXCk1dHXqQ0DoklTd8NiOV3mXoF6qMFmgc
doSBMnQmv/VU9H1Q+TcVYy0EW6xW7BPffyJ/rG2lpeqGg2PduMlAqaUB/qChXfLK
Ll8+0QS3W6ImJ2seu7FxNyWKgvLyMmO8/8r6EfFX2sZl1P8gkS1KsVmGKNr1YtOI
+XBc7oZUnqgTMs/e4v4lQAWQIsLsiPXo+ciMP65Ky/uXbdVKAezN+2kVCP+rCE17
dfkursuGzJ8vT6ptH4O9wMtdL7kPHsP6qQ8XZvBZLEI2KiOaaMOfHCpMIwkfIj6C
rGT1j5+dA3/HPJZz8lpgnbi2I1ULrC/UpP5SkkdTfNEAiCanfQpS/jI+EV3EvwtH
sFeXpLjV8h2TI0FZ7vPn5NGlTJyqEPBy7yxShYpolwW1Wk5ynFnO+m9EHWujfUXH
kgIOfx8l1COWZqkT976uk/80q33XmwfPDqQQOvF9cjYPQutYGnyNztvfuPtm8e4q
fNDa3URxSi7nBpdc5zgRoDVefj5sJHlcm+JgRkFRBIX8LrIAOS5juk7txcjS05p2
ZfnHRPQJNdX1AeGMr00kztbw6TzKqZy832OraLOKI0Two6MfdyI2k560mcMetLR+
aXekrsUVzUFQyl/efqYy+kvTnQ21pBUWGCoWrr5CBIr6Mig8ACPbywaNrTz6++97
9ddNJ6JjIXLLEwWCuC4UPvbTOhUOLr23hcTeDEqqy70W7n7bn+AJOVsfnIiMLpMd
SzyJnVYZJkq6wbjyEmsgV7rlP/jaZEzczLNODZ6aFR0P7gmGzz1PClST3OBdLDUB
+Z6HBgC6wkq1il3iQS1Prd67m4zUb1UMTzJ12gahVYrgvaCHPQ9v7091Aw/XpFJM
tIAvwwXcEuDliLCJyG65ZfAkV5Bc5nYL2/OMmnaaO8M/z/qJieYTtd7Zws5YhtRn
gha7933WgPZ8dkR5JRnIMDh84dM2eeVFIrhJwT5kuQLGAx6dgGCxDewlIqFVlBWb
ighunR7JOozOOpoHferJ4SDIuUBlns5p1Y8wBIH1XNzDdFA4N4Mrt6+jEIxkSYIg
ml8cYDkF0nd0FMB3hmP651RfD0DUn6Pw44P1TN1q0Ep9BqLljOtRbGoUafcGtAFe
xudhAO1ByJbG0WvWKLxubM4Eh3FW+gjSs2oStGH3yH0UQvRD7n/99AuY3Q+Xdh61
WZjsYqbWUzAT1uOoW3FhMxHog9hnGBe9Ihg+jBLJLenBf5pFemYYKKCOWCXfWtZ/
TxyWpgx+YbepGOWoxLmJMnc96/zte6D2ykkLTzVbFNmxYP5zERCPgwS8n0GYMqSF
hAz9/7JzsDo2uw5fsBWb5KfSS1vPj3gcY+qegRTDe9zX9O4WiyN/V+JUHrqVEaHU
mG+Crjo/7PDAFeSoOvCUtGeF3FJ7hy6lkw0LyNcMyi1pRNon7XMuc2Q0/7uzZGMB
ZMjC7SynRji2gRXl5i0J47m2iy0NC34pX9CWW+eDkfwjKktPHzCN/DtzqVRonpXY
AXepqctdknj3hX7DWV6rQd6+Z+EHHd4tbmTkvVWSSnZAfl2bll25Y+kLcLYtBL6q
ZrQ/IyVEbDTL6vT9B7wi4debPZrH1BlJj3Zahg9oK7jSBycPKzDHzpX/EFRKPx9l
WgeGR5BWj9+URORMjHuI6IYVE3NhEYqgezZyWPRb5uBY8a8YTvFV5x0wY1+nidcp
JIiZONzbmSGZ7aA5Nw7dwFE9JnO/hAdC30Dhmy9ptTmlyEqIRsBZfJm/bSQJOzF8
e9SZ4JGfmRY7egcMTaO65wRUFkv1cpe829poOzkya3ZZ6KFQT0ECLFmamg5KAgEw
uU00R1t9HXmrf904Jn/JlWQCzzqb5mATVj4LQwOSk7R81E4pNVsT+0nkwoTfmmPz
kZSIgAxdIrLlD/5ZPPpFXpKQVWyCspJVWG5Yak/tdBJlgmjoI+jedF7ZaN5hmPES
eLFNocIwEasrN4Ukf05SEezB10xhutkMY+DT8kKvMeLf61nq3LayU0qtJbh8pYKt
b+QshSeHh7oPako39GixjmeBsyTwmL7mN8R1bI1uhkP7uv9hn7OmhiNuUB1OTcHJ
7Ypno5k8zPNmaVeYjT/7h0XH+CqtLPU4+qqKedOgU1+I97JCKD+5HWLusDHe2oxK
VTEFWOohggOP1WBInNEz8yR3l0U2ExFwIi9vz1z1u42qBiZW55GsIeClJYvysvX/
SQNvxISkxYeR+sTmrdZvxWp74ElkVUnAJWnd8Z3KxVk=
`protect END_PROTECTED