-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
x8qs0kQyPYZf/uS7Cp2gzx+UwIbTEzZEK59MTeMvJBqB99tSIqO89DbbZpbi6Q3dNKidibvaeBAz
iwhOeQS919Hiq2h818mGFVVRL/aWkXZpTdyoSY0KensNiyGY8Uz06Co52olPyEh5zDIeKuL06X6z
P/3TXQmle1Wd87ckjNLMRTfjYz99gKtCGoaBg95bfk5niBpZ/aX/0tUUqP/m9SvBhf2862KBdin3
GV9hTwzVQKDMMkOxj9BGf+m+LH8Bba5d5RZrETpDEvwGRrV+ANu4j0zb6w+NzbPMre3wkiGgWlbh
MgCa9bZq4JY5Yrj/rz6ZBaLnGUQzHUP11wTisw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9440)
`protect data_block
5VoSYwjqLejoTHdKCnL0w8tSYvsFTTmL2yUN4aRC/KiaiCNVosCTmCoxq77s6KP2jIQ7uU0mT3uB
a0HlwIfibUKh+Vun75oTEQxveic1KMtnEV7E0UXG39jdO7r42C6L+Szz6WAheYGOCNAfBBMBmNSF
B+lXCPt4KV4qdDGTOzN4n6g4Dk5msU99mFh+tyad+msGh9Gi5tG/babyCV33fMolL/DJ0Gocdwqa
Vvib7xVdPh2iEX9fRQbccV8mwrCFdtvJhHa+Az7Mz14KOmr5QqA5Vfaf2EK441C6eBVJzaOHp9Mg
9nMoz7fuzpuNZ3LfJi/7KJsrCi1FT0oPlQAPxYZpRJr8c+ydXaiffCchXSRuO2b3cA0sDj460qWc
5R8pYxtRxLplukFgYx0GvDALAgBdnmX1gU1ygCuzvO0zUp2eoY/ER0huSbotQ6GsPJiO0VAfNOtE
u3XAJs539BYUbpTisXG1bhLYZ/t+MemOOrIarflBs5nHUpebyqDL9Zf/0x87u3ezmRIMugjrQHN9
UTdMJ4xkDTJdkQVbDIEIEPW6Yr3eYmJmBE78LwPLf/9RhXz3mPgNC3tri6Oihi/lR/N0pixyc30H
JODcdnywXMVH6GoYJyGY4vAoJeLu4RE7v5A3R3wVHmKmdYNo/SGD2Z6GeGsxwh+MoKaS/Ts9LYI8
N6WKt2JY3ghmXfNNcDaBUIPKC1tTozsqOTiKfnl1DsmBg2ANIM5XAkYg+4oQqJWT0QRR+SQPVfok
w6PQTSazQulUas/CCPrBg19PBJEnuMItUuy7ynY/mMX6OhyxUsGP6HCxLOuiHk1Zfc/90Vk6xm0m
yuX/5nlgo/YlAnxVsvbfANss1U/Spb9IEmW1zbuoXTtbc8IY30bYsy220kfHEIIu1GbcbUzkPKmK
yMNbZGEYsmJU2mDcsIUpu4xRlzpcCqUjeoIGCyl8vtK6i0HrqouCDQRRg+hhtb7M+nEmuq3CrXD2
U7CeTZC3tCJp1BiHRT99SfgQdQIag5riYUc+F8tZLEp+IegqWod8oB5oPlMQIUDG7dKT9mAKRwN6
PKhBziIsLwgckKcRj4WJStCHChRaI0qVPyGTJIJrGZTqwVdyQEabSzB++9Byv6QfVswPqsMMo3+G
IZhBMGHvpsT57irjYaAbD3r8n3XXgqF2MJogA4xptti0ZCMXYU1neE8nDxObUfy3rnp9D2kc3SXn
OrNBVua/XwI59WVsTToCe8VNQzUschFXj9zVWfMRg3H70lMJZn/PE9tGdjN7uTu7sLcuPB217uo9
4uO+B+1R9wIvK8OQUH8ixW4tEm4Fn7I3lT9quwhxDqaSECj6c9opnhtTO5UlDTcb+aOJ5aqGPsVp
jptwTxvlWbJqGu6eOMrpIuS2pkz8dSR6szLzrJT3frEurPDi9wAO+tc4DruGZnBB/weNmjJtXVtk
TJzA/qqQTAyUggJuYg/UITzt6KiQ8Dn72isFtYJTYJCIFPKC3AUuNYAqTCWei0Vj6O2KfZY21SUi
5u4l/eMFPRUjyfsO+SAYkiocVVhBLo+fGih85wijQx3kzCMsntYySkSGFcIVb6OG64/LGRvD3Wp+
TJkC5OWZlDc7py2CdqW5kDNrkxHUNNesrd9fPYlLQbkzDiTJQAXZiF8ZSYcc5I5Nk5NEDxs9AStQ
3dpJVSAMNv6hU1X0zlmQETyNhD5fkLXKS0ZjpxVXlbuCaVz1XWn+P0pTuZjAmfpqNkIT2CGXiwka
h2nqj80Bg3wS3Wmcw8NknXa67MLAC2zt1fuF/EtEiX19m8SzJKK6oY/Ik7ACl718gILFT7Tv6pAb
qOl5kt5vKuH1trxGzH7MAWsY4WvCmJCdFVgdAxSpg0xxLn9K9R92h9hH4udJOhVX5h4GRfN3nwTi
VO/a3CJQmJcNcQjvfHuiSowDZBN+C4iJY+pf3v1/klnPjG7CWbQo/O9eFztaws9wa3ZFu4vC/+XL
l063DkRqprWKbhVJwD/nFueMP45D+1Iv8IDjNJx/qygXaSwqAAqm+tTbwonkJW2phb4ap9/VWkCi
BmFMHWVdCrhsDGGSW4GpNONjw0GZsY1T+RY9mB8ZutQlVmIO7+jQZ/uAkkEi4dMHPqtVvGovhtLG
ri+dmcNPMooMwtwhJzwqI3KuKkNPMrHQ0xJNgIqDQQ6Dw1iY71/Qb4qISW5e3Pf4KisEefbzTBXz
U56kIYlPZPJztCKzHkFKFK8zKGBDNKoKdwOLoDsL9AtP4T/5rh9ZfiII9FiRtL5jHleKcY8/Vbsm
AFqgOBur60LKqS9H/r5ZhhU9De+wRCpbp5ASTW6S0sKTjHsDcUOCSupF4MVP0sH1meFFq/ItUnP8
lN85YfXLpaTcnIOrNpG3638u8qqaWpO93ROyw8Ey6cS9cbk/P0NXNmJhpDlkzDifAu3t8LsdPOZa
RvnsOBCQFTOJURaPVw4Mv7VctVm0XfQwcFwpL5TD2f4bqxvCUpYVu1bt5lrM5JSoa8Xw7gJhqp7T
OYKXV3e3ESstyfS/qSNW8v9HcLrGR0As2aKysV0QwCsOtWgx8ZRzpGt1ARIzQ5DbyfvbERAHlOaZ
QRaSpBaE5S+CFgQacduDSyN1U4XFxFdJ8vaqg7iC8Mcz0VZVOHqWdKrmumYovwL/Ycx4ta1Txm7j
y4Usp+3NFJmIf0M1NM88/cLo1vgDUpCBPuXYIRVSmPgoQra9OAiDHZw7SNyETrSVzsMC554CzCi2
wPL5GZJ1ZzHVbC66WiLmjaw5REw5e5/+/opP6AOz7EEEA1PEi0f4UV0gcOUEyI5YO3DDaVZPH6YG
iAqxhjE78g2rvtiiAsRk6JSiiRe2HcI0Mp7QQO2AVqBS1yGFcyySJymtj6MJmK4PZ2v5b4271HaL
a3HFC+0gn6TINt+UhUYe7CztUDu1/QhxG/9TdQlE+ZsRYT/j7urabR3SuCxqNTwm89+HPF67s53q
tio1+VniGo0pQGUWoRgbHYru8AT8hY22PXrBABrTuQ07ssk6Xb5cq+V9y93QQboLOaA2+j4q9PGY
guAG7M2GbmymnrCm5cKXVnUILmxJNxI5DGPRggT8xcZG6w2cA07rrnUQghOeXNeN7h56etU7ELcy
SrlsdZtgrWrKBtygedUo2bMMGNNvuz5tOSE0/C28oeDrrmLFzSkWq/a754EaJ/84AmRuhSX26R4F
ArdeUvZ7Zchq29xtGHLEgun35juqLjfQhA4D0fFPigtkFwmu3uHPZKLcgu74Uq7mvGjv8raC5a6y
uEu6dpJYUDCqUwFge9wUJzxbWr7GBuR7yWIe9d2tx3R+74oOrW+Dqa6BwgEPENXHBsK5bLfZqjbI
f5vxNVyCE/6+q+zLuqSPQC9IgETqGVbXwzekPhDU1ffWkQ9Nk67qoFWjYHo+qrlU9/FG0k0YMW9V
2QZSroyqX1rPwhl+kzwStjqQI3VRZfsDzZ5/DW5QHz8ADcqXY65/H/oYx7+L3uXdN4tTed9e4Cy8
Xyoq0J9Npd1gOovd40WCWTzBCmtvde6c9bz+0GGOeGZ5QNK7nm6FtWcFyVyXCv+5OChJfLz4swYa
gaRfxkEFOrzzASrpkReBa2hROn9Q8uX8NzSXF8qDupErW/J6OsBNlwof5h73eefMvp64xRWXRg2k
bXXOV4SgZtv21jSdkdqAequvyISh0WInwP2pzRTHjGhc1CFpsa5ll5cPL92cqwxsJsZhWnXgDnC7
MktpFVWPvCm98QGGWcQXr6j9kyOKEzNYKwgOWCSiWv8OwJCcPuxlnTzdd71sVG+tVW2o9xT5yIxD
c9rHi8T9AJt+9gBCICHrX60amri7kxBRoAhVdrA5deP1l58HJmvvThthCOQRnmJ0LhKbrqtnY1Kw
2kmoGz+DM6ZBZiiGNKn8s+Be/AhvFTPrSRwChiWoNqKUhNvSmUL/a4mQjTehY3g003SgdZH46RHb
KmQUohR+Iu83vQRfglhoOrmguODVk5+G/TspABrSJb9jIJvj6+yoaDajNKCsmReRmeXrIAcIYVkg
DL085gSJdJzpVm7jb0XEHBbN1DiKc06g8SYd2tujgTdibULR5jEi6MNrDdSRU0k6gBbXFScBuVPZ
oYXI2GNssYKy9FCG9GBbjYiC6L/SFioTKDlNQIexhZyCcEJ3jrPtJSgWw5V+HIOKFlguCwl1VrjF
pNc+ODJA+GSigdLCoLtcwh5mlB+z2W90AMy9EB4SJ8MVtdpqTk5THYYHYee2qBp+Oc9F5zSlA95e
nOBJTwSbrXyNGASFVD0U2iFH69Zcyt61dduSeHj3EIR8AFo6nrfCa6eRDHrylBVhrjdx339HR8Qn
27P0oF7b+gXntqVqmBVHPG7/O6Y9+wAMa78loRq7J2QcsTlh8TcWj7dOvruxkbclJJ5zxVJRKWJD
E9rx8G07XvNGwV0HCophVw20Emy8fRMQdrfigOnL+hiBdcmJEzmrVoIAU50ugrGgcvlDMST98Rjv
2SyfRwW07YF0nGwsnI2QO6KDQ/wquGWW4clFp5vam7JS7ro5A0hiXCRdA+09DqFAhUbIQ4lCYaDD
A7YjZCbS+Ejc5DhDnFR8DkjBVbZCPqLl6cSjRnY0+IRpkJfxD258n0NikNcVQ5/8v7mj0GV29a/3
71jT4GTfnZhVSeqfdlr1iTvrpD63r28S6ph5G+hJpt6J1GJmg5GY9FlPM5/fAoMXb8YZ3P1vr31o
LiSm0s4U1DOLs01UF9zpo/T7kzwjp/9ORjpD+lyQLnkWHA5aN8fQYcmTRGuZfVA0swIn7rk87bd7
52TjPs6GwiJOi08IqUyhbnqCIFk6KwlHm9KX1IPf/klGap5h+zTNtqxnd7NWQPIvjHVhUedJCyr4
LsPrZjgPU/lbQucgyS3AkWgAfGNfnotSrHfRnD1gIINYQqC1tcZpVZ9SHHYa1vmb2trFwFhveC6f
DIZNDTdIyvSDjAMyyLX/K6u+HklgvVnXuliKcKtPqF2jIQgP5C9jcWfrVQwaIDq1tOuNSK5tzhUd
UDY6yQUUDov9WCLtQIK2VzFQ9uOlbFoZ/bGQalVm+shUdvLMxymlN8cgbf0FN5BXW/FcxKD1qwaq
ZLQWpbiRCyUcwMVxoA/iEmbCz9RSWLTyZib37WJFxGmbFFjPDn9vCYTD9s8Xj1ikXHgZA3umUCAF
iVXjCGbHui4I+9ufuTXLwlnqHACSEoAZsJZZSDxXr98Gq12V8svPLSltylenVVIsoWBwBigTBYgb
ZOdR0/nirUlO0vNpQuAZowuIisw0ZHrf57MId6bwP2u3DqKDpE7fPHORwPmKuDU60WNSp8EikA4a
MHlVu26vHUuDcpKkRPTeFR0PwSCJbNhaC+3DDrVYoVBFY/1DobqVGQzZ1/ZyiKaPBWgWqxe75j04
Hnp93j36qu7SIuV3bil4cPRTg5SgunyN2OZ8eM9EnaoNK1+5ylJisvYLuGPUJhY938Kdi16wYrN7
pfIiXM232Da7ohEVWVox00NFFsSl3MMmHBLHJOLxisgOflANW6KF0PGQpg0zrr6xfrwksRq5xGgY
iTMv/2lkZB5PbolmvQKNyIMPRJGvpbNVKTGi8jyIgiID9HmTsxe43hU5ajjs+Oz40NVM/mnx+5VH
inG0bwG+4Eehx76wr8JQNbLvrh92p3dzTy/LeP+YWppPZq+bXwD0qGdp6Ns086lsMXWTOKHVTozq
6uxnSmWbBjq1himUkGh8Aw9QGnoOda8REUcCErnLkYRT2O7dgCd1TX7UqbQ+ij0HTQb3NyCJS8N+
FFPnInxiK2V9vZukpc10muu4SzSAPvAJlccDFh5h/4bCW9ftewixHxFYlmc7xssxM+CtCFO3SN0y
0vdGTAKKROX4ueD2cYrDUMIlQfHF/I1c7LZfNpmO2B/VgFY4uVrCHkbAQnk02EdESR43INK5gFW8
5ksIrp8at4NCPcSMW8CVJBzAHtPTb2YaRsjrPnDdiH3NHwZcTfntwH4iCOJZB66CULJPI771/QY5
NQnY+8PzP6AgBYSqBh588lfmxe0QM6RLb2BruS3NaH6E9hFlg4Q6A/o1J0bQyJXOASegxn+X0Anh
X8pLvkIOSOtHcj7pkf11hs6YdiW0vcF8HUp3hnHYi5fr1ncjanlkiqEzr9JNOtcovj0NCZb0Cor+
rR1eeGCRYBeCEQbvypUjL12Ho8n4fNh076tMreHaOboqJRrCON+34zk05M6DxTR0rrF20R9uWwRE
t3GHKKmk7xgi12yQS7ex+nytLhKKpd4i5AlbECrF5xDbJc69Zl7TZtOjoKA9woJpJUYmT3PIv5GH
894keGMyP/Oz2zERMUOg3MCs7ML/3/LY8Xt4Vb/4wrIgoEvaydnXwuC6CLF9ejskmvMaWxZhVvy7
d4cX16dN0u4rGyoR879qw0DCCXYWAT5wG+Z25fc6B5XwPLsA53g0bOjdBylG9YNDpF/XwQVbpzGV
ZndPn+oZrOIUH/hJ0rE7wqMYugHD6Bj7d+imJvSD59FJbydRUb+T0sP+RtNLGSUXte4R+KE931JL
iaU/o/DDyjMWolw4FdSC4mZf4pj2CUUUWu7/OWrjeb8Z2XAT9uQvAbhs/jLShrcWc9dQVtroBlVQ
+2xwHaJRoEdvmPFAPks4yraZvuMw7F0pPTRHYaRnqgSwZ2s1VWQSHCGc4JU4MY/EmxvTv2dMFBXu
B0iJbk5X748tQA2j7pI6jM+acHl4mxzatXXVXm7B7YbVV87imyGvkVUMK1chpuo7ZhpQ7OCZnn6f
BwhzOQuKlCGwbDFGKRRSZsri8Npco0jUTxftB7XHiI9fzx7MHm8VXYuXep7mG1S5XU/6B6f4oIaT
g2n1SXB/SvheRiMmFivg2O3AI87mKAx7T3Pav+F+WnpGX2VaWr+mmp3gkJsbZMcJXJ/avusEskmO
QMGFxrpV1B+8TIfQCx7ffpI+9JSLSNUiheOPC2PlCLTB7xPhC24mjl3Mw8ZjqlpT5tujswznCq4N
G00doEiHhWsXwQ3lY7+aQPN6Am2sg+PDnVMooz90UUecRcvl8R4fJb3FvE6bq+AOyawmBHR9B7yf
QgbcZKQArDpmogm5di+v9niulKlK7MMPygD9fsTrQxDUd0CvOvJpoXuWbbuHkkVz5djaFWB/tOhp
t1RKMhNNWQha46z0MJTGOzc8QcoswKwDN/KpJHYnd/YlGidvaiNlBwWzqBYb/bK8wRIFwrtdFkns
4MWvdb3jHpgMkhlsbXMeB9NaLVloYItaz6fYqJlcIkZF2h8ZZKZPQAglbOHVag7PbcoXlFfiWtGx
ETw4H3aP68g1vNpAEUGhW6Qv0WC2bW6qnAA9aN+vlV3gqbbcRzfp4ZKsk9Kkcsod+oiIZp8DOL+6
9B8dcyHM5ykaZ6HqrY2SZ9J/pQRghorNw5ixxH+5NkenJlphAF6bGRzXH9eGouSxT5HW1wPZVeRg
alIO/SWALKJhV80rPGuGY+woi8u6tkCcw/YOKBevfUm42ie8SD/cU921vkGOwiarRz55toccZDG1
cvSgmreMtY9LczHyoK4lQRh8+9cPjUCCL+8MZHN0bTJid36wLTKIWPvC9puKY9A+JCZ7gPcSEUiE
5F7gERh/hreqQ8d6KU9+B5h87Ta3LCz4Aiz48SriZ2FLc1EYTWaOJNUvYTU5sSqnrd4uF2FVlyuH
1+D6gdVRBpvTMi2gjNYssOggkRfg5DQDSSQtOhZO6pDtQXarCp3T+AbL1bo1dRSYTQBrxaKwDVzo
ocKj/hYoH3aKqnRLAvEEKmnVXCHsHdfhphcGj/+rnJ1LbyPLPD8MO7E2TZgjLjTWJvOcE+S8Uc0q
lweC6Lew0FwW0g1jnA26Hq1zjbPttVyLsIG77BArsbgaOQbbVzlCLSVIfRT23IZhrtSlPmc9rxv5
GAD5yu5+Vcw1t5YZm+/xfVrZGj+UFW7j+0iC7qK8/HXZdpqiEpE4VqTJF/asyPnTql1uF8VsGC3E
yUJzD4J7NMAxLEqq5FGyP8350aIewWfhNQsvmrR44dGYJ/9OSSfYryaoqi5O/A4IhCP/4q4BP/+t
rGQAY2h9bKGk2Qb1a9t8k8qIkTq0lOuJ0NaqCodAlrpvH8VnEpj6+jVUZqpZNBZrn8W/JJvqKAwp
tU71w1v8RawgFxAE5ykGsyyJoiRLMPomIY67+Rsig0ol2xjPUt0FngVWR9SWIjPb0UGDBEzV3HfE
Hvl56eewdhMZc5niysX3kwy424XP+kwXECtd5dbmB/mp0UDQwbrouDctq0KspiOwNHGCs02ZuCAb
pr4JvB20DPOImQbm5nkMN/kxzkVzYv0CvBEJUoZEylypEhLlCnAzRfaUNgvhJsN8MQog5wU2e55J
ZEKvd3MZn34LbNGtgcbQ2ypJzKS23F2fpEHt4woBZpv+GAjwAWyyKRg8cQs/CZUNvBKdiDnrGgMa
o26C0MlUqIDEvzycQz2HyHH1QkiQNwS2yaweVA9GsCGxCCc/UBsxVRAWfzM5lzsympKpR+XruEzL
BRE7yBrzlE38LGaanrEtE3JtPBJrzhyLRwae6xYCUwoU/Rptgs4Zz+VQavqooBGLwUo5uQMhe1yp
8L60SyLYkUMjFaDrlgCEj9Dk5dtYtLe3i+d7RaaRAQa5nCbSMKFPRIs9FZWCq7qFQSWTKRCA/Ko1
6vCYvO1p0hhRRo2lQvaO9gMtUvgpwm9OJjFGqNpANsfJb36XWNVRllR88pUG/vaEaQRlEqUOruV5
DT/I6WY2Tbl5iE/gEALSJN2VHoFEYxsHIUDJqkeE70fQpa0FpHHzbzbF1N5jDbhjYjmEt4SjHwOK
4El6kl9k8qtBI00zhI7YjoETIOmqUmRKwpEytyNgxtzzQjcXh1m+rZXgoChbzl0E+r3jmQH5gJRC
OzvyXUNFNLc09Djujs7b44kjC5tuhUHwvzK8zMu3zN3hFDcsUxttSWBwauoCqy4ZSZxO1GUbmdUW
4lLu6/niYvcm4C8/S1SyUL94/nDxJWODyL0nd2ePuRCBWIb9h/3SzAj5enYF2fldniX+r1vhP6VE
rAZ4GLlm011l8/qJCNt7BpsXujZRjdh/gyR3YL/GU0S0eYs3LxTPVEbmuq1w+KYL/GXArqg70vG7
4ThSoOf4GQQkZc5OaV/HrGTsfNEhbXir1MmMO4DSR9/OQ29Kdg3YasJ2mP59PMEMoPCZAfXTUN9x
FZkxmfXgjTB0ebG4Bp5PAzhVBRFIS6x7kOE3EY5WrPB9MriioHNVzTQSUQ6SvUl/VaKB/n9OfZkg
zDowFWBOMned4ca8yEB9D3DdrRsWWa15hastbIi0YqLrSN3rBSoIu/lEz2S06IZEB40wpkouGVy6
5i+zBQKdwBgkLAGvNZvJzHVpliCXuI7gXgqTdaDlrcbf4GVciNYcqSZIyK/ditc7pPGo3mBnAWzd
AbvLh+xW7G4J3NxTSh7UQauUwsXE4MxOvMTqZw9DpMzAV8CfPtxFVGFEfgCqk4aqW2o/NAyQjcJx
wvAZExSyH/zBQ8RnszMhWv+k/0Jur5EIgHBu4o236Fg8JEv3joCh20wHQI0PTQ188IxrprqJVGxc
tOcvxTP7+HOtjtFi8l3kyVMxeRAq9woSUDxWeSTt3IEvBYK9JQoq7Z8GMOnzlTpbZFUm9ewkSLG2
4R9gLCWerOyppa9jJbGDtCPiZ2/Img652EN0MPhlJkzhJEJDNNu6Zp7At/Lck9bUn1sNO2ecuc9e
qhVDCmTna4ZDyYYQ2muE+LXWLO9BgcV2Yq1V8yoaCiSeHDSvFgExYcuGvV2fxLHm7uqO9qeJrhYM
9Cc1x0nTiaCuRUNpcjVZupDdJbct8qZcHV1J/XXCvlB82oJu7nFxIyAnjyDECtOe5cchKqoGQfF3
xW7B73IqGPRZveb5Ef+T9t9OIDviFethSF8fnagoYreTRH9yh3Ylc+mUoLcgCcnUOM8R4BDbIA8T
diX0rRdO7teRGIbiEpRYhQCJh06HAoE1q2x36J/C5LWaboBoeMHcbz0z9cbo88gwR70Cuvqq7GLV
bKIO0GWmhEOttO6Uy50mxr+DtarEEw2bfqLQmeRwEGn7b20k+GcTdtVqa7CixgwlV2NCYoqThjEf
AXestk2aNcN4hkW30SqXwexeCq39FxqPUN37Zn6Ovf1y1St8Z5XHhoDjbO9NcU/926RPXtDHURkF
/hp8o/FZWbPDRNVS4grZ47PyCpFmN7y0nIxjwud+j5uxgumlDmLiiWnycDJHOjgsJBAnz+221yV7
6+Zzwea7j3axTEUeZoHSTnjZZ2dZ71f8xURsH1SN4f/95okoEeiBTV7X9YGjTYcQCcjB+PzvoXXT
rSdUfLcHC3nl5FDNc2sYL64ztGPhflbWIK+zi2fXN4i8YRC0BxnVXAmpVb4P1L0h5GsucBkjguMl
5LQZLJg2U+TF8r7fsW/MoKcsCSLDwhcFQnv42q0yWdl6XFSg61i7iG4nrq9paInQ4En5N5ZT4MFH
cyziSRmr8Pz43W9Z0SBXpts+hdhPCg7ps76Q39Vn1KxnYD6SU9Kg2JXWJaR0VNuq8gyRKTe/dQNC
9aD1ICr5ruwB804UMs6TDpJrwyPJZAWQ1zD225tTjk0h9vpjblr+4a56eWvF8K9yjpMLKno4HStc
P2rAwI/jJfY3Zsx6ZkmHDRMkFLRdBPuXPrXSz1w+Bp4QkcWZw8uiEBUq0Mb0N9JRaiIZDp4QJ1KB
k//MsvaJlBB4C6fxn+P0n+6m9szSFfkwClgxPGBivxMI/Z4JKrMwPja0bfodZUCbjCgu58ug3Lzl
Acz051iPVY4m1gLmbLFM+uqt7B/R62lIKX9m2t1/mWC1KdSwjQ49agxOWORyeijTo4IKulkLhoj5
UqFzQnGHD592TOAZOz/X6GmXOZMv+tVzAxEtQipl2hYVbrrRh9SNpQnDoIVhs9LFaClG5aDuUH9m
bLzWGTe8MAVj8YJ7+aaJObXXZVWZcy4iPaR7l285z2e8yo86do7gEOpKlhLKUFFduZQyuuAv59jv
eES3TfCrUQGU3wZmhzMc/KR9K5kXWxSfACtJppy2NMhalD6Afg7PUyT88FSncGoZfWl0FfnwfyYN
vXsMINBKre8S2muoG+09sJQnf5kjTiWJxQbsiFd0yMZWHWvE65UfEXJneuwmX2bB3D7u7EQRz8xe
0at0Kmn0qnIGfQEyZU4qW9wd78d6rWw31ytELdvHiWdtW/Ia+v1Vi++5II28lWmaszpQ5EL/bLhP
xJqCLyFCKrF13f+zd8RotGLIZjqj0b0KT6yRnrATLrxEyT5tN+R9WgFVqQAEWWkzgtbm+Nk9ZuAa
ddqXGSXELXxC6mFIQc4JcILkr+xkDiHteUpYUaxNpWecqC7jSSxuiLNiNxeTGHWDymcNEF7/77lV
uRePygvGu8xc+T4IHvTnX4R5FHwqmk2oN4Z6XdtNe1/yU2wufWE7VmymL5kAkt/Bc9pMWvy/UEez
wBOYDGqrEU0mGirLdneuAzUZkXa/+lcKIuuoMXIhRUlBrjFdAi5F5sN+LVTYBfDHyhvfSj7LjbOS
7C5RGd0szzs269glzSWJVjpWeWv57cB2xlw0RUXhyEulBxNa5+a4yZ3oA/gzE5bRlEeETsLHpWLC
fmcDFTtJuKETYTPo7Pb8SnSTGxLxLnkeydF10WiWxelbnu+wBjbRFqWZM+SRiA9aaWxSToBDKtE8
UYUv45AhV8AP4XA2q/BqIsG1SWPFHpHQMgOWjiyZ8kESRuztYOpX1vJsISSmNPs0OekZ0g9MguFP
eARe9OfCx1cT3qj97ar/HusgsiSU4meCgX2fHapsi9uOPstgAYG8t80CRkx50UDxJjoNht3wflFC
p7tn6t/HEN9my/m6AlYC6Vm4fc5n3jeFxAcdxVGrO/nEEQcRR1l3bmc4N5q60x3s/r4ItUfx4hfl
7su55xGu5ZlSVufzwUCwUtBdCSbv80lyjDxPL1vfTI8QwpfiFxAYI567balRH/yjseoeM08UKdPA
ezXuiZO3VZfnNjSyMAtby8h9P4bKj3Tr3KQ3UTkHiRRxPLdsj5jKQ/NOOcn2tlvCYnM7ouui33K9
+7kz4ZK/5o+cfTBm8EwfHX4GgVfwUcXUAN5zKYHXt0nFLvzIV4J2e5ea8dYiFT5v5FwQbRmUJzBi
SoGZnR8ioAYminx27KPYFjtnt8PW2lgJv0ZmfAbTLSmZn5dRt44+ksazF0MYinQCh9CD4In1zd/l
d2AvCSy3u2iC0vE9PPJhAAM6atfueXLtkGlyoUSEWIY73xPjNdbuHRVsju5O9yi4xLYkqoZ47Nyd
Qepztp2u+Gn6/dLvHDkGHAEAAfIDdqI2wSTca2sFhCwFl+uDjqGMmjjpoXnCkSOgfyoeEt92izWy
TIBdju9p0CQv09LRSoJpFbPDUz4X4dx5XAKbOiK83Y1M2rI0rdpPQCEQAa26m8DgLog+xPRzs6jx
jxI/YQlIH2lv68+Phu/GDIK6GRZWWVegyRCTJO3nRk95rEF2P9UQ3kvth+xSPJjHkcPUfaumjXq4
h/FSeFEgqDG/Nl1Ef/5MPiMmaZ2dQZfMDfrYYk6lJJf9qA4=
`protect end_protected
