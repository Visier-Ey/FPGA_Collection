-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
iDMc68+YOrDAd0pGlyiYJ+iG/GSLWiUMhlbtrJ8qa8rj3sxkHHzN/lTa+dOkNl9jJkf99i/ukzp0
OvTzZPMDIJXgK8anhib1gPzba78bzEEk96dZra70/NPB0K1jeKETyLGY8siBU5CrOYyJTDIsM4Ms
Jcw8LDMS5r6yS46/TejD9Yw5SQEUwRTRqiDemcGAL4/RLM379jRW1mRyriso9H148jRQuCiVDDfV
iLqh/ojo+JqoVdzzXp+c6u0M0FXt08GI11ITlyaLOOY1wYU/qj5rB2RmiX/29uVpm9B9Gz3lMZRj
8XiWTGiVAfVj/uXAh6rueM1ISTBdPPyNxRzzHA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4176)
`protect data_block
NiKDroYdkxWvmwxOBWMcbUfjAQ49YGjJ17Jt41l6k9+gw3EAjQ1ekE07qBqzxZTGCGuZ1UqSHdVI
nnZ8utP+QGCqBXfUcGifs8BYYSBg1ZrFqi/TPYoFFD3m/VLptpYPsLVy5YNlL0ktPF2Rr8GSO8jj
DosWRpQ4R8E+eRQbm6HqcNRqzBHRgXvvTdauIKzZKsLWHrQNBaC/XJ8/UzB+qVK/7St/BED74dpt
DcxI8LmzGAd0ulj4cyzhHhytKLMxB7pG09znitI61ttYFkcUPvdl36cCvS0mcP57fgmJRuTirCRv
6YtZOd6zQmWtnZOb3NMXCqeiWmW7Ys+1FIc8dYJ3zFdJI8SbFmDfaJNM4m8zKTN2lA2/tgeA69we
VvPNN7X+CRy1/aroGIkugSa55s6FKpsU/YW7YmzYPdjIfcbWEhxIZZqGcKZNvZUHqUa16ER9O1El
89Rj61t4WxyhYAypv25MR7p3qY/vWjeD/Mjvlayd7cfHvnmecq1g/Ho3Tsnl68EmJlJvR/5iwL6c
PrqLzLAnkdKYRpdzGg7z0m7I6FrqJIblvMOHEgHMn1m8aF5lMQo7ak20J9RxGHzjw9GpF0zSQegZ
4tBwym032zKwa5oVETNmoMUgHjhrGVKnkQaisFOZeUX3E6i/tjVP+LJL7NM4PFco4EmdwwPjbJi4
zE2e4TdJJr+Vj7FqtZc6WPkeb4bztZ4/JhIF+Bg8FYPRyhMES02SL3y/gYCxKhKC0gfnqLxT3/Qs
gfobOPrNsx7WtHBdVdQ0/J24FpUFLw43fF8cvI05ON1tYYQy1eHXHRrh4S6b2KDnYgXbiQKYA6cC
aRcJterDK3zBZ5WlB6D+lKIQPt9EkUHQ1txNs4VjTY3e8eUQ9L9TJiRH79QIrTuzA5+Ef5uMFmK2
MZGZSGuJnvw4PXAcaxDfRG58yd27XHPCg7JJk48qp4N8Rn5GoA6FH2vB89p7coPbDdXiRQf3Mihn
7p4c+3zsm2ZkoscEubacAqEesQICkEVboKnGK0qb+wXrYa0cMHbjT3gRuNlI61IrqHMenrbWZrOG
ZRmVjMYkWUGoeUEfxu2EGUhQlR8KAxwWZahBsK+oRj7Yq1homHAat9zUhGmFxfNWIdxfqEIxWEwJ
cKa68c3rOpusUpVG7SGgVblzFb0hHl0Bu4ocKIIzwQRDMY6cP3le6qK85IT31a5qo4hNIHsWQ7UH
i3Mkv+CuivY3G6yjpvobDzkJXwviPVr17qTH/jY/0OQCUrO/FhUBEcv/qI6dRM3N3sM8llFrjQg/
Yx54HZH+SAon1qevBHN9EtNXGQa5Ka+fnhAJqe0+j4OlvQ4kIs7HBjXNxiwbqeaUmZuMjSU8Bd+4
Gthla0BPYsiW3tVkF1eazk/bKTKEGjer66VVmFZFjnonba8tQONHeMW0XyMmambXv9qa/Lxun0s5
Ya66yWpKfy6Gakd5+jB13orL4QpmU1empP76+h3bL2IWcAhi6l/in46obq9lF/4iwnZSaofRq8D7
islMdU83R2U6y9dx2TpIFbF492nY6TGnzAAfobt68skzRcOBDSLln9HGHpY/QAYF+TuoEGh8TFYx
yEWZE3n8AK+ijvU3ynWlePoiyV+myfGcueUUuPw+ZAheypuLLwWvkpUTkHkL8SVvR7l8ofl5zd6c
BfqstgAc/DRxGSaaYBOv4kphlgGoaE29vUVuvm6kpP76409J1L2+wqj7XRp5jHfG15zRDeFEkzpP
hVn8V+o16YqKx6t5GoRgMfM9OKXTvomYweOpuISaQSTZ0UAfVCAydYQlWwMIDUn2dsPupok4pRDV
DSDvu/kNMXmpmRG8REWCQvhcclSpqx4y6Of/e7LFgBf2yw85YgjX7xbXCDZAqEEjVJPK2/LYUNoT
vlFckqHrVe8yZf2Nzc+Dz+6c2YBwWwU54EwZaB4xdAmI4aUcmi/z/ifPC5VQ+Uyj3XtBariJ7IMn
WertbFF4Q4MpsO9E7hEXsa3boj2dB6gDMwqgZYNUAKJGbyjX0qyzzYDoBzOIomU5n15sbYDH2kGQ
JFTJY0mkTKvXiUOBSHzbYWm2Hu6rAAi4dcts/Q4NCt6m7z05kzG2kRbhymfM4oZLVq+Irrbp+wBA
XEmIUdfnWPcFNIJxwKb3prlQh6R0jz1eMD+mfQ2hmQNqaY1OLdv5yva9XwAF4hdsfsyVjtwY+6uQ
R8ucgAbwHJXEF9EMTEvoP2vhAblHoIi1pu1M/Tiir+F3a9YIN43Spj5XhgQsE3epr4E/+LwR/PXz
lvPLFbi4wzei7Z4fn+XWko+kxD+RTMH3OTFxZ7nlrSCRWxpSTjVSlUEFAhuBzok9s0D6IyaGw2AS
1droGFYvKPaQoxDvzAa81Fn8W4GIF4z4IDc+4OftFjXu6Rv1U+x3Q1zIkmzICOf87ttYMwXrDn1F
AXREJZa6JthiIV0Q+kfuMTSzKivdoRxRE0xF2Sw8XQmhG2gF5y9t3WGuBuvu/yIoeSgOlqztKKqd
FalfrEIkLXl/LCJlS+XDxvmC31ZhzOByJBvz2tnINNAbG4i+j+mV31A2P8u31WFuHrNSHOYgIpx+
qUAmpdgs8UWLBwUtkhtGUT9FXdI6dSk+GI3rdq6aVZt+ijZsCeyMFp4JlIbnznC/AB86mP+jHonl
B1oijgunTAIMUi/Kp45gemrvu+jHKn4IrJmwI+qxxDQPvROp4JAzoCC8eec+AgAzN7k920IXm4ok
91J7MrfbJxXWVANXqmvm257aGPXkb5HleDfGX5ERTum4S2YPqYTGBS29E9tbVkqYHZkw1ouZVALE
xopW5p2U6pd5hOSoEMy+NDI6pqJUW7v8/x7b9wqSIzLIAAVm7wtVPBdoqRYKRw5LHP0boQAZ/9zQ
WzU7Thv2MTL73KaAOEjpsgCHxgc+OwBD+UDNWiFXlNIyZuQWgPypsqRIrC23PejeKDc2sAuvqnKB
yZZFUFxhPRXRN6wA+OC7HhGmw4drcyMLLkt8JDVG8SXIR4K/xwyRN/CHEx2jvqb7OPZTuYvrjOv7
COaAY+EPGcxnMxyH3nARcpqKAW6iBr2Wrl6gh4Xe66ct6jtpy/n0Om+OKSG/vJ80xmpobWDsnvwa
lWvBtQAgD9SHBJ0pAh1yElkmgEzguXwjSsA4YUasWtTVDvfYN+0KTt9caa+MXHEFa/pX8w90z3S8
12FQ6LUD4ewjV1LcPI4ViBrTZvR4txv/EcGIPYZl5g8OMf6JzaaVaTZVDmuoMBruBrCWZvfbiLlR
nMwXF8o9mRZ3DWexu5cH/W0ytUztUuxf3JyxvjpbSsQ9KflgVVLnySPmhTDcET8u7IyfCYRKJ3y+
mQtnrMS9vEyenuUSM8LMeb0lug6ySPF+hIlcOJru7NEroUc3Yrz+y8ovg2VVsAjZLrQ5xDEMeAct
ng6pziL6Gn+ZIEVq+z4BBUWsvqVu6xY+z0AMqJLVu0L3JSciVm90uQm908bmmQa9BM+UmyuaZcwF
/DL+hzgrl6DngaDqNOVi3X+aG/c2WA8lBQOsqMBwZn/T734mpICff1hEXW7hEwAwRoZaSgFOPukJ
5HN8OcnaC+AmZz0wuocOxmKlXcJ+/mjInuUivESXpOVKCLZRX4eHN9wNWbJvLYaBCgdTEWoZYoYV
FrbNlI6cfDt/KstybxMo/agqD2RYb4Sr2gK8v580BLtP5jROkug9foAc5L8gSeuDZCnuEGwoUt2+
LKY54ojn2V534yh7LsEt4GRP8OKvo2YI7SVIFl2OR1aXdJH7zvtCKY+tEIpwjXfEMXUqsuua3vCG
QRbsjQ+RwVBj0+jwlWHwweA1upsPY+Vkvi80Seh+miNy58TOVdNfvNeC843enG3zkoUnPEz2FdeD
RMVDbncOeI6zVl6k9vhTSmKohEq84XjFzJlRspFWVrCk2+Y4CHfs3s+YWM68JmzCUyo77jcLcQ7r
94XulllaodnR0sPsCOcj+Z1hGSQuzsRTHJL9i7K62yp6HEs+F4QmyRffHasIjYUG4Ay7KnNqyvca
WWY2QF8uZLPEeQBMmuN/bDHQp4Rz2t79zs2R7paAvrrAPllduK2ry1nzCexKI2fSRo2CMXCEyl7L
WRxSThQMH88od8ljFXKP0u3kqmu8nVJljdqZV5KL6qcYic1t0fZITqTQIC4c6DgQajIKbdGxMKRQ
xVry7wqaPwXeg9CWXWHiZY5WYUCy0NV3MhmQ3Ap6V+8cvMp9mtGsdAYq7Sq5hpbEoBrS9PioxDlh
ZK9S/kq3p2uwBzcaFq2R1nFCEtz2Fpd5pUIG2CAREIhYbU5jprQrpv+z5lKsJMI2Re6nV3bKxC7B
/17r9AX3mECkFudFWPO5NoSni67/lkDOFpDOwji+AIbSO5lEvlnPZwiLs2zZd26MimMcMxv9xC8B
LI93V4c1NRGnKuab7tD8IlQysrficYLp4Dbsc2R4KK63XuUxPSNYviKsYOVFNXCCtA16vu85pcol
Qjbj+Iaz2iqUYrec0qveOc866Kn81kh/vWowertEAbi+rfWuJLiMInSmiB8YZCwWAmuHLpICOsI3
sIeImhyxRUnpsPpcLxySJSl/3ax8M3S33dJ2YxboU6AZVo2N5rnblPDIlXBKYzm4Jrmti8fi9r/L
6PQOuINxW1dQ2/6wagcyjNkNxGByIFZDj04pOQh0WxQYKqqHnCuH6ypF9wlHruBOPbWY5q9kZ9dl
C4JjIujR9IEvVKfroSJZqKiyHkl+oae0YJNwZMDQ1HVU+2ZCn9mfthY+QsTOYJP207+nu3nKKKb7
uwVyi8VIqr13Sh714sEUKvHfTt6qtbOb8FHYZ0EtxCGYOfaQ1jPTtwjuJnHYi+OiqhdIQPadbVFV
6Sa0V7Ef99L82G+onjA4PbnB4McO5fL4zHgdhmXzwZj4Lwtm+Qb08TYL6nPcDcDApCFZXsM4bNKH
EAz7QV9n+eWIV7Wg3hLQVWDeb1M9k73DqdW6HMvaAyKilxmqzqAWZjCxTQzw3tNpG1tsxhIWZJ03
apQKU+60WulegczGTGDF2RLSVvA2Bvf3+6bJ2w5Y9OxHEQj1h2JmBHiFBlnkYUKaMK0a2ZRiidn6
yUOiIa51Lb8xKyAQyv3Hni5VOjvF2/sSRs1rkNXnmEWmSyW4+4UcvQgAeX37dZBNp5ax4PbBt0iA
Rnyq+fpy5rz6Atvb+b6XuPlaOWTpGdaGS0/Qhx5eZ7dXl9CvmC0McUU+A/A1/Ypzrt9SSebqfK4f
nic1E75iai/m5+SXZnM9IR6mDEKyGhwhQrmtTaXGcVRfZBRZ/6idZGDlmybWJ+nqumjo8ThzDK2i
9Q+AHr2rZ15qu5FN38j37ygQCld8d5p14q0mhvwT1EK0EFK78JDZmNSme44C7Brs0xLQvC7W59qC
1A/U6U62Kd5jrmraKSpiDBv3ESJfiGdPu3R4Q17itfdkJpso9Ivsm8NeK6uKWKtIePNG7sntDoI/
CvZeE2QGHkCSi5XzN0qehn8RBtObtx7QI9Xx7OA8xMASR+WClRMGsquALq8/M/xLwYJ5WqS/Aty0
ZEKcUofUDlo+PnSpZQEG
`protect end_protected
