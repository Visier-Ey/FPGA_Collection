-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
--pragma protect begin_protected
--pragma protect encrypt_agent="NCPROTECT"
--pragma protect encrypt_agent_info="Encrypted using API"
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
--pragma protect key_method=RSA
--pragma protect key_block
pSmc+USrg0cROKhaYmMtUrVkpxU3lffOEuoIXBh6zxwA1rVRSmvxNLr/O6ERrssJ
KToF3ZQkIwL0Mu08yn0izignsxUJ/yvtdggOx3cm0K/aY5WD9lMHkvrZYjGkyeuq
YEOKuQr+r3VVC2lJYxvsA3UjIGqz2KZSxbuf1dY1MlzyeD8xeBqJihE1MQyLRNCg
dmAgQt3ZbMLZG0s31lKqtO/VAmKTCHmoEayeUU03TkebXUMjlsbugV76+MOhm2g8
KGtJ6i7rd1B7E2qrA5JBJb+Z6YAYI84phbgygTmQwnD/3d7mvPLwuYxfnI1E8nB8
TmxIDFIy76aaWh886elV+g==
--pragma protect end_key_block
--pragma protect digest_block
Xm6KGfrAebk2gSnmUMbJ9jj6Q6I=
--pragma protect end_digest_block
--pragma protect data_block
3ee5jClTt5h6akXayKAu5qgFQA3PVZd/6gohhE0BpiGyQxTgjT6KbYo2tgaZaVAn
3a86KaMoYnMMGryyjHZ3EK2/iZ9T3fqnP9ZghjgwiTfLkvCr0eo9hpMxeUu2yGm+
l+8RJ+C/PcY2ZWlaONTv4mxdEgAOWFHTZVEExT3ZvzRo5f4jelH92xhmkFDsVxuG
OYhuvOboS74ri6KIUTJjEiXURjzwkGFX9LXHH590ROb5p+G3jJFabGlRZMhIRAFG
IWYbYPhA2rtP8tPed0zns/2ThqZ8gBq/IJSZjSstegfbkKfDgw9XI4Isu7ukz9+D
cRQAF3KgGvGPzB9Sta4UpIpwJ7kxNds75uGgoXwPW7dP6cGJbESWM5f3CXoglll/
HOFXAxqoyqC8pbKzOlVz7LpEH3VSimMuGgqMWij98BCUKuRaTy/L2I3HmphDbw4U
tbZm1G/Kws0PzGgrbBfSJy3C4zM0R2dogc+BgUMP1zLhwxcZ7xnqfLoewzaL4lqb
lgl9fQRLj0+unSeOZvXgMO9YKUleFMyrZUk9MOa6yuAz/6ZqcNDhpylOu60rxeU0
L/45ZbNfMKCBH6BdS+Crk5SHu/YM5I4n9+IFwC90qqthiVjf/MOkUtl+rwM8bhVV
YPu12Vbpl85R14atW6ESWrFw2vET0Vv0sWrMaM6kVcsYkQtaP1PlqqR+9VFZsSbF
+aFQmMEJv3lvPFfcN8OyO0f+3Bo2I1CAlo2JVIHmXYO5K4NMr08t7XbSn2jY1jDK
hgXao/VGsWkkfyKeqF+KUVH4+7GGD5Jd3oU24IsoV8f2OSQY/6/GHwUTTsaTiPKJ
gJ0qyzHpyz2nD2vMH3F0gEhNJYgbwcL0iug4P4cb3IyNrpfv5W6bpeV/Cnqy4/Pq
kGoybzULJkcfq3lUuZiy8wYshkMd2piTneTmTFwzc+qKhIlwTZMh1gJblVpIeA6F
CrIyd5WrDyKjfk0mB1zmue91r7kAZupNYW0fUuYpI7R+7gqBw7hR/ids5XFdvdMC
Jt/gYilmZLu6CEYy2BCbU/HN+phjLc6pReeymjRYRXp/ln1JcxCFnYbmU2fcJSaS
6nV2HjutzBOjqZKhc6AHpLh66TerMVAapGOfSPX2c/S32i8KT0w2npWGBli76gaH
JAwFcVKOxH/2ck43Tu+CH6OsG69Grz4hIKxomlpm2RTk3+QMOPYdK+/2C+lFLjBN
HnYsXmd0wAVWRjyjawZbwyrkr1NrYqtoRzDKmVpObiNRPb2LS1WNI/PZMUtv3d1D
tpcmJvkvMVleLj1g8XZ+7TFhDhlIacH25Cpj7NQfYiOg3rAdpNAnzwB6DCxva7Fh
J9HSl1lcz0rtc8qoDASwPH5d2XGWyNHfKryK/ncA+oaDb175n3B3eQm2gtt/6eIG
9uDfMkDf6CHJp8T4Rl+7phzLRcVi+hRLp3/y56ragncVxmrfLmC3ipY0eboyGQaD
wAe980RlwounGbI1mdYEutWyrkQvzdk69eKch3vmVQ+Xvgk0AKh2YzsjF6uEYW4U
xwszd36A8xxViIc2wdagaRpNJACtNexTg5uTmnaVtSYFYxpRG4YO0OlJqQA2rZN8
TG2lyGZHWXAeVXxRtYZi8qQl9+xE/Oa9GSCbB2VtzgKSBQzbEEGSVFefsl/RcOen
nkxUpsRAZzLGvrfQLQ1m1ksjIDVLPkugZA7IFFKrAn5bfWc2+xGL8dN5kneN2P+p
q/XdEnffqDR6Q4bIIp16u5BBD39X/RWXpZwunvUYhvCeOcKyuVSIMPHFnpIR6/3s
e3wokLu3FAyDGmil4ImjsR3KIgQXejoL9EId24nTawcCNRtxqxznq6Pd5XN2emVy
wUxHRtKgHD8Y3HwARZjKNs3mIP1K+Ki0nEblppc0RALz0Dr2LdC4D+a92IznZVXv
eiAUvZmjlRv4xbqUDQpJw23N8d0gtrMNUo+U1JRw0RIpG75APO0v9PcYlpJzIt49
9D1yBDr3WJalysWcc2sTrivtabnV67rLJHxaor0HcdQ5FuQNstuZ2viNZZ1fWLZ9
De7bZhDFG8f6+pcaE8MJhotUB8SOm6JosivEECELK/K3x5plaVQcxTcJvRyRgYjh
tSd/DMmIlJUyGNb8/h4GGxYh+35JPgmSGkQAPGSnfwbEKquK3KEavNlMoixgUU0B
kE+pY6OqyFxBXSILawbEFX8NYCT573bT9YZpGxGgxM6YIOnAVw1hYBvGTRY35Z6Q
+3lwQJQVmRXikXbAitX2V7FZliA1FilDhXOUHugU7HPDSIGuS5ph7knuNtAXLRvK
bLR1nKi278rwlKn04eUm9WiBpDhnOY44BgBJbvi6CUGOlj+hYOwERnG/RT4r5GNh
MA6EGJqKYKaqujn773BkYCnFw8ucGwDtxcJiHv/0HlHRFwTdgoRclUQY0c1MZZcD
r3ywxXopLkJO2i+zDhr/9Hb054lAw4HzlmtDZY2Hy/FMKjJovrIBPur7q7RR2q0b
tACOZInMWsJ4wiryJUpye46mVVTomnOuZ5kbrxUUsNssEYeN+33nVr59XJzZPmMk
8c5KaQDYiOnbo0Tpi9tCvM8W0wOVY+G5ipCMva3Fj4Pj2DR38E1DHHdMTUada7mP
l+2QR3nq8aYD+bB4eXzwna1xhzS42Qa1NBSKzZ3koh6uCcPWK0gQXx/2M7rncrpj
2ZiU+grKjt3BOhlj2f6vZRqOfWOBmr0xlX/Mj0PAA2nt9qGJ+hnf9YXtmZeYK1/b
107yZXbQ2l7HbVP+jvLEWCXgI5WYmJ1IO2+jHKgUpiDZtRfGql8ztXd+aDf8X1ot
cUQSN8UJSDajDPFuqEann+LlCYChti9toOpTEjgPl+YCzmzs7s5L0meq+wwax69Y
dxMNfHcYbGguzvudkcjtSVJDiptnFazEUee5ntSI2W8UPYOajvS0+xqLno3EgCuM
5tSQ7WMiAhP/cP47yzW9/kovTySYuxpK6HhRUS1bFo9xstn4zwGI0F20gtPuka0U
SYq8k/tR64U1APVUFCG6gL+Tth1itkAg9nhFQrdSixL9zyKWVV7dtJqqj+aT8q8M
fEtv6avk4ljG5JNJxDV2j1TJDz5kmj2HD9BYSY1y5VGRGX3VA6LB/q8RmZ7s1Lux
CSsBH3JfR8Zrma+q5Ksc5wWqp5kgsO95nOdIaVKIdoXII7TcTcbJzb464KvMImzN
t6ZMRNArmgYZ7tCnTlbo+otXGJQbzqmcZl/z7YBgmF4a18Fg3l+UEE/fOmsn1e2z
peSMA0cMcgZ0xgsIqvwY2VQBfp13XVnPkXIpbe1B0KmuOpINRhg2HDHc+cscTlcF
onDnkJBORoMbpzoNFCDOlAyDAKmi6e4vQmXEVOSPPIdnWuNW08LS5VhQeYpT1KiY
jYUI4BByeyopnpVjMufIh4lMyhCxiuQoaNroI6UdjFYtgk5xLzDOq6fAKnaF9eml
dogq5ATeNMGJVqfCk+jRPS4DngVCJkObMfWQ1SN8nn8fDwX/VtAN0vCBjucJyC6M
ejCqJmUIxj5YGw3nI9rABrphVAJqQA6Mf2cfIvuxiObBPx0a7MvhAnY52RMjRh8b
LxPWEUq3NeDafu+Tbs6ZygVdE5KDGkkvBMaadF6T+p2mJxYbSgSzlIxSAwdv0fi3
iPgqgANSdsaKu4oEn9/Lyv1NUYTGm4qRBh6zhglebhYNdeAnkDXHA8cHVgvcAXZG
N6CGI9OR3LcclL9WHQCUc6ibIeDMN7DlFwCtn3lrwoL8DLQRFZeMfWg9ywNwAhuT
wjgcnJjRyw+z59mfjNaV4Sd7bSPzBpc/huqPEkPYGEbTn/4zPhtMj7vj7jJZSFNF
KMwYA/tzq0WZAtdHMf3Bo260GWwF+/jx0BrQkqGsrvdUNowpCLPHT4QlzC6rlJP9
xprw4wY1jE9vITw57nH0akCcoMKSmlHzHOMofs1R1CmlNtYnOhphZD+SRTW0nCTS
grflu0ZEBtN7zAr600QJwG1NIN7u8MuAVU+z34hK3NhPWURWk548zu6NwklveIxI
V90fZEGkgIyUlR8CJUhdj/OBWghjFUTfGkppejkxp5xddso/4xZMSF+96RTuDKg5
gwfH/VQEaXd7aWRyttHEsiSunbkZSazMviGct/f6+ihIAatI45x7UaBl8AHBRjwT
yDYwQlwi5bKCKkEvPviNavizv0uqTJB41Pw0B+SjzARKa/ylcAX/nxNY3nc3nVTn
FYBFX59lA9RxfRP/9Eae7BQW8UW0qR+KqU6tdvgDLpfvQtsTA6zhESB9hLy/opSm
wsCCqAKE69yClu1J1blOf97l5bfE4PWpzVIPawuhwvgfiQxe9LLAo17JHpk8HYe3
nNUp6SHxrUOGUPRHvD07v2nsy6Vo10pLkhTWTssX5CO66xY9YHZogFTSNnY9lNW6
hV7tQIRNEcA+BaR6G2rrN4awjE2Dsg3J7VbyWMVmryQNW+49K/EJnZPq5T3wr4Gw
QuEBgAlUdL8WuFGpUq+a9CKI6Q1NEAwDA0q1iUhp6+EAwczR1q3Oqf27aNGBG2dL
HnfeBBPc5vlwYUwTqjORINu38x2c9rO9sSX4X3dNUlsiJSOoTT5Wah1hmAaTgZQm
h1W2AAC6diH85cMjb4B9Mqxk5ZrCM8XJzDgixJuzoatb2/zdkKZitxUyuC6eDhkT
1vBBDUh/BeK77sCg+bMw6EBGGIBwOREqnGDI4LSpoSd/47KqZxuURI1glF3Jc8Sx
Ov56Ky9gZFi1FSvx8gGnLg/xaovqPXy1aXTYyHz5p1tuPYN5v1yiX0SCJV8M/LQ5
dGUfffH6tDr4EJkCqGNKiKtB9HwNJ2vhTCQ5b7RBCQDKQcC3j/yFMiF3RVochT5Z
n7D2gGVi68AA9wOXRH052BcpDdoYzoYUGLPwKHRiugWYtcXOgnbHp/A3HmqaQ+ha
xxA6lUOADf/vWwRHlGfhuU2MRtzwjeiJ5UUqyrdPmA5HRu3ZcP7Tw+Xn40P9nscr
FYkt4EI/Aq13L6bULXtUehELDcWeDI3KzH5SGtd5ec7veXGprT3SAN0PJW5AwPMC
4Cu6ocImpuRX+mBkFElhl/pOSdl974SKOHoK4v+fT6L2KjNgpi+z5h5w7KMBD2Ae
Ci/lbTG/Mdkc+7I7GDvxVlzuiAG849GbYQgfFUXyn2Y3XgMpHsIXr47V7LRLZOjL
pzAgUhAoPRBUm8AA+yioE0Aj9rexKOOrPLv6atkUzLvZsTjvhXNLoOHDRJEd5bJ6
L18nvXqmN97BgSFdohhsKzmAaKbvr8Bl/lB4IgJJgzIillTDgjaykps/kWL004fZ
sKtU9KrqhSOyLhP0VuoPKbeOyQEc0wflz7MMPlTmMB+oGUIb2ihxeDXP5T//0i+v
gQyFicl2+noS5JtXYbBy8mTOOjHyAX2MxLetNtEjzUttg5lnUIBTYUoRMGb9KqzF
8EeFfi0gOCVPgn8p89d2SWg1IMALqxg1RJDbmyuxlN2cMxXjzLHLF+eh1itrLu3t
ZAES+urO79/r2zRu7OW19gWhTHDep+KVRgkEmj7MVcvrS8wOHD8vJPnYCCWa8Pcn
N2EhTDp83wzhJstQFLknEQAnGhxJJlitkyTMBeafAm3A6OYghw0YjJuqw1Ay9FiY
8H1kLZs8Y48pXdUYvPuqJLXk68/hk3RNbyR2MhEscZaIDfzUU9jnsZf8upxKQUJF
JyKGfkSI0UU4gvRi4TS0m1jQrPIPWHQJ0aAzPeA/zZTZb1qZr7Ae4lgx72qU1DWy
prCb1lgXZ9vwuZ/OavRGNY077XBjJJSVvzXPn2NXONUcLSsMYF9x6/RnSMqvujA+
/3+gafvpjz3Vjsve8qElq1/5yARUrhO/7tlqpsNwEj2yDMhDmkJ0400cEss0UCZW
Y7bFVavCC9xeFKZkKKFg9HSwyDe2VRTHDXruvjyVE4wWU+EL2C0YsWDSqa76zons
dHGPExYOJkxswBtgo8uESHYAsMBbaIJWBf76i33mxjKhOn7/D8AqgcCjlLKZHYwn
xAk3q1aJnzN5ge/zmBxszv9fcgpIlovaJK5iHsPLrRTZvR7DXLR6Ze2Egk4PjGQf
HXYOtnc1b5YTjVxLH+EVoEbo60Bmwi7MgZtE7z/7Owos9wAWluWKrl9d8IMXe3eo
TbHprIx/+z1s3I0HLw8D+v4WF7v50omyY90iODAZfQYySIrQOvi2t5AZ+AOQFHTI
HaJyYQMk3GyXx5I/Jcv8EKISgsLx5Ng8dxXm4u/uTPGdOOgpbISk5yJdwxKThjfu
0KHSaGCvC3io5Cov+BlAhZBlyOaZlFgtBTqvm1qceZh+eaZ5eDLUEewzvTNDRnGz
IoOxPr4UkjuCWBBn0tWe1QVT21xjZksU1PrWZFm2eXNz4qQPbiaCXyeZGUijLton
rA2/y747Ey/wZMz9azEg4JdMLvQMBpfUHtGJjFh2BMFKTt7FSSjvaq9sck1XHDIK
YzOA5oLRXSKs7IzNkvSXFCp/wQn4S/K3QdSos0Hgo1mb/AJfk2csWFOwEDPDQXg1
zhNCS01gStnLoSsT8/UCn85i2313nxCkDq9Qgh5lteh8kGVCFY7pyEdkhS5tIRib
vmuc9EtioBVdpvozc1E0R2jZxbWRqRxplIQQZd5VV4RGo1P0R62nfxjXpiCJtWpq
qLYybNgx98dZoML0SV0Ovpxl4d+R51VuPCoyxXhuH7bvCA8zSiPCw4itKcty7Xtg
NwopLh/SgSQZTw/ARAJg42yYFkCiJ6GkB7qAlA6sqP9ne9C7nI5cJq1bdeQl4yYs
v08tuGRn78TyJoS749xAInFbJDGrcsAB4xSVDK2uWJu3dXyt3nQRWI9peobCCQxd
pVhhyibrQn4Lqh/8rd5E55nPkzVxQEG9Np53oLLzZrPjmOHmFgHNI9SUG8jPnxFk
y+tgxYcVkFYVFg5jm5hdPIvCceKYt6krfKB/Jm5UoBA3w9ATurRj1/EGOseQcnhs
+nN/hVoAK43L9Jdb1W71clovLdrj07D1WzfwhD7ZmyK08runNZ3F7u3l3KzgzMHR
TjuSpSodehzzi3tATFK86UGrJiHXzHjeWHTs+yZ1SGfUsZWC/6J8sH7zb6tKDJTv
K8S3kOT5IrA8aQV04HnADRP4nt0QgftywqPUCtXmyOVihuWRvjGdlA5vUxAhQpWs
V8rX33z8fRiMncyueHX4Tz7dS+DHF4Wt7SEm6tkxFHPlA56aqOvB/3BmIQ0F/zi9
eY5ISJ+U/nci0RlsYrlOS3Bp+vyqzW8vbc1XabfytvK3WhKNrokWPZ1PvxOyuMyu
Nu7VB7kCGWjge4qejLYZfBtbbH8V2i+IyzrxysUchr189vdt/5IgEnBfyGR5l41G
wJ/2NKpTgi9QYSvjOhrxaupLWuNmNIunkqtn7i7eRYt4WJSq/xwWaQAzpQO2Awfg
9YlTaXxW53OX174hJCugr5nm1zWlehKSPX8cK51UBaETeZF4wJ6mHW/Sc9Jq22Rp
saxCmUyPm8Pvko0uefDqaIW0js0UFTzzbzFL/CwugrpYgBzh/L9I2CXDU5RM7Fdu
n5gb7FPfn4WK51uB5XQoL6WNwf+wl/oz+RzbvLMTi2Vtn1VSRHctIZT9aKv3Jf9C
ErA+kRMB2kFDO5Sp+7IRnat7YWyOb6ExOOHAohAl/LDf3W/rrtlNuJhUSRApwibg
QN6AKG2UlU2snDwUPoOOHDJP64maj+9cQqD69OM5uG68DRMEf6oPQWROzl+WgieX
cfhaCQy4H95dcbcoHKruTZ6cXmiPQ6xfFEAO69xJ9JFniGQvsbPGlEbbRZ0BCzLe
qoDy10KMSQG4LyrWQLsAB2pSZZKyvrD5e/K+TfWrn0v9UbodbB9PomW+9rFGRP7s
3QXPhFOBjE7172xbDj+gD2wdPcORvbRApMObFhKeqCbjQu6p3TUTy3RPfXFPpnx7
i0cSF6M0FQQeklTW34mzOOr0jwD3K6NPBVc6+UYc+akFLcyA+Z1ebjaGqc5spOqC
iS8KfcP/DKAEnVsKvae1wLa5AkZ0FmbsOGXHcHTlRr1Gs44zLkh3y1VnqVS7yFUm
m+8rSK1M/NSQWW6glynZdGkFRQPQsQHwIBRkmrS0FWq8HW/jKLhS+wRCUlOQp4ss
ZGL7HDy/GLuNDZ18D5ZDhCJKIjofMcmSLR/AGf6mOv9mVEBBRmkeD6q6VC/a20Nd
pIlppJoMg1mtDU/e4ZBv+GUm+zHVei+QN2GZPIAuskiK8R6OPKNNu6/hr3ETW1LU
S3fYfcjIy0kgxse8k9VCLUagpQIUpkEAMxDSfR2SRZV3A0FB8NuxA8+7XvvPD6+6
eTSfZoFpdqijyYX6pa5VoR2ppAbcoilH7PCEb56aOoDjRMzVPtTev2dUzHYYMh9/
sWXuqt758xfHC7ZuGi99dDY2PMAXzhTyEGRFiewWveRWfB1pU8VJlcNWhveefZow
Q26VAjDd3Z2r0P6lpfpFrmlzqAVBkbch6VKJ1rOQO0EqhyeKaOaK8ONGdEOs6m1y
xKhqXvsNiIEycxrD4nPxcQnaBTpIJSdRjpnYn5d7KDC7n9zcSFzohRlO2OiGKAbM
Cj8dUrsop5WKw/92awqPjpqRf0DWZiEvWhJyt5xDCZ7oBMB9yv7Bb5omTRMsiOFw
l+uIEoJ1sfx3Vl9t48GbbIYk2Bwi7wjsG0PfXT9HZoOM6uwXusoH97hPCBux+0Wo
o7d4pI6nWprixjEATJfZStDjPw9ITh0uc7FGac012K88FvSVv6nqFpe+os5IxyVK
nmxNOyBL/hTSO1KEhJ0paiwApmzxomwvwRq+SH2ehC73Q2qhTBebrqdrXEHXjcEv
ZrGWRmu/O1Us4YSSJh5q4k5gLFs4c1oloY5mumgVGItr4lWSgbS0mhslmFH0xQlO
7EHmydlEs98v10gccXOm0kzlkglfzllJXHuklnGzfKRuTWf3CKBfAI70W29eL2n6
NqfwLUkgWL/f9w2nC76tkkgJMIj51sgjMEfoFnv0b4MLOLZS7fUS31U3v/PD2D/M
G8ssu06O1qwKnv1E1i7KgT33s+9PN/hRGbqxblFvIquhF1U3FUdiA9ds//i4Z87f
7yHo/DM6EQY+bFKy+oZ0+bE3mOVNzhUfmr+9FoM2rzH4DxxjVIN3dKgv2h9CHq1I
yK4x86AWBwoC6WVa1+YBDUokoI5LAS6sM32iDIvcWZQe5lEuxcw2it+5KS8PEHm1
1lXVtVEcsjuOivyGP2NRj4MEVlMLc8ppmjtsO8vkFzveIRec/Y6vaFwgqDSmdZ3t
8VWgkf0reR+hdABwmkIW9hkwsv07QbnNrTz0KX+sBylMF6fcVPf6udeUW42dX2ro
XpRRyiIT6bIHnUWUMayJhXe0xoB60PAZ9cyA1ZWVwEmnmxg7uRBpVD5DCOof9PGm
H+TaMR+/EloRT+IPl2+MciwrhCTiP4u2HoNT0ahrz+UmCoehipK0/hlGV8WlHBse
gktSeKWdmlV3ob+LLFduYlK5NqLpMFYjJfvQWml3NZB8tBIXEt482MIDJXJtpQnl
zTs3aLypq2o3yOqT8N77e/CF1zeSfgTidFHWlfAWyLmUpV2RqcTYtWNBK5C6iyEm
jAtFqarP71whAt8CB0/dBSRs8OnIYvShSckTnBWkjKh6sa19jmgORh3u8Qlvzkxs
LgW6kj8SxfMK3a6nSgAQwAT4DN6+uwFEn9/d58urMS2+M/58zvD1aInLIqXZvoCz
l4D7C1vzfTh8Ua5g7w+esV3So88zD+0lDQLCBtwd7+7vcAXRoUExZ/8X6WQKcngA
a5tgkn/A3kZPTfOIsQWBU6QgI9nAtbJUb0rPUeP/VWn3eFPSKYYkJRTw1zU//WLY
yAJXO5mK9Zecm5vjRCNK7k+/wyVTN1BLUmf81aH7vD4807E17MiyaTgDnRw0YN51
aMS13i9JbWmkfrpI5vQQEg9OHCvqI2JRI5MRvDvw19DJzz+Xg+Yai8blmpPd6Qvn
qwnKtiWvbHLQcLwe0XlNwKVI/U6a408ki1lSiOQmkxKwHl+O4VMH/VGtaIPowBvY
FM4afPXDprhTevpM65GbyWoPTKehDPaye7cYLpekJyT0VA/lw8FyAiKjIiJ7J+b3
Tjz1wrF/JmT8/pJFmG9b4OaqqfTTxtYFo/GUzpnYvLAGJmSJsjubTMnGw3IioJvq
OZYfl8q3GBLYCpZRrfcsgVQh3lCtr871vFAJeL390bC/4Ptu7f3mJegsuVU6YwmE
MGIZuDKPAG49G9/sHCN8jYYpUoo18oID4oagmGGoxh/37vFYAVPxYJM76pwoDx71
CBw2SuFyCXTVz1r4hTQoDgBbYF+mF986QeBIqQk0iY3o5EKOzdAOY61TqKYtcDUd
H5UE2FcSKbMRLaVpBCHe7oCOFIiYo1zjq+sL9MyG3LDzvDuwbB0LTEqBVmTpOoFa
QZk+WMi3R6JNfMFvrSgWuHmpiYdw2YFwaTtepy05BuAw3Q4OFx017HnpbsjNVTxX
48hvY960Ag/pQnXD1PtmciIUdSD1WgLbuBfNnWLib6tXbM1auJYpX4sxwrzLV8PP
IgeWEaUEu/PCndBZc5vEaw==
--pragma protect end_data_block
--pragma protect digest_block
Ipz0tSaoqsds7/pcXTtOjgAQ3vs=
--pragma protect end_digest_block
--pragma protect end_protected
