��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���Z��?��1*w�k\�d��T6�c`@h��S3���u��څ�6+���p"��i�]Ω���-��s�i��>��m9�h�������Y�d�S|�B$EdB��Fm�a�6\�I�&��� �l��J� �|�SϳU�Y�r����1h�G��ɓ�mg{�����4kLK`k��{������8�B�dۥ�,�"��� �j�Tq��D0�ۿ�I��nK� -VcJ�FS�؍�[�|�T��f�V�-51�@2\Ϛ�5P�W��;*i�/3S�mÌ�	�!��$�/��j
����n���3��ص]j��@k܈�`�D� ���%�B`N�0G��޶�� ٌ̞� ���đ�w(��}�b��,LG��O*�!v�`w��˕GFP9�Ԓ�6��a���4�b��`�[ظ��~2��z�����*���}8��9��BwJW���q�������|�l�m<B�R6v������?�U��� ��T`��P��ɳL�S��� �pl����_��'�'�0�#�E���㨵�DLB�;}$u�F@d�ޏir�yW�x|J.�k�T@�B�Ə�jM���:�U�I�F/ۊd�5���Si���$9F��KU#z���zj�oT�Z����B#^�����SO�m���{����/\'�Rs9���9⃳�%��V�2�%�шݬ�Z{�Z�����{ۊ"xB,�nP�#��>����e&{���[�S������}����
�[����B��.z�������ܔ�7�p�݂$��*W�&��dd	6<Gz��,��JƁ#,�k�(.*�{�sbs�%���.\���?l�M�.�'!���Ts�����Mt~rA��U��%���xi7�80� �P�7���7^��p8�X�eSSG�EQ]Bd�Wؼ����9�}Ѯ�Au���'���N��f2\��g3�'���L�"[�,�UbiPBB�����+dq,a+B����E$���Y�I� �	�Y���kuUR�����(eV^���Tt�BA���A���DC$�qQ�rW�5�������C�M���<-�d<�[o|�3��]����H%��6s�3��[�ܞ�U|�oq�n�{�ǋ����:@<ؐ��T<Ϯ������.�r�SH�A���4����Z0��6^��A5��'=�fS��L��^�D��ͩ0��*�!�]�̻G�th�>�?%��4�/�ER�(���H��=��Rgl����L#�@t��@�jrї����jP�ޮ�4�[�+t�7<*���B�(�s�����T�Ln�f��8b��.�L,����3Ʌ*�B�=���������T/1�}�i?%�:|.���o�4�E�m���/X~�]sRWɗ�4D\s�S`�
q5����?65o��M�w�x��V�'�_�H��לּ��?�M��
;�&{J��ƚ�YX�-���:���3RÆ�`��D�$�$������G�u��a��ﶭF�Vj��O��}o��)J�n�x����';��OQ�܍��G�$�jL�!�j:h��F� ��/�Ĉgk�n�M�fj�6����e'犦�̟��C 
&���G�y	�U�!\��I�a�l�����鉆��Ʀ�ï��?G� ��='��6��a#��)�����+QB�C���
d���_�K�F��Lt�e�c���5�mk��>LY�VedI��.��� mFN(^�oJ��$|l ӵ�����I��i�JF�ʙ6/!2�HwT��f��N�X�6�>�g�ݽ�� ;M��H�Z�![�����$U��ȚV���.�|������`�\D,��1G>:�oh�]�~��*we�K)�<Ǎc&C��ZC�z%T��9������ݚ;ό[5s\�"̡���|Ǥ \#�n��͵����~�� �J>�9;%��Yc�=s8ҁ���Ma�W&}����uwt#��^�o�)⾾&���o��(��dB 6]��i$k�:s(Hk;,�-C��dzb�����"K�8�=#W��$�[�O\X�.}A��=��SO�u���n�|,�Q75���y4ͧ���12ev^�y�U�eҒY�H�s��I`zj}a�	��u�bo^�������2o;'�yQ�hlMFq����