��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���d�v����0�i�=\��A��?��� (��1_B�f�	�Ѻ+|n��y��Q4�]�aY�����*2�y%����>��������K������ �
�D��z�z��C�y�B����
_�U��hkF<�~x�ܕ�c�&@xAMhֈ���z�	D�ɴ�$����/{҄hx�3�C�[�a8y��x�y��#sA�+q�d��"��W�~`I��|�t`�Eu{1_�v�1�8p��c�}O[���	"N͖@�؅ʬ�̇l�:&хu�=gPQ��̠����8d�'�a6ʷ�ŝ~�͇-o�&8�}�`/b)Zmxf���n5V��3~��)��sv����㴎��C8��#k��Og�j?ʍ�O�f��}̷}.E���݈�M(��a(�q9��!ė�z9wc�Y����7J;y*��B��p��{�!�� �P͈��)��(7{�B*��IOV0:�K��`G�B̼�+Jw^2�TFԾ32-P8'#�"o�}���a'�)31�k���JxN�6Ck�g/H��o���c�����fe*A��7�8� ���ݨ� _�����%��=�=�C����I�{It�J���W��N�������.��%���׏rV����r#k�.,t����Zi��>�6]�1#Qq)z��v
�O�It�C|���\��!��_p���j�C<$�!".�D��{�C�����n���FMw�L/��Cj:�]c�:��L���y���}_b��R��Cm.����/�|��J�����)$UY��H�Eʂ�ԞO�����H��8�h����`Ox��7X,	�{��8^ɲ)���u��Ge�?�kY����8�G���>HO(H[��� 0��\rŞ�*����֔s�Ùe����5�
	2�,�y1��6��q�>iڱ
��,�$�dp4�����n� 9��kC}T���q5$C|��-j�_�OHHK�� �h"z)��儮 ����)��˛%��N��:�N 0�����5'�����k��.'�����;3zI���v�"��O�yȀ���ކ� �A?#�n����0��46��]��DO� Yh����<b��{��d>�G�@(�=�D�X�����Z@��.��@��e��R�b��Y(��<��T��Io(���q�p��I����<Z�T��9�ς��'�[�Ba�Ag~R���3H�|�7�_'dy+#,K\��4�m��tHn������t��Q�<��KZ7��8F��	�xd�A����4�@﹏������>������
v0��c�6w�����=����w�`�)�<)�Y8a���M�|�9�5����L~�T��-}���LY�>������,B���ā/֜ t���g�	������ZP�9B�1Dg��'v���b$�U�s�G����c��w�(u���T�r��͵��*{�����g�>ɏօ`����)����\��W��\�L���n�y{�L�7A�7�{�x~�<�ာ�X)�X4wC�`^`��ex1�@�mE��GרÅ�NFTYkl�b!�A��M#�U#m�peNoEb������;~%6�m�0I��7�Bp5n�G��Whs+�>Y*m�qu�o�sN�{kǷI��ѻ*����j>��j�H��|�g���A�[J�L ,���.��v��ֵ��
,l��Εªq��ϟ1�/e��f%�R�,-����.o+t�eE�^Ĩ�KhA1-�lݻv5�v��QD<���@����n��I�>�����W�C���6���XPl����Q1ɖF͍��*������&��/
8��p���{�W7����7e�ԑ 0���n��T�ݍٺrd�I����L��#ӻc��Uy@[L����QVXV2#˨��T���r���� ��8E�k?�ќ���;�������X�B�<�򔿧����|P�ҍ���d�:8�V�Ed�Q̲~m�$����>�D����ӟ]8�����hK�FMώ§��$�.�A��\����Q[��^�[�y��C�v��'����%�������>�~s���ZD6�똰�t���ix���z`��Q��FM�a�H,�g\����A�����z�B���K7w�I�Q�Et�WV����1l4�G�F\����֞_���q��EIu��҇��J%��M�m1�d!LM�N'�/�l_�RY1%AO����4C�k�)d;[s6šm���u� �a��Ǽl�[^ʀcV������{�)č�wL��!�#@��(o��֐�9��zu���ە��L��t������J��\dSh��~7��N�4�#���������`� �
�e���{ǯ�=��(�v_��F��k9<U��٭=�A�F��$nW�%�
N���*�M�����/}�Lp�J�y⑱�\����1«��=��RlՂ^��z���X!�"�Z���Y�9���_v�XW�ѭSFP��ۀ[�ɿўb��rƌ��;	,*Z QX�X$���O�k��]��p5ڼ�*}�	(�+�����6�@i�-�p=����Fr�V^O��+�O	mUATo�� "�K����s7�hHl葢�\J(e�w�L�n���#���i�˯^���İ?�c=�}�1�7�"�	�_���Wb�E��#<�OVlmJ�Q�ƀl�O��T%8Ǩ!�r�/N��qc�bq�2���5W~(��4U���]�y-`��'0��ۓ��l�B�5gz��<��o=�m��aw>qf�������Np��'� lB�@��Z�T-E�N�<		&�5�.A���:d<24�#\�vܠ�?�0%ldВ1�)��"���6���'~����+b��!m9��^6j�g�|cI5��\��$��S�.�&�k�g��I��
�ſ݃��AGx����� ^H]lh���� �*����J��C���R����Q8I�]w�T7�Xs��n�d=����\yں��L���A�BXY��Uo����Ȇ�����5 �}Q���N'���1qhF_t�X�ɛ}�9��(�	�o�wI�`3�	د�T�V`��=K�}t-��ؗ�:��Z���QЙ$:k)Bu�K�N�5�����	������ k �	�t�=�8�O\*CR,oB��u0�K�Ø��@2�os���]1y0/=ԣ���>y�t��?K��:!�aǯ�ȳ�(�����Zk�C��0u�5��_�|����P�_v��޹W&@�dA�`Z��%���'àq��ѷ�K��	�o~��Џ��۫|���J������Z4��7��խ��J�Ͻ�{`kB�S3�O�[�e�t��R�>7���iv���+��T��<>��?0���QZ��i�S#l�F��6H�jKX��jeT���UOC/�ܖm��EI��W����d#���7 ��'��QDy��,�]��1�u1*�Pak��zsN���w >,Tׁ4E��{y�A:�8�r�΋�LBn�Q����'�٧;�2������~E4)�.V��,���;��~>��ê�7����n�X3�K�cŖH�8�����o�9���&%����l�T|��V��p>3Y�?P�A��Id2���D���o3-�O� �L���u`PR���mv��ȟq�0�ძm���K�QR7,����g�>�$l?�<~8�9�vL'� �zgΛw��3h*?dB�qbD��A�7��3 �\�i���J�$��.Hn:��Yt�����86!V�c?{8�g�5�V$K:.#�G��,����ؿ0�:�"p��Z���>{�J��h�N�g���N������z�� ��		��%��o^i�rx7�Tΐ��rt;ץ\���h��}��=(�PE���s*� �u!������vz�ߜJ�����l�x��q��7Hkx��6�s�V��>�1�Ѥ��`�%MO;^�?�"}A�����mRRT��$�3�:IZ�7j�R�s�E��H7 B���2�sB�|`��Tа׌E�5릺y�]���ʒ��)��v������x�r�2�G���y����ω������� r����������|�D�Q��jkC��#�O�I^�j�W�m�f�<���Q���f�����E�xFfuZ����#���6F��|F��8��"P��,�nq;';l�?���G!�ţn.���}��r���'ak��֙ ��'�"��]�� �s,/� z��u��`�":���R�42�۠����pl����O�1�D����μ�J�bz/� RG�}ga�����a���\�o ?�"X��I�<O4$�Z�g?y�)��*Wg>;h86b�땼��IӋ�̴���;�%̫t�䡈]u'���Qp@�I�� 
�����{�5�OT}��e�>����G�/d���XCޣ��RXx�S�хŖ�o<�\��j@X�&�;y��M��uiK�F��y¾|�N��2^ۂ���ݚ�0�ç���  '<\j�^=q����,�g�O*-�n�u��6�������o��������w�߻4������vz�ÔVN�w�tA!m7C���7{����^=D��h����o>���;�ں��"q�:f�����XN�_E�����tˬuُ�殞�S��w�����;�-�p�	���H�$��<�������tJdP.a-]�V���$wب?λ�&�	�*�m`:�?�y7e�|zvr����c��Q���a:6�LH����ݐw'cST��Mᶙ����~���Pm�ȹe�l~���x�%�G�K�#��bJ,����8��e��FqQ�-��*6ƒZC��B�.��/�r=r5�SF�y��_�Ҩ���wɆ[)���*WO����"���=����0P��U��~x*eC'�_%�͖GA�}�S@�����Hީ6���-��ND/�^��F�Fe̦ך�
>G^��J�х@�׭�k��m]�kf*�I�h&L��Ȱa�6ݘSŃ��H�h)�`���}7�}\X\���A\�FT�o�>%�jKV+v��o9��e����T[=ҿ����fbS�
����:�W�[���F�%�6���/�W/����� �(��m��HUo�� �]8>jPX���I�ͦ��:����%�b�[��n�a�CE�.��Gt�����T�/��kX:����(�����V�I<� �+��4���G�@�� 	-{��h~�����d��
c�?�y(���n([�%Y��
�Y���:�S�!�Ȁ������� �)��0�Sk\���h�ID30��RD��<��"E�#0��Ě,~8Q7��vLo܋��m�K��{Jv�ge�(M���R�w*�T�D��Q�_&�8��bO2}��֌%��H�d_
0R�6���r�`:���'uZÀSpъ>�R`����;�X���i\��~1n��ǟR���&)`g�ˀ]���{POb\��mO"��6� ��(���y`��
���@��@���*���ЫO���2)�I�XGb�=���mcofbwc�Ⱞ^�ø0Z!�%:�E�}`.�®`8�WL��?�K���W�K7�k��^J�`�z}yO�t���WP:V ��%�h́��+-_�Q�+�*I���L�ӈ4�G��Yl�?�z-M���0Q̏�$&��yc�� 7�ՐǺ1�#d��޲�1��P�EO�G[-�`ѽD\i���D$�������nҊ�Y"�����U5�UA�:~=v^ �ޏ�є�a��"�����ޥ�/2��#a�j�.�[)�����&	�7��HV�KN+41
�=I�R�b~��1�>o6��^���l��}h��b1��S3?[x�<Vq���V�:�N���o��WQ1Zc��[3�$C/�V�=m#oM)�����G{��0��r�3�R��{�C.�y�B@n��
^a0[n��z�L}ۛ��G�Yyؔ�*�K!���o/q�n�4x�rn��S�����%��4LD�_��ӻos5���T}=����F
�I�%O:|1!h&�̄rG��%���z�� �8�����n��W_�%:���oB��	�v#�\Ж�a���&Cp�Y>J<�pR�z.RY���(�]PzY�!�_D�'j�(���4b
�~ʙk�@`۩�X�裸�y�i<f����~ʹ�C=�-��YΛm���-�{o����^]�  NHŇ
킓�j��1cD3(dw���`�³� �4�Hd><a[Z[|FG��b��K�_&�0��B�W���@<������(>Q�et��,f��P�p[�!{ gy��},��]��Ô�t@!�ȗ����|�q�%�%t�խ8�E�QY7IV��^��Ts
�k��K�(^�?��P�P�ӱ�B��A&1����W�fe=О^�h��H}'ш�aw�7���b���U�<(OZWe��z�P�8�QB��F��s0�����@���!O�nШ�zJ�dwg3������Os�n�s��〜��$L��$�\��H2ȆL��g����Gy����.��mU�����Ŝ�Za�[͚wzm�kA�RG�����3-�'�E~�
Myi�r��a6y��������(�$4p��?�*{S��|>F��<�Hp�Q��1����3�*9���v�����zc�\W����Ck70��f�{�\X��Ƨ̝�7��+/(	,���+��~͢{VYk!5�A����Y��yjj��T�ibr�%�c`�������@b*�έ�7��ڭ���I�'៻/c��_���D�#�D�������V������BK	��T����3�>��(�=����q>;i�b�NR�ݫU
_%	F��C_W�F�vI�� �r��W�sɛ���?(��MP�����n�q>�y�(����[T[���@�R�ջ���r���[%Y#��M�H��,�G��	
�݂Z�V���%��[j�7�I�#������@Fe���l=C�1r(�ss_� �U�e[���D�y����
�n2_%]f��c�~M�+��C��ʠU��QN��_��ׅ��G���p�K�o�&�|����E�x8e�x������_�O`��M闗���' �Ԭ����NL�Oa�O��l�R���\?�2�11�n����  T��'�K�ѱ���x>�O/qW��������P������ �	C��G|rq�4����|x	!��e���;!�)�]�'%<* 5��;ΨJĿ^��*�:�Q��	ɑ��·�[�`:Z��G��*LI��W�h(b�N�k$NC�R�5dX8� �۸���.����:T5'^/����@��+Ǎh,VD���heέ�-{^C�3�o�i���BK����s�?�We��Ŷ?;v7�(8���p�P�pXyNT"4�W����r���!���>�hY�QRa��޵�a6�By�� �$z%;�����w�?�߆�쏴Y��O0%�m뺡A�,\�U(jݩc��m�����	�Gc����� W��_#pw�t#TY���TZr��0�%$6,����úʋSC��-�D�eE�w+%(��V����q�J����xN�X�����ZK�� ����aj�P˳Of�V�[<*F�I?N���v_p&���xO�?I�`Ƒ�3�B^e]ʻ�@0�-�l��Ae�v�D�d5*{�KJO^ ����y��WM<��ԏ� �;񌵸�a�	�L���6�p����g�\G萵O����=�ۜ�&ч��]���j��𫀌떿1:����ϱ+\�Ӓ�^u�"J���+�T0�5�РsW���h�B	 Y�ӈJ���҉@^b,�W�]�.�:--��� ��˩Ox�ֆ���`����ҕ��N����	e��V���	9ס"n�L}/<V��ζ�?4�+:?��dm�����-��ض��5����Dy�^��]`��A����*��ڼ��.��A�T_{P�p6�+�ém��nD�n���������@a�y����vK$O��j$��V,)��҅�:�<-A��	�39ڥ�?A'n��/�2��׶@�=�TB�g�N��1Q�A!�?Ԩ�3�3b�cJ��]�~��/�e_��{���k����H$�yq��aC�̿����W:��9��w�<A��%��u�֡b���r� F9%�j��H��D:�z���3d��y��pFâϰ	���B�~�,P����n�V�7��U��u?2��fyc.�k{�fx�Ud�%?���L�N�d�<���o���i�x��T���K��}_�(G����A-�c�`�b�Jҏf��+���c�O�Ѫ{���ɻ瓵��U�8%��1��O���ߨ�)��i�ll��]��E_��v�׸lP��+�胐Xe}u�G��,ݵ<�8��?G�Yln��ص(�$�s)L�W���yq��Q��
��c?ʵ$l���4�P��ܦ�U1����0(yx9=�'��2�L��Z�ԫ��s�3�q��Emy��b
�֌PiC��[���b���B��9]۫�P.���]�L��a��s�i'�1kT�d�52�oj����6��3Ͷ��i��:N�1=���Q�{&��v#<=�h�.Q����}Ҙo�l�ЊF>�ga��$;��q�G+��^�	���a�-$.af���
Yyh
�#��~��Ci�'k�WK���+�)ug�}�h�PNS$�>-ͳw�{�1���d~�U��| ��xy�ʜ�Ji�h��ߥ�ʾ�X�yG����AMc�j�D��p�V�����e��,0�O���i(���x��{�Sղω M�c�^^M:�?���4���Pl
��[�OV����d�}��b�f��_`$bZ9s6�^��U [�G�J�T�>�ڼ���r�DgĒ��_��49�Ly��W'�� Q>�~M�/V	]?'��P����)i��"}Ϗ1� 8ɑ���iz�M��[Ӊ�m��5�-\]@���x
�/��K茰�n�� \���p�����G�S�hЁ'�	�,�f-YLUܟ��������E��%G�PM�A(��ߢ�J��Gߓ��Y�;�yr���$�|��� �u�T�ן��ć�a�	�F����h+^��� ����YA��E��(�W�ES~CVS�	�c"�,�|$nrf�:̻Q��,�1����Y�9�_���	��������:�c�-k�xƠ�e�=#K^��������ȃ�(�(V1n,�������@�A�}	��,_"�k��	���?���c��:��]�Ʊ�}m�>
����K�9�~�s�_+G:Ù&}J�Ėf�S�q>s����oy�p���A��Ri��Ͼ�	�ћ8x�ʏ�Q3Ί�2��j����o[v��9����ج}F��s��]�~'J��恐�{ 2"%�*�T��Bb�W�h�6��ʌ��7p�����2��Mh�L���b �\�%8n�|���3�b��.���H��O����JA�mh�DI�#�"�E;���K1 Z0�W���x+&�wytHe��5q�(JkT؟?�!����|:g�����}���JY��
�;6S$��D�(��}�2,(���N�s��Doi�h��4lQfݹ�������;U	��V�t����y3����acO�e����(�-w���=�E ��~ܲNZ[g�v�}ah-�ڊ�;��7�@�҈�����q�X+�i����"r��=�gI�-c���B�����ݙ~�zO�G���RBS3�R��}�)��Q� ��`=ۻYy��$��r�%�"mO|9i-/��-�^����Q�d{��S�cJ�ͅ2�!�D�aR�/�G�3StϷ���NF�y����vϱa��Ȧ��'7�����-����~���i�L��%Е��Wj�IP��ғt��s�� �o�vm�@��E�x7)��P�S��0Y�߻�;��a������¿����U4$��O�����D�b�����L�ªnŊ�sl�\B)���0��U�<��K������Ĥ��K�pьYE�%�GWc~.U
E���A��<��!Y�j�{7���@�4p;���k�}�(˚�`���.�y=J���4׋�\�2�'=i�A��{0�׹�j���h$�b��L��_��F�T��xRFb�Q�}v[�g4�bV�!��PZ�8zva�*�h -wQ4ʺ@|�]0Bp1GէU�F���ǆ�Cu_�]=�ve����6(�Z$�0|b=-�����{NyJ���z	����,�ll�?�V�����]`�9w�ҽ�_?��Ў7j�g.8/}�~�����M7ʻ��Ѣdb��m�.E���E���\q�Ihsq�iM?np�)87���T��7��qd�OP����J�燛d�`��(��0��1�V[0>�֒mH��f#-i��ގ�!|-����K<Х��1f��q�	[�1>�٬ٽ+ᷜ3n3�!&�p��_�s\t=n�r�0�Z`�4�N�=��J-ʄ��I���6]h���K�T
��O�kt��&,���ts��W�D~�F �#�w�c�J�nd$0lS�`0�斑��swBx[�U�������n!
笪�gV^�"�������H�����&�������W]������;��e]$�%�9҈t'�c��+�E梔#�M!�<�CRB�㞥���	z�V�!w�0]1��!!�#���F�[@��`��륦u�,�f_o����V�*�{g�&���˥Z�n��S�hj����p�j_���Dқ��z^/j��D*@հ��:�t׈���p����}�d�ׇ�kAzL^�r�)[����yl<���q�t��b��
����j?�F�`!%^���B�l1�rd��N�@����z���W�ӳl�h|���[X�?�a�x���F�b��Yn���8b��u+��s
� �y`s:cI���:
�C�2��j�Ŏ#"��_v'%y�nR#1�?��
�m� �t.��R�#��+�#>��(l��;�=�M3���h��f��#5̦����ˤ��._��	 X��C��/tJ$A?�K�H<b�hކ&�:�k���/�CU����8�����hF���[�rx+|%"��_S�cpǗd�jC�q��v�˅�T9��O��rEpL�R��:sdY�����,��1�+�	�KD�ǔ�Թ�e� zN{�2R*|sj<8�{(*����t�&~;��Y.L���/}5P����:��>X�r��.�|	N������J����g���!�Hv2�l��;qwb'�hn��)Ν�&KY�����L,`��\�#���-To�~{��°׷w��0_)���_��+]'b�UD\`D���ʱ�C���eu;ms�!����L��X��؇��[(Abc9��.m�Y5��exX�ڥ�L*����'��3)(xЫ�����2���Ҟa�{mYj8�7��:����X(s�O��#R�6`��۾R^��|�l�WAUg�����mZthQ�z���E����*S��������G��13�ZG�쏍tX�J0b���^�%u�-�A�(��ǽm �{9�������p�`K�W������v�)e=���m��	+���fbdWlm���㦐Q
m��=�Fy�cX����ߋrx���V��������RZ&ӜߍK�F)񉣣V���P�ve��^������v����P�	}^/��v��zJ͹�)Y����5a�.�M��e�.U��u����}Y��8��}T�iv��-"�eA�/��Qyr�z઀Un�N�m\3\>���a~ "�SP��B)�(�]�چk��hUsi��X�ló]��4���A����ʴ�oŝ���\s[��"�:��I͚�E4v�j6�+�����:�����]6���\�6U�?�Y�#�aBف@؁(KfpP3���$Q��H�Sh�Zd�܂�T��c4�2�`P�r{��v�aZ�����Q�Ȇm��<Lw{�h���԰�Z{�[
��XRǬ���C���p�2$J  ��̦Y.w�?�����	��-, ;�'�NP��̟,/����v�0z�+��3���a�\
�l�ۡ����<�ǆ����<�8��0Pl7h�.��A=W��k��j���)�PJ���G�����V%��mfBB�H'Zf�LnkW�$~�Efɕ�%NB�G=S��8.�t���(W�R�{5ڄf�kPw�O�(��(�B�:���'�Hy-�k��Ƶ�T��^��-�~�b���,���F�=օZ�S�&v�諘U�Yk'���n��"�Ij~K4��i���v�5��}��$�m� �zC$�c_���Uv����|��"E�Zf�9�w�'�J�	��w��T�3���x�N^���!��iE���VS[!����J����9�i�@ �g��Q��^W�6�z�i����vd'���EMJN2�CՇ�Gɵ������n%�訅� }f���EJ�� �9�)0������D�v�'-��i-nGXǫ�=HFW���RCb�^\]�x��}��	�2�?�Լqs��[�(�L��Κ`v��B!�J�v�����Ҩ~�d�\L���$<���ҹp̻��`���bC���!�"˄�ch�$�I̊dC�j�ƻř�� �7x1�][iܔ %�ؑ�y���xѻ7�Z������ۙ#��ƴ-}�����ĆZ��C�9����*ز���\Y���� F�ӎPW��3�����n��.y�=LA�B�������r����9�S�\���5K��t0!�fpԩ�]w�l[n�cѴ�� O�F�Oe�f6��x���{�߂f�K��z5#�r�?�fb�y��
wj)��=Y2:��Yt,�Z]�f�?R�&6�`���|`����3��ئ֣�������*��f��f������N W�o���Kɛ���ͣ�:�$@���fƞo�%�I4߁D��j>Ԭ؟�c�SxH������-����&0����y:����/���R�xU!'��Q�rT©�yt�����ާ�YiV�6���Q�H�t�@��,c����/r�	;t�KN���mJ4O���b�0h�{q��)�TCg9��2����+���#�)!e�^�A�+}�H�!ѧ�I����6� ����R�7i/����8Ȓ�{	�.Q2f�[�ܚ�&U׼;�},Q�=K��T����f�mcoX��Oz�It��"W&MJ��`�m���������L���D���m����}���*&��t��a��lX=�4ias�?k��!��-����C�t_�~�0�#�$x�7���S1��	W���Μ-�-�CRT{�1�48y<������G�����x��y)F�i�O�X5�� 	6���	�ƥ�B�}o�S��Wk��S�r����W	�p-n�X�6/�˫���[�E!x�]��|f2V�d����w�}ap��H1Fl��0��F�PNd����9��_j���ğ�\���Eߩ�ol(�"�6�U���9�4�{�ү�RG�P��$a)�eQL:?�@m�J�c���6�͇�U�&:�9S�?��֓H$7�[¬M(������K�{�wM���1����/�
��ǃ�\~���$��}�؂���
�ܻ���J���t\8̄���(ֲ�v��8�ЊX��|�`�`�pfH�3w�lz��hO7
}e�e�A���q�>�4��۷�C�؅CW�2@aq�]���O2�����.�B�e˟_����[���t��h��	��@O���<��""b/p�U�|�����F�ݸ���}��^DW�\���x]{�{]i�DQ/��ۥ��`?����^��)���QUe=�'�'�l���T��������Rѫ��k[	��D��yho��Y6%r�8��%N!��8Æ�N��O��L���">���8��������=Y?�����EKҊ Ȉ͍���Z-�!�[�z��l.n+��l����-d���yR��� qR��bU"eC\�	e��	'����Ν[��eaY��a�����i��x(�IN�#�+���d�:����kůQ�k����(z�{@�V�<K/N���ήnv�B>y�
�n�ޝKאFE�I�������wo���Oh���������M�:�&��,�7ue�p*����#u�d�(��d�!��Ki����Z��|)�V���]�< ���gmR�J���_:��g�V�Eu����� ���zmH<�#��!�aq54�n��!-�:��ꧾ���G�3���(M?���H�U�c�@�E"���/��{��-s���L�𻫇�/�B�s�ט~��~E�I]_~R�;�y=f�Xߖ���@}kĎ�a���ٝ�v�ø��
��e�~a#�Ҟ��+����N+�U�aP��ꠘ���x2��n��I�|o�ˋ>�DN��C"ZB�V�/$k{���@���C#�K�x[A��k�Y��ϫ�4��)���g)(J��~����_�$PL��(�1O���J:� ��u�f�_��3��K^M��� ��̿ WU߃���f��
9������ ���cr�2��H�B��|��,���)�]�m]�����g������%b���\6آ�^�ڪ�X������ª��pO�-;��aU)z�9������p1����b$I7�?^4���Np)dX��qg�qzYrQ����w��{��*�~r���͗㸀��;����L�!I$�I.%���߼�y�יx'� �gI@1B�c�'RB�&�.�t�Oi�Ѫ���mn!��ăǨsj�p���{�� |�=ׇ섣E��g�e���*�s�#�`�#�Єf��g��tV�׆i����!7�a�=^����ȝr/�Q� ��y����B�� =:�{Z;$�(����3�)����ƅ�.���QW�#�0:Xw\� jݪ˃��y�16j{q*-"[�P����(��g�:᤹K��sm ����}i����q��`���@1{Qz;Vv���:ʷ�A�)�^c��Y}�澨�������B���dE����1O�MQu��u����E�] M/��������-�O��Z~�c�,�e�DX�K���ŧ���� ��д�Le�-ļ�B_�����$Sr�K�����mm~f�r=j�QI_��@��_�t@`��f�������x)�[�=�G�⯽?��	,%��P�q���b`_i��nr�^�����M�4b��7�.+N�����c* 
�1�Ư��ʼ�\��k����`�nh_��t�5�qoD��p�扔Y	.��,E���˓Jy���r����3�@�^��,j�V�"�2���eh��[!�H�w+�2�)gyAx�z_�8��)usfU'��|۶����Sg�^���T�)�bN�/i�>\���+,ƨ.YTl� �Gp����.�hq�כnl���*X���T��v��iF�q�z�+�C���J����(�ǻ�o<���ҁ+u����z`�DN�^�MV��P�����
A��i�>M��1�u2��n�8�c@<͢j�%��L��($o�P�8S���k�	JZ^K����&Ӷ��d<�-分{7J����8R��A}�PϬ =�����ҥq;=D��	�� �9#ةlH� ���RsW�u�$��x~��z�Y@G(H���'�V�X�Փ����˫�v)�[p�l�}zh�݆a��沕N��XM�xԅ��H��$f�yҺ5,t��(��uᲰ�X����|H��#z*>�z����]
񷳡�Bf��&,��f[%�G�sT4R���*
t�(��3��4��t��$���t2�btJ�u+�B�Y��J���q���F�Z���6g<�1`CZ���L$PjN	���uk\.2L��=�Sw��niZ}��<�����8�� 4��,vr_���lʤ�-d�>lDtVճ�������NY�姺�|���@�� /gw��}���J������}�66*�jL�+�����0��(��8ʿu+�R<Z�;j�2����koi8׀�>�"�L�+}V��'n�?�d�Qͪ.�����F�jDFI�� �����$;�z��_W�i���n��]�V�t�&�˭�9:e���S��̅{R�������4�"z�2_b#���@E��5������30���u���X�i�� ��c�?��0wٻh��o63�sB�\��M>�Yv�	ŋ�P�p�C�KY���	`��-��r��xw��ס��XL�ʭ;;m~�lЦz�L�Ι���_��y��Z�-f�u_| 1끞"����<$)�Q�c�<|E�IR�s6H��q[_N2��vԼ�o��w��f���C ~*o��'�ψ��j�8�\9G���RU�N�*<݅u�J��ވ
x÷H'�8������I"٨�*ˀ[˄�-��<�f+�,�FN� (���?��En�q���=+�(d��;7
�R�<J�PJ�59�y��7�$�n�V�~?�aU���
#ֳl��=E�c��	>����y'�vG�7 ����ip�n߻���D���	��~�W�*L�v��F<O�A�Z9�ۿ��\t��A�g�#�u�GW�2�3�ˊ�~]-4MI0���m�ҟ����T[�\���jХ�n�o�FN�o�VB��\�4��A��ي�<�n�P�c�g�8 �ϻ��z��si�ԛd�=��Ofl|O�U�
ʋ?��Aw�pֈhކ
e�&�����z�#�=5R=�_�����BN7=z_T�Nb7��7i���zIw<��UKfAO�N�a�l���"*��*'sv4�f�m*�s����ܣ�TuHڋ3]�*q"�rs�u�p�7�IG�tp��$�?K�q�s2���G��;��,�H�DY�{�6���H�n�{�Fw�h�j����p��0-��rM��Q� �4	��\npҽ <�Oj&�8t'�
G�Eim/�y�:%A�⦡m��WY�rt<Nko0?�%jDL��H�u��B��r��lV�d�wީ�Ad��U����
���oُ���,����n�%߾��@k��
���s�6��d��T���k��J��+�c�Ջ��~A	����b�����`\�%Y�PQ�v�w�!�����H�D�!9��\�y�.���)��$�R��d������aCNS4�-`��	RM19�Ȯ#ʖ�I��V�GY* ��~�g�އ۫���%�{)bLDy�
f���-.���꣙P�a�^�b�~���T�L��;Lks��D�����7? �0���}M���^�{jw����I��C�$g�
]�_s1kw����������V����L%eU�JP�e��2b�K���`� ]uU�kܿ�9F�5�_>���46V�9ȳٳ��hm�a�T�>��+�@�e�
�6ˋ+�zs��#��:<'��o���Cܿm���Y�b��W�f�<����Zd`x$Ǳpo���E�艒�U�$cfU*r��{՟�䯄��YRy@������ynC�t��'q�W��4:�O+C��s�N2��XV�_81K��byx-UI�I{3�0��c��!�j�$M �ip���di�]m�	?&���0S|�ĔUO�ѭR�#���!+pNu�~l-�����g��|Jua���s���&��!���>o�Qf(\ �ڨe���Ôz<	�Ti��)/:o����'�'\H�.O������ù<%���4PX�z.Xhc�3��O������N���N�"�j��]�b	t����0���������{����r�Y�莾�]2��r�����y7ȼG��Z?n��k�6��6���������Oa��Rg NM8���G�r�V̍0'��nq��v�P��v:�c�º�X&q�QW0$�����(7�ɍՠ�(|:W+��㼯�T6��.3q�A~&�Rd,�﯑��g�+,+�D�U����緊ߨZ0�V�'��I�ʰ��*_}��w-���`�o�CJ��Xeu)J���`��Cr�'FxR?����k@�u�S�Cu��쭫g�ظy6���͎bW	�)��xg�h]4�h��9R�Le;a�\/MD����pQ�����'&P/����{=�"�n�zm�b��Y�pns����A�P�!�s$�1-��"�mJ��ٳ���FFg	�@�!��]Q/B�X�����cX<A������v�?s6f_H:� 6�g��H���>�F:@u��.A@�#�FZ��&/i_���kh���F�s6y�?s`}x��n�J9:�a��JL �3�iP�d7&C���u����	��8��	[�'r��& E7�ْD樄+�j+���9I�z�=��"�d�rNR��Yyێ�j�Z);����XԘ��va�A�Q�t^����ӫ���ғ2��2�(�M�
����qo����i#�s�]-�I��l#�_bT&��gXmB(~��+qS���X�^6TV�b���S�R��l��"�Do��w}�,�����������-�HڅE�~��7�1�É��9亄[��d*B�Tk��A�I��2_�����Ǽ&�D{|ɜ��Y�=|!FOҍ��}�͙%�U���zV��X;J��t�Mw-�?��.6�X!U�ME~0g6�3�"I��C9H���a�kL:i
�ׁڙ�+�/Q2��l��[\�Y��̨$�6y�F�w��w\+҄�U���*��<����v��X�6Z�ů���� �`�Y?\�cwTukz�P�e��C�/&�
�J����|O�D���Nw1��HBȽꇤy�9�q�j%Fze��{4��g����5o��s/]������OZ��Jk˗_�hٟ�m_�����K�M�/ʩ?%5mR���RI`d,T�F��!e쮲%4�H�Q�	n����^l�	��}i�VzX���˪�b��a{\Е+m�5/>$�������)��|am��bM��U�X�����P����\ ������Iw���;HM��\�Ll��d��Ţ �ߡ��u��J;�d4ģX���{���Y=Y���X|��;�l��A��c"[|�]�Da4�Wx�'B��Nr]��*��W����������_�tϭ+9�P9y����R+j�/P97���+rS*� g���j,����j�0	LԒ��F2�6M�٠Z1i�[t��x�Α��?���^��Gx���"B���"nI Y� �θ���_9l9�.'X��DS��"�4�޿�ڍ� ���4=�fSd����僮�>�>rmӮ��6`�S��0�{g�\��f�ָ�����G1@�״(7L\�hĝr�T���k�4Kh�]���tt�R�O�I���f!ÇNhyg}��e�gӻ.��gv��ah@�v�lA��z����P��.Iw�%G�#��[�dKl!�����!'"#M�k%gŞ��D}R훕�I�5��7��|�<DȖ��p+�hy����7W�-Dx�R�G����a&��GϏ���#`M�c/�=P�/�^���Q�o{P9V;ꄕ����2h7v��`��<�D��؂�6%��#���-�W�<fYK�_��y&���1) c<8��c7qh ��������&���:�C�z%x�:��֜�h�^
��Ok��x��#\���ҷ����#k+��s5#����+F] ���V�B玌=�*�#� ��&�P�)g�f���$u������ڟ����Ը����Tr�����>�eW�F�B�q�;�/G�3��VED����f%��ԍ��E������w-�˼���^E<�]=҉N�а��&��<g��8�k7�%�Q�R-GiE?������;����mG�#Ws���~�3���c��E�����l��{��Rf�S��`�f@�aG����Q �r ��I�dFAq��2�WAn5���-�'�����s��x��U����	y	����X�}L���Jv{8R�����]|2��C�4�����.2��8sҙ�g��./4���:ˢS���7�}�>5n�w���A���C7G@����H�c�	"	�����~ßEgv�������|�t�[}�(V�����?/c	�M�m�C����gE����yΖ���Lx;�\����;*��3�������r���Hqq�i�G��e�k����\RJt�&"�=������(2��x��{z(U0|
ha����;w�n�Q�A���`��̒P&asַ�����u�� Ug*�\��)*�僡O���$���U��Hs��؆-L��
�ĽY��n����yI\}�F���I�~����9���U��5��"����&����9db�z|�0�K<t��*���ߡ�����<�1m�LȺo)�u��)x��v�����R�.��T_�j`�"��?�*�]I�]x��69;���w�����iS������E^(-m����a]�,M�P�p��Y��Z����ml�̞�Ȱ>y��dc2��-Sþ��c{�Kx2+|A�-`���Q��;�cM�2��(E�EB��|�m���ֆ�N��R���:xK�4���T�T��
h"���?ˁ>4��e���(Lk�?G`(� �/ͦ���Л4ʧeI5ŖQ�ODAX;�?p��3'/
�F8�4qi�j�5��W�,p�QF��C$"�������/G��塞ui���h��������Θ��֪+r���:�K�$rA��\��J�mu��i��h���^`b�k����m�p��U<���M���f�7aj ��]��o��1= :)3{��� ���gwȡ�Y@C�7�;�����f�W ����0*�+��;�@�;s�A��w�-����Պ���;ܐ�R'Ej��H����fG}�ƈa���-5s9���MC���M3�"�E{
};�bN(Xc.�j�bM�ǬO�&�s4��͔���=;p�0�U�n�y�Kȋž�{�0'�h>PP֮V�
-<� 7� 2O�$�,�p�}ט���$�B����V]���	5rW#�z�yf~(nǔ�o�O�j$�Af
����i�<G�=49s��+�"�Tp�9��K�Ug#A{�EtF&�՗���-�����}��]NQp��)~�
4��\�6^_[B��ŕ�z!&nc�^��oA���f�J�#ٹyK2O��PK������bk���l N����(I�[ݮ��@r�QO����T���w}P��4{ �<�l���_�y�?�߷�R��]���E���G7_!+Z.9�$t4�f��h2�=���+��b��ùO������	��t�*T8}�\Pф�l���g$���Q���q�_,�W��&s�X,�G�ٗ��Y۝����۾Q)G�/�VB8�h�~Y�Z��-j�:=F�Yi��P.���#� IBc��c�v���O 