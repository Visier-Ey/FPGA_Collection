��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���J�l����9C���%[@ ���vK�G%H5��ۙB3aԯ�g�!�
�:��JN�>k� t3�[r|������D�����P����gbY:���Ռ�N߷+��͒�P�v�_�?�e~`�\R	@���@i�Ց_�a,S��f�z0��.�� �-\"q�I*I�R����yjڰ��v�`9�����,B��tg�Xb�?ưn�픇��y�ߠ�7�S�ޞ��#yF�v-5e91�&�7�u%\�=oB�\`��F��4��0NM;<����r�˃���GH+�}��+��z��q��2��Eg�� �����)j�FXs����!u��o�0(T�ri�����H����0��kF���:���/U�D���uiT��D�Xcύ�_����*�p
S�!��rǧ�����%?m��x:����'�qGxܨm��<����S2ZwK�%�׏�}�B@��J�n��.��L�c����� ¡��݊뜚Ť��X[{�췫�Ҁ'��5*�0�����&�C����[b��<�u�wF��X���M_�+�g�՟�ܗt�NQJe�A�,X��\����ASwTg����&�����[�3����m.v�B�u�C�9.�KT�C�_u ��{gz��X��Y!� �qX��j��uī����١�Z�0�e�N��@չ�`x��1�h`���,�eb���f���t����M�O������`����6�m����{��֎���Q�L�3��;���FV�H���T �z��i��9���g*�ϯ�^%�Vo#����0���n/�ٷ��[R��ٱJ�۰<mՈ�s�@baۓ�=�[����&���e���̮E= �XG_aΓ��9q~�X�Ջ hL�l��X�xj�<M�(I ,�;v�O2����|h�5*��YP�J���DKR�_��=�ƛS��m���_SZg��g��'�pf��R�w�S�#�:3'��R:Qmj�	B�4�?mÀ&���?�մ��4`��M�����7��)���-&�eWb�lG�X��0��Vq&��X�,���9ͨ]�׊�$ɰ5�[��~y��8&ْ�o���s����e�˥�5��䱦
�$ 䚣B< ��'
���1霑�;3����k�Eִ
x`����?F����c*�&m̛��8���!��孟p��Ѱ��xRۻ��{�� ��d&�VX� ��?�C=�C{���5��ƿ�<~�j��.PQ��1�/gRY��r�/�N�Tۑpu�|�	g�?��u��\ ��� �O��)�4q�P}89��|�����ǣ@m]c���o,s��~OC�t�Iz��(�̽�n�;'�kר8u狾��2�4�8�P�=&�?^a�l�,�{�@`M�xק6#d�zɧ�H�^1�VoA�h���u
F�GD��-����#�9?��~������7v��o��}[7��@��qK6�`�wv!׮�E"[P��,��4ŕ�@��Sb�u@���1қ%��htlns֊�����p�k�J�G���S��d�Ĭ]��zL�ex�Qb3UX�d�I��d�>c�ԯ����,ϼW�p�@���KW���}�	3��)����T������_n�n�S���gi��X�|�5�\W���W����$����d��[ڄ�"a�|"�E-m*��Sȥ��m�Ƣ�g+ߵ�m�s"�ǇZx�;l�f�Hea��q|=l�"c+vk�Zv�F= �ʙ�+��W��o?�%-�"���\;�9��u�c>kV��5���˨�~ǇDo=���] ᢽ��ن��HJj���5����u`&�$�?r�g��]?���x�H��pP�[��a��N覱}���_�ƯN��`Z;q1�P�]�pv�l����0~��.>�\LΠ�����Nn���q����J.�p����D��5�IRl�r}L�͎!��x�v�кpx�����O��?��-w$["�Sw� �b�;����{�@>�f
�%�SN/:��l,O�h��gY9�O މU_aZ�Rd�އu䩍�1э:P�|fb���[/g�_�jz�p��ֻ!M})&Wʍ����������4*�LZ�)^XNDҎ�"��Ҝ�%y(�K��7����qO�51��8��Hݎ! ����uK�y>z	G ��,4��R�?��zJ<R��bi[�d����D$u��ʵsT\��/�ζy�,��"�;���/�N�aW���h�������J'��Dq_fڮ��Ki��f����Bԓ�^�PԹQܗ��V�pJ�[Il�</��N�;<T��6k$R�
ύ�n1�H{LD�� �tzy`W51��n\�%PY�ʤ%�ri?X�`2��~�k���$\Gk
�Z����2��ذQ��G�`XDT{���=u�M���:_�W<���oRb	�����@/Vn��|V�_�[��t�dB�*�ko%~�}�` /����B���.W��V\ \'E��7���j�zɤ9�ңB�:��=�[��>�GC�Qc!Z0�Z&Ƽ�����h�$H�=�ve\����?��
T�����*H�@��o��*�_��E^']��a� �.6
�xm	�
B:k���\ÿ"D��g�R�!�ȡd֓1����E�~���	r��me>����OA�k��K��+� �h�LT��ì4�H��f祥�5]_��	���L���Ԗ9��[@��\ܦi�b*'pm�Ƌ{�:��5g5/��V�7A�ף޼�p�P��9��B_3|��VlĞ"�J��W��:H�젿�qD��x�MJ��66Z�!Y�Q��xi2�$XD惣_d@���&�gK��O�����##�u�Ŕni�  �aX|)`�B���0FܐX_�Lmΰ�	���I�(���`<u�.������{Q����|g��~��� cBJ)�B��Ǌ_�9r��<��3m���l:+�CW)�r ����=䤆�� DjOX�H�qg���xW����t�g��w�"���8���r�b�&�Tٯ���n
2���ƫ�<�2 M}��\����˸bmᄟމ��:p�R7�h��E_���ϟb�B�r7}[� %u�)�Z$�3M�g�k����/3Z����M<��٠),O�if��M�GpHQ��DN̈́gHq�db륔?��#�%
$��y��6��:n?e�u�'#~wc�.�Wv���]Qo���n3�#��f�.��b������f�y���]��s8Cv�,(���/��b3��C�ɻ��PrYe{�.��iR3��q|�}/�9{�GBBtm%��w��‘�E
X�)hO:K��C,����ʃ���ϯ���D|`�y}�y^3hN�a���w-Kt��'Z]r:J�z�B�=�m�W���^�}J�,�4������Å�p�A
�
mQ]jb�]�?{���N���rt���+���ey�G�p��Yg&دVd��A����i�U� ;�����]�Ⓓ4�"Ro,�aX:��9P�@fE�x�a8+i��0�u���j-����G�:�}��ɵ�E!�jw�Q��V"H���J�������^W�Vk�n�-�JR#FNa Q�y��bf����2"�����:x)Y�Ε����t��\�2:b�b>���?l�4��3���BW+���v��V��	�'�T`�[Ǧ��k�i|("L`k�u ��g�Wf��dbC��7���}kN(����Bݷ�����2��BG��eV�H��V�˶�,��|ĬC�^� ��r���i�Q���[�*����-�Pai�X
��S/����Y����a/%?i�a�F���b��P�������.E�9:Q�U"k��ۄ.�c;�)��y�I��k��m?y�2�")0H��u�4���K���z���\9{���.�� ���.�7o��>��A��q���kZg	AC$C������8�G�
e$�A��o	���p�QH�*,E!���y��vQ���bw��bC�d'�0�E��:�����݇id�o��/�5SdH�G�<g%�i�Y�b���;�QO8����[���W���&q��v�#F��'S�"�h���o������I���`0n����B�H	v_�o ���|��?$T�P S�tw2^�s�*Mj�!J�x�=��Az<bۧ��z��i�QW�3�k��ࣛ@�z��4!T�`���յ�a}�r��ͱ������|��a�b�`��RS_Kx��[H	�`����B���M�g1"��� �춌J����������$_�΢ z\�W�������������ҩ�\'�=Ӛk5��ro��DH���l��~�@�k���a��{���P2����0k��	��*0łƾ_4����J<O*��w���}2ͅ@�;p����J��L��`U�l@��z7��\&!��� 0�S1�`a4˱k`O��!�
��^;P��0RƦ7a��R"�3����ݴ�%�����@_��է.�_�bA^�2�-�j8Ǉ\��@��&�p.Ya��4H���N&q�_�c��������#c���`�/�p9���C+�0�>x�H��4��PN��K����<_`M`~��s?N.}hK݅��[��`6�X�pt�+������86Y4���/ۜ�Qw�j��w
��i)�Z���
��%`�A�U��;��R(��݂^�aZ��m�7?�#���ǿ_���+�"��1���Tw.���S�b��'�4.�]i{L<U�P{?2/�G��X�:Pb�Nf
����쏒����U)}i���on)��5�Ͻ��cTT]�.qFްc'PE4z &�b�2��������B�Yơt��H T�Ҩ�8�q9X�X}��!�}��k�l�A��7^�ɇ�E�������o�W@�٬��jD%��I#R�����,C[�	+��K�����9��pJ�)�}-����I�z���F��ף?�6H-u���?�t ���Ψ`�uڝ}�r!��f�J�
��5b����p��]�	bM����cv�|h)�b�nd�ќ@ �BQ} ƥ�=�����Ѻ1�9�]�Ԅ��Ҥ�/v!p���~��'Љ"C�r���Y�����H�Q���"`�Q�.6.4R�dW'w��agQ>��k���p$�����y�@;��Z�����\�U2� 6�Mo��e�7���y� 9(Fp� G=��W$3�����ܒ<)T�:�7dێ	�������H�ƪ�J�-Kw��(�Y:<�	�������<�i �W�C����ë1�H&�Ũ�ao������t�t��.��f�������G�PՅ�O�vPs�HP���aQ�J�Xzǯ��� *bm��l�*�ӹ���ٜ�]�/^J�N��0Ӌ�b
F�ݦm��rX��Ø3�O�! �����0wh��r/�Yw�X��718%\����І>TLZ�1�~�˖)'�}��M�'��]+��#
�K�����{�`��=�I��ւ�b<UjlX�yK��H�8�MsZ��.'�����&�L��g�+VCò��־ZN��d#k�!�%%��MЭ�4O-���=@�8��h�2>��rЀ�ॄ��D�(�%����$k��1��Y8�FI:��c�a������v4���/������[�PuF��r�"'T���W���U�tDc���q��ɫ���c�r��Y���fΣ(��FC�G��E;��ߤ%�����]Z�w�L-)���1)H�G+?�5�K/6u)��	�])�[��'ێ�3!E��@�=����(�E�G��e�����w%��l�����q �Q�_�ꋏ֥�w%�#m��wbCsA&�=d�A�)�܁0�v�-�?�։�:�l�U���_6�j�I���'_F6���ƶ�b�h�s�����K�a����g������E��ٟ"��,�?\/�W�[�SUAs(2���iz��J{�8�5�Z��"cem�� �M�?Y*XG��$=7
�����nD��� ��X�c��~����2�yl�(�3��*l�:^�3����@�z�¯�w�Ү��U^}�k���i��R�+>�2�~za�Ė� ��ٽ�/}�]��[f{A��
�����,��Jԣӈ���mzh*S�!8�cH����+�;bf/�_��@4*m:qn�5w��&�v��픿�z9�����5	΋ ��%���IЛ�,v7�� <c-]j���9�z�����f����:#�m�)�h��^"J�p��e�����������k��\Nrencә�4��i�:���.~�Ŷ��B����!��k�����cvTr�y�Q��<�B*D?D����?a��X1S$։_?�ۖ+Үm� ��16�\~��یM��&�.���T��$�{��B&jks_�R��
���dä��&�K1E�X��3+[���֥5X�l���'67��E%.����8L��ɷ��"��w��6�v���;�ђ���{Bv�U|�	�p��A�j6	ja�ӯ���C|ݯ`r��6�_�[tV��.�F팚V_q����e����,�0TP�n^e�ԡ"�hğ,�݇3�3�)�׉�B��>�0;s],(S}g;�%K��Gd�=�%��� ���:;�@3oH�;�K��C��*�>og4 c�N��ʏ��2�0�����|�U���c�X��y�!_c�WQYG���Y��ӥL�q	�
g~(����)�at��7�tfj���9�He���W=�֯p$�'�U��e8Ps���7F���Tp��:�l<!��,�ùY3�ie��8y/i���6��_