-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
--pragma protect begin_protected
--pragma protect encrypt_agent="NCPROTECT"
--pragma protect encrypt_agent_info="Encrypted using API"
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
--pragma protect key_method=RSA
--pragma protect key_block
QPBZqsFwPu3DGb9//Ml4/dseRKkryPMUZVdkfvSE0HzvY2gkm2JNDCRPzzlP2nQr
EJ3/8/yC7yeX8fP7gUss0RlBWzpw2QRt7RTfSPJhBy1MgbXC+uArFtOI+db4mY3e
cfRcX9i0bydFATD5q3s6TgWfKlQ3XZ13EaFl3FtTb7bNUzYLNpC9bCWQOxBgaEcy
XFBx0mNe3SecIWtKd3KVH8f3K7EGWKL7jHQT7Gjr1Cg+opMnnKYBNTN3a+E2d3Zt
33QLtlQYfToGPwnI1eICvk22bcLSpzIBT4dlrleqpNHRzfBY+CxTOeiBbrsEWA4+
XMK0tU6mo9yJ47U0/57e8A==
--pragma protect end_key_block
--pragma protect digest_block
Q4CAWzP6f4oSmqxQ12DvUNKDMAQ=
--pragma protect end_digest_block
--pragma protect data_block
jL5Gro4lfkaHqM5SRBOKH1sxrPrQdiNZb6SO6go/+L+1u2tZvOcv/hVmpEephLRd
0mb0kOj/AMueC60/qU1fobOukND8kCHIrou4CQ8GmVMgvJKFptCwYIswTTeE3TZ2
WlK9g5wbBeJ3X8jQoG2piJTRzCOjP10A24vHgwvJ9V89yikmFC9ghVIsHAOYnbj7
9xLdiOc4d/xetllLGghBGVMlE7Am6C4SvByaKNEg12R2sGdBySIBbniSJKlV8AQs
8sOZJZl2hre06UeQmXhuGHoGpvZx7atW/XfvqTwS7DZImZxDz8/i8pfEXeJpKmQD
Uwb0cVIPV4VklRNojh+p5qcgsfx0Ab89BqoGsNaOT80JK6yX9CXd6i+wjwsRExt9
n8tvkPxhXZAd1Zx5QLMcjvxy6cP/Nc/48RV+hygEKQs2RQx19i3+kkCbk4m6S1/7
77Q0xe0y0/zrx6x6HobX/bFsa5+6+FNO7ILlt+qUDUz9XlTieboDI4khYaXfTGBH
zsbdbe1avfr7vuICLHLkedNb23/LtfJB+dbONDTjTthbx2fm45OEgbBNvAuvdPW+
dPimKZ1NXo1ydHk1Tp0bv3PndbaN+yRirRod1/Uv0Pw3Aq3798Ze6qjHIHx+AdK7
p/lvpOviOQX17cziFEDgghLA2jJ7x2pQ+Qxbn7ZFYgyXifODyQgI5SkWlr+q/4Dd
0jcMwWE37l2Z1oxiTYwyazvvLnGachsDS+xs25Esg5FI4u/In+QdEUX8uNIbE7rM
OEMDY9sO3AP4d0Uhkpf2/yIohQW/bvPkBGmUKws/SM//6khJE2HSwJEWS+RALfzR
oqAtfCOwLRMCekc5Xw53yBynNUeSU3aao/mVfosIlx5slIBmKxPsbOTnold/X7cP
5Uek+kH4XE/ErKZOjDTNaTfnPJD9+k75TdIw9HTkTx+lRFJAH9VW5mIUJaOa9vXt
8EDZTi1wJwjls20Wmsj0RO15makwadfoWcGeEV/v2kl6d+hodj1VYR2q9OQo0hxs
5yaHV8P98xJ9GhSNDba7MUldNUsoawy1pP5QkCo4Jp2TChVkn1jAxDtb37E5BcTT
ghJys2zlyJy6mpjGguoZwFzPrQExZpW/sqIcrC8654bL0oCYz+ZK9ZgFMNpIFmzk
T56Di5iyZL6p+7AlT5uyR2m7XSO1N+AC9NQOZ4bm95aXB2Mee92lM1nCIiqJEaZR
ypd+1vEES4M1lLrwPcXLa8pWUSsZmw1Bb+lQ0K4MR0UEReQlmOZuAJ8uO62HiM6G
H/lOXEK2TZWoX4CSY0LP7hqjs+T2Rse35sI5rXsMnvdPZ9rLdQggvg1GrZVqCrVM
cCN0fcEqGcaAacF6PyqeIyxjwiJEA9v2oytSwADd54Ys/Uzd+HeIfPMylE+97vfr
F7WLFn6n491RqfUUxD7Z+BizODAcafvgTN85/4Loq4mMoi/zvyBBS0UW+d+HY0gQ
FSdTNDmPcY1E6znInDPgyxhanbCEit/Ixv8Jys1593M1xMUUy7CshdKlxqj0tN0w
SquAqyZ6IVyo0S2IKME8XGwnN3TWTT+N2cI0FwlmlQXmxzX9RAzPnuhZ9Lb/4YGZ
OwaXU5YJfuXODpocWdopCwcUDm/S8TJ+SBwE2Ls4lRPvtptkLm5FoxYzKqtWLh5Q
2htAVFvwmVLlPnEFptQtJMG8bNwC/Bt8KPveanKRcnpZ7jkQTuNIMBSsIxDCojpN
rQopP839ly1PAsDiSpCXICD8lZx6JINwZXuJ/N4/aMLRWrgV3Pio+yDUN6uFYLJn
T197Am4pR22U1oGF582i8xE/VPdTTsf42Wpx2227TlP3BW/SoF5sUybJevnf2oXz
sOvhOBFCzxR6yBKdR4sQ8l3jfnvISPQEak/DavEy3SyuMGU9nNRcSLXjLnQQqI59
ZogmByeH6IshM7qUL8z6tn5OA2a2CwiFqrqnWw0Jb2EWtfeco/0VtC2g2IYgiHQa
toQIjpOZPWqBF40UusajBjzrTT8e4Mp1iDZ752+gENHrFIadqj3zY482Cp/vUhxp
nSivI7Llp6zP/vNLTaDueRSo6+3wvYP7522rQ3nLF02v6lWcJfRcex4DNo68rcxJ
Nxaiu2q7gE+VLchLYyyuxC10xSkkT37VDecFFx/9D+TIDhFdyEuw8vjrNmULybqK
iTNLrKTgaJUFBixqIhwu19iNJ3zzdWarbRqIGz0dc5H0Nx2XqU0Q7a9MPBHXesdl
VivKlK3zzNJsq5kKn9n0Ox7ooyBckynTLUyd5nKsWgNHnIDoqQavlm35hxQqbDdw
0zkCYqxPaOe44lBxLJlD+qSv3s+3FgqPdSPIbnVZC1/sjRrQqrH9a6LvNcgWyGkm
czQ38Z/VYKyMVrH2/LKyx/wX6nZvcvpqvd3BDmAlgS5EEPeuP3LpSCNiu2+vxkHY
jZrourPmby7LWYWoXY8VXVClS/n/ELGf6/JVIyiSRP6NSWICUWlINQgQPKsloNlB
3Z94d5hYdqjxPHxtvywXTFwHp//yz6Az6hPneg46/M2eCnboFzw1YFVrGF5ND4bU
CQgXVX6cL8kV0pB8s8OpPdl0q3mRPB9KjMaU2AMDcAwvYfK0bODFGWOGWDMpDXIh
8yj9jkgmEytSKha/TSgD8iA0NBcrCg9jW82qkmljzAihorE2RGfqwkEc/SoORVhJ
kroEGuxq4iSUM35fUMM9+USkDV5KE5cyFFey334biW5TujaqoigRo05NtP/l9O+o
wD7J4Wx2zW86MxKfx0bqH40ArWmJ7kEGiYPQTI+FWTCuNNKEQVVnfoZDOn+KhKTR
GZASIBVp2KPn4wud4Ubp7yLo132HAQW9t7UY9Vg2oMxkdPPHlYiwId+n0rLOc6TC
026sTKSXsAHJldg5uScUTeok1+t+WwkwrZsqigVrVl7SrRyj6zcWYL8Q9YujGfGU
Us3w2dklIA1kVLk7JVHRojauFnQuwRvStxda8RERF19VqIoLvoHL2s9PPlnaXv4+
GSD8m79nlfDqAg+2npGOIkJVAukElmipbL/3zk5MI7TgNc3UO/6wor7zsurHcehm
WMQrV4c0JhOSp36Ur2wyeslBAhnozFv4tYDggKM/Xks78O2NH8Dy/Sf3kmtFcfCD
wFrlEqeCtvcmY1YVguYjOIUKtxQbWStslqI+V9oHcJWx5SooMMBjRqr1eDBK9aq0
HreHi4Zo4A9uYLaGM4NN1gYNyIlZBXnVAgB39XZjsmPT6X7f9pYxZCJtjeNth8eT
NMkOHYxewHOuJCqgGFgZYUbTS2vBtatRcgSvEudv55orhLfRxBXJc0Dy6yMAgCpW
pRC5HlCqdql3Zk6q8jIBQHboQXni1BQMRSOoPzzKLBQdZqKP4r497+ebo8vorj+2
SGYb7NZTWJ2WfefkPaIKADTlL4k1/FkzPbcOEV9ercHeaYxcAN5P6MwwhTQCh5A2
941oP2Gr0UpL9Dus/sDVu7w06aOc92DtCbKNyPxwBKoKIPPxL/mKDjRVRn5FVLNx
9yU0BiktzTfp743hABGi+rWimmSQTDa87S7RK2KkEAVbhL30l2Am2RAvLIRXHgfk
RJpsU3D+4niGPRq5B3L8ssVqtQKi4l10N5+wTg/zGgJ+DEQDUb8oBjqi+liydnXo
eHJOeBgvwMoarmeTSycpPvJCF+h+Ax22at80UfqJem6ozkNvQ+q5uUol0usmB+X8
RGn3JguRjkr5CLb9Jubj5P3yPgSSMGx0ojbJGrbs4CwIYSVh5Mx4BnKIa9FOMxO/
ZkvkFnnTmPlc97wntBpc3/ny98vR19CBEv3s7j4neHIjiXXC+QaIeoWG2T4/Ouo8
wWOiLOO905H4E+5h3nmQgR0mITOvK5j1G/iBk6jQWfsAtV4l8yRp5Nk0ZXYF7zPh
jO77whVZX5oKAvGfLlPqJcfNcSPwwgPIkYU005iHsx2n9N36r8YUGRLke54XlFe9
4RSPu7oZe3cA6QyvB2YU6D1PIK1GZYLWhyu+5+djn6vjunBqBMa7z49iU814hl26
Bzr3iUuWdSry5Ydjy7Tcqf48L+PbhuJ94y5IVnQ1++SqThBDn0iMoXKs8uax46Pn
AhK2+kXnsYkRmD8q3yISpa5wcwQ1vVfJU0wXajJsGQcmsuQ5y1COBUhF7D+TPVDv
3wsGgtgEyIZ+RwaTOunGE5z1b3HBc/+eut2eUhxXfJkY0MXeTkvbm4QA/vljcXwF
O/i3MrtoOlYY20JvIZzqu4laOC7LEClvvq4zhGqV9ZvLJwtaaGhYF6ihdDaN1rYN
MMw40GAiy32Hw6fBaD0Xc8a2W/B9zQP3nJ9oBsl5OJMbD2kMhcLeuB9DfQUHQrvq
X1uge15EJ1kCIzNJcoW5DHGjsemMZZFOAoAPV8koSH9XrhaQAdC22ScPejBD5Il2
AP00xpdpQxJWoyNsEPns3mmZlS1Bj+EGlRizj56vWBcQwwCaXtgfmeHJKbiV9Cgm
gpuV07HhHH0bOBh75K1dUDSDvNF9He5l5XlnmVu/Hqw9CC5oFtBoPG5Vh3PMSBiK
C2MH7akvMKTHU05RFBPtWrMuoxNxX0QqfbjXJLhmivX2EbA+ZpGoXfJSkjXi2gdz
XepvBybXb3Cql3aP1ZntbmXgqXnYsuxtntRIdjF44bMOsj57dTwkJ9DevgnJPS6p
S0VSDzyIYkVycwxAiFf8BBqI+oAdzaIj7G4INcRcnQBA8ghnJMJ0iryc5GptIgwe
7Aw/+A2lfbSwNZTvq03CJuDQlxRSitStHWp6cQxP0PbzD3oWMX7f8Jutzkxuo7Ds
T7856AvPHwF3rV2yTXWlEQXeqAXjRXF5BUjFf8lXtPWxisbt37PTGv/SDcIkXs6L
sSuoWNrFpOlpw1A49A5aRPlrZ8aH6+JK4YYWXC4BleWv6cvtSfXsfSbt0OQgHOj5
0cFERdU6dR4IroFfXkUwrgd09LKXrhILx1JcOkL34+4b3ifPw3/Di7ojQkj2GxgW
EtRQr10XxGKMCKy3dxy3HmP97wwdJDHJ0pWEQUWxIZ1EX7Gi+QhM9O8GWuAYbkS4
HHrSH0pgoJNmw0raWjGEMtwf0YvE55FsvaNCnp2GlPEaL86dWs+iojZgFV4XdxRn
afKTPCn9M7po8WCalctNXSIw0iRwcEVjXqaTT6U/OhwmsiWN/Fcko0gtCAOwVYDD
T+kmPiCTyzNXu2kAn/Pg8S+FKoa5FOiYCiupOPz5g01UgDiRKcEd/KnXkKHF49+Z
BpsrbJNT90VsGiHeWHxD9xcf0Mft1y3ZmXb+Gr3irJ9Une51l+hsV/XCIdJk2HOR
QKWLfS8BJYTsyr9EBkb85OOwOYUBsGXuNYas6zW7kgkXqIMFWx0S/lvWKW0cPTb8
XzcBWGzTaEldAJZRIbUluPeQqo5j7dHYbwD0nOZd0nVE474smU4psV4xxKZ0b3Jo
oG+97gwlEFjLRIknuwOFuGC2Npn3QLLZopLIy8g50KsU/0gqDoJDT+lbI5qoKRP6
KEnsyLT0MO5dHK/hEvm17n7WKTH48cs8jg1P9XzmFC27lVUJXNd/n+AGM5XElok4
4OgllMsqCr6YnyHpdT3ZEocPzEZzbcfDSL2CHqZC3R+6zD8Wkhm/QZrItbOwfOdl
IJuZnsMm0aTT3LflxN8cfXYBa8875krFPFhy2HrlAUPNQqV1Ktmf1x0JeyLDr0Z2
yTkRSg3uqMlnM4DOvvlzSPWn3GAzj5iKYj5Q/ZXVOzgQmtDEjv1aSYnmQ8Kij2x1
OyoiG7V0MypzztCxKSpZr0zyTG0aXjUbmrlcBf52p9fN9NZhpFz9OajI+qRWjSJO
aFQlECPbx05RqhzRXWffKFCSCBBf/9oyQSfuSOGi4qVtgLYa+3b+FHakC9uuUL2k
4FYlRznEuej8a/CZWLvM+Kv2pybuuL4qlC+Z2Xyodl/8OwelfrPl3c94JZiCOqE3
u9Em28qTpLTMrdPfDpFoNAb9hl9P6kZ9+XNCOR7zv71ZEtm9D8/eh/AUIdDniKG/
Ov4DKF2ox/a3UDP+BZr06yH0pgTEIJcllV38Owyw+UK12aVM2u4yvR9O+XcyE6Tq
quyuobGLJwYabQIvqsbcZuqdMYmwRpR0SE+xoYzvZ1c1Xxan++cqSoeDn55lcElI
nJqetrCNxZjjhsS3f1t4JOLF6TXkBkBsGEBM+7Hj2pg=
--pragma protect end_data_block
--pragma protect digest_block
KByG1aGFiwAMIGf4YBWRsMXfpPw=
--pragma protect end_digest_block
--pragma protect end_protected
