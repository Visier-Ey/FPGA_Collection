-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
oMXWXw3hc/KdZQKXOp6vqR635Hva2nlpOUcJ1EGSoT2YzaNTAVpBNITnaNKaPfW+
6ZOstvcT7rHebAwLUof5ZyPlbnZYAtiiQpopYyKWBvc40qiXQhra+Yw+HWc71FA4
o0IVyRuyaw+PiCUBedq0MB/nc/CzLmo9V/hL8Znc2VA=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 43972)

`protect DATA_BLOCK
1c7cVYmumBRM37f/8cKWi2Votbs5XeJncfnveWW90ce3b+uaEFqbj/Ts8lyOUnav
1ErmAF/YIEAjrX8N29NpYA0Xfg+O0m95vbQkP9LCDrC7lkwy0qexDQfuhtLCjQVA
uSm04IXZB2kOPziMee9puoiBrggpTcMvHDpqprqtJ55R8d01fOPXpwMgY/dLNaH8
BDJ+oiqpOR0rjk6jBecD8gIWF8A6UvNEsqPvnxM6K1v5JIucTghY/vVNWMTcYntK
4xwNxvt624odokFQs+5Mx7afhTJxu2EIouytlGfFYD5nQBvrto+zZfUXlBbnaNmU
SZmiQB1OvGauSnD5HjyH2SZOqtDVvlwce2CTA//fqFuEDorY4+m7pW+c1Nn9RKww
a+rkzgSUzXg0AVIP28hzrzfUubH2F2O2aNOpoNtNCjne1DphUTbkIqonhCHedsib
VMoUfaAP3PWEKqEEYHZwVuIiZwa/PLPCUiBfmQAezCK674YDkKn7CFB2feCKudYG
EZjBHEdmmTor1SHkBw8Jy5JvzvP2sjWQOn7oy3OuWmAuMXymslrRJBje9guGUYxA
9bzK7e0SyHEbfQ4A6IRh28rgunUt/LTZj902YVlH8qbZGOW2rWWgjrfWhEHZnVWp
pZ2jKjahaeu/n9t0rpQ76ebAK82egG6DunRmn2HuWnSgCoWyHUDaR5zsfXRyB130
V2KprEme++fDImKbyKtNHlcWTjbMvD4dbRFqiG84ZpT9lWeuY+Ticgc6X7NN6dil
su/K+OXZytZ3JOzz9pW/NsiOJEdpviDNOcasTdmS5KGDpndm1S2M/JzkU7n0PyuB
gjDXZZX974Dug6QtyOZ42fAOAolm+p7dQBp06H5YApX8bigVVm+0vsn6QVSj4dM5
w/K8m17PZUwnQ4+hUQlVMXAG0VglizcqB/zR2B9alMHsRDWB0FRuqED/y6cqQfpo
SNwpcm+XITy0qAhui8whKIdEu5zdBRy4b8uEj6X5RMUU8PVLnUbbuzcsgLFWZs7y
X39zTVlgZQAu868kErrXz/WKK2dpA0ay97MT0Wt14v8gRkge1NbHn01L3MlyqMDk
IQFpx4jKQvHCIlEadj9VHbqizY1KwY5QrogFhiaFbA7Ks564pD8YjE3XMq8cJd20
4Pqk7gfkkXLHiu39udOqO7C7Y+gznUDIeT5Q6oKqticLck2MXICiwRcAqi7z23D2
5cPXikdyi5VtToWw3yah9TH47aLflkulduhVO0HuUNOV6vXvX6HF4d34n7JtVFAe
6sODmL0jxYCPNtTgK5BzylN9LNK3bsKGuWo/Nw2qx0rgC6V5S9+IVxw3eI/STIxc
54PJ8aYSsGwTLtoCf6t2/nWM19cA72rPQGF8zAfsJUdHoBPiAXMHsJN1MrMZ288W
e0UrLo7R0Yv8V/aeOQVXoNJFHkIj5gqAbX/I/BZW+3L5O5zFSRWg55MpTaXb+erH
Sg0mhUk8IBMM/nkwtg1bG/MRi1HTosAsg49EI6A/j1MZKSicZlT9t7WDrPcB0cT9
H76rfnpDfEdJ4pXl4QTnQShz2nrkTRasr1Ei1hev1SX+x/aH/fXTldL7GxUN5Vd7
vncXhcLboWLPfd/rGCBnhXAqmnhzLh3sqEV09aAhtJTOy9EyvxMPYZcmV5S8PDCd
KYJUGcnU97G9dcsCRfE9J8VMhGrJRNzuui/f8rjLEXyitZkJgB5u2LdCpPbOnE0d
ZmpAbs9eEuOWkKDJ2F2Ps2ZmZeg63IIae0zblBP137BHp2dcX8wvEcHFcPiV3XBE
YWWX8+O3FCnUkBj/zkFbgL1WLZ8o4YZGa+sS8270NcY45xrtOcn6v7SsSlPPB/Uj
mQT3rXkUXg00cnGihMqbyTMzyZVWyvAdCZ28dm38VqRT4wpFtQktkfduDp9Ycp5m
/lMKcwNu1MMw6MOTZWM/PEcdtVlrBMENE7bihueWGZlp6FES938mj+sHQccrNg/0
Z8pXTB8q0Gk4WwEwgyPlvDAvS4VWXvmNSkhZ4KB+taTFbEwi7llPhygVeu6jqrIk
AME25/MVZYX5OvO1nzWpsPJunBCAdavOQlLKhn8l5RU8zvyAhyM/x74th8PoyYX8
K+aqe2fOQ7eGvVdLzikjWFwXjes3pwFvQr824hfUkwd9EyNwQqdD7MJr1Go55byn
SoBFia2Ui2ME6r8sFvnAYlsIUZnOlFrFi5O4zQGCfJh2BkfB8OGSfJTD1rBBpTJJ
lRy8bEAAiAYH/vu/EcCaMBlt/BYpF9PoXCKD2zrf/cQKOi1dChsnE52DDj5r6ANk
Bzf0Cn6BRpzBCLcDxodypt4fL7FnjVnQXC2jn61HMSEXjBcNAxwO9GQ+sdp39AbR
TXdIFAXlj49dMqmJMagGvx+OBYJJDz2VYeGLhLLIK+gc5PTwzKqP/kS/q8Yc6yhk
bOwifCBQHwfxJzM1TsfbhgHrRRz8CfDZU789Lbyr9MDmybUXRk/16u+bXCq4N7eP
d5z5scx06TV5oziEv7KLR6fcUkaeKg+NeLB3k8EqmcZ7nna3/10K35M1L9QGJS65
lfFpjOYQUac1yMuSQBK+GEu+HmumjQhNsuU598kQb1Gh+K5gBNWLHfB6+cjgjqTX
+fEFXYIoQDOFEferFUNjEMXp9BzVcpGqSL5e3YR+mRXWumqgArtESpJzzRcgtIfD
VAz0oYBCyKRVurVwnK5QLYNDJqByPXjfBUvWqNTYpp7RIrR4abNdCATEyiAtRqAi
55CV7h+vbQaL+0f+mcGboOUthA6nDBMSfzQexrbNeiHFxxqjhWUY3VvFLALsKPs/
krA9xB1daIfIBsoEbVIgJxij+7hj9/9lHN21DE7KnQ06LEibjXiFb1UutrTXa5aT
pTVSxF4uC1VRY4KG+SbRk/d0spuOPgzdRrBskdOTjO/3tqPaDdmQK81RQEEvVjBE
X9AjLgUt5etyoGz00zu4/5BaJP5Buy/n7WclUAIop1C7QOd7t6q9Vfl4y0nt1wvL
rkR0DaIh5WP//0yAk5pU9kve5GKvIoaq5okXpQxWebnOGsGTuDn8C8hCgmpzCZD+
LYXinaKm/tcGf5BuTn4buyz1CLQk4jMGej5yVntagShquL9lJeWBH8fPLBJRfodw
boWv1GvHx2FgFrh28YLDBRUikFkQA1D3jq2TypbsF5T5Qw2kvJz4PiWdQ5er276w
G9i3EyeoSXCUMweeH0Vaft9YjJsJObPj06I5Y/akuebSi3/ZhUTdWXTsQ9rRI2AG
dEWkIiid9aLOYCq11VoncUJsJ2IQp1RUQp44B+qamtaXXIU6b9HDbKaQw3rY7gj3
cVbO2FucL5MH6gUcYqKfAovkG6nr7arumrG4RPxTsrploKKIx5QBW1Otm3gviVz2
2EL9O2pHXVz741DC2hssDau4lTwHgfSxcJf734ri88GkuqbwnW1wCxTizwSOG5QO
Fpz8daHA7ItCx/gemhclzMFG0aKJKJir66rOpErg+0jYipvz7iOjue0kA1AiUTBN
r8/WhYeIHyF+QO32te5JRkEqWSxz3TqNSRUri4x2rhsfKJ4jmSyVBEuntNT8MRDD
uQUZUCwllnnlfG68oKic+j9j9C1DrWeox7VX3UY6VrGH9UjgsBbfCNnBP3BTIeLe
epLG332m+AyYaB+ZhpHL5nplw4+phLsncB3ISpBIggNMfDN/E8kymeZSGScWVbfX
JivxCWobxbTcTHV9+UApBD2uoiw08H9IPCtNAqGOY3/MTo1fyc2OxIYLE8wqJc9I
ICvaQkzK0+5x7podo/V2lObdvDp+GGtICrTdU96TGEwQf617opcaLlMfw5lGIn31
UL+kwqCGrCVA8GZhTIhPMrpdiwWhjmhZ82VIsM3DTU37H2jMKS4SON0wsGhZSC2d
usXNuMwjLif6Vk0wXHrt+Z6vJ6mgcQd916uBDyKsSjqQG/N6mo0aqfHTZne5mGZE
Xzl4R81T6RI8BU8smss1aNG27es7CtPHOO8RTCdcoZXqeCBG3He1sU3wZ0kzXd/A
nsmMs6bQGp52lAC5TuO1AcEXRXZPBNlu5OHuFzJ2mLsJvYu7IE6iqZtlen0Q0Vm4
LlHiTr+ZhbMTn03NXd+lKNv7UxYAmQIJt1V+U939QLLtNXsSVFnkgGJgBIBaGAu1
1QkKS+UeitVVY8HQUe/cjlcrt+d/FeAJaDa6OdyhQ29jJzDFpki/3K+RRv2mrixL
U1fvOsodNwhtUwa4ZLnjInsuy+nxLTK8URglzT/6gLabM6n22J34hhbtFo7hO8G0
lnjfHKQEqVkLAKuAPW76uW/q6979GwmyWwZa/+NUWgqb4dzJaxAX8bGNXT9DuGaQ
ZxoupCLC3tfpjZi5Z7apDpsYHUgBXLf+FToes3cU2PM+leXEo82aLzwLLy4p6tZA
fA9KBenQMdMd4Ecg9+Sckfe5IgDeN5woyixw+6yjvy7t3u0n+vbEXN01/soBG8p3
N8Ov3XCIMW9so4OoBNu0SlcuZT4Ks4PPf+3LKbKifUJrkPx1PDhRFMoCP/wSoTnY
/l/8DLSW1uW3b3VyR2rryKb82p6N4QRN1yqt/bZO88CZOUw8QxFBnFuhYqi3q8PR
X9mKwSZAZLoZfpGOSvqi2wJXQ3NPiAUQMoQGfd1aOdYoDio4Feqdra3n5xMzMatl
BTj3sW1EhWiFWQx07aVov6+nsTRBBG0Wx8mFNSOmhieQ2+5+Ljix2AN4HywwjAS0
w0mxEFQcbcsjv1BcPaKmNKgpqdWrLGroc2//N9qAZyAQfod7yWSH5ncoM+1d0Sea
XR0gsjQyfH5/2otU9tSgCzX/UrfwsYJaMqPtmVfNM0lsb8AFd0MWwGBPnFcIla/9
V3cWPY7OxVarBR/YXink18nK0+xHPILnyfLM9XQyuyYrRHoDDaiPjfrTD+9Kn+SN
31Xzs4LJkGhfzIJKq2KKuTH78oE3GQBcUGVuN5jnbw89urtu5cHDZ1SqCRXY6wyz
lBsGknSB08fjQ+ZkKDqst+oiyc2dy15Ad8T+yVuIUnjTewptd8vG7G8RfsvAIKO8
JV4VRmUG3HNNgNSUJ10q6E9bc2KyeXeRI6V9KA2dI/EuFe28Q/DRLcpGEfi41vS8
PktCHFoOE+SJTeL4eprJmM82ylJAM4a8T1/xSqrGGEA47PQqGs8LlvIWlRGA0WXF
X2/QZNBe2H+14+f1/4X3Tldbf03L5tQlRS5Q4hQhJF6eDq/Hb/9UupVwCeiH8MUC
VG29pbSEgpJex2p0XWq4/jC2HWhINjdVZ6UE4Nl14vZZn7J6QTa3dFnrbS8lXfUm
9wfJImrzOqc0vUy5sR0of14cOIjMPRuvMwxB/0TxQpnzpr+y66ywc4zYUNWl7/wA
c+Do3k5tvm2d50sNzELp1kpMRAZv3RhbIZaTbcOB5cNNtibcAvfCEfmvLRq/nxPX
gN3MNI7C8/MlLJmU81mlkD2gG0vYzhYD8F8TvDBKpUHdu19inON6plRVv3WrEv84
bRvDAQ5bdzJ/Ga89PUohUZpj/yve4szRivtNGVFVkefoSnfc8Zg3JWEnAnRVE842
6keDk97ZDH4AK27yZz/U99vHmelMJPy9OUEKTMBzW7qKV1YGeFuJFX4bk6mBRCIJ
0K7EjpS0+7dWR9k4uBBCxEr42uvKdhHWm952WjneEdgADbm0J25AMKzlUmq3oEVJ
N5C6z0NFvOany27d2sUVTu4haqMNONEZkoYm5IZAhdDT20T/6S13obEeOQaDHYzw
ehGa5vTyFQWkd6erDGy4Y8v8jG9snQCshO+QXkyZ/aw50GLnxiysaD9IMnQLzOrb
fjgunsBqwCTTfTx4IKDl8TRcl7jOH/C6kw5H9DmqZLDRYNB+PXMEUO4ajHa3BPaJ
zIR2R7Sjdbf1uU6Fvo9S5RhLXD/yxYEmcdaZfpn3gHhxk9RpLM9LThjBmwBb4YnP
UYaAfuE0gtlgQ7wo3TKqsKCW/ZJX8PkBp9SlZawDnzC4VR1SAVfzhNW8HUMKXop/
FyvyJzgEVUsymL4vzsZYfFol97/Ho49A/EqisNjqHFgL9ZMBvr2gVj7dJvqnKEJ6
7MJjuAkgyh8vK1xkQT5R1bQVSA7gw2SU25SzNmxJKuIfosKiT7SNNkVP2pVF/KD2
Ha6fg14Ksiqrke/I4cfFH7BNiU3WwRTnWY4mAgcltvz61WT2FQ4Cqko1/Fkba9VS
mPwJSZ3PqhEj/ggezhfInHMzHfSRpEPhjDfOhXmVehDB3D90r8s1A8o0VocrBmmn
fY6Fb9ZCEPcOJE+JpJZY742Gea1F4AL0geHEJ8QsFqtC91syJB/RKVdWiHDy+7Ud
bLUwJEwVRS+ul9Vcu+11DAbxhGgt7X/W+CZHyExVu53Zavab+T7S/gmrmNTjzSGK
Bp8c4j+9gzqQwAjQjjsVptXqklC4T44JHrkD4DStJ+/99OVMC6cIuiZoU30HbAmE
CR6NhbAacF/Vm4JgnNWtYU67CEtDDrcv1mmbXcFLw2zFvEtUPu53rstMbL1+xDEu
XKPXW/y2+hurJmPxX7apL4KfxvE+ToLmWZNYOmPuLEayK6obFh00Ln+t+tLqqqFL
Zyu/GnRHZTQ/Ryu3E+D0zOuYGlRJfJwDcky/wYEWdv5l32s5XXj/c7Joea4V4ExS
ki7f/YsdQjXzvHhICQu+yoThXBub8oyG1ONblOZBJdl71ddnZXPdP3Aauaf33BAK
thTS63Gf6Gti2CyXFxf7RCWVplQMQC1ZDzEXziB94j1aWawqDBl1rq/Kt0k7pUKF
ySG2OA+SJXcrBTKB4lUvlUfAUvaNgXE+sO+KEv4MS5RNGs1xHbnMBZ5HqUxybtf/
Vo3ULShI4xGBb/MjHPuPrTyR9x4OVOTtZ/e2CBdaaoqcWwAKOWWq1IwX5oDzPZ0H
zkXPYZtHA3i5DZ2ioMddzw/MXC0aosSDQRBv/hkCA2eM+Zm+JBibKmQe99pN3UkS
e2rN6sJBwLhiHlXGQztEEjdk9+jC1TR9KI9Fzwq7JOkuHUVwx/ZZ3ROxQ2s+hdm2
vZtJjKiCyruqh3hx7jDvmD9evBlZ3iL34qKpYBYVA3V5Ice5Zsd9N9ipajAgCqn8
ISQ+Sxn9f5IJf6uc++5x19iZnwCxxU9Et/d4iOefinDoRZAERSHqrBrLk+AR4wOD
WAnuQK8gXwW0Jv4CUWDJJvI5RDE93PN7ZWr1HuyECdqCPyiq01xDhW0S6O3DZ+kR
i9n6SOxw9hitBeb1Cyp48pONCOpUotNWnQoa+/m8cHzCBqg7v+caX5xRifVwVBRh
11aqQ5sewGZ5L0du7WCbzoOMxy35YvdRr45Xd70Z4srOAY6wzdqmIf9TjRaV8ZWT
ossFA4rz/zbOZjTbrauPjuwfs3HP0R9jfsHuO+WPmTYEylkU98dQbkLfLymNIDHH
dlMmLh5Z4REVek0lfRNJrI4tPL9G1BueWXyhNiBODeFboUcImLIEg0ymSlDloHla
MgQhE/i5Abemv8V7dVe1VsI87St/xYDvoFYIdhPigeq2+bgYZCYiKVSYfrlN1zOu
nmCic8sPFV+srn02S60CbHDrVZHIVkUKV/n9t6lUl5/pzGjYoM6aav0esI3Nkr+N
FBTekiYBSMi1M4ydq0Mktj4lubCDwlkifeWiNZD+P6FVUlSb5YoB9M01Yf0tHmzh
wkQUEEL4QAbec60zwhmqmIOEMU01/1M0YGsq4qX7bGifrG6ViyFl7pdjV2B1SRvZ
D1TbgcDD9m0XYjmCvPNQf61t1dDl1sWil/ChrsgisCr/9Et1RUs7HoRpMivrRS5h
nAZll8J1o9z3NJqBsbUQ6wJIzmAkLSa4BrD5cR6pRz7TiQtXjhs0AaCE4kXXfh/U
RxzAwyv8bpQG/MDzq+rOAZzrEGSXiZDKUG93vXVq9XfiU+jpdfHlTvjt425bs6Wy
JQwzK/pdzQY1hFZozogrOjcsRs3kVxJgktBMEu8FUDugRLBcrJoyyz+KOBKotZzG
eD/Y4+ZuHjrRv6YsHERIUkx465OmifS+83wHhWBVVwz5m4F4hXPXXlh6XHutL0q8
m0qnzG9jTcXoaMexvqEuXwtO3R66yAO/sPdzN6HPjrVEYMWamuAjCgwBAYRSlfF2
BrgnfksPn9Mbv+AxG/tuu8iidPRIUc/IB8b+FMJ30dHAzRywQGGlwgnEAVb99FpC
Btg703lbe/gLa1xoqbI9U7EkJ10hsYnNYpmk2inmArFA0imTZ+FEgHSHQySeUwrp
j3DTocu1/ddHl7ZpsAikG754CHJfWVgaEeqcZ0TPSbJ37zVLY7CVRs42lqrw1JRy
c6iMJFAsckgU0RZxwwxziOgYvlveKEGAoDByN4IntWRNTbVBAvVc2DDxCSUn2vMx
wYUfpQXtpsUmvPAcO32o3HpjyqcNBaXrC5Xyo0gd8cV4yAhgtoVnRIjCX+p7JGS+
my5c+XNnm5Pb7tiAKnneFZE1SLzGfzfxBXTRrcAMyoaucqb/kgYfy3YrubuDoAMB
er4jpZWAN3AHcNN5JYYN4/jWJLbyYIbqbVPZU/OSBzT2lBBckm4E50M0PWfY6NeZ
Ba6MrjPJAF8sjH3lmBMdxFJikl4jmrdvGYb38ikLGS5Ze9eJmucgIdQ1XNQQtQs0
UD4epoL7TmIZD6oUwDYtwKVpYyb8TulOhX3DEb5bW0zxeEL880EHg9Fx8J/uXtRW
m5kLo5s0QXnvDIVuj4fX9tKIG3rhVMWdLERKPuwLjdfeE6e4qlZjF594LivVghR0
VEKZ0IgVmXJ6Gg49KkzuvYN5rRQHE6sxxsys1SqBAOy7OfVvhKlQw+2gzHzX4LmD
ctiF44PIz7apWQ+zx01wpOP1LPJLj6gwvoJDAsRWDu2W4/2M0yyyg2xZ9Ih6rLD8
Iqt5XzyPMJXP+0zRNXcTrCTrtQFQBBTsDjH+W0hd16TN2yDJ0rIKGny5o2wmLskD
5+2n9TDW6KOPWTYWKa5x7MeHbjCoE/69kGdY0mWY4hWg9OjrGMLuAPmoW3TtnxG5
warxSa4HlTrHpB1RLvRcr+J5iSIGij4tzpvpfTo7GUMs3EdLqtqtbkk2qiPPHpt3
NjZcnwh4XbFgYA1MdsdqYcXrtxTfKfPy5LwS5qmFrkU0DSSlOEGO1YFzw+8ZrLYA
1hFZmA5orElYU4rppbYSuixXTblzsHCpBOUoD5JVIYY5/Xh6hc1Hbn97DNqUsAkt
doxkBV02AANpDIOJSKNvVkkHEouVfBSp25hfdOv+r9qcLZyPZGL/KwDvvqLQPNMA
ltw53VkDShh8YFQA1TFlO5lUyQ0mj99U2VYx3JoJfq+AVCqkj9XtZ40BAZTbezsx
+7awcoz1fMc1zBmfjfDyErqfyBP7+niKAKOoHL6YxEsHMXeLEPZIjMiYOhqJ66sE
NUW7Hzf7juWJillX1rhczKXTq80PBAICUa+xavJqoW/dyoZUrJC7wqBNrU3g7p58
JroIekhRREQR+xUYl7XOHxLhMfSZq46D7GAaYmI5VcA6kJIgP4+/JmwUCBUySCds
slsS1GOkPWHSG84jprumbkof0mDyCYP/fwvadbuR9UmWdU8X0QM7SAzm9qXjIoos
WF6jVm1Fu37XA+A110glia7JgwDTiUM1TfGOguDrBRYhJYuNPVO20mRut0D5as6r
cW0sNDYUN3IKElKzVFWrTMLYh4sMIi/2dYr6syf8Jdumg4rbNKhUjB9ZUkDDU3N1
q3y23U/KmIsPq4hFjPCfgXsv3OsuLUnq8ZkyeWycMc48WQhYa1Or1jnmuwYhBgcu
xtmUwrpz4EhUsNSACdaDp84nERncW1QyWWsfGfQNZ7x0w1Haaut41P1x1GQQ8d0c
7lqCGmXic33MJF3Ck3LbuQGvs20fobcGjQfN3ddFBvzAxidt+DRTvRqN3ZHTAuBY
McLYCvjFljl8cd4gq7XX1hIWpVqIc2oXh3s9Pm6w/508L0OYNI1UmiWSk6WDiqdf
fZwROi3wd/1FqGmDsfw6Qg3hufC2I3Q133weIXJxmqKY67ExGqlNo79UVrsZM9s5
p73GKGWJPhSwmsKA+Q/0nmw50Ve4Tn6eP29IofNd1Fn8JAGa7yOK3OMgNne038QC
iM+gr8V0XAvlCTh+LOcC6ywzHEbMxML/TL1S3Gf1eVlwFcoYfCAJzsT/P8osanfW
So7qlEexrJIZdJC0I4K609tWdBrGzT7rvy8zKm1ChflYb518M+bb+tnTCoSeuRHl
QangInPvEIlpgATE6ahofkjObwYr51qW9t0A3PfzA8/YIHi7U8/p6wR9GD1Q4y6F
zmT4q3iDXjqcFxcLzzGnd9HN8X3yGmGAb8ZjOaVU5MnmjLKpTTimscyyDX6YKrSS
v3dC6Sn1j75XYvRg95ZdMhETr3xSVvbyPQmOV1p/CwR9W27XZ0m9uy+8fWroHHmC
UQIslTgnb1EDZ03zyTflwcHRqoxZNLLfUdQqp3WLzZEOMevM8t8lHHAUNIO+JZIW
cbBFR73ARIfQLrorQxhDIsrW5/zTjchJp/WavYga72dsRXBVJ0jIb0rML39lOWsI
6wH19McxJ3XhCWC/sNxY4YmO/Cr/ZzhjHmfegaRCVLhjxuaAz1HbS6sZE3t170YF
gVOQnWkvpyjZNILU2vJVvw8lMjA/43iRBxweXGCt8V2PsiGzZ5QG4RNi/Xk1lhME
73QFPolv3zedS1xkkIau80Bw9e/tbkegVTmcHDFIaro4hR2VyBwB5Md849NjKEPv
nPrUArqdf8W05kmknWKfpsjMC8Okohic6Z57X4CsNDFWk1cniRmeM9xCYPq3UjrG
TiJBM3M0fK07v0c4BdvVMlPMT10BUyDy8V0Us9q1Zw4Y+jJ6JSWf+yUa45lP7FBz
hXn/1Fr3+J7QK1ImhzZOnfWd3C4dqCAh/BVFv03HC0KMXNnHQFfG7bVwyU1HW999
OXFc/Z+89XrqAr6dS9LHu9LCT4hSdgciNVhdp1ix9u8vSO2z8QaSAcHCHW1alisI
5A+8EqNdymbygM9geOtEHIQK77v1UhIYWBnrYw5BC/2SOFebU/d+xB97lnEWOKYL
rVhdqujlR5bIKubiCyn2SCwJNOwVR05acaHuo/3ZVrYP4ou3nmwDMpNZp7DxEySS
HtMuYeRCsnUy+AvvDNQ0Ag6ee5anK9ZAjx+JRN3XUF9RbHdt8HbKwDgPFcW9jUUm
Zd4CjqX0814x0cvRq2qkd+bwJ72XrNwZB8lF1EI9Oehte0/f33lBw/iwRh54ywYw
w45Sg2k41xwJG18wQfSSpDuccWE63e+o0qCvbpGfYQSGLxQGVaQ5VRglxIRMSbE8
MtX9ivwQ3mHN7D9aaNGSW2BfewHVy0d/4BhclVAh6opd8N2ls79Na383BUf0CFFQ
6DDo3shDlyrzqBu4E/7aGOA3sGZgvUfZoDrQJ1BXpOoYXVpL+L09sf6oYnltwiDQ
ehss+jZyJcooz5V3KsVG+xFIxdtjIA3x9QEJ36T3zKTwfiDuWdjMeW1T2z8s5E3w
a8tZlrMpsKMrPe6IK7vitOqDfbvh+gUBCaVNc6+n1NnXLC4iNXZbWrhSHCK8xqGU
wFeLH7ntbuuBGComwcIJoHS279gJ6rbY1TEvoBo4IDQB2ERK0n3MvwbsIQbVbxwi
ukmka1ktlvfHzwDKuUXLSHK/Lw2AzJW5b79+GH49fJp1pTJhHPAVz9a3F/VJ9D8J
IkJ2dEdxextJG2/ht9fJTYw/9INbyLmJT9RdSmowIahzm3iQ2ug5P3Uh1pzu5Mu5
YsrnkmsoWUVB8cKmoXj8D3JnyCE5QAGDPTolfE06Eo755K2vVMRIWbmXlT95YO5d
/ceN/FllWaODRzfiFhYo3zz575K53YM9x7UdVEabp7pguHu5xi86ZKXbDuz+DFYf
XHKSLxCk6qY7Paq0uwAbfMh0jcC+SDHqlkypPF6lpF7hHFpjR5rVau34X+pXA7RU
bi2UUkmymTdJ5jhm5+1XjlfW4FbTroosWgxm+NUpxMalv0sQgkj2uxzRk9K3KL0l
D21kpmm1I02VWJL6UKz/rsFH+WPljIvHLraYC00YkhZnOz/ZRYGuo5R7uTGJ+eF2
AR0c9CsPLQMBRuCs9eq+0+PDflKTkC3ydP90LOvNgwvHfL1dGe+aytKapd79uj6O
AZJdNDcPXJDamf2yVoXtjd239QLBOBGRxKvf5PO54LpZF9dqS0mLeIxYY3JewLNe
DPwG0frHcUdd65Q3tWhV4OziwCcIrB574lnD1Rfs8SpTWWNHKoeEFRM64CLNqGWQ
SauAT6X1K6zvNKORx5Xa7rbxDSEN/znt/dT2gh1xoyCRPKpKlRB5ZM4OPon/vTXW
SdxE13SUBau+ONXbLJU4GbeQ8GjoUtQv905V5qel1O6f2JQOyZXzweYe3bJMa8ni
A6CEfwbjXtD5Z6UNB1yJjhloiA+190YJmN4CphMdvLkQGonPPl5snT9NakbgEAKl
pzYCyMsFQXqYu6BrV7Gwmy5wlYxAe0iZzZi28xM0CcvUqVKKWajEN83dzdOEk8Kn
RyYi3OHyy3XuF+SWy27sadFx4o63ET40mB1zyIIfR4CuAPGMcGBD4gXbEB14g8DA
oaGNyrC8HQkLUBgSxKtQC+hJYj6fFeboHmKIgJDbkdMnnjP1VVc/H2rmkiE9Rrys
DiACBdyIy5XFXV0P4uc7hT2OdFajJ2JFL3NffizEmHaIgTsjaHzaABf6mcsf7LD6
xpeqnqW1xl9sWeb1o2OQIhAUoFvP62Bn+6TKLffuhF92UeR/F0oamNSZ2z9egNkX
xY0EAgJ4PjolJ7NHv/2F7dj2xSIduy8ZVs5DlJugLtt3hNcUckRPLoT6Jb1lhs91
9BusAkQhXcgq19rUroZIRH6xxkQCiaffrUpizmWX2gifHWLalAsrMzg3con4rohs
ZFZhVdQt2t24dGvRhhURp/uJbj3DKIfjSob2r0HUSWzIc7wChw2uQa5iaJG7u1RE
ZUGX8v9yg54puMckQai8bEQ7X/N9QEG9O6tSb9OItlu98qOO/H4IWr7Egis0mV9F
y8NzfDLprHG/l53leUxctRQekVwYG68RJ4TwFzajkHA3uD8itG40Yh/pjPE4d6Vg
sM0qd8iCQORo/uVPSnrpE2Uw+CMDFZHM3tn6Z1x1oB3NSUk12Smry4/3UB0EvaGC
0PKRlpoTLbUfjOpCp1eOFk1Y8uWE5X+u04GDWr55NITX5VgCpYOqeTrBU0QKDYHE
f60OAvy7Wzxu+kQmSUz49RH1QUh56bNkALI5LpUOwv1RSZ7AakYSdtOVMzCLVk4e
JYZo7v0jEdF0jsKZPdnfTQ6dCvCN+nZhFrWyuOmSA9GYb0lRkzeZ6nflstcnPUc1
QVot99PRTydZRwvPDxpNIb4xXMOClUR5tJIZywh6akt4DYt2BEWScQYnmH32vIhj
BUw/zTzGStx6ukcXX9NicQ1Om0quu1ezFn2f+Kjd6mIdoY3Tq1xpXoq1z3NMWNav
RB7mLG8XmI/vcfsuDBpR1zexjOjcxsE/6IJWHNokHf/ivxc4/MXtrQBso47q/dTF
VXaLmJ3bslwgVsT3DVTvYduzumlkST1+ykSGlIwOqssVQxtrh4etwDDZmkLp8lqG
9CkDnHyQdtKv41hgKTW6BMuuH4SNn2NrWHMNnjgUoDABf513CEc4KgOueSV2fgUj
KKQbncrYfSZFBKz2LuimbnBZ4zXH2va8LD2D9hdJ4Mehwum3r46ln1q5dln/2bt8
YdeGVZFkjK2qzeheXH3QxhVM3NqCQR5ABqjbu2B8GJQDXG3sLFXuz0BIBn6jPiJJ
19/yVnnx2epg8sjef9htH4NVpDCFWw/a0TcclI7g/hZz5/6iwEjExaN4XXBTs2iD
6zDyfCwSGAcnxhgL20Q73lJyi+3F/bej6ejGOXegNcbZA10emY9Iyi+Dah7G52nm
YYAdiPBYbDbxxXqOddE8vJRsPPbABWgrvjsLnQNme6w1i3heEFuCrLwG4aCFEEEd
9/e2lzGsGu9XgX84AuMlGQ8Cm3tUe/WNNJRhrOLmEC5/Vf1JTWa7a1coMpz8l4nE
24+wLwk4n5pz06r9PDj6Khf901nNWdL2qb/a7jjzxsWnWfd2vr++JsN63qBvDkPN
oFYSrCI5Dl7TLgz3cSo6eAhWppEV26U5dIiZoJ/kgI2O8HNE3jMsMDMYicSxhJOP
llr+jg8N18DGyDlVf8qxberYeW+jsoOjZak0AiQNfBe5H+vZpEuXymp45xNMcNkC
2Tg0R/YPCs2GkyH4wkoAEFH0u+MXjnl/KQIvIlFakmKgADd4Py5HVvcvsr73DhnF
6SHfl+Z3jXJ9BbkzrfSSWjpxUUyaFXSBb0rzEX4pVnvNpwwQ31esslaZyfKdo25U
aZt66BYvlbv12UeM2R0Uvhi2SSi+eAX0rABBr2oSFmowM+OTMkN9KATruH+U5JQE
io6VbPK43wUuc2wRR43EaIVRTIFFOQMhkGz2DH1bDE/OZYVhsG84vqzhF7pyGnVq
kKNmXi4ZWOnmMqBYKS+SY7gIu8oYro+/qdYVFY+Lm1b6JNFXTyuWF2jFzHmbT3gx
OQ3B4wV1NbtGwpFgkdH0oGdh5vcJN4m2z436DzDsIBy6zIoyASPodxGcTZoq7n3h
OOsMCIYHLzv3sbxr1L3zCu0j6cmfwdpeUif7k06t61XZqbnFRaei7/r7tyUdIesE
5fL3vIbCuSFdFLtRgmSdoUfvvqHKYSaHu4yTxVGZa8bLHxx5bcCJzqqDipRFRKZ2
rkvVNiCG+zZAwT9VTQm1G/zWnDi2SKUfkYWpYPpwuhTsfCJpRP45UZQhi00Gx38/
TPi8U90IoDRjUdRrWDyUzitMjJH6ad2t4iTFTB4ZOGiEgyfs3hRjHluaQhBNdZNj
oMu3qV3AkSh7ZsG1N9OcYhvRO6IbveSTHTwMB9juAia/C2Lm30KWABoeepT11qTF
WogMoLwGnlC6cVOzCgP36KZwD7yJXcebuLlLPDX0QvvlXf+ZC+nAUa28RJagpDJK
q5c4GhVdFIFwxS3XamCzwKut49PkvqQMn9540gYYkDI8fo95jpTu+oNfCNym+Auq
mDLMl3ZdFP3QCZxo1Wugj/qsuC4m/T1M8wufQIvNcwaLRcPlAZnUCEeRazzLXFxC
lr9dXvpI+MFwEazORIhOg9irD8I5Foa2PhmZHEso8CGNl7lBgLhAMkE62E+nyCms
0e6ZuDu67IPg3I5fAUiP1RbAWef1UbwsBOuENk095moMsunm05hJh4A9sDngAwVC
inkIYs2QX8qepdI8+nYQHxy/Nd8lG0YwIYjda0khzVXcbJxyYDf48y+vVIczRdrB
K5rRZEedkasMXAvMg/GrArbKX0cIyaR06mO4yV/RPB3FM/FQJzqRObjoDybFAk07
L9M2E4vbJDp6x71PX6t46RxJaNnMBEqb9aOJ1rb5IcUz5vCxZYUs0buwwQGDQp9l
e0FFPGT3pOXnfgFoqoVlqxhuUZ6ELRny9cTQBlI6eKUi0nT1r9LFaeUvjgwqOHE/
0Ks7ZMkhDpSfCydTQwF6/1HQvuC6JYLkDUS+WIeMx/89M6R28/xzXwSQNfAmL9u8
5Xsuz2sy9t9tEmkvO4JWV1ti2oGlZ1VR1LyXt9OapaHbP5N8OdmSQh6Te9cAF8kg
Q7AvX8w05VvCZOiu0zYzlBtqfpxMEHdD79jABwN9P9IpobV/z9h1gSYvzspRXwOp
mn9shL+s4vMg0JE8pK2B/b2zZ93wQE33w40Htv/MdSg0Sn95y/Afu9VKG6GYaqkw
JTko2rooQDpMR47GGlZKCqlWJJ4TKLEAfVrnnVb9Eqnu67H2cdDVWlNNXRqxG3q0
RNDU3A79aVjn/GueNwbTbxGhZOwuzUec8b5+OxNy5ycw0VgFtLyQxA6c0Az4P9yi
Ljvj1z1uWhxI49Kv4OnKUzVkOvYBnejbHzSd1vkfc/Z3o/Fq46B/l7dKF3xdGx1z
t4f3ownX/97DA+g3gT7OeZPzs0Xj11d5TPpWpVJJQq/3k/X02Mc6FvAQZPUo/fbp
c5ahQtegm1pGxDk+3/c0/u9nP5cOuCycWACevH37R6EBiJ+NeMpuMD280nA1FW2O
iiSFLb9CqckCErZdREcDQ+rlA3D52GIszo0jnJBvuvTH/bcBEuc7peC5SYeI88bI
CtJerAumWIRFek9Uy88K75VL/dXoaL6XJYVdZz8uYxn97JlJ7Ig1t1ZmLRbbLQzr
ol1uz8UT/G4g+6RxSLmkY3+CtIhYfx1EjIe5355MyH1DImlJ6jYkQ8G5YWh7qtev
htptOmk7An9iNkCtkPJbR9nq1l3IygNREKhJEARLpOjp9twseuTh2SWPBGYRFN5C
x371/UouiAonrSdAUY+UgPMcTWRMNR3UQRj+gGdAgOuDAWRzRCN32GsX3FX3y0eP
cYRb71vPK27cr992pUMVRwNuQBlMcIuDD+oHEFdAi+0CAnElWAi6QAnHd4Rt3cUW
hjtEKQWjmpluRKttnrtqTw9OJgqftCkrKpt9G9uOxqmcuovrzD4mlSuCuCT0LV2O
7KtsD5/kb6jJu0QN8IbZ0fK2cMD8dnj5MoukaHdEiNbkJ9BYkhSKqkjXl4JX/F3s
zDaQa8ig4/0DpPyawUsyWt/l0JBu2i7dMXNgtPjQG22HIisAiHNY3kN+7KCpk8jD
PIgZ853dcupdPAkIni4dWkO7fttPAhzlhw7WqPsi24Hx9rBHCtMQUkp83+Z7FUGs
c0WNMsiklX++lBbNK2y7GyJblIPqbCFDGC/hShay8kwvnnOt2UXImFCTdDnIfNel
idCemFy7rowHzmdJIo4f6uO45JX35f+42r/uXJLAU5s2yCUIRBC6GhxvJMyt0RM+
3j/TYOj/an/ey9SHALM1dhNQltb6QWrMxZ8mcJ03v6M1DVhuQBwSsJ1hD+v/wg2L
Nkn0fN9kE9sGfH5p8vxiiPBWltsA9mJQ/MAPJW2ib8xLV0QsLUvkyKq76Q8iyp4W
D6vJm/Ht7GVhhG8rf0jtuaK3D0vpkck34GgV2Neq5ZFhFFekNDpKlH3d3Oy1ReBW
oGhAst26Y6bnrMoTLnS6/6fiCnxwb4TZRAAadKJVrehAD1KlYph468vgERu7lQNR
TqYsyIoq06NVcmBxaogzJsgMJDfWuFq7GuETQftKT6uq8tbWxVdaXWnFbzRy/Q62
YORBydJ5fNr49pmtvwgFlAmJ7fxXT/XEPMlG3kExk85kBoxQAc09sZHm8hLehHmR
VLxlJ1rYjqsKJb1jQaVtmOjvdB/JxFQznFeRKwCmZR6MAxxiID6HRIAHuNhEpZg9
JGycTiW8rLWnNKALUYkYM/osyP6wCryTolVNOrxwGmkNAwBd6p+0RVSlf8ybcmhl
/HuqXQwc6p2uceL99rKbhXDUfvgvvfR1YCzXPtBCRK8xp4PlPYYYnG6C6EVSactF
81TIMB0zZkGqJ8y+GN8dRBNrkeg6LVGa6kgnA/QnJT1U7b7h0UBkDYxVaXse8kei
4hKAf24QS+Wswm/0+EaI9+K9hY2hn3prOiWW60B1eBDK3CJHlTO0MUhVg32DspAx
X9/+XqF/szG9I2TF93vpPme6MfkMFjZyygSwq2TiI0f2dYE1TA3gIxDaQpx+IwlK
vAnKGZvlb1v/4ZJldmvzEVOOJYpO8qeccly//s1/+MdyCD4jyiWXSnkKaxEZtLsM
1WGGU54Pf0ak+q1u1Paztg/zc2YVjyAPOLtqSM5A4pYKZ5quHrL/BQE7HMnONany
uQUici53YA6bqtdw9ILiHcuZrNUOvolv7glH9HSiE9Aa10vL7Dmt5WBrP0xvVdDj
jh5v+Chn/JQm92tCfKWYVoS5eKCpxDcA4G/VLo6cB1mY6Ypk5vYi4wbkbTZFvuHX
DbQ6sZu1BjMSRmFXgt88ZRqjRTmw8sruBtASaxNe8kx5K3aVQRD0UOmUkODPvzLR
kqom9V05tW7ugMZRgdlFBAAEq8IBNXA7AtUeMgQjRtI0Bavb0vLPCZHCW8CVA6WS
FH1BB7ZRq0T5v4/TtwLLeg/X9ocsZByfnNCPKTEw4w7uG+wz7knpjPVXugxfwtqK
R3FBzSV4488Z6lMYDWBd5hukjapDoithbemwYGaWgXYvbCCuj5jqpLA1NjP4B4jh
KyJ4DnCgUZ9f/6zwC23c/MaMxydzyDa7EMee7pigdww4fGsmOaccnIAUfpGq8dsK
usWO7zHjHQhjg6g4eogWZ7RPdyo3Tg3D/doUYIIlQfQ/G2ZtzGdHPPUdpfy2+Ldv
1s5wFYcos/2FwSH41C0d6N7r57XEvY8a0amu2u5ZIQFdPp+E45zqtckjI/7fhAv9
WJzvIbqPf4H7cZ0pSIn4mzrzsGEQ96VZjvneEMg6qJLyr88IRdxPTEWDsNvrjmyj
WOh6sRfL4ZYLSBjqJT/YpkcpcYTnC8uY2o0LGSXOoMVcfVfvb64rEsRg2ogEInRQ
PbPdGfaDzfe4/FcT4FuAZgDE5fl4W9tJe1Bzitvj248HxXbhJaGgpZt62+4j8h79
0gRPCXRwfKbY6BxZvsvYfGRy0hCDPxpWxQ3MuXa6i2iOVgn1l2ALsDkt+RjykRcN
AFdWlbmHxxk1wkBgzDojYzWhOCdEjika3Y6FG4SlLppWFox1iyEzitljA/7n+K6b
zvPECRxDAm63Wnph0CcfDlXyUZqXZ11u/cft0NXHD13QII3eHPXFDKq2UlFA8IQ5
X7rwFTBLjso8TXofsPyTicq4t+L2A9B1mDfW4zvstUUzAFE8/4UYo2QLB7d2UMax
rKsBKCl6OkJUxPLHTOdLzbRAbiJnklMi1lgVZh2bH87FCpcCVGPr5012Fx/B7fDK
uE3gvrUdjBvYSKAlA96QQiVwbFPkQBFcwjTHiGPZj7peJXs6ItnVvEWaiD3CX/Id
HXSgjS12g1OaBjcPyM3TaS0aq1Sg0UE0SpB/vkor7KbCkaaqAmWEcIvMhfFQbEXD
433ZhEpiqYpGoK9dA2TsgKWnEUtBIIG64P8yBNXZ2tfJniQosIqndt7WPDcnskVK
yoBqHDUq08xivs4hV59UGmvRGBUlDCb4+3a+oN/vS0pV50bhZvjZ/AVr7Mqzd4TX
lSySGqnmIH0Zlqwg2idvkk93QlDsguTP3xj/aKVG0QUfC4Jbib1059MAucF8bDm1
3NDsuQYXrXBm/ZocnMMgX/q2Rfzf8TGBjiD0PVrUEleA7rHIcxphjwv80gt+LiV5
KukWpnSL+rRUsGM9Slh1vy9/XhT5ZbJsjbNAxjLhMRSVpUTaQeRzGqIG4vW+qY0r
wd4yfeDa/N22zYpgHu6brPxtOJFsZGWlQYDevdASmzOeiwVXkp5balYEtqLL2xFL
Iaj0TwQPdSPiMI1VMrCSWji3nmaAV9oTlA4sPjUEyo8q2p4jcOtU3oNQfv6Ibaw9
gmX/cBJIoTiZlPsh9ITPSueXryrk5p6OjwOu72248NELx3YZmBS628FYYdwb7E+S
dHfdoBhGIgHhF3R/dCZqC6iJpxauIH26XG39ZOZJpw+eiIigC7tcxJDI289G/EpO
N4k0tYMx8eNveCK7s5R2pvQ5CXHWNQny0RGI1FxiAM/YD2tgqLgrkz3/im2/cVA8
cdmtHy6u6q/6oJmEoX+iJWCQEyM5af/PMwKhY+AqGPfj3F0FjGMUxcjDXjkO5LKM
1ovExZh89OAsTGE1dnqlpsDqfWUCbhQLQp+UsInBZqiFhygrIo5pv1MNfr9CA0+D
j4lp0EFJaeGjQHvqpsJJGGicpRXI6IyGonva31ciK6HQJ7Th804/8LpiCNL10grO
6rZLINKJPiMwaUA9/612ias8ukGLMoGUW+itr3qv8sJ58/E35b9+wYGSjQalMEwZ
d/A22Ihyvlf6bQXnHUoaEJPv8nRXPjaGq3AkogSIidU+rkJaONxnjRYIrwilVJ86
1lYEYXJo1gl6MKlrQ9+TDS+G7DA3aB20eJWFIlox97VeXaym9QyBFeo4jjKehwec
tkEIw1tSVs1NAY3B7U/+cUWLvRNuGXriKPcwApwhrlMrfAnLdaONtQ28KUZ8QX8E
8MPMN2wbvTV4UxHApjMuzTQgfj/W1Jar0PjKeNq3oH5ZWViiRLib4j8CRYpXRku+
KjQnuRyk8xMOmZSX1KpXY7gEGUbQTFXLUupDbuV2qraZWoh3sn3lzQjF90NGVx55
4Z/NFo5OU2cysIsbj3p3KklbxmL5sfxt7K4L6SMI8vbwYUBfRovin/NnAHE34m/9
vMUNATYsHgfselagDdnu3z7GRNvjWQjlh0jLwIVZI9bg9xZvvtLvl7HN4MC8yLHB
2pDyZNXNUDzTIApQkjuei2bnYsGkM882JeWIcdb9yt8dKkcEbY79lVLgvO5xlenP
7LCpTPNukp+961D5dOFbAjmda6OjpHVmdS7V/7178bsja/xvC5c/5j35g6DksWUL
oGURk2P4sFhBJAHBaeOgdqg7hsx19+bhf4w5bW5F9CdswJwPc5DLog5aPJkW3L1d
X/xF4sRLsZJgX6DOUpjFJOK+/dUcM3C+EE1+dHnX5GB6yWbU4NcohkWZw1at0RDH
Rl68Z65/Mc4kPzxU159xJrh3zIeA1Wkpi9I8vowimopLZuFj6VQCshtuhkbJRv9d
xDSWN2B+6O6kHALHtcBrz2ZyCiHfbBumasLs2GRMiVB2sK91EOZuYeHYQ3tmlZYa
3lsOd2n+5FcyicBOL5M3CZ3LftvvCFdGD6OS0aBkjoHD+GeFzeyPSuxxlt+rPK8C
xuh6dTJTxTV96BDnv5Nv0W5qIG284LEV+h0rFbegHoo6nZXIwFciuCwSYlgKN21r
0z8vqZEzUok6zqCpax1eqLq3tTQ+udRvdMh4TQBfSIOEeUIpnSwF4V6r87k+Uohv
DM4fKjpY0qEvwj/o/kYNckR9TRr/aAqK2599kGUMBzJ9KGC12mf1rPiwLg71O2aR
d0QAQt851JX3B1lAssHTsqbDepmlG2CnfVeRcyEyP2L+1IWCVmOqmN35ZfWzvKMQ
atz3uY8gh3G4m3f1v9bcW95OrJaWXikZXBT7p981jklsrHp3vaHp4i0LiP3J05j4
vWPW+su6AFHPoYcUqDUyuCq9XiRKR23+PlZ6V/S0AU22um5GXFYmWwMXRWSGv+ST
2zxBTVzYDq1TkTl7sB2GY0Yu0CBe0QUsWBb561zlFPIJDgqkDZaCMFpm3P7HFuuW
oqp0U9SxFJIpxrq6cw0M2+3i0WEfuFTewLi9H/JvrISNwlAAenhZkqNzgoCMesFk
Z7kUmgw+lz/sMyLNX6aftuz+iDd9Z7ecaoFkCZSpXy39Bn5BAsGk5jwBwlb49s8Q
HSjSMujJtBpAI8fdd7TdMioYMvYmanePOFKS1o/cmCQlAJo3AoJpNpLYNjUYovkC
ihzIR6Mw+44adRiYSS1x86XOZ59Qp5dFeNuwIuQboVFy0NW9Dry3FQxF3AYSumJ0
m98s4BL5aCiP6cHd3uD4YlEdyeWMyaM5gFsgb//Jvs6KdiGK2bX2tx8xpcVjQHRH
d8WQuEDXplbIAsRJXIH9l+v0ez8mo1U8c2ZEDiQDTTJb4BS1nufMrWmss1vfJC+2
2/QxrLwdjh8zSg0DLmZ2ehG4aXfGvGiEeSKMQRYgEk3I0QDdtabIbGtbOOuv4o56
p5g5klXVJ0WuYSNZhyU5MbiEI/2/r9/W5+Hy25HPwkFd2h0Ruk1ud1+ihS2e8GdY
GBjkmEa1LhtPEGDgmEExTVmZHKao9STyw1Y8zMKw6Vkv2ehiZ3P7GUpLx73kKDRS
L3/IKVoCy3HrNzJ1Oijuo+jTFCXxG646+X7rZpE7rrd8LXU6MQON1S4Gr/6WzkCC
cd92TwBKccFMAWR7BO6zvWli+1V8XoDvTpdLkXmSglbk0wrIIZAvVAgN50IFV+nV
j72eoA7yeeF1SFhpmyR9FokFWDoMYxruRzfBjcr9EeKsYbwTkQ/JoO5W2VI6P1Av
jxqAkQwpjv0phfYKuvbHuiXPPnZxEmbBHu2QeqwY5mwtaArxnOXozId+Dm0w+WIg
u72DUAoeeZEyrsqVT5szBqGj7cXkvvWvmcCGWfEhuX+wW5G9eMEYxMISynbuoCxU
lzVQbBvsjWQwTYeSsBC8oYZKcy++ILCeBjk3ZYzbRtOEfl4pANRQo670Ky3TDcrE
F6+G7QCVXO54v9UK4Ze5YAan6PcZhJ35w4bczZIXClZPn4HfqyD0uGi66SbVDn1h
gWYYsM02Il4S9T94vezz4+282/RK7+c8jtHTOXIfggkcz6GFxB39s1QHEQlq1n7g
qVsZI4gIGKjvkj0Ga6aUoHM/z3gUVFwm9wZhvqPbgjejjbgugEyyKYMmpINXt1KX
JmCNsrcdcj/m2dU8eEQt3vbiv2dufa5vilLUWY4jgoTeWkk7bJaPpq1yY3SwG2Km
z7/qi7fzsf5IdCKj/PXKpNqlfC5/I+eXEDdhPKAWoFOAsbIsF2ivwXGw3XRaYvEe
kDJVT5omdAU/4OMripll3A5x0WcSpmzvjIXbYk0SGLQ2zz79sDLD19yNTMtGQHHQ
LMw8xNU/QPAwSMJ/VsQ023u4NScPtBqEt/S7LzjRVc8iPN7gEc4O3SvZXmz9b75v
w2JmoRFOgS4W8gQDdyLGwYlxQtOuRXjPqPWoF5mK2fzXHH1lb8YAfS12M4fizOaP
gtX3uCnOMLIUSs6UQ01+oW+ytvcdiFORjyxCga23wUf51siX3n85HM++uUKH16QP
cstlfWqU5CLFS10e9N8cehb8WxtxQUaPCajAVzs5SHu+KTsbAaxDVFmCKLh09CBx
bwt13lHReS7/KiG/xRdbWNmgjzjsdKvhfsx90lB3DUQBXAqdMJbAPm5Awaqt9FvH
NutYfUsBGdWzwLZNIEOrO6qnjR2XC4biB1/bVURofi+aSzsGtAX513dLTH4rRRdS
YaVW1ackTCgj0vfN6CIT+nzr6WZN5Y8SJmyPNkPlmf5W1efEixjRTz3WhiSBsM2i
t5R7yTTGLV2fxvlc/qWm9hWZEcskpnYK8rH+1uCtuI5Mhc02UfobYGoLxZMhj4BI
/Y6MRG9eXj6j/gnXOQhbDIqt46QQr5Z/IHeCoEJVZTC4W9PcW0ht2zexbJIHn3au
f/ZzKWic0rqd7GvqZMFf5Px7qrYmOOcp2aZxpy1CyIlHv3V0xlpN8WCVINWhzc4P
+Hq3MDOUGiD/41F33UHFycgDFYx9Mv/77+nGxK9BidJa3v1nXEDFXuCHKNttE8GI
mmgorlwQHCfSOoCHmD3hQLAAEYsFOeqL7vEHtn6ymqUpovLe76ZyiXkFC07I5zl5
NNpqovRxxrIPHSib6cA2Db9EN0b4z7Z/Y7MCO50BVj3Cybg/Wb1PeU/O2VWgwoGM
j3MvF3nbPXWfBTudndzLj27u4oXsSgUGWudLaapi1O/KXGaLW4hhYVXUVXcOpIwi
85SKKGoJ4Aizjng8MS37o20r8CAl/rzXPbh7rkdq7MzTE9ZCtpbx4Jjxhuodbd93
lbb63m7v1j/CsN/UdKhjZxdM3t1YHuMHNMIYB9TRZ8z7L7B9uYBVmfExVSP2mRBI
BsEtM/S+ykl/+Xq0xbu7uzl5FP0C47wRPOCS9nV8PsMfN1yNPYllQFvrlTMyaIz0
Quz4XhxGdI61yOmVPZijabhAsPKP4Rf6N8zfppHoaNQeF6jWLeS1m4+irEvyS/gU
RIBpQTNzbqlCIzzOtcoVE6vdldFtiBkISw0+/zsFJXbDQk2S+iyKQITGkbH8z8hg
c9o5GrsUlH5k1j0JbgQGK+ITin4/HU04ljmA6rSt/QA2K9/a/fkGKB+cQjYYNosu
rwJ4ASIVR6FNtv7uXkXfQBvRgiP+kUJfJ1oUkBVS6R/dA9Z1pbcKK+OpULymqBoB
T/30sGYcOWY/0CqIzMTzv9a7lTJ3pupREH5U7zaEe8QeBy2kprHSl+8jd/V2idZG
aPcwQ35aLuijLyKQzujjOqH9hd+vODthLzUSda6QbjyEQpJZBADFhbHz+O/cZWpt
iYP6iY+Y8l3C0DldsSyfKfvRq53GxRt/61GQJqfvAKfjJ5ULdXE7ER66my7gWEib
3O4kBMy//iF5U4rDTgpXyD8ATj5LEX+ra3bAiO/pyLYCCz3Zn2ZBiwTS2ic62qZ4
zkZcaOH62/26AEgQo+DuN1al8TiGoIOfPGkeNPChbCgCMP/sTMf34nNfeglyE7nT
KAYuZWO616KMYXUR4NiSmuZ+HplBslHTj3XeWQQjjDMwCTkfoXXOop1NCcwH5gLc
uh60zpOD6sGgJstP4IUpikLkliCFAT3ixZGEVMWlkWBY7ZstYxJ6d5gS2OE3GS33
ImPrYo+xa8+bgLg+/20Gi9wKsP17JR/erV5eWZte/yahjvY8Pb8p+wOxZG2rvw3m
LNjNmsYLm5+BcllsGC1EkdicxQH1ZzfVzlqG8phionAqzKdLCbGgZG+K4/Lxydlu
Pm7HKxuLravxAumrF7FiXNvdmwORXJxkFq5FAVXeJf9fZi06MjP31OHIya1CyPGW
9uzOgIjha4SzS1s3Q8Dlg2tesJFfFvDwA/SiF/l1BcCUho3FjwCLPV4KtBjCsgQz
6T8UjT5jvS9muo1aaKFmZHSA5wWY5bMcQIw0pkpWwhR6vW0GmxLzCS2v4SKfZBnJ
kSGRMYXPsnBWh0qFrbVoyTuXpjSh3hdn/CaBKrrtKumphLnMgXi2gGDxiTJEyFk4
DHdIRqO2ThtfbHOtBBBbzoah13O7pnXeUJo4kWAG0S8DO0zKrAd01k9oHr68PDwK
KL61R88ATg7dHxEBkAp+hrZ9VJCXxWYsIaio0Avjw6Byw+yP9PIbk/fJfwDpaj0b
R2EObTmKfjVLFVy5ANFbH5cs396OdW1VbvLweZ2MZClRRUMThiguR+1Tb6gl0O4C
z2pkt9TcjcNGEuND20RCqvvsWoyHRhIr/hAUtuEn5r3Q2xgPx2gstVN/7LBrlFus
ekKIIU8c7eNsEVe2CsmpanFBFgVh7lBO8pbxygrZNsjL6xVKTxQv5ifIBDfkeK2T
cY+gE0a7xv6GF/l40dsZXRWs03k0d1As8M9W1UERwZo1SL7knqLDZj5/sYp6Ctfb
owGI1A75LCISHTyE0EVnflV7QmTIhOZ6PRPe6jKQOzzMoBqMZvjZiYCeXSuY4QRm
GLbPPaY2JN9+NDjzwQ6lAnUayr5iLsyNTMwuibYXXn4GNlwf3K4McATJ8Sis/VI/
b+VmEhK2k82K5YKTsEDpeE8Vvcpt9psBTmS9P86z3birCkGkRSznLzyo5HqZ8KUd
QmAGE+0p3X+EyVgZeGoczsvjmubuTpNIdWmmNHt9kQMAnJH3piSnydrPKlyOlMiV
YXjoVDrEuycGfW4aZSDnbttD4xuYeE5xwREbTgTSVrfQZBl//8+ltyp7JRPDf9ZY
H2xu1FJUmfj7tAfThIv74ah1MbQ4uy7hkbf3ZEKgHTbgXfoB5829nSBZ4c2SxSGB
E7rmPmZWKxfz9wkkQ7HvVF2ljICAnlSQ4zNoZBLAdz1+WFTgMu29x62b3lUbzFZ0
qfFqJdeAuvdGzeMhN7KvD6dd6wIOZitwakD4pM61Dbed2hv9JpKXY3JjCqvs+Til
Fu+i+Ti6RZ0+f8IECtGa360CYL4e9SgG+YIE00WvKgCEpA2tfQYp5QTEVCby7+ef
xmCs58GJARQgmW0sV0+eRIRak7ppt8masmKjR85Pk7399WsT71bQIciXkVW0q9ex
i284dIqYTTS6cYh6c+t3bHqJT/xhGvad0SCNw4MrQgyFjhrc/H63eg4FefsMdia2
VVSjuUFhcG1j9dchlPEjBFlj1snjao4TePh+/dmzWiSYWqYCCL/CL0GZ6HH6rdXJ
O/mkwdLUEBetE6Wy21RXjwmeaoA4Sa8Z51JiBhjprutImNitaKQ1/sNDkD6Hnc5T
/bqbcSE+eJZcnzBS56mZFTd1q5fN1MWPjGl4dJ++I0HBFGvTlIR2l+0F49Pidhqw
bRDn1Z/NUaovGP76zOL2J+Rc6bt3pGNGCGM2muYo1ss0lsS4IvpvtXs8ZG0eUSLj
5B/w7+E1wQ8kX0fol95YMDIXRYtH9/rSEjx8Kup/IFjZOS8rKEVZ5eju0WUQV3Mt
ixJ5wV8QgWsx7I95EsXcxcblVVxzQFIfncCLGi9xHZD+62p/FuA3iT3Uyh4tyfTv
CWQX4+aCKNgU9b7F95x+RA33TQzPVxGT5nPSxt4agGpKmXiNwbLGQ/KXEUSWdCHt
Lu/hwt2Xvn2HQ+67rFs+aHfrAZP8eB97bqJVaUUyhrKFD6fk+kNqiCgQCprR/YsN
AThBOwb9dHmAiZlprkN3g+0VhoMqRHlvWrsBLHjI37JQwAsQihIlxFV2GX8INOVp
TA1yGujIRywIcOQBBSCb0gXdLjNN8r3n6kf1H9fEZ6MuTribVLOunt/1FoLCdUR8
SN2SSQhddoTbbz1TP/X4GFvrFRcmgSQsC1pdnjz4jtqbrdVVP40fTOLl5LaQUjhI
vPq4S/79QzlXEqYTvNMqh5FVpYo5P+AJrA3OqRwPY9kN07CyLVlXQ0YZT0VUbrjc
yajqpwHvdvqzf424kaot/DQ1heNkU4ZBRrKDX5bVxqG1weR0cBndsTKvJJjyoo/F
bH5rgrAK1c64RQ2s24vcFjL4xLW3nvbJOisyPWcfcpQOuP/Q73A/EkrpYwKx5fJE
qjMH0ZJPc4VYbkjUgF9yAvJZ4Ea/5eI+a4kmn1NXPDVeUvHy9f5YiQjuF3t4RCk3
TCFyDbxWNDS4mkG64g+utkPb+4zR3s7SILZuQ1s3l1ANqWR+w1ucAzkEFiA3t6oB
Q21KLKqgT6prhu1tNhh4Z6Qdal+tttsLRC/S7m+kkq3q4IfpAH7ww6O4MHMVoSxy
H8V0ABCbIU3VwKTxv3HbtcRtkZ4Djx0KFr9GIxu0FV6MVP6yl2FD041ag3Kw/e4y
ITGLodnlGMA2A/VCJEz8DLuEAPI4dcdMoQvjH9SyKZV++hQT5RnpDNFsFZFM4DoR
TnX9GMc9t4g3MFoftwVN9oGIpKp3sHfRCIfmzFbR4j/8m0pk3A0sRsjzlasJVUcy
9S9xp8Av7WGpBIrbe4USNnwzV61kuC5MxCuz8aU/Cu7puxEqIaP4XD8K8hhNJjZF
NYGTquNGTWH+Auw7J++2q3sCNDGY27HvG6xsETTPXo62BAJ+B3xcZxsQpf2SaviO
1rVW/f6OLV71jh+VXePGS1Tu+UVapVlWlDWH9JJWt2GxJ6Q8kdWc2LZoivACMGFh
wR/wfnEdGaMnv8DOTiPI6Ar4hcyLlyM7VIjyAOTA7iVkePlJnRcrNhJxE0nNFQ2j
He2m9thnlK3cgE6P972HopyEeaRly9WhwMypS16vzZg/nenAGRd5bxgzM6rkjT9p
0zBt72zWH+WY5Gcb/pBVJUGuk1Ok1LkJY0Eo5fqtr1WUtK03oQEc1xKRzFZzWZn0
YZvCqNXcE2/NLjfra7BDqP1ZoYYWYV/BvVMygoAajB4DnAR9owkzeceU/I0U8x6S
weIj/iI7G2f7pME+JtpO1tkjvvBOIOIomazjgkdb9SVSUimawoDPeWN8pH8oF1FU
o6qdFXmFg1SSGF5RJZ35uBPo6uFuDFZAGgbYR7ehORSCRXMisjr225fO+vXCXCsD
6XzLeaSSkaWUKFC+t3jmcEnPp0tOWhlsNCIU3c/F6s5WtWyZGUw7Cn7Pgp53c8uD
E5i8TM2FikBdobysi/p+rM76XzlbQJZNs8p+8XGvXI8Y/E1hESDTaxQr96WYZbk4
B8VXB96pTSs6nwCKzW6yMWEKWZonvpqR3kKaWYu6wBnNujmVTlSKP8k4eSA12v3G
HQlXyBHagtAMtZYN6aM/4E9FoAMwRAhQzApT5rwbdK6WXtfAyUIyD6+3oGVncewE
sOxTyCIoDBkAtFR7BDRnY601akzugfYeT1UMNr6I8ebpQ4qmKDPxFZSlOHWHEPpW
h++3df/TL8St54Q6mnXpg4JekS71b0SFHknO0ZjuPKgVa7JTA+EeJsd2rMz5bMaW
lNyJljYNvFntoYv9x4QIQYAWdLzvq/3m0y4PcLlTeEiXLnaGE3/69sajDjCcikpw
LnAgffRtBLrIVyXXgspTSGa+9aW3fQ11ad7cpUiD2jqZWL2TSgxakkNTLeIPPCAs
jB9KGBcsLWKZm7929A01e81/VZIvng+Dg/dyqC4x+ptdaaA2uJJyBnNU0e4KlEf4
p0jtSmVgYbbYoMCz1Ror6afGTMY/se2PReS0g14Pa0eZV9Xfa7Qw1s+fX3u6USFi
Yx0+mn/3YZA6e4D1c3soAMoL9N7+Gm6kkPTJB3OZRKQ8OkXXfjFKIcU4IGvTYj3P
yq7Y4tk6hOp5yfxFetkg4q5OD8t1O4B0W6snBpICC+VzDlM60gpXqCq2gRfo7e1p
XMSZk7BfP6fXssXILgJcwP7JvSteH14alNSx3beGQbLniEsayt2VDK1Yb5x4gGif
etb4vNfRm/1fZ/lZx0W1RmXr5xU5a+9S1/GkznciQt06drktJw8qzKN57S58B/A5
ZhT4Yb5a6CO/qZ09XE+mKJQTX9Ygfa9ePNdiVsTNKYGe+NU4DoOPYHLq3EJ/1bxT
xz0vvSHOmdDmaCExbU8QJt33lwcS0kJ0rlhsRu1BoFK1t4hr055UE70WrWilE0eB
TjDFXP2Fsy6BQv4P33VZtKz05Clljugj3SLzR0jrWkQfFDb1N1LrkKehgSLjYkiM
sHhht1y/vd37bY1zYRthOp+DwfzNVquh/XVQ/lsIYhGr9R2CUz7/a7d0OkcEu3eO
466f/fATD8QF4A+UYEjyMsBcGTHgtqa+qTTm3vCX6Fr3VXGEypWxkP4EZshEWEE1
om0VDjC2eD3Z9oyApcVfMuQp5uVtkZFGdHKUL1IpfCNBe9rG6PrgwksE9V8dgzPy
kL1p7bltFL55Y2txvWw88uj+i6C1lHutKIKYvcyq6PCf5JX1pyfoxb5L4A75CYEI
u4yu0m1VBBXY5TSBIFPOtbU3Gr2si3qReN8m139+J45bEeeO2eQ8dzQtjohcvZIV
iTlfqdnbe2g6Yw5BTbOqeSBysbIGFHarEAXT37sKq34GMxAXkwLCwJhQQ6SEBi7s
e6O/R6loVaDXu6sSvpkjJ1I805MaobiQxLFBgK5NWd25RXBSmO0KWXxOQPVQ8rZe
O6f+nm8RNs9xlRaUZjkMcfu2kVquE7Rh/TL8kwGsByGcK5NfKyoYxmU98w+usTjG
z1RVuRY5/c2MVsOt9fLj4BYDEFt6RV1xif8NO8Unw1auqjm+Y1x7l/Rh4irHVQkp
yO/NFqF7JTTDnSn4IYarxPZR3popWI+8A0XuQ+WMdp0WMTIpDicu+v8OmbmiUwS2
9r67gfwZweQkKtVnZAiWVESJwYy2FjXDXJhpE64R3GB8hs7sF/vXlOILlY9jTE0/
gZzj9M9UYOhybzu/lslimxTUuQKUlqymnxeoXljiQ2R1HFAfDcHSt6ONJWFM8jbo
mIIMmOd37FSilKS5TCopu0ve/Oa2E1/dkPt+pkBSg7jTQn2BU69//SP3f4WNhNCQ
79OskzwQD+fNBmp9Q5j38joB6+rQcyBH3jxpKBQCu2Qjy8cqd8GQA2Iv373OEFeG
bNff1IMVeyJB+i5l/OeNrkbvRcsrdUrwtV901OZA6AnwtZiLCpn9V77lN7a/RV8d
7PW2aDqsWlVpwndiSXUrcIGyMwWdu21BaOV44MSY5J5+u8io+GE2kqoeubyd1t0x
R8fPdNZRW/CTORp6jx1LjHn08btZzeL5vN+fak0POrrl3W7hZ8Ae+C++cGFs0bEb
6IFUoVEksZvhubQywHQaAgXKdSox6HRH8DSE8j4fMljLi1DL+46rdjYL8Ke4hKa+
hra4RD/UTy0jcO8hhf6tlSRKa0D+/nTyWdGNBYwlyZKFFcI1HXKxYDUEqDvJcwu3
P+kbpJzbK/T/wLFo8/v2IagIfahX9/PIRT2ksXGJeUNjQB0werpMVAVxy8orkUL/
nvBDzisH6UHehXl9w26iyZsi9iBj5Q2nXugvXFEWfa+L/SZj+2PgFC1egP5Lravy
i6n2Mgq8QIwGywp1oBkE3358NxTnehAOIH1bQOHL5kJMk2LGHHiX/miC44BMSKk0
cGeFAfohzaXAa/1olHZ/fzejBUYrcNJHKotG/ne6YbjfPUgOFIlfrHBtF2mbgsY3
hamNhVC9BkM8RkEX7HyGLlmPa0VlOmJtTjAL5t+vnWAL+QAWvZqdtGEhJ+DIa2Jn
fq3kPzNxSOVyhTWklc9mPKcQ09JsgJHXD5gdIx3sc823KQRJJTA/BkmOncxKrA+4
hhDNrxFmkwnJPdWPvUm8038Bv3EKGRyl9My7fjf1wB01csA5Asqn4wV6Auk04ftV
PvCnQkwLgevk9KW8SpgNp1t8nhrtHnHIrdHUm7NpefQmgzWLK2m1u6fTCaMHzZCf
P70FialhQS+oGHfo2dRTaSlgKOoj2LUWKaPwK1Vys5M+xcOdPVXWhJIZ/KAb8sRT
ZQDCbZdl/OqcqdMmi7e0iInP4pOV8eycEQy+fSGaVBofbNejJfEkTbK7Ej2+mObd
iMRialBK8debMRZX0t0LCa5OvsrIxPXIswnQ7Z9tCqwAhWQWFz1JSt0g6I9LkdkS
Z8W/Ily5nQS3IJ+8mauraII1mGpUISQFWSlkqxQtgoTQnT0OPLlY9QxvdwvRmwU+
i59CXy0LLOJpjFF9ykbr3ZvERyYtYSlL5O34IclPVpnlcPOWIISL3BXG5lX9ZhDU
3gH9Z5iCGgzQNP/LmN77xk4Cq7JErV21W9ypJQyAVhUFzDOORYXyy2LdW7WoOZhJ
Mg54YxlRrrUPdKtwB9mSZzNjV/aNeomwQJ1wJlrhpULFOuzuUAY3G3fWg1UApIdw
A8xLAeyYORWN0KxQJrSoBxs5nafjXOWiqbCmwEjABxSFO2ZuTXAyW/ClIbw+q99h
7nmNz8jSpz/40GY1eDMr3lqoC9fuUEI4TXHAJAn0vZxHrznHnNNZ+oxwtAuzlkJP
5fhyz3nVOxxX5vG5MZyNtgLiY+GC+iExW8UXJDo76qIpwKwUv5iUXElNA5eUcxTz
HJ0E7WfVe9QY8v5VKOYc2tbEaT1hBPELhzywqZlpn72VYGFDfO7g0Sz96hQvtp1O
tGzBCwekFqiUm7QzStruwTsZqUPETKpUkqvaa3cyIW2lv+TnCv7kgYYVOpwFm9mP
OhbBI/jmd0/Fp4CQ+entKNr7iQt2fcaCsFxWSCLMpz19kKiALYDjQPc5RA0N5EtP
mKWGWmhFUPL8EnApmUR5Ee8dxs66QR5KHRlyBe0xvZoQBxFnuX6vDICQn9qhuD53
xFXpCZRyWXIDIaE7ftotjw1/jtJBxPzVvh1ktmhD/GOQfewlOLTi4D6zK27ySE/3
wTcWmU8QJJiGFHpMxieShiXyEg2zAkAL/EEdUk7Or5O1mdRmeZGtojyD7vIYr6ZF
H12zWiJ4myzk7v9LIc7DvAfK1TBkcEXVIPzLVX9s8voXtTp77ZhmH0a2yYGTnXtu
oEcfAMzRpGOL2MyvDWPGttLI85CmqnfxoUFw60Mr+e/ZoDWYj9QVXxSZGy978M9/
DjcwCJDi8McYmVItYPsjRctYWJOonxg7p3USOQGiWq4SLM1+OvSXL/S9OzKrokHo
ag8E2Hu5fhJOg53c0DhSD9kTfcSqGa/rqWiY1i68g0OblHi+dmRAjwOfEzMAdcsi
SQwMJkVWvvwck5dXRJLhIRftwwGjD7FXZGYw0PGsUup9KKx60sl7hqkCIUL5/F4p
AeC6GehMnel3Zi7jm8DYTR93GX4ctMRhpgKTKibrW+LjcvzvojdUHwlGNcjCT0wA
6e9NfkfQMFw7F4nnkU18qmjZbL+85MY+JRG0SAXMZOvlE5Mg8IQx+IrQ6XDjwhJq
uu2SC8KJLR3+/P9HfiN7KTo+tZp0WAFPh1HZFsdAsnMPztqgN4KJPZTusdD55eB1
0Zre5aKTzrLWHz1zXmDutyGWrYbe8DSuUXcZ4ElgH539wW9Bb0CpakMGOdSj6CIn
I1As3oAeGgdP9TjDuT9WpoxeC5WdTI//wOA8sa13LX92BbNHMYhavPD8mT77ac86
G/RLobs7nqGekTH3OYqBgoewcXsWz3C3dMe7DDJ6sl0XGTAYFVMow3d2dDoi3xTd
g1oJC3jvfXuSgSZ/GF5/5Eh0MCVECZsMvhkF0i5veC/zye67q2X+iaCTB5sbOysm
sNIJRimgj+38z182lHAG8qN+Utz1J6yJ15SsyXHZ/LgLz2We9BzU5WdRz8wzEzlJ
9eFRjRujTkZnS5P/lE2mXqPhs5vRuRD70OYxNswK4M5ovAD/pjaXAcOr9ZYe55tp
sNvNxWGUle6rPz+JO5KR/w3JUeDOo8RXdQ/qgmHQx2eISInmHgH7WYKwRabxVOXg
/8aqnZzUa5AEuQQpVdvDQmz23ZKkrzd2ISY3eBMtUhzeVwk2pSIqNjcc/SEI9nG8
Li/NuQCw/Ye5PvwimzBjSWLPTVkgu87kYhPTia/cuydN2FJoZSirHaaQKEZg9TqX
z7l1kLeYpqsymCP0z+7fzIGBkWhz2wzMiu0puNAUGEP7xgzza9NA/uk9cmObnQZS
Gvo+kvbBmIk3nDmsmF8ox4M/jlfD4UzjYSaudm5+oL+DwURRUwdxWBDJg5eW9C6h
diDNb5eGkzqQsqBZgIXtuIXEtR42tdahhPmufLSk5ghyA3QsWpOHAovCezoLoMtk
K8K70fOOfRBNc4Cf8+NKBiS8HAo7fpW6tIZFfLTxJyPbGMXON0sv0z53CcdJznEN
TD5OuVG36VjKtrEd43zglL8Q/QVPfvVdS0dQjzl2g/JLtqMTAD0o44tjmmVp44W8
Ga4p9X2dtsGQPPOYGe/JxywIx9Y1vtuBAlLFpRpym1h8TIqO7H/oOeO+O66FLzfX
1Gbs9Y4x+eDoUTtikAVMmnUmICZAzuROPQSS0I2Fse+VpYFlnT597mF9405XfXLt
he/deumYJXt9FUCha9sQ4ULISGnMeDc9twQhc4NwKfDtoPpxYsXW1+6psB1m1dhz
k1F+v+j3sLdlT4S1GEepmp5WGCfQ8rlvORsUO4WzpTvCOeoeXxPoh7OB8JEj8V/B
ro+D3DZOBkr5adQ5UaHhCUfuhmqT33bJI6+MUEAhX5fJ6guHLBBr/IQeS53n5dXr
Gs9kDYgCLMyxF9XrIk0Bwu8OJRmQu+Ms0fAoHmE47Bi+IGULUbCa6W9UQb3F8tBS
IAD0dwZlrAVvtwZXjuPLG6CxgRtxsxjRylBNep2j489GAm8ZSj4LL9Jn/dlwGRs/
8FXXC1rcLO665L5uxi5lpCq3dDU897mosozupLvNpY52b7bPtugyjW1iG9aPPKq/
QD+ZkaQVJSY1lkU9XI0BJZpwJL4aV4bwYLD0RFiDIpFtTsCoOGDww8O7TTXL0S8P
q12SVQ9vQ4bPDKFEQ1MSXA+Eeguo2DJIX6BCm+zY7i/enerBL3BMtyoUbQD7t+Tv
m2heevEASjx/bfGpJmD3EFm8kf0jzvwOli/62B+3wqX6m3LtaKU9uxfjFSXiac8g
VAKad4aVaiGNcHqBt1YlaCaMF1GBVmv23ND2QcwclDafHYIV/qysUzGciCn/NNDU
ryYGSYdKx5bnc9kQEkrWaAy1IBL/cVw9uc/JqOHsi3x833SIJM1OOrzMekLii05x
DCa4zUKFWLHK2VVAZ4wHpgnJicsAvn7XvAL97LBNIJl2jJD+y29+xRMaewEacVvk
wuiCtxcTuPecrktuklA4GlpiblllAaIPWSdqMdbimoSKnNDwFt0M2EAIiMkVtvr9
i7W5GsMbGTb51Ye62TV3jYK0F04rBOPuWKtaV7esHzdduOJF2jngbZ0dxvqVnph2
k7NC9V+Q/gbZVmzva/on/hNtcvDuibac+N9ResWVhqQ2CUwJU/A02QZ0pWEWAWid
utZBxfglZ2Dkb7Skmq45u4OH8HGTRJtbvqLPqkB9Dhm8ArrE0jurHsSgGnSJSjd2
1fBMmUKGdTr6tE8tTowvvLE9YCy4wrxZtd/KeIwJJF5mACuJDDc/cihu0N2PLCx1
mVg1fbxzMfv/6w3JJtt2YZpg3zi7xXibLr7cmai3juKVsmeZrUMQggjF131Scz0i
HfT9SkbNx1RS5juMAq2+00RpIww/Q2U77/wFyXGKeO0wuyfB/zkhHuH1fhOcNWML
FOM6uV/GeGeUIWM70amvgHLCu+gXKNkQplDlBvwwZGLgWAJUVMkxA8hI7e1dEj3I
UBAtVnLMCh0mx76A1O7OWb0RbbD4XPi6LFig8pdcIVysNlqc7avhtAkOrzsAUiI6
X7nmN/V4DTc1cQtRlf+KPJjfcMMcoHjapM1rrYNip4BMCL9e9mDekNW8OqeF09lA
CIWry/TmVMSeDDthpJgF34efCAfEdvByYtlomndU5Tl8el3+cyuUBiTLBqPh5eYc
4pRtwhGUne1oEfQv5x56BR1FUzyZVe5LMc9MTeoC3vU7LGPy3O39nojxqZcrbxqk
MgGcrDfQFt+Se5zEqrEgDJvRurC4HdTfvqJKu9rSj+U8sjuA4BgdqHi1QZ7LkkSV
fD23WfvaWyKFBu1mPqyZpiKgIVaDfEo9JtMbpZcvZTFsrEWf7zdprxAWUQEwaVDH
f0RUjp7ltqQmWV2uEZNLRZde2Usmoz4zCAHe4PK+7+ee7lqd2cVujVd9b2ZRd9ir
jvKgwGJm/S9r8kumOlSktcsDSDy3qrpXdcGeAKGFIxAK5C/2MEBpI2XreHWRBX2U
Rh4XvGPp7AmzW0O3hdc62XtiFldgREL8AG4xdG02x24RCAC1VsCSvtlZhOUkTiLq
GkIHqeiErdAhEJrlkvrYG2vNFqExM1fj3zKKi3R3Y5VCHvYdVdVLDBn0ZqL2t0NS
KKQXskldubbNxMPnsVoAsqrKpzm15i6UYAX20fgwGk1d8ui3qFhqiqVi9HDjlPKn
96fveV6y12oROONFN6+AYTDSuTpMqCAu++0ISPa7lMhqNcjSh7uXndps6nWSNyie
/0uBhbvGJG2PHh1l7RjZ6OP+IzTpCgWSNtUMrp5pMZMg9EsRQX1ZfrjY+rrsaYgm
GyKnW/6WAPHir5uaV6lyrTL5ju6mAwhdWOfoY0rpEQu3oyqYvYp3pWVdVH7hnSu2
zaQsDE30uGzV47c125QGyHrHFWP9uUFjb2SbA3ar0Wc0yi+tqmV0O4Nt99ECKKNX
ZVYsQnqryUegOZ7r2d2MNTOl0pEeVmmedEIhhew9ojzyK+0nP1ke5TF2JvCWkcde
SVMty23lbm01ntqTVBwXWszKAN2M2YCEI3kzC2266dpY9v0ThGoPM3ftTWyqdov5
SUK5BMKG1SY0fZP58oGe3UiA/BtyUEAthNxekf1n86PCQ+SheoGB/ZZ2CwtTSCWS
KBlKAeGe8UMmTnShgKMXb92MHOGDhswn1ysjn7QqnAuE2iUwWE9nIHvB57fL1rDA
HbvT8Hzxhd3m4stOr81vZJw7SXUEyX0HcKh5/BZeEnxnNWStaPs54tN7wvRNf4oE
XaU3fOxxJjmu0akHeF/UavUEIOON476q8+/UHD41uwvnqJHj6gTlZveUc8wiMn2L
C42GYz8Ua8I3/6p/Ek9pRe7Fq2eMTVxdzJPMyZ2Wpb40Ksr5snskrF2spSYuGYP0
G3qM0fGOVHvxD0qCi1d6jdOnXOQ5oNT71YyPN8Tgj/D9ARsGSjEkVqt1tDtxlb6r
+HkPE3PgqKNBE4S+u31hy8nZ0qLQyMa4qiCFFoWxRPVCYMpvGYI0BhowOMRMDUsa
4cn7/kivEHCi0RXJbtmyUq46CxdChArI0Zd+BQiDL+E9hRqKj1pT8Ax7poANOsXt
RPyUe6UkmZs3vPUr588EpXIRcOgyKvHVdeitbUbz0Yuj48QkRsUOyLJtvH29DWoz
/+TZ+22bkf0s1eG4epLFexYdnzu7Z0VxmqwExC8XlyiH93tOoBCF+S0ftu2yVLcE
hpSQRMjuvSm8fP8WUevidZmpCHQv3rlr1nNTHiaSjnWhGHKXppMqzOG4ERX1rjTa
1XW9jv2gjE4GOzF80HeDfAzV8YY/NsA0PxkEvW2+ZNsASUE3+PoIhcv6d22yplVo
Jh/606am7Zpe3ZeYjzlEdZmAE57UFJp8U2ibQlLOC//VG9BSDK2Pn/ATj60aSP2R
+glRJExgrQAEEgClKERD1kY/cNjbVEW1RzDPwoc3M0fO7UONtYkHsJIYXHk6GcDZ
3bV6l9ukcQpivOGYHj9qBVn1QjE+xIrFuZBcZ+G3nieIhfNCCBI6XAtym3sEddTZ
w7+/1ehWZRKzPE1a3wq3KTjrY8QMVR4IHINiqUfN90p6Txphz4Kp4KiKyZ0uSPIO
KV9p7GJ6nzRT3AmlkP09UWHnUT4Bd7VxWuXLBMZS0x7XzNnu62NsOB1ezzJnsbxQ
bE3rapfHgv/qiIqPrqhXtt+MN2ntPNatQuEi82Zalb+FGqpqIKsqrOyCmWr5ogtr
T2wWEiJqiBEAvFH+O3ALkIw6wI1pxy9nxXZ70KUyZhr9e1i/QdmPrUXfmApGnvcW
AMUqGXFk16zwouPEn+KZFL62ZoS4ro/nbcnGJ9Gu+fj1lsILlxgefMvdwUzXnniP
M7JmWe7Ou+VqWjLNs5+jJAhGQxiuvjH4oQZy42On+cbPTg11lar+CdTjas9K1HN4
PHTzZd5Tneq8LVwOXJ/RNa58nIW/VTc3q1UBoP5BZvvtV0bBIG1S9q+/9GukIuul
7YYZ/L23Nq3D6hwfW887kioHBAtJ8HO/5MpgMlwyxr0dqOb1vB/MBvWeI4ydZIbr
KmIFsunVPtUK0RK5mSMLjdSlweaWTNrh7Kl3XgxQf+rRUdMJloV7soYXI7CsRffP
hfF9ED0DNHtsaE6BHXrkdQfgbhr0OpwcKV3sVQrcbosevofw8bjYgFhcrLK6ZhnC
uHEyua0Vth9JHSGauBwnoDc2LuDjGjsAWDSOvY0u5/CBD+86XCqvLIc6GRtslqEG
zviHkId9T4OF5Q6akZtXQVCiBIjtULHCDDOU9F0HrDp7kgDNgJzH+BDBFRe9oHrF
Jy8JIeVHeJOIRCHvFwSrQRnHcXHdap82iBcc3Dkvw3j3XPRsJmSashtCU12zoOWh
zqLXB7tFTwSyFqGqayG8NMLMIkFfA8/phqk9pUIxMPYXzSSbwnFz72UOnrzUBwUg
sjvYIRB7VgTD7CzM3uyZtFOv7dutQ97DIGtg4AkT/HrfmViT2wSg+qBLnw0Xk5Ok
Jdd570uh0Px5VtOywQoG11uBLC6UYbjFXxGgbgy6OkBUtygvA+YkRLANdchAoEr4
vmHy58+tZM89nDvsZeybYl7NP3v1N4YJxgPaunGvsJQaKZZGIH9aA4iE5UQ42fLL
UbyjgcsoIjN8xwEP06QnTk7XLX5T4xwNq/hPS8r0P49Xu+z/FxUHUohp/4ZngDDj
hMG+aqfdL64yjxW9rUf/h8+UIzB78WW2DIduwg38rtRk7GbsYORLntxOM96V3yPU
yDOSmC48ujPA6FRdQdvPgNEuPvM0tV84hHsIzvkWeT7kXPnqv+5yjdW+4fnYP1hs
fiSXuGqDb+Z2r30bhKT6aur8Dg9mRba/5/Iqza7+Ut3dlnsUFQYb/WBiO7Agccm/
khqs+C80UgESBrjzhXW7MYahgFIZDaI3x/31s4sW0mcxOKjQwECWk2O5synZrWy4
jrwksKlAUOFDKcqeh6rohIZTrFgtI+8O5giKfAJWIk0zuDrMrGVtMdrzbPGvRP2h
h7Tw3UxdiYQaYNgtvOaHA5DkiUWzwj0iuMPtVsjLpN4fuWU7/rZEseAmqgkJXErt
oJ4wfbHVOez6scDWaUfoUhg4BE83eunHg84t3HrmuAFYetfR6MfFsW/RR1MU5soG
nKFkujMtKU9dOystFdyaVRfpluZvIOBTRGAM3qo7h+AUL4KbBq+kzJ2am/30xPxF
k0pxYUtlAOIivS9YikmLlid3aSnIp9g7+TBzY79fIr4+lPGWDCStiMUcJwkdmlS9
JuJJQXSgvIsoEJReSHGVYaUS0rSJsUl7f3erSf7elHBSccek494w7S7mLvgrQPgv
9ccP2LllxpdDdEogsZRLQRchWFbaAtmi8i2SXPsS06DWv70PY3BswtEhnt/z+b+r
9wRWQ5j5S5st6p9pDpS2ui0CTqZ+Try6yF6MTF2Df8KQOv92bY090wujndrdxbga
3bh1gj4iL8pUnStA8HGNUFHCFRSHY7XTxSKfIo5FK/d6QMB5G3OntB/rLeOLA5P8
qEMiQDc0ZvRR8Fo44ila9ml82LB6myp3RhmkRlXOEMMsl40if+gNsJlfaZFbDOmk
J3Vmy5efyq7LqqVucxY8t6JLbFmuucbrKFllGq5o0p6xkyLAaSMtdPXNaEt6rJqP
5H84FYbUalwo039rbAITX5yCGV0saH8df7gxJf+a/9IiNCwOd04/cHg32qsFzFqT
a8Qo40s1gmnggbpQwVS6PGuER5GMBFgN0Ux+grZFG4dLxMAYEKs4fwzIi4AFw311
3qe5CrGunMPih2m/3yT5Qt9rtNe/4Iy6tMRtjmWZtVdy7nb2HooYl60jvjCWarSh
43WfLpW2k2cXsBioFjTZvyRdivP5ae99lG64brQejAH/UjHgXk0VAlZ7u/mFL6Zf
INs5rkfyhFlLfMHLWhMo75b4JoVitwiauOHXdPOQ+49ieRKozmCc3JdzEO5HlxUS
Nr2ifwtWK965sGwVeQh9aeOg/65AGlnNoN0Kaw3a/AF53LOQ2KtEIPZm67+gMFK0
N4E7ANMbGUoQmB/OoblylWFc4WUYV5HkHvg530AC6ePLsD57INh/vqgh/Wj0gS5p
cemV5FqB3KsCeCeztW6l9UOlK77jf/Xfl/jlGrMk22rfVorByIMpJTZb7dXNIsgc
a1D9rAT/AlPFTPpUULGr4+lntGeKmx8a/0YfhxvD11Hg/6K2BUmsNPwRzbBsiw15
8oKyXFCFpbWXVPk4fp9PP5mnsR9K6UPnG/oiEI83knRLOV5GnabPstyod3Cc4Rix
v+wOtPKTLC7UKuWwSK8NKM6p/f44/Yk8Rx+nrha3gMN76VoUaiaY2aLV49RzD5Ol
B3eXbnv1m9sjC8yZ9E/L20QFlO35PTuiP2MwbEoPVEIvpecubFRbcbE/OPzA5Bbx
UClxSKl+3rA97OgUyC5/quyBtpTH6haj1D4asuqQs158FORkCvIkE658jZ1gaKoF
i4kGmUyU3+ez0GilXlC6D8em/TAnIbH+dI3ZegZmDMX6mrBfIJKnpKKhUFWiABhg
njrOFxH9Nb2/tl1PqFrtsgMHdZP2nqFSLtPczIsOZoz/Fv/wVnQSkbTKN7hdsouY
oniKe+dnR2ZvkQRRUZzjCZnYlmF7+xeorNvZpaBxnPgaXXoQD5U16kK2HqPPPSzH
ZmkQFURl+59IPZEDp5lKho5mDJvlnzAg4c/hrlTZGEiGAtsdqzopSSmXyXfKhOLB
teqjZZhaBhKfQSYzyccIKo75ky7MxWRo4eV0mvr6TjfDBvfZR2TWCXnn/fLa4two
2d7liybBVD7XaXMAxE6PPilPyWyH5FD2SSJeGqEVBiduA5jzme2AY5sjlFB7hpix
TWO/LuyNVRNIJyN4zugRuZTmDH6zSeulmgJTClUQ0BimKEwuvOEbFMEVOgirqTgY
6Cn9kWGlt9mJeVczE9eSdsIsl6eYJdCroCZEqWcsul3ClAvU3SckYUSL8bl07tZs
b5Z88tvoTJq7Gz2HbjATMPJYLasCyZpBR7UlgVigdE+2cGr2nm4XhkKZxAwcwFLo
qOc3ZDLD/jpS/9lgvAJZ8dF7+1yoLRgxlpVk7OAKThY7cghPTvLQV86Gn4YHE6db
P+YJFloHssVFUIo00gB6eE6XHmjVtegq7nqiztaFLybCChnceQERvEMFbOsPTTzl
AdnElGrT7qFrniFZal7YUrMq9cOli3E8TagpKnygBrpxQ67tzO02eRGjDjvEySUm
aGFKg659fYboZs+siha8ouVqXWuVXA4tP1bCtSJSsBA2vFqSM4074g6Q5o1mUI8+
sTv/gXuc8JX2nSl0fmB4g906XsJLLYr6HluVVh2zcTjxcWdO3MjND462TWDgSE9T
aLPKRo7vUvriU9e5bcKfNKTnGfOv4D4NyFebdytaOyddkSfg3Opvktmzh/0Ipt/Z
JZZ1+x9xKd2BYCejil5NDZlAYFGJkU5CkjT8DCCoAIQhNj05o+EM20p+HHn85gyJ
M/ZZt0EczSZBsHsqaYgdb1xZaG7z5W+CCH8pjsSZQgri5pASu3jhywOlFDWOhWbt
F6uv59TrG9Zwc2nfwcZ8Ez2u71dOvaI63CyHsaDIWSaTehYcNOrHg1sO0142K73C
iIUYUY+FyDbdDasHeWCmY7MFLebQSl/hdd6ivRASxoOt14ua66g7INdPGCkgBeUc
lF9/FCWbQlaeh3Uvv5x5SusbgJhx6oZ9WVypaVA0YhS7SVfXpzmWD45ItZoSCnoJ
iwa7A7mbjSArRp66fp+Riw21qjg7FDdaOtEvbQotP2sThP3XmlVig2Bzbv/L8sam
t4z8a+KxlTVQhfcidNAJVGvF0whSoaU4FOuO8cdQF3kv7TleChyRQCiWmZh2Io9E
g8ki59WJzjd2SgVY0EolT2K4ZLZL+QARspaCk2TEdjJRwpUEDCRMVWbfmFRix3Hz
dmqojsOlgVxpzbbF1Iy7VyqiayVjgdmrqMY4KEP9LcO/L/NIaZmjuc8h6FQSAb9y
HuP8wrZGEws5YW/gh9WjhZfc7g6e5zAQ+/v6f+jr3EjtxRBb36ZG0ONfFyTIHE+k
t9U9IhlX3LVxqO+Peqtl9vzY1Fk5/j+ye+Zpzk4rph9kZArJhHfUCXp8jXSWxnqV
kfptQI5+i2CQin4j2Q16kCgGvUpWvpCsjnMu9N+yjbs+Arh9/KMyfG5z2sxP3528
lvFzM1qVLO2LqpikU8VHk1tIC58aNajjwviRBiE3DorbmwJ/hZxfbVQkS/ZdpryN
KAFEtux9FEdKmf7nyGZhdltdFe3aKTfq5hYRfizB3mylLrdHMo89SWeh14eJjHjp
v0j9F4PgZQ6XMnYDmfs3JIUEFaHGGwMPbDKq/9JZQTV9PGtZT3YlSHSudN3B/TWq
gSSOouSZoT8hWfYZjZyPNGBq4kmk/R9y8s4wY9TcSJo711P9IRcmcqbSbHp1AS7z
oiXRA0RFXnyZzgdtEB1+U8sce4FF/7Gn5KR6+q3BKyuKtjmCv8EqIjwSajFkX0X/
8tEzKRpfap2rt5MEeHYraJRbkhOkyOIJKra9kUr0nYgED337qHitfJFLVtAqu1O6
v5fha3eyLIJkNz9SIvBnBf+CajQB2jItoufotzE0QzZkaizkV40KaXf+TBwhXj1G
/Afl45Oze4Fq3GEjrqtTBGoWXgwa/V14YoptU7YnNAAWkYRoOrwgAQsAGOo3G5e4
Zl2skpwcVXEAkdKnwL7OMqPPqs/3bi1CUA/p5BvRN3yzwiOnsYP5hFbpJydd42UB
pjNvIQt6WamlQAw0OWpqqUUpxqcLyL0uo/yvQTCCnH7+csQmhPq2zViKzMXLaAx6
+tihAybJESTOoLD/VlwLgYAL5CK5um+p6Lou0x04ZqJV1Pwg8tXty75os3fSBfPx
new8OSdKsaXHDe5mTJRhKKxRhNAQFAAKRicgFpPWNu5YbGN8FyeTypoTZ5ctAeqP
b74EMOiC/BogC31oPaNh/XHMuCbFLq5PSx1UWIXkahEdURy68R3yk7XDHqe7kaPO
KOd9ZN+r6mEdVqpa7gTq+fo6ed3E/cXt5b9JJCV8dvyJyO2kSnVIEQrgL49YGAcE
OFhLtRkkH854jR9Z6k7HIbVuYyKEu5g3C+ShNb1BeculDT/2lWInZmFuzdogbdWX
rKhc17ODsIwF2Oz26Ws8j41/8YJz3jM4x1cfJHrVAbaVvIF5yAmN4ZfPWnpEvRJO
nW6onOH92M1L9ZOg2WqCFwXjbII0QDJc1UKl9/uRIgHkz0iMm3uOD7jzCYomZ7P5
6Zs44so1zFAsrh0cifw14ppVOAyTbmV7SeFZ2hD8+uwDawgxncfWDkM6YW/FOkaM
Nm1ZLo2TB3Z0+TF3fXtqh09tV8hqr/mwo7d9FyUvcYZP2J6txLNeEtswfvPVPXSb
l1kG4flgxyCvfy431GGmgtM9s7nz1SeSzN2F7M/hyddnRWTc2lszIZtxamGjjHuA
e0pTfDtdfYeOwFMm8dluwqxYku4NjMILFrrYk46awvPnSmPfR4YvOjY+dVuX48sx
7Wb0irDiSLxFRcqw1dgVEu4UDG9HiRlOWtepXwb3DPwubFwv07K+3HsZze7YzT90
AmQmQrYixalSad8+9BgepmMbEd15p1jf44OH2fLRkpyPGSKsCnz6Xw2N1fKe68EC
sXnZ0y1qejKPABXbGcigxRPp9ZHColGC9CYprK7N2JS8VUKe1ECtAcG5RKyAXDAp
rIUpMy0Wgg9gSAKCugCfXiyUyJw3be8+s+nosQmoubO1lHGwbZlt4INF/SxJ857+
FF0Zayne5AcBqnmFBzyiJ9TIYUW8M6WKxfzbYd7+hnNIn1nsMCxMgA8vCwE+U/AA
8BVUp8TzBLZTQApPLfnEoeCes/Zh/ncsBpLL3ya4Nm+koBm3Srmr7qEk7cdABT0z
cNAIw63+ZZ29E6WVrBXOikqSg1wkdQogEMrzN/PjWhddvMN5y4g4bQf+3tAD7vr/
o5m2HB05w+0B5Uqwsix+4k3MKjWmN/vAx3pP6eqCnFPN90x5Pskf6rS9f/pV7Yok
EXrZ6evxkQwBWCBi/Y4Yb93/rZq5vy806l+UWrr88pQdN4QIGfAZHVQM99+ybG/x
Qe0x+gxoL2FZQWoLpyYCxkQSqs7ENwxN/O+7zdCRbFv3z1fH5q1lsSKlxLZ8gml4
8o1KVIc5NBr1ZethosVNt5l+U2BROzGZj7cBXldkU3AgmQvH6QKVQPsijB0/NqFg
OwJn8q5EoP1bKCxAYdW2iDQ+2nd2MZGbkJ2L8903sZx+2uKPNXkl6lNCK/Fvw0tF
a+3oEoHQ5mNMgBJ3vmLq9O57EOQ0dcp7v/R/9JZ/OCaEfd7FR09ycQQoNXy5+OzW
VN1MDJFTVjTmYrbtnjANtaw6uD0y/2/TK+09m5NmYvvtguBDVB5uIwfdrqliNZ5V
qB2P0aQRn9FUBXFktOT4UfnT/TMTmacFSR/XXL2aFLp6VkBjmyrTmF5uy6+v8e+K
3EyGhFdNGMD9LS/AgFvDuHdxEET7u3Ti8/hxsOVnFUvuQ1lqcigFYbGetFXdhtve
TPrVxKWMYjM1UGp/MRAyP2fNthUOtFSyy9nZJKBXlgFTLrsazJXqlPXrj9xOhK19
YZbvFor5y50Ktwqw90CZ0XjjfWVNuHTUTkodH0yU+DnD36fNUsC/4HF7Hl9UJPbL
nbfyDdUfpJ1SpbtoADqJ5OW6Jih+cvW0ZP39QQ9Oe3koAUhTI048N65ChYFqRRhH
tcbXeLm95Y49ucpAc4LGhHh71CdjIs9U0UYbE4ESaP7mRwJjr4msM+A+SF+HHdeX
Ywc2byhS6KTpfG6FjjI4Wdd3b8QYsFk25irTQW7ivV6dNKIkGfctfHWta26scrbK
c0HA31PukSN8yQWp4NjEK+b+KA0ogiG8ytWDA3ncNUWHFjw1zo62jTBV4mRED6bW
Pfw7iAZhLqllUMT6hU80xob9VLVpV8WEjkdL4vevD10PMun2RaptR5SKdn9QNRFh
frt59q7/jkHukHJnNZzVfIsDPOT9U71k099SunOh4axlkA4kXM4SSEnNtMBg5VjQ
ExXa1eiwYsGjgIch9/wHAo0Zs0aTcFH/A5WR0VNY29bpfNC1xhyfZt9mncxihb+G
LkK/k55DuicAbKCkaTd5xPcKMvurZuXnSQTsTVRtsO5FWJHQ5X4B01pNYNZWifJe
ru1FQoYpdmbWceK53V9uY7CIVDKdES0x+1d+CiSyEkbogHFSQOBJ4vUNBTJFiC1F
y7lSqtl5Vnoy6nUy5u63zPyQwzs0XjOrgiZLv/I05u3pgiz6mz/cTA5pmnr4NSxu
2VfcgjjI4fxMX3Nus5MlHTobhxK0qsabuOALHm9o/wwLyPgEqrR6Lf+T3D17e2+y
Bie57wECwYD7indFsXIC6L+bbYm6JLrYcvd8rPAAiOhsGgh5Fk3D/mc/dY5gx8aQ
o6xhnZGhRONVQw4VfntrghlZxoj34CAnAGWEey2hZPwESvogExDptvaxjtYX+FKZ
AeMkxrVtP7i1CDf1EmJRYf9VZ/AiBeqvW80GfQyCLWEXGQ+moz5d1x6yeSWfC599
v9KKEzfVuy8nzhij+RWVRs0Iij7PT0Rgt4wQHZPh6l8ILpOyUkJz096eEsoNYzXH
JvC1Z2KYbHaAaBVcbQ2bqhxCQAdJreUFb7UqxMN7auXZOglmg+rFOYZpk2A0UrmF
l+GitcLksLdgVxozKHmjcgWrzEw1nLK8Ir5LRC/ZsChQ/Nm7vB9UMNNyy9aQoJpN
VGBicyJ5G7vsXPyVG3gHpO9kW5li53rMK9z5QhLV0B/vq48wG+8HHm6/xcMZvL5V
V2q1xKdIchsLxOCcivCONOWzP0VM83AEJ61jCXQ5FuCViUKYH84KjKezMdBSNREN
H8qJKgE7om6ud9iIM7SnYIgFvQeQXaQ4doFb3SqFtAWe3rbXmE8/rwAS0w7h09Au
hWaMAwqZJFejRbTHI1UXKl6N2TgnKphMmdLg/M+yKjrIZoxgv7YcL4KNQLkE176p
tqrAWHGHvGB0AqU779aGZVTHOjn8HWJ+Fzsv/OqvHgvTIqEg/Z2A8JdbdMRMmBIu
tuY61scAhfzLsCT60Ongr1Vz5e5Db0daww6/Qg6qq0/SwwRHb6XHqoEcPS743NYN
us+iYCif0hq0AZhBUbpXPgePZxKkxiAIt2zkOkM0vmw5a7PFPAdlDWQxKWBNxuv2
zprfN1/CTsD5trkuespUt6Np/5472bcDvohpO3g4qWVWtDMRU5goYWSmPyg/YACM
z+IaSvAEzrSBvBPUJHxIlFjm8XbbU1oJDwoZY+s3w6A0kN1Mz4vxBJvtiplGFdiW
t3AzROUAYRSftFjPyyNzZ1i4CxUahSRZgQQw9yUz+K5zHlFo5FLHhulhO3iBZrlt
dbYRiTMzOoqZioBpimyNv7MS4pGI0046OfvICvmhYWe4jLZjNn2MEKiM7Wi4d4Gn
Sa0AW1CfYWgzvUUhpiCejvyJbwXw4caWmMP6yFoTTmtXYoo9VPARjTB4JfhIadE/
BDZq2iZggYA9tasXCyQqXWINnrJfpxEqTSd566VCVk7MKS5ei/ToMR3RmwQUM05z
NrtYdPBhuvwe7aiFA3KqT+Xeu2g7COUSlWG/ZKNW1MVwayoSaLLPA4yTp8n8XrEv
iN3VlRQB2eyX+cxhDzAOlsouWeR/Gw/cFzL/CJtlQ5/wtpAebkuAI1I8Jf3sJSp6
zu95aj+ETyWiRll65pP70EtePVn/o9BJKtbm7Gd9daehautEPKEPZI/8Y3fttjmZ
HXFmP+qvK87De/ES+la/n5Z1dngtWZWEBaJdsYGSHi89JVGfynK0b2oHYBemYKFt
gDTXRIVaF7d6Sn3KTvXhid5y8EXj48uMoAsN9f2MNl9fhOygXtbVBQy70sGFAa+C
uU/YdXKDs7F58wHI/tAvyn8pREBhF8reOoDx43HLttlv2CvSKrr23GiYilYZgFOI
XE1qJbSVVx8NQH644IsGHtR2DzrEHX3373pwqHnx9B6GNu1iIJzmyTGTmOcJKFSf
ErraWDM4TnGOa7pHXZyaQxEvoUhM+qDzmC9uuWX6kWlCEh1HyfLvmactGCnV0hrN
GLElUm8iHEGrieSc4jNTPz1a7NWt9uUneAeXuhHDTZ3oM4H96oC4trJmdN1VzUDC
EN1SZZE7oJxr7IXv91pslljFC6ZYqt6BRwaen8ETnECYewq8ahYmVas0GiaZIO9b
aauR2FtF/YfW6jc0EHCPRBUuRgvn1jVqDPQj++VBXTMaCf5lmkyrSqYtlenXuUfy
h8fIenm+xEXetC5AWd71wY11f6B3fJkk2pCvKoIjszXt9I58xkraTUzJ+obQOWbS
yHpqCIKF+k5pcwMQYE7hrw5CvqXBKm8ewPm05fQDi3ZvtBFvbOwsobsO3nUkJB8B
QYC7jWdwJYB5irww6/q8M7N5dwBpZPznkynFD/WXa3VG3VCpe8icqr+c+8dxRtBy
axmY1znuw6m+M7yveshAj/qo2z/x4qDNvrpTWKolMpoW7mT1BSxhgoPSHGbjTWsu
w8aSo4eKq9Xfn1QbzjolRUnsx1DpuquZg6b2hUVkFyEy6gyDAgIWM4lFUnc306Hb
yrE2NvVHjYfJyOpjxKnrgq16ty2VYxtmLbnxl4b6WHqs1bCSP33PG2l9Neov8Arg
aEflkk4y5EBkFXCK0alF+uhyHj/PaQqJcVUwF3lEqum3fsYPhVfe0tQnzEkGsLEr
RdVXdHipzvM7vs2CApB3nMVGCwze5Tek1R9TWyXtz5cP7Mdm9h7b5Bgr/lL/pqXK
W5Uk0TqOBCOSIz6QTx+YSWR75/qvWlcR4v5V8auPs/lAF6w98BzwPPjKGeWpTktH
DCKriedf81hZcAToLEqpXZViq+DVu6UMstmqxlCeqbS91ArqL8B214sz5aBflI9N
2+NZV3GyIkpqnPni2oYMNGNqgEXgh23ojbdIS4rYG/TXgE804ENZOOgZY82qdNVc
yC0A58Eid9bYy/pDX8soGvBVQyfcYF5HQjvdvtdvG6eU2X4MhCJOz6f4EBuzWj43
BxFo4S/KLcv3hGBzgGcc4NiUNK0gomUo20cmqIJGwScwgWue88phUwIcA2MVbV+W
592l8di/eB9/3IZexVbQcOOLBdAiOPzm9krZxeluvP6v/YT7fr2sBPIBkYFAAc6i
poP9kWswZqEql4c8pqNm8IuEAUbrRWPyMEWenacdny6m3d9178Z3k3ZoYsXZUVgK
Sfu10VWSR5eOEH0NMvyjH1DYVt68OJj527LubjT1rfdvY2TQpfOiGKxmyMG8Uwzb
Eo7vWiVAXnwaqmiRtNej9YkSW0EHWQC/LI4nPCrWzSavCDeUHcCDRtFbU93sfzj8
91X6M9SgAwUvaJmqxBFkmbdEJgaSGhUS4qxgobntSs9ZJWk/oT2S0IEPieWiQUne
37Eq87VveLXNvDJFzigVLI2OPBoNFQRYMHwwH9c9nMeJ4duCREABdbSXWDQVI2ya
EDPw6VzZzgh+eS+95ooU7IGskrRNbRyGTAun1ZIchnpNhITqiXslK/CY8gkN5ATg
ruOVlwhRXBj8ln1OkyJCyZKeIRBAKml212+SrX385x+uKvOMAalrLR5VenDuD8Ys
oTz4DevHuXHREZntz6YZXJO/Gixh2M2tFmOJFhRxEIqdorfNpcSDIL7PTp5wMgXO
5PwbBbFgPJ9weK6KoFT5425DyEgjxaSMUe63yGabRMNh7uT/DLZQPpRnmgK6lfOQ
9QTGys7tB+l70StynLlkXUWLjD5o/TZ7nWV6fHHxp/i5b537z2q4UqDHzcqq9Gnm
O556ScQIvjT2LfbRRJQqvyOtMdPEMJEpDAGyZbZUYXi6hIcKCMvPgf9CwxAcXa0N
99tRSqyZmPMDGu+ZHwiZyampc0ByZDWgbjORUO8VXUbuXh25hGgFqoOtpfeGcNDM
jZknSz8XHePneOsQAFSPjZRn2nE3I1AtRfAYMjZNqFxuG66hx7/K6K+gBMHHOfAz
7aijBQkyjrRjKsbGWb+K82kXNKa1rRaHQo9YNGEAjGxGuc1ATC5wZXAHZIg47v5o
L1fJP/ej2wpUFefyeNd5BztqDojSPVXPYlG0IRH/k1hofVYJBuK4AZUoCL+1CHBz
cvi2nWEUW9Bm8QCDoVjj7GOv90KwoG6N5lYx57HTpHnQdVp3JhtYJRVHzKMnRm6a
uKvicv4LTkEWO0D5n1EQ1uSxQFMVIB1REyaGDdctIDE0JWkoRaFGLH8wW5Prhu1l
d4uhI+ZRjcuU4YrXEmpkegAHpBi1i2hykraNEFdcllILz4libSFwNkk1qgLU3Fae
SweaL8qhw3PMFnl0LUKwaLmpuVS2HkxHBiQRiASVxF3yARwjsN6wfz6bTbJGrWOZ
5GuOuP42WOOF0NnUPvrCFWEhK8IxGYEHof3H82rkr6udWh1r79h7HQ7MK7D8K/DG
L9LP67LwtPub6Wk9xL5JZFhldnpQ+ljXfa3TgKgs6AZEfg/XA6mZc7tmMgxSmNVe
hSUpz1hD8jjQUSdyv86TJqwiPqXuKqAE9CJINz1OCRphgO52KR1twS35D3kTrp/t
p5yumMK2kfPm1tW6HdhH4BocBGl5tUFGWQANNI8Y5gORkTTIGU3WciAC7iFUMcPe
IMqrR7+8fz7fFvs2XQ4wg4/0S16Zaza7nwWVZl5mRiDQeIDcYRYNE7+VN23BgsS5
hWaccjt4UZ9qt8O8sAilc7x4HPnLqVkxoUDDUFuh4FQpxufJVgoIPh7hDLpp2KPs
hOJk+GPfOGzuEV7U14MJWBx8zi4JfiQ/l/XabJfvC3Bw58BUarl0NywNL07DXnds
27p8Wfs6lHNkQ7a0MXJ/WlQgE+Qh6u/7VtJqgGMkPsKepnbUXv/4menHD9M455Im
Q2lucPG+gdV896LLM6c73WcQyB/CvHQ0rTtZf08aWCbCDbupK9Y0OmynCIUQ1grS
B+ZQaJ8OETIO8pRsB7cErrRMzmv8a92RbAYW1bamVUdX3WjC01ktjyy2X6v3RqPv
6xeo0smWqB7vkqbCcgRAI3QHRC+z34n6KNS7WDZBW3bnnk++n18uey3cqBJnLJsc
dSwyUI6yhtfaIQPiVKKrTNgKYg0hBZCvOwqfDLToc5caayhD9+1kY3muQU3U0Qtt
lfbIvQM+FFWn591aUN7Mew2q/u7Mco8VM3DcReRzH0O+MkahgeGQfpuXRWpmQzK2
EVEa2Ls092Qcijd8tLAMX8CLVZKAd7tt3bVhKBSW1DxXGgZiJ/Wl86QSNXC8P6JN
tKzmRc8101GIOFekmdLcoILLiADXgWPusoyEG48x31s6+xkHb+Ttrp0qutAZx2jc
XW4X64dIfd7eFz9Fg5dcpF2yXrjEe64PP1JAgJti6u1wj9dygaBT3T42Wi4hkxKd
UNdCNiP5x01FNf39M3FUooBTUHvmAckkcAMBDENQ3uqHs+Ga11NeyZ+Zx2ju3BaR
AiH2aXkpzdujTwMHOJG0wjpqAFdP8UkPPdnDjmOEpSrm3l+mwy4X6aMwQKcVwdcQ
t7uoP9sf7TwPXk++cPB0ub/3WMPsOa0dq3FhqKmRdQuIS1uPugJ+U2P5wF3h5CCL
o4+8bWzSmEYeYTQXAUxWMuuRjA9aHEsZvKFIsbe2cgviXxpmZ4SARROC8uS9duds
eqHsmQIMs+TuPnawBzJBMb5Qq0TWMV9o1hENlD475Gj3CI/8qWarm6fvblQfKD4p
sBdeIyTI14mUSu6cvWzeL5xlcBvNhkiswNbJtjwgE5/eHw0iOEe3D5uavU3mKpML
3o7d9ZrcspdRNsvV016H5ut5RUc2wts//ZH69ZcDWvKv6k88p13lSkkfnYfHFF7I
jNa5bHBBO62wb1DkOnctkhbS2mEo+GVzewq9NuwawyjhV8PddbaSBahBKazVJns+
8vMLoCPyXDOnQ9QF6/DKuZ3dzJ3saoBN4V0B0yvJlRCjjnb/OGP+qgE1EqCfsdfm
9cWaKktZIKFKdb1qarkb2ipUcLVD1TNw40OeX3b3fgW2AQOdSa5Czu975pXeh88W
NhMGwhKTTvPTDXAtS9Z2moCbc1jSJaDVoUfHbwq4xgQYhWenWZ4c/Xk2TjDHLDlQ
U32PuJCrF9NTc+3Pr7C1g6qrNY8bjCb/YAle0/11X5YAPeQ1GyhmZcTJlTHWRif5
riOVaEkNnMra6C6uIbvoF3fHhZgZmz2JDSJx9S5YGYv/loX5u3mS0GXhbH/wJNl8
C82jFzI2dLaRjy+sBSHyj8ypfe8Re7prpRQEIcl0s45YoGYE8Q1toCiKcP8NX1pP
dKnHOO0zgbWP+IOCo9/FC54ANWxi/l5WcGP2fvu0kBu5pzK5zxy5iN5B+qvYbeCs
rpMNA+Vms7bTPdi2aTdbZu/Bf8PVeEyo9IlL9fASrc8MR5d19YmJvjPsKY5zeYKj
rA2uQhDMGrhDevuTfa4881cuuDoFUEG8QqClH83JKWn+++W+sNfOgf/gB/ep8dZg
Aj2XR7XY11HTM5Mkut5TnBsIZOfjFqUw/SAOeDqjTcX8b5a6xEjVN99UkaA9XaJ1
GaF1X+gXD/Z5NfGteooNFR2KW5OUrD0gr+0xW+gMftDx/Ait3wn5TuVgoJQ1IRMB
ktZuQcXtgHUuL7hvdN1btrKF6SycSTiyzigclNanRPlTiWqtlm6m3TCHWwY6nPRU
Kzdcox22t0TvqGuc0xYjibuhLy/gD7A/ZyaHbnUgHj6D4YJkMyN4ZL58mIJZOr0m
60+Fo6+4z9IrYdLGqe7mCis/1LFlGP/+VBoSpkfBK03hEo5MFIpGIJy8hSjyPhuA
B60T9SxdrweNFsv5YRYkUJJ5jqzeS50wRXd4Xat8jIo/Oj9o8CHjFK88rOy+oVTB
42qd9w2hVXpwQGtQzz+0MD2BAekegeAq03nILYDVc9qFFcxKh7kfl0AuAL4DCKS/
gWclb7A5MDtCeEwTULAF+BkAjTukZft4RufheFNg+tRnQpIxy7WmlO2M8ykLqsE+
PgEg6mxjedgsJlPm5ZJmLPyJPXqtXku9ta1kf9pgwuFgz/LmXa3AbIS4zw0YXzpJ
+HdayxYTtuhSb8q0X1pdxBijJAYfOWA2ls3Xf7VyqJS3kSXU/qL4eaX/91NsPtzb
VY5diAsaDoat4qIkC2TNfdCzz1ZGlYWXJyJvMTyrMYtWJaYajUjm0F7qiMGIiC54
k6556Y2HAhxJMGA1NT8HszO7Q28OOlN7bqm+2E1YfOsdeNUYNgH0QjCMdu9KnHu+
zbB9aNbcMnPldB4F//kev1V+h2aGwd00WBvxUwyYbUIMwjX6OG9SDUQJSgCrLuRk
MwRm6UcFz3eCpmcgXofa8E+rShyUJaZl1XCro2zcffVTbSVTGtLHLG9lcBDDLW+P
tIne8Oj6DwZKp4T0Loro1DxjLShGz9xnrK4KAVmO41m9Wkq//jDSbO66SP/yr4H6
eobxgTN2VyT9MFLM5YyhChEL+Pr5rsqZBj+TBypSnKyOFUfiUqHboj2G9IXL+iXU
9+yVr4FP8OQ1j4ru8w3yMsuLDsl2/TZmgMTxzuBdMm+OiO/eEl5x22IXm7Wwv2u2
vnFBoGKZsWcjPLOZl3WHnSEN2lL5HeJUHkV7Q9XbZZI4IPxWQVKAE/wQ6AmriIMk
VNzIUHJBSBGvGh088skQidRsTRg7UO+n+B4IoxJ6z3p9ukVgFbQQ/7IEs0Qwr20+
93bBIP2tPKcipx1GWnBb7+UfiDQsZ05mYYlsG0+r6kfTI/lRa5zS8WlV7Z/Q3zaH
W8FKiQjUV60poXM5nCc4xlbENQpwLXPsn1w3lbUktTh+iz5Tyjc1GR16FkH3eED/
/Vm5z33kr73euYXr51t8qQDLhm53asYlUT/Y4kfniHbzzc6Jzmf8QFi7MkZ/+oZQ
XRbSYaC73sVFb6I54p2G+FM2w/M2pYb8E6Wu+8L2OcoQG4dLyxTwdlFbUCKFpy8d
JTyawPX41hW8Ng5GNQeIrfXiC8xLdbnewy1D3+huntUUONMCkqvEqMTqBLx2ULGU
svYjMKfhkpT8dw93c5SZYyAGt+5oUtS3Osc6RdY94GKbgDzFARVyV+ZEFmuGC9g/
n6J75mxPb6WzsqjuvS4fu8RKm4tPy6gR//3mToMUnrbp47KJSx6hmZo+Cks0hPky
J6+oBQlIWfIsduHoelZKcejBbQ1Qku08Y9cYOLGYVGBme/+209ZZIU6JbVO2undY
U+sSby9rKemS3+BLpp2GfvzeriEZPdUEs2cNpYUU+w5D5gxJ9MqX/g5TIWPEUYhF
zJ+o01J/iornRkQ/xSNNcE0MBRjxmFTBhQdwu+SBGuBEUlaeA7LVzqwAzHBepnLh
ThO8e1iYLmH3J/Wv9OQ1YDv2yqPfqq9QIh5l3jdyvCIe3MS5C5GY9lFeAf63pOzr
aTiQRVts9eeA5sB2j3P7hZk95WKcgErHE04NxiazEAMiSYmHDPjQ0fJhg/s+9cVG
mTRye7b/c6rYmlZjze1fzloVJms8prTfDP406K605sKH6XtxmtaSKhmb9Z+MIr5I
WFDXCptv467NV72QchqaNB3yx2c46n+25hHBkZM8LBJmrrceTVpawuOBPl2tBK5P
HWWMbtGm20/v4QkuJ9AWjhVkyRDyxGLcjXOiAfcvfdKVG1JY81aqYumPxe74uB82
P3dhAUdhpgyF8P2m6x2cBU2z+7Msn8ml3gyOXKAzDIJayli2Gc0YKPuq9ejeqZVR
6Vjnzawes5DQIlosTdQtmolsUVbZQ5rf2WrqS2GHJBz/A7kDtmmpMf09iqrcqZ1b
aYY+2HgJHO5w7EdTw8eV4jafASpTc8vi1G/n4nFDY5dYpB4MCUoUro7HjQ6mg9UX
0p1e4SnkJ2pBeGkmlkvHSOzKLGUwlHX6gGrsgqRCWSCzKC7lpHEgOVghEOxo2Qk7
XTf2CJRp3mU72ig1WmkpsyatN+J2fgHEpaPYHSlJAUZg9Wy2qt1k+kFe2UI0bS+6
GlE8YX9ZQf0ezgJZrmShcof0X47PfgWMJfa8B4WkfnBgerSwB9hMzg3nG6CMfm90
U3uIF0bII4vBt8LLIax/dGsK7REq+Fw7gnkWKFb74f2Y9UTEXGq0QDcZ4TPMTHRp
/rYwU0LdAMM0Qey5JyKhatMs+ajgcjTm7/MO7GKAfoMsg/gp3Y4GWEjkl0NFk1jQ
qYPwXoRjpSLPA2pPqPaEEUWxafhlu7vb0LdORcuqnFTfInjgFyPSNjwtLKQ9Lf8w
SpmAcmr0IKDise1YX8M8hTNMJAHO5VnLrTVfyw61Diaww5CjtVRbCvVtoL1OQnb/
SgPcJiI2a9NPjZTHpUsH89nyPqiplcq5sBOKcnmcDBxWHjxAHdtCx+NSbLHEgCRb
P8ply9t3YvoRaPyOQF3unGMzn3HeBuWDmFmL7EnSl5YSJQoqI7gXkpD9q7/CDPpX
gGgzOjCfNbbo6O7qhq2bKJzJs88wQG3rCj+oZKdNKf2goWa8udiXQkvUIH21HJPI
BQ9mTFH2A1X5fFTh5s5zuYlBtIH2H4qLMHqilTTbE/CEtgEwVjBcwLg0xzmOKtKk
xfLZS9Lvk/KsTbBGluhit6zUvDHYlFsbm4uL65uR8pvPBw1kANrS715KXQ4k0U5f
+j/HaWz0LXECbHM8j3x/r9zYAGkexROxKP87d7q/ZtAOXYI/Fz9FfsFcABY1G26s
AdghieIrtW8wxk/exGmEo1tjTbqACuOa08tlcdlBqmpquQJir2eTY0J04oIVozzV
2uf926b1N/M9WzT2kDRBlmFgUpmqjPNZg6V4sNR+W2cEmvL5aWQ4BygTF89EN/92
fSxLhuPjzQiocmZQaUGWx5pP5zyeUlZ9N12V6mrJhnOEc598PoadLxiEqUtL6rZj
JP5KR1fGuU5LDi0j1nzGAOczyK4JFnjTnh2zK/CvQw4y1tQvgt3Qm9+ffXM1B8J5
aGzPZrMFGtKQrLkIRMbC5JS3l/0MzKiv0JvqoxciS/dn3DCSJq77DThGDFknJSJD
4mWx9mlrL2JNLfHcqWE0hE4pF7A9dSHhP0nBN1oYj+RCEzYONz5+zLu0q+GlbiSk
VOcz4IFWxWQKq27i4c+OyAfV8VKxGG3icnGMxNHJVrfb89EZhLfJW6WwhqzaVjBy
ZDn5D5vCNFp1RV50FRQpDelzXkkk9uIg0fFA+bN16zbMYaQ5qNiOxZpMuszojicK
xpOHbpF4ZtDQSk4+Qf084jpT0lCIHbJPsSWNglJztpsKHw/Ze2XLFK+GEdZaxyUV
y9aEscV7Sz6mO0LzSIazCbzRK2btfyXWLKeNWFyi5gm5I9JW5+n6fxGW4+LhdqYo
zQhji6Fx5zzWE2I7M1gxgCq9qkYEyQ1QgQYeM7T29eiNlXFpcyURNV8zsOSLg2S7
g3iDdBSSGql4ujix8vs1WzLHP5nG6oG4DZAQoM/4/8qJ6aT6jrP+667kSXSV7pCD
Vk+4knws0gXTDSRgAGVJkiuhZvnZKwtguOipFojXo2HgWWYv6SA3OOtIxtKUwHG9
NZgj5diK2NBUO6cmubKB+dY3noGUgs9dJLMXXANUENe7M+ZSePHBiw5aRRnVnCFv
7CsxTribai+0WtdiEjCss+fPSHLC5nCgM7kaEu0RRoqi6WJGx5Zc5yLnIVmQ743V
1O6KhxYG34Hxd0OMaBRn2ZwL+NK2wwNraaL3e8+IVMoRAiBqo+D5Xvo2Z7tXCYzM
jA1pVm1vbw4cXkWolat8lHUxy798Ih0KxE9kuVOTFWlRrOWpWULHSe+FdCYUfCFV
J7ZJWDPormu6zlq5+uZdhhsStHfZWfGliMtfsiVQUDpzzOO+uaTKhHmCFzufiQrH
T2Q/0HRMEX+KELKKZViuogLLxcRx0NuVILDqol7worYdiDhAGwgqQZoITtz6uS5b
+U8HEuY0rbiK18QHf/dTnCD+cFgLVK16+vl0ZMqfSsrb4vjmz0CLVKbluH5xMi3F
j5CpmDfWJaGLA0qTWB4Di4LroTuBjJKNldYUb9ddRfPaHEJjFh4IGGVuw/Pw8nAM
EA/FFfiDYMJivNfi8hDyg2DuLrqvTRcN4tRoc71RJAeDYOHTkNZlItl9NQxIkMuJ
cG8hCLXv/8oLCs6bRjoA/AwksFuKeF9gpc7f9ki5MxWF4rEoQ3b0REir+nJj80jb
siv6Z1WEnuMtXnKJfVegBiWrw0uyXa234YIV9oLNlthkHK3OUZUr38yNaNMwlr9z
OEcvAV7dh20uRj8mmso0UGOareKjdzq8/DBYUwb7bzgkdoa89ib9ChtD2dm5CmDx
Cb/LYAZMoDKYz6ySSCJPWAtwIYfQWXBGp1sWbk/lc1qHrWyJ5I9PSIwc7EVs2MY7
YKsk/CJ47nXWRUmjim/a1YBbDmm82wTFZ65WzZf3ywezd1D9C1kx3qgkuIpEflnp
yzStU8e1cmdkiX7J+Wh4AxV7Gy6TV3BtW721VckslLqIBHXlpzcVhjrzSVj3osqs
L1CA1x77nE+8LaAY6vyfsYbdXzVve7zAiGTboADZqLS3UFdeYohA5WLptmtxQSIq
bFNC4d91lEeDAVYucNj1X0iBL49lYrKI1JRui8SvrRyb6BwwRB7ae1CtIm2haOAF
g73dYdJB5t8nC2Ia7BhHV7RyNch/s2wt/FPrKi7MYhfH+2vF14E8QcP05HixSypG
027OmdO460grgptCY1CUjj0w4vNXvE1l8QRO8knBABWZ4wsBXACQYvwow9nukaYS
/jtNSYmVLssk8zgaXkP6dXYwyqIYpy+4ciTjYlzYS2o1rJvR7jL3jhUP+9rwt3J2
S/2Uo10MCTtjIGQh3wrmXUk4SLtRbaJI5XKVI1cYBFRsjvf5ML/iLplZ5XRv7Tds
QoZ3KTFNbfQhZvFkxPm32Yfci3qCMUfDXa7wwrNCGudh8KYcYmi4HhvbDv2x2cRl
itdlEASE+nuqaCXKroYtgwy3QeL218GVvgUldn5i3owyW3bTMJyUZd8XwtHusNwI
Tcm44xQXfgx+suqSEGbheTUnnrVYV7Pg6of5Rw1XAV6WH6jypBQ6rWbYBrUVUNxw
mKMyunrLy3iaxgQ5ayvW0jrp2Q0NAOQ4wQNTR2oaEjV6JLL8tWQKKFsnJBA+zP+W
6etZdz0NRLGTUYR6vftbRPZNJHqRxneGgWerHs8+VBGEzxlLZ9ejH9eOq6ITPhr+
uUVLGQIRTVsXJS5B/6I7TmAPoRDfj9ToUJkSNPPUeC2LO4DCZjkxc8KcUkDNVge1
4aLnr96tDakBfa/VPdk8Dsa4eBigIx+ZrtFZ72u5LW3IBBU+jVzKUSrWdmThrWvw
6rwFT0NF0NipupECpzNQ5M8AKg0MlsVqNVkad+qOZbA3Pntxemo6aF5vwjqH5qvJ
cPfvXgwiSJbISIgvD1w7dzOkHWlP4z9lku2Mevn+GkDb1vvw+M2wkJAHUVtc5EdV
X9bIY2j3F+6o4SAyIn6b8z0j5sSGJUVKj6WunPfL16p2Yh9J0kPbNQ6cSxtiaI4N
jGD8QSaJgXVUVH5n3usfNNspH2s/8hEAuovjx+ZcUSsEZs+SgombyEAJv0vDzJ3e
4bim2vl4ghFRi255K0LTDLuzl+AI4iYj0EXYjwIcrzjfir6+HHKlx3ixbwzpd61A
FRJ05wyJ9pCUEhnfGH2t3zx/nzl6ONE2dlPWFpj+zS+fPBWxf29toftk8a2IoZn0
ZU+xCMKPbUBJCyBeDmm1UuqzScQ9tVpjE83tToozXvlYRmaFygknPS2hsPx26t+v
5aiuYU+/fwXaJ4/Kq/LK02mCxgCF+R2liVc5dcm9bUSACLJT5xKlCABbYu3S0161
Ho20p8yQQ8vD14inUdpLGMrf2xBZ+IQTSHnNCMxsPOj46U+lks+ypSo74XOgTuqM
HqtVBPAjRODgq7itmtpzmvHhgEoua3Qaji7iU+FUFLqjnNqnOQb3g5Oc9ovzJ2ir
Jro8yBkC9QKGejbunBj0ibk2ylCb4rUY206T5FfCEc+VoDZ9QZ2kKWtCpLAWdQCJ
QAYFYJhBfWmbHQFQ9hxKOOxxlLPnINga3vubOt9ActvwD1+9XxuGRv2OseeAWfEX
bR5aiw90gAc279Hg9fcFsDpqG8NdWciVDn7vR3CYnTxLYO5g0lf/UICqqrDgd2se
CpLtk9Ljbfc2Fo9Qb/VrPKoHHBr4dkf5SgVGOWsBdCk6dhz/7tyaGVq/Dn+b3NNa
wERenCUuyt1cO7ZFsWAdmn63VetzcGAhRHyQQ1EHONV7FrW4boN2SVVof57q5Hw2
uTXMtWMHrVBjAPh0fdil5GgYu4JYUMBK3hPsxGky4EraVjy/D3BfFIH3vskStxa+
stFC58XIjv/vAiXUiOgYrJC4hAXxL8T2Sp3IOiCZ2DyPeT6ayS0d0YA9CT6TmWZt
3DDFh7G//g514LFwaugg9kEyayOvJg3sOmTHWSxI8fs9UqstDIQCBtWcnzV6yd+3
7jQ/GYgnGs+MUb6DEKRETdAU3BID3PTtBpCxYuvVVKErtv64smtDmz5e6usygNQk
KZv7/QqctfF+QzjWExSVGxzCIuokTPWg5GvDR0nAm3ZQ6+iXnNQ04SVXHo4DiHDP
WYsSzn6cIOCMNrTbyLCApGbL17guGifmtWpLDCw/kmio7qqKd8/FSz6cz6pxjaya
/qJYMsVoryI9UgR8DGqhyGhIJQyf2fvk1LlRh/7COomWzHQoP/P9xa2OPBOfhTna
/ppaSmpjaBC0aiKVlBFqpy5uRwUduqlLBqAIeKuL1tdzf/qDK44TSJ/oRm7QWo4p
Lyv/QOciR3tge5ZORC0zD6mCAxEWykzCWYkLNpvo7tumN6xGHDx0n5LbYM5lJzXs
j7qqN2og57CF5iqPS8lTJJfRRpjXPux4hMmd2ATW2aVMqOTxh6uTsEnXzu3sCm3E
y0HJrDr5UPcmNlvc9GkHwaCiCvnGrAXl7wZpli0NKuRRa0qKLdgE3s/G8YZotV2u
lYlU77STE/LkBW4EW3ZUftyq82m7TWG5hsCp1zAc4dWYoKAvRdK3rF3vg8H3otgQ
sSs8LqZ0iCgTuC0rA3IQYc5el4jaT+wCiQ8X7oVYjgoA7IHD3PeXugYSGDZMpsIs
H3FEbwWgrfUOjFvNBHwoVZvhX8EHySbnwpKYi64mDDYJO1LC6TlbueasgU2Ef7EZ
SHVuMS2EQK915FdTpDdsBZpzaM3JZRPXjcv9+LhaYUxwCumy23bX08UrFv64XKaf
nqQ5uo7zLCc/27lqkaKPGzqlUwPadNfCYg+rS2+TuzlaU6SH76RJul6UGeLMKU4A
LkSJb/spYeQa0Jft4UhnYo+OcHNLhoF+1UXew7yVYMC4deLAysKH8F0J+DInkil4
sDlYH1txoEKExrtSJb+OL2IB+IiOIgLKTPgEZFVZJHQOTtDj5Q2x/pOVPmBPzD21
zq2ahwJdnNxuwssj7D6ZJqMnkx+Ct0CcY/XWyrHb8EhzrbiyWZNJC7UaFKz7M4yv
/kPbuctoPFLByJ4uQAYsp2sQdyo6z77nApOojroyLdW5193Abr9AkCeSSD7WPN3N
1FiWq3PKgbMSdAG+vQ9hfysRUfmyqAttBPE0hLEDHiPompw4qY4978tmiijaG+/V
HKsz7GPrj/woILdTx0lgRXiMkjEkS22uM0GRJWgdkMWFDZCfo6n9vWUVwVnFGilK
HclUBGHim2n8aQuk8v+q16oUoRxQN+x6SQy2FaOu0bU=
`protect END_PROTECTED