-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
aCmzSzJqpv/9JWvg/jfkc9l7JDh5yePfAfYMVk8td6eKUHv8uHv5qUKeo0syJGeY
Ug91+EY8gF8bM5CjNmj8Yb4HPXb0JQYOEZaYFzFPSE/302MNwjir+9+NDvVhIz+2
u/y1zPfP1qhfumAr2ElYZQQViBfqxvDD45p7oO9EM8o=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 23375)

`protect DATA_BLOCK
iiyfdcQc4srCaufll6NGN+ZvCxf9QQaC/T6edsW7kk32CmqAMZhDbsdPwKD0/KP1
w3Y5D/A774mRRiO29feIu5Vc5C37ibLrgw+oWBMc17V5HBiZG4Q5dBhOgodzkdYS
GlgfSFfgIXf6QzvexomWzFaCPx0SAFALJte29DOAMI5/JWyrUDDKzjo4hI878vOG
MmEmkZuNLsIqKA/9waSqnkFeGvK8PG2uaIUfYknp1EU++CUniR09Sus5ZgfsSPur
mvTvRhuUz1jDEwLiLUTWOsXN3gT3dGxgcjtu1CSl9SaMOSlhrK6ncyK3uMn3/9vy
2b0ZFvxTrWcpCXyR0bClhGLtCZfAq4gcry4BBeAvVSEi9SaqnKVDvp+koRtmBKxq
R2dCdufyDkRjqmSJhdUvqqh3J9jQy30WXKSlZf1IfwQBujFLN34rkAljYqEd+w/y
l+6q0xEYl91PEkOFMfyl0I1d98zGYmBJGLpRRlkBSKtAIQkGiZKdDCZsXTMKXPJ4
2d+q5YZRH2YVjJQYxEgxhIQcV2NT4c6KuwBxOHykxCMQgJ9wXpl/DkEMVuHjnrOL
U53dkmyqhIUP+u7BuODqqWL1tfCOdCgN4eJUZGWM00b6EGby3BSLXXKgZmE+NJqB
M1XT3et3kM5Sb/kzUBV35w6QhHoCINK+fTHIywHwcLNli/NmKEMg8mgx34014/Bk
VIo+au6OMzzdUsabhTKhPpqcM5W7P5bz12r5cF71P4gz+3v1Ao+/JQ5C+sDZatkx
+7kyvnHDTdJSBO7/up/P7K+gNqTViZXhZ9cnkr5EDQD3Mw19Rg1RxtehE2EVXctH
BSfdxqHTpV/3sRMFI6N+m9Y2o2F3Z+ACfKi2ICKpo/XHdnPDkdPMAD7uivvzWxPA
mRW/3hpyWT+ZDcYRIEQmNeAHmd8KOjyGIrjGg3NvCVyHG2V3XdxOKJF1SrnEojOV
ndc73DjVu0rEi8WP6pSlcvSxCrXUz/BAWqAPQPpOsufvmZY4kO0aPiWqfa17X2pV
sd+XNAL+Qwjr3Ds8DtcUCj/7r/hK65iMbZiyHoqS9sC3gF1hfDQ4MAeovOGQvdue
QNWM2NbXYsY67+03wdGQ4wJuAUugOT15rps6sBnUH0mcqKHE4NiziWYqHedAxb+x
iEKdVy9+hjmX997QSKg8xV3/2W45mZvdyaHhPlxuuyJalmG35zCg7kY2jD7DZO4h
Oi/9J+Etz9gO3hBjl1qEc7LLnPcGNJBC0VCZVp3h+yJYFXqFE/UKGQFXMEC66eCN
Q0l2jULIZulNpwVMehqudvVJiqgQvIGBrjzrxIlV3q13GR3Ei2x3NfD6wQDt4vgy
FUwGShUXiJ651oRSvhWncO+8vQcJwxHxnntvvDJtAmStPltHETEOP/Uzohx/7Svv
IBv7zEgsIdBLKfjhA9LbpVx+Rze+VltoarRLhfTJnSMVEv0f91ut5HQY0oXklDs3
Zii2X9MitbrxIxKaCeWDWdKLrhmIb44LyBq7GJTa3/k6c1+bmovsFm+w9WxZa0cB
W9ywcwHRiQ2gT5s7S/4MAC7JrjBOBXAc6aoo2zM73qMPCKeIG4s7xH23hcPjV/Pw
srngprEvE36ArlGBzCwnbUDGqBTAg85UtN0EJsUD1XATansTS9jH/5xdNYrMbc0E
R3DGIrsa7Cx8x4+9vDwE1sygoCIVrP6rtbra3H05hP27in33yVZJv/iErBAP2qnE
dIbCAlMdfOIoBjnhvLtx5WFQeQ6moqvP4ieJA3DKqKwwyY0gJ1kIEqkJMuzinkR7
khRS7WPcK/fN+UOtGb3i33jmDq7UrxscrfjToRdTXYdMK6hjmMRpxBB1UyCB5le7
o/r5nT0B5ccOEAxB8NDlBAEpoBgoCNWrgsP4ot//BsDZ/8hF9ahXuR/qG0YSmTmA
Cytd4Avcd39wmTS5ajqf9UhJtCILF9pT9RMojhrNgF66QgbNQtpqSsm4t5M/O17W
q0QFkKkisWRkTvMHXtjA2T30nfA6wzc9HPi7PjLgQP1lRrD5ia/8IliilTsc2Hog
zUBbJg9ziHIgJ4JJpKslQ7q6qfBNK2P3L9d5h4hWqyaadOkZFCeUrhwnDg+ZEChk
bPs4/ZQc6Q0VDFkYjDocVXgS9gXUenUQd5VBsSeqYSMrV/rGwWZ87f1yrhPP3m+f
keCaaXC1GOZjZekaLMM/9QiVF/WN293sZwXR/o6mc6tm1ebaNw5kT5eXbs4uBFjA
bml7iOZVMotVR3UBgfMYTlO3MenEOVenupnGRApRdcFEbLqo0YEHuJyVRDGmtGTI
sRPdzrWN3leozS5jypjzsWhMvslxYmVR4gy2EWIOjlbmFIHe0DGQazZhuekPRDlh
tfFzZPEBngY2/iMQ2uGhmjuFcP0KYYDcosc7bavV79kb9p8qLnv0ox9zZVh3cpfK
vEx+0gyTC9++i55n2ArdSma+4Nj7F1Oyd3rAqkRqZeYahu+UkYF+GhmWLgPd8IQa
V46ZvYetLsGPoLrUo07d37zGUtdZYblrBAi1v7Kpto/VuUnnq34rPhrsd1SNpsqx
3GB/JMtMduA0RY82xrmkltbqHStQRhMm9ku2Y3KyOlwbXqA69KxfiJDwD35Z5Z2a
kDSwnPCJzn9a4o5r8tDQOmgX7Con24DeQZwEy1UjN+HMS0RtBHNRkvh3BBMJpT2N
HdKWPIxniWfZ23/ZmGChKCqWJXueLd9oLJpLAdcOQBXxsNYmyXo/H/Y51AiPW5mJ
4ACpyMQlMsOV0nGbFVF8OEyVhPiJlTHxfkxeXrfrj5ugJdYroaFcs7hWvo7akZ7r
b3pdVnTMrXolk6Se61Bbh998sIbo5YOcNQgBNQPnfLQsnkz3Xb4oa5dQEeLk5Jy7
hgH9ZZH1+3C0ugXRkaQQ93nKxON37Vh7bJLcpVN8Ff+xI/LCICOe5PKBVabiFsYz
WKP//1SDSX0A+kW8s4gv+qgyXs8srNxucZLO8u9wUYV5K9eToq99WadfwETcgvJy
7DZe9OYqp1iVj+C7xl6YeYWKAqccpgbvWhR+5RzRtiKTTM35PpfGLdx6eJQ6Uzxd
1Nw4zo/GCa5j0o1DUGu+oIk8IZJ5p0AbLj5vLanSUDcOxIVZdXpzJW26BcVnU3Wx
RARXsTvrrcOctvOMmn027cLRoTWXGC2YQhXJKWlh9axxa+kHN93gfvZtpNOaVrdm
DyzvdEeEOA52WJKmBNcQocH2itOoOoIS5rib7spKCBCfE1pLgPe5NEpQKxn/ZFE3
2ct7oyU2krUjkmdFC6nKldEuo2El9YMgC06+LKsdE86bkfSPwTg6SegUHIca8wjR
yvtBWK8b7hpMeOPTtapBGJsIUNNcsuVskTdDdEV+I4kS9lOMZFmVlkHwvaTeaoS7
hh3yMBwjQ1u3rbQeg/Jej/NrroN+R4GKtQItU6AzXKxtL6KCdxyXRibM/trTkTaI
aYnSNV2lAYDeUQQ8GoJNzuJeDDdzE93cGUEfiKLMSK+DObRUL2qHfpMXBeU/sb+s
6x81d7OuDni056GeoNTM5Vs8uRroO0I6oBluPs+ILT23Ma+tL9kQn88IiqrDML+8
puFn7seOTb6xJgkeoV/A12S5u29RVdlgI/TOzK+ktnBrYTzHKrvVzVXFKBUqLGw4
5cpV6C+XdwnN1Y2LsrGMQAH+JEnUiR5fv66D8yFbvw4ncEv0y4k66ezS+Us2hR27
rPOIMvASV30n5irWjcVRp5Vs4j9I2/dz49Svas15iWq2eaR83RynctJJgAHF6uia
VRDH4o761F4EiTlnuyMypP1W5nIjDLGgC5RDeocYdzPODOLKpn4A2qvtpmJ95s/M
Ury0lnECQZsB0pjKYTSTTqErvHy4SrtZ8jQDeJ+JaP/4/giA90T3D8Nx6LQp2TIk
1vRZ9ZbvgJpOHuPza2IuaeMY1BT4No+hvTFUkvpupwQU0/ktrkbF5omMJnlMEzy2
XYbekJG4RdUC3M3ZiH5ugDjBuOyegVyI+cUNEuAXec/gbuG7zxjtetRLG/Q/sn06
VfET5YuMyRvWWAiulE7xmldSHPeh7lWOMNixCyiwwMviFolcwycOeBtMW8YPKRYF
66cIVKI+VvHwWTTrjDJP+BP6PX6j6LemKbesgOZM8j3Ijc6P5ITOoOvsNjXzXPU2
3Ng0iEEr8PPnEK6rxSoKrv8PbHaEs2pwQ8fkpK6MAFAv/SKG8cBzTFxs5dQdB+z2
Bowx0w9Tz5jbpIB2m4U5XjFm7sV622GjFIu1zyZUHe8k6Jj/wiGgGhOi4U5K4ZvR
zRTPWTMrByBDt+mmRetjlas9GGU2bkQq6CAG/1yzCH9MVZy9WSFGGMEqUHQtnqiN
RoNvtPn5hOkX7u0TFcDywUcgVQG6axiy7x3wbgVIh7Nmp/mvBKroEUK71ThFg1Hd
sLw7FnWQHLqaZqy7t1K1qK5LiWALTj/jZI/+wak58LV6SLT+DtPNfbbniKzlntWc
tJZGVvD3r48AfK7vIHCkPavyyCd32ouqbECUUp0KtJiqdOP5haebO0W7r8AvbuEF
3GX+tDc3HkISCi3gtKhPF8eb2a2OB+6n6FxJs8Ph6Fw9kLJzKF+ou3yYK2b1wQNc
OqB0ySrIZUS5cjmW3Ocu9xRzm19uRJXnilaKmqJKJJZNXpaC5DPcWpleHwiCMGPl
4tTBvQlqKcCe0YQCvGc5jNpLapxipdk7ODBgJR6N03KswxNVkxeXNzInvoZ6VYCF
3xXQRyWrklC4PnZRUu6+RTsjMmyrwZ+8pI3ymeO4Gq0ZyZSJZ2rlBIWqukOOeF36
DwxN+xm9AqNfwzJJvpigeZ8RMolY/zLzct9AR4cACT+lB+cPORwq8KH7Cg3UZVCm
1rV8TFoHvbG5UUrMFJNO24J21KdEVqtyzIy6FVBt+mJK6FeFyul7Q5Kj+XIhqThY
AKJ4g3NOY4b/+bY33l6cP5hPaIgNmeZn/eqIAdGTJnZvBEwpbU1IFe/qzaeZlGG1
Wt/grYFlDb7QtOMCegT33lz9dwxR/iJ/dTOzsDr6TVMJ7uT3nZWkNYmViKf3ZSFR
iO9HRk7YLV1s+fO9VTZVQ1DOAWz59ohtWUYTkxIp+73D6YyupKoC4JAXNfjhy3up
HSip8P56nHCn3NX/1YPmvms86iNYTfuxxu5DazD2xM170B25QIMzEY9vjM1opO8w
DL5lTFWtT6Yp7tpByAnsoohuH97vCXND4Ycj+lObcY0ZCGSzChNB3M2Ynvsa1m0d
ON0s3ITj/OgLFx/AnmzuQkU254FMVwyG+pH+5AjaB6zJ7QcLbJHolpX/Z6o2eQD7
cbxG2y0/91pm+ERyfCu8NKNs3JBT3PDm18MWzxhK54uEky0XrYTTaVQ7H+iV6oij
HFnFhYNNdoDxbDZCfprFxC0NCsahe083O64C/hdgGbQhYEqey6QAF5m0nb3bZ8bM
2X2vZlxnGap43wHoE3UptPoqQaw8W2DVB0Rn2eFk2S2kR3UWOBChrEZo4nsgf6dZ
ZBdTCkdQy1Yi2JP+tcVhMGfus2Tp4u+vsC0hrOaAvFqMl4VHT2tMLPRo95btAvNZ
/4vXDqyNkBHRyUwwqSnCRChkhXDhl48CzlBWEQoDX4UlE5xeXDn5V9MgnX/MdVBl
vBC3iNb8WehOyuni+tp8TAs1LSyfD35kaQGZyAhJS+DfcsVwOZn4W0YzJl/MKTVX
UW2s3v4yFQsNC2Ywqa657T4aEd1zPNeINl/C/i8JTG0QS6x8GOl0byeB4udb89Yt
cmA2kZH7eeDcOHcgeUdHx12iKxSXOU+JciZQpZ6kXFop3DxYFGHGCqPAS8Jo+DmT
BFM9+S+XAfGIh+2ARyp+Z/M3OdmhDAQ728q0VHiSN1tns6HJNkf2tpkNHAmohOr/
CakDRg0dKJYpWJOh48c1BMEhkfrw+PvBh/vM5yOshUjKBmZMAMu1Doq4YYW0iDlp
1JucYSFeOiB33WRVUqrgo5EjtcreFo66IcfBVF4Au5aqWSk2Dj21SMMqm/0WJnDv
NHzqKa7T10ss6xhcbnVzmUULgIfllaza/A1iztLzTbweRpyZXqYXCekKD7T/M6Ft
bDVmQyyQ0qCS05H4fbPFxQl3fKgGsacXqD5NCQyuvk8hhBpRsFJSZ2ZXbe2aPqRJ
vh5vMu3Aa1GleP2IwWDYM1mquPxLL8TbzleR0E+pq62skhxHGUGw3gEmO6spB/wk
Z+fIPQ7N4hEK9OwM5xPcUVKAObgEBFVULK0oCwQY7IJOGTYHtGTfag0OV+Lg4seK
84A75/+h11l/jqrUlyeYti7I/LD4hq2nsGWJviCDZ5AxB43iAM88zRz6VXozm8UL
3c12sRSVIFETBUwuGlIcOALz7rUpddfNR14GQHN6VG6I4pdR2fJhI0ptQ6K9tK7Y
v3Uo1tJt3IgLH96VYxEWV3RvWQ59LegIVHTvr9CqyQjh8ZIdamZVi8NLuh4DPYAE
+0Ppj0ligRkji4+E3G3K/5F4KaRPbB0WdOldvRzQbHvlpC8t5o4tvyGAYKJX+UQX
QOZuyKmCIiPuMLgmPW49jRw7NDFFj1tFbj1jEUz5gyJzlljm71tToKT3fWZEn8RY
VXN+nFAnkCKXsfaIi/c2S22C45Dq75b1ZYF8pMzCg3zWvzxim87H9xNCPn0Z+v7y
okLezyV78SzkA4NjZ0NLhQdzJ+ITdiAnXz+oTZnhFMwAcCRHsR6jPjXQk2c0dMRz
Rb1AZU8vVlu4p81ClJssMBrLaaY+21HSdn7Z477aQsByWv2s8dYzyVz3rqDyaN7z
ENB5N3Myq6Q0KLWGXEgsOWYwuNPCBdHThEFDK9RYTF597MpTYHkit+6D4CUKnA7M
T1B6XrJidPGsCrKKXCecEn4ciPlU/Ssg9eo2rvo48+dwum20LpS3SiYsBiovLHyh
HdMKRADBxEX1dU2VrIyf4D8foL+lCrmWwI2SQ+4QeXarymKf+uoNtTgcmPvxNz7j
23/eW8DEaV17eLMCeUVNquRlk6siT5A90q765hcvOldjqqjquWMOM9yhMrpkVAGS
oM3Fyldnbp8aK/MN8rGPEX8ZTZvz7V2T2qsxMsytgnhlsqy3JBO5Xehgii2ivr9L
ctXNaw8/6LB0VYGdYpCdSfaZyeD1twB62xvQ4qxelJI1YkJXtsQmJzkup9fUzytd
hT2KR6C4pgF+3ya6KLSGGWpVHPA82Z2HPX3pSE3Lx7BjOhxp8DMBaTkuvkmc1Frp
MFQi8LBRaLz8lRSakqwDv86WVfI/wK16O+DA482/E4sPU+5NNuBT3S4wzo/EY7La
ySmgLcElivQk7Rf/ec5Fd258by1qwEFqnNHzzLtW+2oXGjJNnN006ABovu39O7P8
o/fIDIVKktUIyR4W3gvuktwp6Krc9Rr6PpLQ2UmePb/avmCAB9aRZaHmXfFO3kNI
xL82cS+Kne9QcES8YxBjSTWQshaoxiH0wGmDXJmHDur+UAVXnYX80LTY+6l2gYfW
8XYCeZH42GAMpCFvz37gu/QA6Ifsfa8tZdgfcREfQGqmc1Vtx0Q8OLRROqUY/7Pe
nVZ5XlZSqMVHqhyZNb1q86rX/T2UwljOMoOVpeYHEUK5tJ2Em6WR9ECvc0jUrBBq
rEXO7/vo34DqESvQpk57PCAPyKDFjirI4+WMoIQKFE49A1Pc1oCG2ZsEX5mj/a+A
o7KkqIDbJXO8DoQKoAvzD7CZPR6/aWJkmpAWVQYCSJnRmxrZu65PLln8xnINytta
liWGV0+11Rj4IMRxRcFUqtZ85nX3Inc/zIDO44jyQUKSEYPCpCCLbJBXD1kmHeRN
dFb1dApHQ+kDPTbz5MZ0y62wgkP1F/1+BAYo0EQnTM13dJve3KYSeNJa/QmhIhB0
r5x5wF8lARwGk9cfldMgLhVrd2OD8yEujPu8fB8Ur/c/QEK75NcnmJ5b4pBgZczY
sX6Lr80Ck8ufSy88J16hz0N0lohEEs4HaEccCbL5Mm9QSk8wtzTOxUPoQPr9L152
VwWorbxe2H2v+1ahPb5lEvyi6iFZ+36n3hCu3zCnu7sB11UrOXpvSbhyyeUbRVFs
fLB1Swee5Yr5ptIGF9Ensz0FeORPqWu7zspD1xhLyyQko2P+OZ6I4A4TSpXLI8cG
8Uj5pHPZ0rvq/BMpwZrexGrFmm1bSWI65d9sfW14qDC53QpS9yeY1ln75Avx+bdn
r93T1WG6wb+tyZvPuR64n2FD1t+uVG2JK6EP6SRq8ZsjQZ1Ruim9yhU5kWJQGgIy
x9sBDuvZaTB1TA3BUY6KbqTfV0tTf3vDkOGDaWNaP74LDLlh5vxlvBUXfG87HoBW
b7Z/7GTAaCfIhash7gFFHEx2dxRZKjNxm2V9fnTr4kVVN/0mOrrdRgg9K209BFH/
cp80fuOxpQSmKEChfmhQge2vRIed8TazKFOExa4J7GrWMW+l/lcrfcScPbDJKQdv
o+c7+jvCS3JzNH2viensn/wCqOGuhW8b4rhzvMZbHRnGRYUlPATOE42g53ByG65j
+YbBXq2RkcKhUZnA0/hClphQ+YQwDZoWtphBlx9tiHAEepfmXwC04CcLvUjQ0Eh/
l1Y4JrsQU0knpnsD9PDkIjeNSVatfpWiJTnvFvEsF9YLc2vQ4zBN7w7lSVBMf8cn
OM7I5vN8N7UlOXriCM9xlhtUjELWeAPGfeSOPly+/+0k0t4J+OGrErPYu4svX3Wp
XgkXiVGXq+ROmJCche7F8xNrWq69or2QUCXkWfmQhliuWIp8wyaAEihRzLoAJeZS
TSh4SpYHiXtzIPVCvYL/cSdemo8N8ufe/vVUiRwu31SqxbZysZwxEHvBpaje2BMq
Oi6eUR/yZcd/V0d3L01mNKt2TaGZojfisdvDHJBj0eIIFEUPn7ahb6ZODsmb7nfT
RvLV5TH8vkT+cuviwXEFjn88yvBCmAojGGBQbCfied8O0Msr4tLACfJNV9ya50ba
gkQWdB4IJvMfbhE7kDPZryWwG5HYFcaW1rG8Xlq0HmY/+1QjAza1600lvtzMs9kB
qWJf4rMq0oS1ZMcAeahupUbpiNJrk2GqLJUULOaN0zKLKXZSMxCCaOauUM9gszv5
GKsWadqKkiCStvQi63jiE484eABuHZgE0+K2sErKMjk92O6fYrKZcNlCl/wDbyQU
o5JN7a4iiwcUrs230EHC1oFtbOOV6/JFUt/bzb+80dLAcma1cPNqCZAjuzld9tQa
Ur60nXye9MJ9IFPNbgfHDvfh6Be9ZOGw9bI7EHe5G9qoXXh5qe2Z9i2QM8yqQNiV
pHPH7Z/TSyJ9jg50M/huvZDIwqQ7pgY20AhMPCGBZg7vr2m1q1q9NeGab1xJdVke
DNIZf2DU4gkvKz4pLOOKYlyEKvh5mXw0V5/cZvVHDAcKYBHJga2TJ2md15zDQtEj
+nUlrLLBKfjmqjulrtlikQQ6G+4tOCcViK97IJe+urVUpgA+BpTgOt8tbzntQYwP
bn4c65r+TnE4vEwlSWpMwFxxITQanJ3eL0utuRujOLeGV2cmbISnoSpAt7w+odP+
io07vttq/LKmi/cWzw4EJ6dONbzGDSuKN8z9N0Z9W8dR3lxzRw97Mta7t/8qKdTv
IAQyNXsmMNCF8qBIoj+d0DzwEJdWdhjrYSXBp2h9GyN+jn7WSVhomMY9XhaSYgy9
+2TN/PRqFn1g4d5eIbbSuqTtUcEU2k9Q/Rpz5F+prN2qSHwxyF44FqT6M4i3int0
AmbNyHVPVdfhGcLraLiSh57XY09PGyww1DJLR+r01SPag9t4e5rTm5E+ZpsoffrQ
lKk+55f7VJD+xmMOifk1y0M+z6u9KNmksrUA0A3IAcfCGO86giaAulMy9muzMWrW
PuP3TfhHUmmc0dbFM4cLuiIiVtvPwVkmn5+uQYoT4ubpZC8pZWn6Sq7+kqLqF0UM
zIxlP2Spv2hSupktvHdVBz5yJtwp0Z2YpTKVhYW2zAK1qFPcldvyjaCjxKV8WAaS
7qnQBDKL/ckf7CuF0Jjt7YQWReSawua/jmk0Y3a3hXMdr6nHMdWokiBXsLk5rQEt
NgojwvvaRW3XkRq6mQRRXm06NdUFy9Utsoju9BvaXCor1ghVGMOtQ0oKAHQgC+1+
FwYdfDDlWH55mj6Gv0kBIf3xBg2o/foOkX1ZLj6L0OqGDGxrpO+jUtPhP0HERmyH
M8kPPvlfyVKHV0QTw03qk5F+/LUgQTZQzR0RUskexfVkLFxiOvlinPcKz6ospzgl
x8v6YGOIu/j9a5nVHJ7aLjK0WXNouF8XEtQwyV/6dTdcPFXrrUh8WNZfY7QCVz9a
tk0zoRkq/nfBTWqH3GHf/fjFskqSC/JeZS6HZRQNtt7OyZHlVmGoidPtIHiX4/V4
du0mhYqOeW++qLe6QRaG7xOjtc235rX0wHMB1lv0HXTCa8ColAqfJSocl/93U7Vc
haKp73UNAYmKgDoxT+5rIi47YI1vBEnYxG1/gUaNurLYvkTxdw2DJ4i+Wmj2I6DF
Ti/Qj48XZLYc3KsWbeOZPL2IxpNjWKQ2zbiBBuDe9cYLEA8+HZ1ZRpYTQ7Xfia3C
oxU9IIpZkSBM2ZEkjhGlL8BnJTZWKrCYZgQgTW9L8tiTUMi4PZEGelrIXnbyX5UY
yf8zbHUyzKEwWtsAhf5mcRvcr8+EGEAUe7bOEzQvmQGzoOPuk/vIicsWEQ+Nk4hN
+okECLH65ipSVQuPSQld2Chv2sEQrX/3jAFZD99BdgoNHNpgyHse2lTMT+H/Tu6f
OtVl3MQTIQdV8tgCuSC90AFhnno4A8GJuBAKURmiBFkUNYq3Z0WZMWXWyi67C/Po
7ZXK8jkfHDpH09WjB9gRC4CRrAXLiWcoLnseIu0Vhga8yH3fAX/zUVuGNsmDZHHG
FhhZTJ62JEMLn2dG+CX/RJIRJurbWtDDO+VAg/dS0xmzi3t155wQn9oZRvhF7H2Y
8955r4hG17DK0jHO15aVNrzihthCfKDFWL7bqvaAOYqzNj/TlVoKBoPO44qcCnZT
vCOeR9XaLzqB4UXZEh77iqWTHQ5OMEcvYjT7OsQtm3kac51Zwh7Hmua437w74M4e
FCRCGY61AANlZY7W9WbmtINlW0oPZQVOL3ipLv2DuOW0kw9NwcfLLbPdGyfwq1r6
VEixh2ki1Bqib+swisKGEy2HoZ4VJLVzyN/FtAqKFRy37/w8rYKwjrP197p4G/vt
ZKiM2w49SHgD+vbyKjkW2BcMlAcrRf0JKT9xK+Rvpb0wveTwVqvZqn21u4qcy0hd
3p1t7Ov4ELJOA8uefzqrMx0QNk/9vqsTrApAeGo2BlIxLyMlh3agaBYRH6TE6qbr
fkjEothuH81g/+Ub8Jh17ZAl4u8Uxy92rANftt21T+wwVRF6M5zad0nxotK26+zs
LM61ufjlYM1e7FeOgjGg2uTbnkfY0/zMuJoSGjs4s5l4XPPWIHVfSbG/si6Z+4eJ
MyGNc4hQL7NDfL7LSdu+qUQncmNe2wsqtfb6Pj5PSv8HFVkIsqY7RxMGY7ymGLoQ
vRryqqmOnQJRNgvXTYUYaJcgnfYR76sNWGy77K5fa3Z6yKOtgRCVL8npAEd2txDa
eGvE1eoV95FUwEqf+r0pOFbmL/5MgRuWeSV9/8fU5ElvzKzrE+PjzNupdWrH6GTb
A6Ziibei1JqJqN0REnZjD0SNY37GatwhD5xHRAmn93KmmAyG21T1eWWP2sS7usdE
QrHVrPbR0nXElAvvfnO0KPQ5VnMSPTY/JLydYuST10F+BEu6pkEOKZnshTFtfKPO
6y98XjiQYAlcn2L/YhoCHjUcFMNvbKzZRi1L8p4d+hRMPu5jFZUuzysSX2kXTfzj
bgJzM6zVfKucs0hS1ySvM3OzRrVKMB/RE56n7P3kQB6QYoW6eJ9NDnA7dj9OPAtS
iCSPIS7YmbJiqFxHeLgBWeec5p8EQPDVGOmMci0caxH/3i+tAucmtoK8vqNQfFor
Eu/J3QZiy5CiklKnWJembiVkyUTXXEdN4sSez7sfUxmrT8UUeyxJlx4pm5KO4vJJ
ao+OIIBBo5T2QNpCCyhdgX+53Gtn3pvJ1EZ6O/mWN7+WSbE/500UV7KTSJmKYacO
7s/wOa9tQIolvRARoZJGE11GaK0aJFPXTNJXtQ2vZ1uJjYHhWchP9ncpZQeC2MMX
jyv9HGdO2rn7tYnfJmqVWeV7sb8OyDrbzG8ai67qs56nA9m6soPLURhIf0BBo20i
no0E39l/AowebJsp1cQRYUnj2GuTcp6qzqOA0HJhr2sbULdblcXLcN49chDqvgsY
QqUbirY3lP53+FBhp2DFjeUWWtFvJIq5vxCBz8/ZdE/xtiwe6xLhZw6bBipgS9Ze
u8ToGsqOhIPkZ4LoEZLGyk8PO+mVSW6ju/9X0q8Msg6sz/Zh26867ZGjM4ucKQyT
AiZXqcIixbGrbwfkD2emEF+Pp6S00J16EXw7OjH79VD5LoSy0bxJ3WUwak3U0i9L
SWXV79j9Yz2xv7fLfl6M0nCBXKetwzIhQ+bShGm9LFLPw7jUTcOlDVNeeJJyDzyc
gWpbV1YZHqa7hV2V9R3i6NZ1qxg7YtouTDrBPqDOpNfavop3tcSY8ocqba3Zs0HR
gmahMu2aPMDZsrNTPesZsm0IkKozxncv1lDGO+1tt2o8IUiFSI7eHLKdLjAYQgHb
+RMEsF8vfUR5gGndQxe5uRP0WtW0YR9U/Jgn6Mb02VGdXxe8SfbuveQKcOZSkYkV
p5Z8LEEoZyStWaYmvKSmBxcPhUpRTvOIIcVYUJa5tw5JTpe7yiQrRc1PB8nqND4Z
zqtjSossSPoteFGwiannd8RK5Og64J02g1djdb12Wq9oPOk3J6clsfZw/4q8p0Mh
dKcPtlkZ5uL7l+1xtV1gJmEwyFD6s6u8ITGUJJaABX9dCrr/4mfQzGZ/LLa2Y8Q+
B7m1ghK1VNa1abit99/VVnjrpNBqUITD9URjIU366XjVeW4zpJiiXecJgt5NJf7H
cfNISk39Eu3QxuQVTSb1wPE6AGWCfoaiGAjpknxVejbB11Iz9Sq6wNF6ojWDNqZ7
szPby/PuiTYoboDAoQR2GZtxwX3NXQsPXm+VQX4D/gGF0GGxE+nropHMo2lPPAOQ
viL3xPwQ9j+fKvln/dUXVmMlU/xyR1gRJVBB80uDM2ooRf1BLHyiXXHDkaA3qQAD
QjGWYbRxtSWu+V3oNouUQ6tlnRKNd3Os69KYSeUwpTZLW5jIFIepBd22LMj64RCS
O76KjBb0u3Un7GQ+4El1HxnnfUiSmimySzdmfoxD4BgaG9BKJjOOFwor5Mq6M259
r2PKRaB+707YzZX7BQ5UoncyJaLoga+w8ZI2sUEMpkl2tQFOMpkqaZZkWhg+LtTB
75PitylGD+LSqlVxqrwI0Eponm43Glc1VbIpnU8qob5F8/C5jDMsFjhM++/xyM+8
mkunLx+rf3MUjdydybHyJ+nqHQrRYa3+zNrVjW1oJEF/4GojkGNsiGp0b836P91r
++mAKr0bsU/8YJE+3OuoY0u8kPUtcXQ0+u6y/yjXy4Uzgrs9jJAeEQv+uCeRYFUM
FHMo1X0ya8weRMyNcsZZL4jKeS914qv3j+cZfMmqHCDtaKUbSDmGATAv6zCuDit6
q9b+BLLcW6J2yB7RIqBWGxptHur9ZE1H8AlFr+Xd0PbkGjWkMmMscB/cRvCDbAhx
zkhiCDHdTnwyw3JvKCQU8jv9clTTRmfHJLoX+khEJ3YlfEZlBzpfU3Xw5tvB33Gl
A0goy+/VxYbGJ9VOGmbtXPvNTC3fO77klFxqZTP6oWkEURAunbc46plzyi5AFvGH
4vwB3RJQq2FFn8bcREuFJZO4sXQcqwqvV6U3UloqFfVdxLsZYq1PZWQn6JvqDX/n
a3lLRiagY/+Zsf6WfvEnyQlTg43K+rSSMIHNf6BNK8hMlXFKft2gG3lWl21Fyy12
GC65Yacvh70S9DdCzwWtEiQs/DzYMogaoaIDS/pRejpYOo0bH+GT3Ot+yukH+0Tu
Qfp+ht1ee7TDRRXeODR4gtWV1QzZ8oAX5JP5LrjydyiPCfAvOu+MKsPqHDRGfJzH
IVKewoVvNo1QdOqM7jne8TBh1yc6z2SZ3Kt/odrVyRMzFk4DelSq2v+uYO+dutmN
WjtKCGYu3nsY3/vAvJsNkOLBmjVOtnF398UUmakA2Iv5iASDlchPCKFbwWriIZvK
sCCeZFOjOQzLspANd4FJ93xyjfozKH9pYcfIzb27JFR6z45Yqv5lAal3EcAQPKlR
mojsewq9tw8IqU51YqxMgiBo+TZnnCTv5Wvl9blWbvzG6yi2fcAP32P8XWAcIH3V
2+9rrlPOYLnSW85lYj4h6wqO/CaRCoBrqQcQODZEWlBQZHIgQgRtGD2YZREvdO9Q
oZSBJFThueuqXdAaXNFsgKo3yiD//JaseNupe23PdE+OFH0Zkb9hsFtWwammStfH
bnClDzW31BN8VSD0IlMr6p3aNcL8yoeEhVWTkCrOeZu5yJl88v9lkFs0QD1aZNM9
NzMTzIbHOQoOefjiC+UehjgP2VHcsbrAbcigijvItyO1V1ZBcycXMoLtyJsWuRoY
32gvveR0O/CR492Wl/1VFAYsv7aiohTOWgJlYX3stRkbzZpkRuqc5588vlD7BcgC
BULMZPel3zKl1/Jpg09L2L3BVEW5D9wkbWEmq2TdultHN4yDxXJd0glytGmojyRx
G1aEM31EsDmqG9qHe9vMFR0NafFOw7easkc9zZP0Xso2RQQglvxqFZDIjSOIcXAm
UGarvEN7Ltdut4pbxsNmZcvrQKhI+OFfXd6KK/UfCTD9mxfaQUXhKrnQp2FI8lZC
L8UYnUqhVkd9PADwKjO9TU+huZLxR3Z05BpQEz3abjm8QMSFsM+pZqCjoGJarSXM
2M2980xE1xBIn6jDUqpinkKpuSNrn+/8aHEdn4aHyiSrwTVqrJWTogndcjM64ZI1
LROJBeahC43WHmXFKaQygsBcrmQTQ0/tZ72nHIqaG6IwJ0ZTVCNPK+miD0lxlN/2
Gdu2Pa3V3o6f+JhB+/5Ur9JUltOXNZNIgmjWAbI4L6Lcmowl3G+wmtdj54nAjG8D
qukgBsVPsNY0jkS5+a70aLaAKZ6ruSM5HIk2Umroh+XDWiXF/M9MO+imUiI+gHfz
q/yeURUircjLgCZJ27jGIWj/CWZuNQ6x64sZdlqPFT2yxKlNUS7X3Z1AQZuWJg54
/KTmls4kq8SkUIvSoAI3RBYIYBI2ooJs8yt9y3yloTsfKeMCpnhzazQZbnpMaH48
fM1npMYIvtwSwOOWF4TjJgUHRnSQHR0fLRMe8zuYL7eHkhwrrez1akc3lykRuVRU
MBS7EEoNMCVIA0J6NDlzGyWXX7lZRVOvoyELmSCVCowHosRiq+B+0ncvs5iM42De
XVtdQznLdv7XA3Lmc2HLOHAl5N/9LllAUZ/Chn4i78ORWHVTL6bJN7CKkexeu3Ly
X+hGVt1D3n5SfmAbDCSEIvQPxuMJbRhPi6n0e67Tn8wH9gJ/XMVvmkROyv3SCBMS
kCmjumjDYP6mnq+5GjaWeIaICgcNoFn3vaNAyVROKczCccvW43h4LbOfzZ80X3ym
y/qI4GyqyfFQ/8QROMlzfldxM2+OMibYGill0uVlu+IyhO/aG74zjnzXq4q0BZaF
UTwODrgmwqS75lVcSjzjzi4K1tHcwN7514HKC9NE1pTORyv47wypK5YauWgaK2wR
dAljCyEroAgL+GfA9m1pa3d/8+jcS9BBZIt8uVCpyDpVmI8A6VeHuNZ4ZeH8Kkiz
XgEWMES1Im51ssKeZgzvpotyPMiUrISAEGqPMYoLzZagM0T5pye8beuLVAmM0OyF
s3lf1iRxYBU/wJCcy+ZtdWbhnFy5gccrBQp2ead5vT64u2QI2k6esWmT3D5C4Zfd
ZZWfiOF8lYC5m8abw1WhEeDpotsFknSY3p65ZJ7CReAw/tRaTJRWJTXOZNoddUP5
X3Vh6vJJpiqCylDWp8pybF6km8auO1dYdhkbExchXO0a7ljjn0GCJhrxSeHxozHG
T+w7LDmsmG1XyxelBu/hHVJnHYuV1z6BX6If4EGIi6OkO+F1+u8EGC24MirM9J63
rWujmyQR6hSp02A3pzBzFKLTUyt+JutmADdrl4BZYybdWfByp+6uN1k9Zl8Y1M2r
JDzKc/MhqjhOidhx35ZLHPRb2KGfK2drRJ1uEB2g663hK0sRgcLUTHMMO+aahFgz
JH19+ggHF2017j38oc1VXdoGJzt0QSConWvNwkkpzKrWsCfrsdQq0Gl2zMOA+1Zw
CywriVUDfwCM5ni3S5reqVMv55WBhgCnqYLWBevwGraCjVjc0p8/A+baIlDQZ+1J
SHIaaa+2OdRMgYzK4a1q4yM1ebElUdmaxx8hBM7Hu5OOeU7HF58DMJAgIsTVId6I
xyWgWKdSptfUSNF8RXhPBbVznBAmo90G37/QHnJpY2qASc6kTekkLWQQqvBCYO75
sAk5+y0Mwasn+vnJYnRS4TdmUwa7vA65XwughIkPc6A7/F/YLapfwygJZe14QtmS
Uj+3iHOCKZe421qYtAdE5Li+yGTobekoAe6eWJTk+ED5XJCBoRU2DVMHPMIGi0SE
eYByOR/X8OwTT52OUKBm8Fm94P2Al9YFztgFEu9s09ZWXsjbWBeShvMOSEP8p548
mgNRvWl7AxRMkK4MMVgqeLqyqB/W1yMXi1FKQQnikh/mkw9e8QZvOtw5xB7Ejveh
YOawU9F/o2h/EzXG1GghDrBnyDdr0M7ICx2B6zTogza5GvRxf6fxfWr9Wbikq9qC
3XAWnaRqojb+7vUrdtDsRzAtmx61lvNBRnA2FuHUmRcrbtunIqRc2KFN2wTQkCOV
hR990yu9jUPdJpCo59sYUvCTuNTh9wyg7vO5Gpks2gSBigg7Fzh70S6pi8NanjAJ
CFYQ1fQr63HgjijA1yM6HyaziDORi2d8Cz458yELQfH/jYH1Kj5RReCYPjdBb/pd
dw+XhKG0tB8cY19sxgINZMvNmk/jw0gV+mas6g5aOnDT5eLfobGZo//26A0kTbX1
qgRokNn6roTEEKIkkECTybyf/PeKUM+tji+f5WIkluaTfdCEw3OpnxTVBNlF1qLo
aCNLKRFU7M7yDrG2McLvqbuAQWIAay5WoPYGDxgiorGPxgL9+U/SQG7ge3wfKrch
NVwjUgZqRULQmk/Wn+lJbKcy9XP6xYZuDn08rqTmrPl8zqHviqMSyHiDNuw5pGi4
NzMBCMd7tH5EAWUr5M2YpygI2rMflcy51k527VSLZna8v2lV1cw7S4jK2cFGJfge
mZlvWdHxEN8DXkQe47MjIf6B0ItagkAAXgYBwkjLF1gHggEHc+9LKVaEVpGvEe47
t9NqaPqXJCFWbKem8ThtaueWWweC3XIliebkIYqqlXeIhrUg8xu3NE5ifNI3MpP4
DghJ1ebdR+Rgo8nV5DIf4bjGkkRhhN4NCWWalGuAhHG0R/GVctX+jtFR9+hr22qx
SWJ4MIFJ3OQGvpZM1/fwx7WX1woc6TfIOO4dt8v6ASKyPrmJlAPfMEX1PXxlbtL1
qlng/ZXQkuQ5Fokl+oalC+TL9TZLdUPW6ucgTC3c1kLUOltJ++LOCezeJ+NqfOmQ
esIRncUxgy7WL/Kerxb+YCCByMGZ+a2nM5n/JzoAA6L47EzSzEcoUEz4MeDCGeit
w4J4t4r520d/PI12A2rmBFEHfOt6TTgbhev2xsHj+ydZHr6sBVTnww1jM5Q1E0Ao
WHbGCtgj/USs6djwnx3VVVQb1vnF9WdaGDekr0jkxc6XCba15+8uFFPNqLtDJ5zL
PJVsmU11GBjodusNWcEDfk+XrqVHypqVX601pzXGp+iYIsR796hwgbPWxOU/srAr
rqP0sE9M96Yz0W4nD8rVUQNcNIh+i3erIWVuhuuD9wVZwWV+Ho+t3OGSG1+zduG+
ATyHXufj8mBTJQcI+1N4rcBUfVo/lzjxETnzrjgq/059TP4jf2xtUzAmbpEAsZum
Y1Nh//Z9+cBDyNWHVEmvoBRTstHEG5VRT1d2lUykltAEUhugqUigneRy9sAPYriw
cCJvSIXP9MYSWvuPup+79SZ5qzmIbkBCdPDt4pYNZESYdC5iTm6Rt0fSAatCnVRN
3pUrZ6EUjc8srdidqEZxwtpj8+dpVby6rLfELFvfpTNfPH5lRKHMlEMUzErxMaue
QRUibwcrs4Mc6jTM4KUs325ScGQR6U6AdGSVYn0UXP5apxas9Yc5944+r5tgNJ9j
wxzEvweeyWuEg8i5YchgFXogV2cb7IodczPgM80JsE/Ib+UGbFaJxIDL/8PGaCDQ
lmpzrgEBXWryXU5FLx/4Ycyqj1uf3f+Y0zw6v/p9aFoJDvN7sqwlVfKOYpaEE/HA
PYokS4P7+f3q8nems8IWaZAFy8G7KTAGcBU1UmQ1OhRCIYHOHuSibwM2tBctAnoE
4aIreZv/I1D0WER6I2fvrNMcil/8mYV/zQKvYzXi17ph+XVR4Eos8XANcKgAlIR9
NFkBTr/41Bv7ybIVr0HKVEy2QMt05Ll2wSb38iOP/pFCDgO9cDv/6ks8vB5Yf/XR
GCqsqOLOLhOQunXQ0YTOekhVpdoWG+Ju/WAGv1XXPMIzQ4+Cm4QwST+nUYMknNIh
GuQ3nXn9F2Lnj9liqBbOe/QjDBjA71yx6fFNZ629nq6HdKy+lFPbi2BADi2+wXEu
EcEu0n53nBltjtuf0n/NoeoaJoQd362342h7BHYZ4qJtwnJVkb2RtTrDMpSEGToa
YOAcWq0vkrE0xy8y0LCZUHMq0rD5rPsZNYCFLai5FV0yM/2gpFttOylxzKZgBk+M
Vv03SXWf+Do1NcFSqTAWc5hd1pVStMqbp5osL1Bz/5DCkA1AwAD0rPUK5/L0DpCK
Pga36r9FcrFtxVKKtisdJc/5zeHD+1Wbu80MXKy6gwiRxMcEMfkm08fExDkDlerW
WGJbdyp4eMagbwvwZ201bunxH1/+lxSspB9eRwkuKGrLS9qgM4a5blz6P2Z1f5IS
W/YoGL/9IQryxxX55EdDrTB6mjqO5ruV1yqrvhWS9cRlo6b8WKiGkileZOsujTw+
3U9pk9/iYEbEFNtRRs7T3jZPw956MjTX88Y05pGXSxX97HI6BW9nQEAJztlPYp0n
K+B6XByiBWnCqroSGVb5lbX/bQXtGp5lq9YDNd5KpAWXT8QrzGCx8cDvqtj0e+6D
DP0iu/O4JBLXDanLvoXLkRsoPgb6jQoSR0Gljtt4kmJN564yCg0K7tnUynFpiKKR
3ZWZZIqw6FIquj3P2YZ9k8qaAQnvKYtLN3q20Uu/lubni3kCqjy7UsUZBiPQ0eRb
jwbXkSGGvqYAOj5yDvpk5zIX1aVrZHVpcmsUe5EzmrWFh3ATQ/awhtxJpkldqJtf
jJvv1LTB90q5g1usM70q/yQrkDdFhnCVWT5fuJshappxq7ESRDVnxz/NfDAqF/S2
LXgITSazMm9/SCXPA5sK11yPLtAzxaXgQcfZfUJycZxEyC3fzrnZ/6sFwnfqtXop
7OfKfiReoUxL/6mEbKSoB/2KE1GkTVbseZZ7WboZFM8AyD2p7DAHaHWnZNn+9vBg
tFK+yPnJgP1NUf+z9DU4y/1rywYCnkLlqXu+w39Z5gTk1yAsiCUpXpnszDUkw9oK
EOQMBzFxt/+4uWMWAuiFHP1azGNR4wsBgrNwTaD4PNQO6BNQ0B9Q9n9vJevPleho
TsXK99sMIrfx81WtmpnQZm0CsYHDK7UduuePBC5kMMMFaiMG6cWQ7OYTQSgHdfXN
SpsIFMBDv/7VP3GvlHJ/9aNaoWFST+tTPT4SJVGdIc6uslIeKW854Uww3dtFItdk
3DuXL+l6fLwL0iuDfKh+Af5vHo6qVhZrJwmE2aBebHhqLm+RFJY0TABFDmv+cLL2
YzX+mzXKiwZKce/sHWuXBFIM4wT0vfxfpG1IP56nQ/WbU4UxfROlXPH6VRNpD4Xt
+GQ8TYR5FRNRMkF7bKftF1o9XiOu8XxME50VXKcj19GUnRbTpnLxD8DOBS79tmDL
o2Zas2a1PjGJZpdisN65vzvV2A/6ZAnkVER6qg/wOg3tNJHTHhuzMNw9hdFxQzYT
i7hSVT4+HrRYRLDdPyGeOD3lOmGp2vs533QcoDPanHnvLrSzxTY9CeSz6a3Lp288
8aaJIKY5NL0UiOCdoCfEfTbY3zwyI+ts8eYMi4L1Pse/DkJ2gKDzBW8hFK3RZyfU
AZnwB1Owpa1EIE3ctW3tTy08qUqMlt6W8bHvQbmBRkBWxhnf8qtEEwW8zyWQk0Gf
r0oC+NAh9Xg58apgbKLHmtWOeQNLD9PsHtvZooU5aUCbKVR52PBtusBId+mKd2Ug
t8iTcwufOKkJAc65w6+y9CexCIrLE6HOx0nqH/BBxLgfkrpoMoZSJCwNXLapdURv
14RTlUAB6wLa4mGhX3RL8sAqhv/UPa3w0mct/a4WebuZyngsQmHUbbrYOlmQAbtM
8REbJDwyJwogdQ+6E/fjJKlhE7IOi+D1PRMsgN6z43YJrWetnIasYjOIbI6rq2mn
/DjQR7uO4gVZnUkg5pEWP6SZU7y17TFKo79ePh3qaME7dlbT6mkDF7mI6muhfF+R
aqLC5iH+BZLEhGznG7f1TGKO7npxH1ASwQYP/SGWJ6dBlUZOg2M+9TpP5wyfRemm
m4KsNwP1fZseI8gm7aHv0Pu4dVUNkpDOkLq+ZChI1PAzxo7zr1sm2RoDOlOaPJ0k
KWD0FtKW9vS5GpKFZTJ7aI5i8RwZAZK8S8Z6hA7H8VMnvEQzdq6ayBNSDVSRCYgW
MJuRucQzrlblK+uNa225un/SFFCDajXoeox1+kah+42DIzGYw/zyBcPNzUrj9KTJ
/uAyHnp2MO4SRSNx8gGcrUV2Ou7CvXCJYyxKg/fkzDfXzQxQFyc6o6PxnwM6ccRa
ImLqjmRxLINMVj36EEUeujCv+HuuHS6+VnXYBRD0PcrM/9VPJRas8j1tnYPf5pva
Q1fM7Np1CoEi2LvZI9QtfM06cPxECT0y1y5Fc+n1I4+lA2PfTjRWeKt78DDbF9L7
aHJu76VZZpFbHig8HNRv80l/0p0zLraWiHgXyaMbus1Y8NLAC/JrVFfnVEU3tz4M
Z389OgdI7f98u66i8lQYy31sCor1W/sEyGaGZuS3AstvLK8gEBr35zkX8tWsjynp
dqQp0+Br7p+yT15tYK+1tx09zdYosf5V8dW5AkQZ+kFcQob5HLoWme3/dI3AzRWh
0Yn9hAe53cXj5jOzrB1eW3QgI4G6HVlqGNN8lRuDcmBNgIEMT6zc+L2OWyKTCAfM
mz6uo2W9xJF3qr2ZGBuk2Fisjthw9w3gTmqXO4YDg7c+Gw4L8uLx8ua7wB4agCRW
JJ2DhRrawoQu/X8/jocF9W57Oe58RYIDHYd6uyvqiA9nEO2QwWKMbBfq7E7NCX38
13HFn7QW+lUP/ibq4+Vk8l/ScM9S/nIZrjgqD2vBZ+uxCYU8MFYJv/i+bi7oerE8
wz7TxaDExjIBj91A0wiHcDp0otdHIDcvPutbySvSaWK8H5PIEwmv4VW6pHy/QJil
IU8qYsisE8eV7uwLbN1rvpr5SmIk726ph7wl5YfdrsAIAUhwH+Osq4UTajMbXhKL
nilu6AlKDgyFsQl3JGTK9yrkPq7tcy7qSXM2MRjYVArUNxMtNXaQwPCj0DdeA6Rt
OzuLpRPxFcUBZoHLe7VqBw9P8pcQNrUKQDXI2YF9bDLp/fCm9BAqPpg2L0QP4WCY
YaD2L1DxTSH8hS61RlZZYvQO644TWGjxMhiumBWCPno6FdDLooweGWfkSBtq1vQK
IIEQeB8oF33jBm+ZL0iVRaP3MTvHywhipIxdc7WARSX3jOMpmpDOaU4CLHvfUMTv
1Y1ZweY3iTtmWOINBLwhQom5Rg7rChy2oQK89W2g8/iynoqO+zFtsFdPQvxhlOzu
/BTnboUObZ+aqayDPNdKyaJAf1wa4dd44Tnq6gZ7yV5ZY5WMROef4nhlWvcYLJXa
EbM2dqRDWRY4JhobSUfQt+zCpR1xOIM8Xg3EHRWqBndpvNF89TUjBN2RX3w3vIWO
icQra9tA3qjVuXa52xiH+lvzDwAhFaNUBNtDiToFZ9w9Dcz3zcAuVYXXADafeb5d
pyrrcZVL8wiIGL73XmAlsLRfXclGMyW0Pdn6f0O0NH7AfZ4G2gSNHXukqlRjhP74
8CGLsrbO5XpxuCbKNQm/4hXYxfdrZQFHFiyrr3QAJd6WfnRofoMLlz6K9oVB6w6V
XU0gJS6ur5cGm1Vaktgyg8lPKl9uIaRHfW5snLcYQTcuToz76HA3H2Vg4sVBLtjX
JX0iqn0EsKDi2Sqart5CPPnHjA8sWhvfItv1mrDapQGp3bKlYZce+LVlKuYjFTxp
rlX6EivO+nCMF8tUhOqXdb9DWu4mbw3f/cXFx7BwctdF6PtevSdmzprZe8KVarMI
iBE5V+8NNQHt3qwm+cBjXIPdmYFsx94m/eMASBkvs6UkmeUDUznJi7ykvBhbnu12
h37EaDzH4d/7JxTjP6hHbaO5P/l1uPLawwG+nmQeMPssKQhScPkl1L4FwCX95tU9
B3Fnv7jHpXB1GEQSQo2hD8M+t1YbvwNtUZuE72UlQ5+DDZpqIXPqMnOlu6BaDqp0
WywW4JL9VuDW6Xwx6FKp0fZG1tu7uGSfgYbyPWGL/qCoeseRkUl7DhDwMdvL6GW7
ZwGNXs5qTLPSDpEr5dxFHoCbbbrlsfTDxP8l0T8VerC84RVAN5FK3zQcZa5i0a7R
D4xgI4C2QjgiJtK3PJdeNZKQ0SYzkvc/nFYmUwq5Fqd+sGO50a6pk4qCDbda2X7w
RE1ILhXUkV0BbY+4qoNBKAuX55zaFw1lQIXL2nlE8IowN6DeV4b30YV4HuvZIf9x
78NGykVQYKZO4+8tzgh5Iu/89llnqv5nNFd/NOQi7JEoBaJjV+E4FvQE5c+vKYdd
kWW2d6885PZsB3BAxdnLXreHTNV/kzq2LamEnRiTxqmUZkZvcS0pidKwVIXD/BCS
5t1VkfvsHL5WVYl3lI6Q+xiiPsNrCwyB69sjOvEs2aRymQWWsqGN0Mq5vQIMxz5f
Ud8SOHKOPaN9DWHd2xXbwstrMZ1wJBrenm4YEgYkEBwpBo4KnuCHYyZDIMdsWGr2
3PgkEg+edF3xUZtmW9AtIjVAQ+zcsJ1LCUWeUNr/8jieteQOU1CiZKpvEUsghfNL
460Bj9TDcohhmMMIMq7DCB97BAuHzZ2pJIsr/ncyZso49/C0mUy9XzyJ3VxxOfRQ
w218CQ2tdbYPziF3XVgqK4mjSooHn+EHpJsIluBIod4pnTbXPeZPb+Zhv7v+Zc8w
gDKfKdUk8l9YgFC0izl4XuHFFLvxitvwXNXdtBRAk/3qDhHeflCW3rufU73z4Mf9
rY7CucM/MyeiieqkME/9g7xGpPk9GLBVXj3hWBxo/I0DJNVs/1ldzVG1QByYk053
i9BTlHJIOPNe1qWeyZRVgdFudyjQ31762OxY2pQYFHAB65udzEocjhOiE68jkGAO
Wytzh0mth7VRVmbdCUo/xD1DVWiVJniLueWfJoHJzfEScP5V6KRfGY+zohRvkdXv
7wEbu7VMZMchjuJfkTrEd5akk6zwaLlZaVbIJAZCS79GHJBX82YaF7eujtY5hjdq
t3Iflu6b86/IdXlV36KRG0wbGi0ZJ0Cp/stfpjRNV9YcgTgdl3skre1uPKCktuu8
2iu1FSFNfl5tkegHaa2E0oAaHRiY3X91XYtOHw66IFGHIS40D10f7l5Eq2F0UXWg
9B1JcQ6NxyG3jK6BvVTof1iGKfwHZRwHg3Jz/acdOuL98tpWAlKGleVmwsgcpr+j
pkuSm/IlIwTuPm22wLLOA8bnewBxiseopZMaC7h0Gn5exihrTzzepZ2K3Dl7K5r9
vmYOf1QvAzVDVsGrJlxng/GtDiTlWI0hXCCSi6ZdjMx00X14kos4QEImMEZLVfzs
a9hsQDNxk5wMG1rMukWyXTSRvJI1YuJB3+l0B+8SlkGodXxj0bBzve1APNf5LeH0
E9F15mmHq/SerCHLcpG/KdX9DoO2loJAVGe0gkezUTe3Vy5Z4wJ0kTuGxJACgpX3
KPE04nzaUK6Mh23PePIgdpM++x2Of59nM1o5nG+w/cKBrUWkTWA8G/QHNVJ2HFrN
G+bIv4HFJEK/XzDQDOLAsyd3WaQJ1JC62F7fZfgmy4rTJWTTRWG8ycplKA64CuFK
jAHd2+o9iZlnxrK4Hxd9PIpWof3Js5xfTrS0y0HUL+8TvoSBG6olOO7J6wr5fmMT
87iC8bw2R+Jp8R8OBQZgh+7RgLQ5KM05pwChQFBtvZ7BJg8Rz2MKBzazXDVd0DJ+
BTzH/AU4Qx0wSXas0oGsJJUGoO4Rf7jutGZhjqlRzzBAVh8XlHc39oivgwM3KGkV
HWhaOWW8qPInbRXSZzfWfy3N30P9E8AyXLlwUcMI/uKN2N3NO2cEnl/Tk1PqEaCN
phLYhwB5as9XxiYXURSxDMkv47zusLwLY0npTN4paAzYhhO4FtQpdsOEaY6cksjC
zljD8jUzZPLTwyhksT4Tf7OqIaZ6E0rwJdxiRfIQLbAhYAZ4o7SxrGf04gRQduJt
+i/u/RPSKWSNQTN+JHO4GA2050zyH9sc2mNFKDe4mZo1o0Q89TQ1tQhccfp30MxE
225KRrSTjZtVTW31lhNrvIgZvqF3dhvORe5TP3u3Hf0XNfg+ZbphW+NMUB9OM6es
srekYFGjCYhkcJ3pE13SdYvvyLXRXFQetvQp7oXuI1yXRMwSKaj7CmfUX59FtT3r
rUMNhqP34yD0C333RCR1IkxFmKkfU9HeUuFZWBY5rU01+nh5uBAf4Rq5Asrfs7Rk
LAqbGwN2nrwsY8vCJVzuoR5sYlUBgHQ97DepQ8o7tXshr7mrYkWWizbCefWWn182
rp4ZAqb4jOVfvYIYf3a0PwXK5EaUiUbdtiZIcOQI+Rhh+yphAC1qyseU8/CwSCzC
YF8V8RBhs/YFYYKHj57TIz3T3rswx+mkUJhX8Ev6tAGS1Uveu7fZSm0lqdPBB486
US6vIBUya7kiAKQtwespWLbvLBPflHtcKIbkEXp4FvbD6IdMKk5HteokHetPxslY
WePdQTOVHVoGC3a+//zoizcbNK4ZG9vxwmg3gPjE51c4U+Vvxbr9RYWqx+HW/ko8
M6e9RvW6Tvm3pWkWyp/7FFzdTy7VTRrc34afVymIFyv3VTVnUbsIfQqukrDQUFqZ
awE2HkuAqkYK63lnEqRo5pTT8U63uAzHbwtxL8HbV01CXjLEGh49iO9ULnm5aBpn
fSxAJDhtJ2acqOmkCJ859ZFLUzQnOu2ouhkIPHeMZ397U3BThv4sjlBoFFhD7PUa
v7C8N9aehOOlqXD14o0GlYXM+df95d2ey58s1ND1+CbuvysTMVu9N+rbSb5FRFGj
kNQT4m/e+zso5h8iYQLo3OvgHlXi9D46Jl26wqApCrYBMj4BnVfa4q7oGAlrr4IM
H77JE9gdHjA8GD6lsrSwVCck4L3CjE3vyCJLh3kHIV6+HCltuO0lzpgUeq9Jp/3r
pDiEh0duh9Hu8aNDEjH2p4bXwEpg/wwq2T2Z787xPRgO/aYDbSTsrvXblVsugADP
AdS/FbhFAF7ciAFeXkzmjdsn3x2RBkRILtumngu2e3sLb4Mic36QGY8TGbo6EIrc
m4XVvRGB4KRemvGFklv3y3HkG3ye6aAFlzoAN4jCpeV7NusTuKErQBp0lR5GwVCt
M3ttmL9yJ57+G/odYZ/tcD5C2YfyUxE4eqguKW/5moGOkZNzFVR0Q4NG3SHBSreq
WdlDa3sW0O66gV/2fFHyz5RlQvwfWHi3WorLTL/FiXSNu7Sqx3WtaFgFx6MBdZGu
+ZeQhuN1yyRWdCqWJHmc5xBzOytqsC8eVuI4vbSKVJ2uec/Mlr400YRhTy9ar+qm
Pv/+IkDH8cRMXTH8bPYgmpnQ0c7Uet6TZr9sHY93dZG6Xzx1HmsedJSpYkPU64kP
7AZZUtEmuAhc8jn5IRL5x5Cdfw/sCwlg1NGtPHzV2RmNfuFkKgPKPERO8ptAkW3Z
o9AefDjXHGQ7klAMPTyhhj1qdNFZcGx3GT+FibYL+1eptenfMAv19QcGaP+i4b7j
RmLWBsZcBDQkayI849MC2WPbSrmG6FawGbgDCCXqgoCsZC8/3cshiLOVDQSJKs06
jvXfxzzhT6Ub/dq+fpjnq7JYaSThYeIyz52P+fbO+nEp2XxVQq3gKnJuonCc6atb
p7rp5Df0ZC/YtGw77BA8kfZoxQuk5RMM8F5IMje8mGQ9YjZkcusnmQRZBnw0Ctj8
p0n0VtzEJ7u/rMe+ZakVzJstLd4pEnrYWLl07R2JSb9pa9xokxXk7EZzIK+Vbzcr
HDmnzFlHfaKp4eEKKCus6OmfFtKCddr6E6YDp0ayWnpgwwPOemcQEb0iYbbssq0O
t5OKPYebHNXUXJhTaCxQip/Qcc6s9OhR/4d0PlRj2JtQDJ70UYN3K7uP4fXZU/TH
sUdoBzYG+gszNBturyHiKZe8Sy3DxszT2vwb90h/MP5fjO0lDgYWoVrgEPij8GCw
6S95BeNReY/xxH/IdPo2NY2N7+ifiJTmAQhnaChLdEjW16myrjNDHTSjuATys5Hm
Nt3Hnb/nn1SEpJsDwTq/8w/LWTAMlRKCvz9sTWRR4cBNUYAchtRoDQGRknpHkbl4
lQYdnXNeacOSi085skNqoQix7ZKgePAUfhT77VimcuzvogM7S1G0FNg9cVbI76uq
6qDbMGIdVSr5lxVHQ9dGBcWQqH7N3/nUqxmrSBgHSMWZWiochQ+oeNjJYAuosgVK
UYYsVnuPvAs4ZFrOnEPrIEg6/zVzM1jrjW6XY5GUfJ1GIcNuNDsT7vJGQzghGnKt
2zStAq0yEg02qty7aDZFJsDrLdd20mEV8aaHjv30iKPoEhGnpn+ycMtM/yweh37u
SVFO82B2vck5q6wXLB+TFun1lFri4BY9YiCj47YHqdBgfq3UCo4yRlj/iH8hIFws
FGDzwi+E2t+58aWfpTQPJqsRCO/mEEAYRiYLbEr3RRW+cl02z+z/ijp2PJMzfiMU
gGR36TS4QR8x6W4gq9N/MHX3cIpGu2C6jlPVjgfJycnvDujlyXW1neeUAet/Zr5f
OCSYQrwmRlwRMfXzvRPtsNaYdUR8WW3DPpNwEapbl7j/DXt60YsYDIMOd/KdCAe8
yOl/HYaXKFv6d/uhGsEyDaJn2DAwPqDZnG7P8OuY1Xio7bRM2mbj10TybJH69l3Q
hKgpEfdQjO9BFJWdUrbay9kFszxm0ct4V7YCY4k5QvwH+CiktkkD5koyPZwRc8Es
Tteef5OuFyhiSCNuNk7+c7VlftsOwrbw79aAw23YLGzNK2RMMN4z5E/qsTp8bSxQ
A9M39uWnHfibKET881wDGZ6ygQVFl40vC19F1DEMMToFIyKDaZdV608TavMZS/aP
ha0zhrq5yfXtW1TsZXsgt3sbxfUVYBzje4+2SENC56dOq2A187OPIZppO1prOQk4
rAQb/NqJq/NiA+t9Frta73HdC8euNo9nvT/4mSwHdQaK3EEJqdmjb+v1D1/VkLXP
HXBKPUtgsT6j58UeKlnrFZ19cyRMZjp4+fr5rzq5zZGMSHc2yjdGPV9lz+kYDarl
OFOq/HJnPjlFDVE9pRWLAyPTAaQDRBisINW6jTmSFBA/shkJPsbof0M/BLal7afx
IMWxMGBeaZPmhEsuW4gB88PcaAn96eXaQPuXcQ2zM8qpCBRSgLFcVpDHfyVudSIF
1gKF3fk0J4i/UgAtfqlCVqSeKhNtTPDvpcIbR69nFw2EqFyO5cFs9eS2XsCK8aES
1XnOWMZYq4kWccofoGkN5mXffTqMZAtRTQqWFJfiaCsnQsICCpPUrKA6wtceX5EJ
vJ4X6HfGlkk8yrhoE8tmHOHkuhR1QnhzMPEKmCD1Wb+HfbSaj8Kj8Dg9RLrzQfkX
C6jXOkPfasmRKOBeHfTUU3irxJuZi2svVB4xNFPv+cLr1xhVo3BJTT5Ay4+qBLS4
m1rT69AMrZVRpZNMfTFp3HO0ILau+a1ttyqm5bzGq1FfT7bbVlT2qFRjxefFXhF+
JLpmRU7iuv6WLHtxQGVnTBTMhIVTsewXvOsIMVYq8n2XKDO1CCRVX5dFaN+lYlCt
uOpbgJwNXJEy4jIvkUk9BkTsp4KGowlFGZfoe2ImbIFs85j1Qaba35nUj6bkfVch
uJjAyj3XGTZqdtKislbL4XRzsn5TkFRkYvvD/OcHvCVyKtbtpj4UyIdC5QWP1/9j
S5jWLPOBbYbbPEThOvRmhCyluKrcVl/H7mTvd102rvr5PeIO9YLzur3gK5M5SU4D
rFz3lOBaC+EYWTPuf60iipDWVAYBv0exn22WLv0bePl0qnTwyWzkyQRpaFfrvDgU
sLEw6JGzRBfomg9oN1ghLYR/gsw3OCnLpyvy8ZphDSvA9eKXn9k8lBoWe8J1Rs1r
GPvxrbtuCaop10DTBWcg88baegtz7KFFxBjDqXSmb4IzMZL+xStjPLgbn1V/w5un
Gm87DxrPSycnpvjvTG+5KGqnp6VFWJEhPHH8tRGnAkW5D0TXaamMdYQ5LCw6t7XH
TTFnenrr+43tRJa1wZjSSxy+DKOm2Mj72azNQ9nRGS0Y7ySIRwUHeVxRnNBKxUMv
YO1xRWIgvEedC7cxMN5+vopgmDjmpQ3BEKqZmEc20HJXGKhvb7so84QM0PWUf6qu
hZ/NIkugL+ZWApgiMhwSajW640tEkopEfgEusemnsox+PeL+QkkSkhvNQI54ggIe
cqNvyr0go8Oh1DzQu8ikktJzHvfmWVXc1cOyOCXVsMmBwmkC/a+L1E2B3OgB6OTi
/+dJtwA3b4K1C1KvuLKKe0FLvPcqmvnFasiH4CKVGMZAaSXj+kbIyxaXPwipDyl2
8hTBiAu3eA3xtWcadxRK7z1Gm5OcTHNH9km4u3C9sFz/W0SrFKQZvYg5pVTv409g
StED3MmnHaTVUjJBeZjaDyy/qnZlG7b14UhQSoD6E4pUsmfsxuocTNoiO0Kh1464
OVShhXmF03foJ0Urr6khzT3DVOYNgc95OE6W8o1sdGDaohqBlVi16cZbq1YweKTL
J09qeGxnVw8T/sO4z+ap6hPNPvbFW7kS2WQ9dnRBdOPVotVPSWwe3Go59c49DgMR
PXhrSXNRGu2GJHgmu/Lgvbx3nXEtK6Shln58Itp4W1J53riHhfGOUYQKgbv30rHH
yDMklIdkdhLI3i1+8zipEr1W2lsA36llLgC4oY0ql9hOACJbjEqZGyvfPylrpgbH
LXgT3vWN050r5klNdBM4jET+WSSfc/RlNItwtjgfaqEpVXrsY5NJdId93qWJgvBH
LI3bMf4RN9jVjM6c6LZuRONzcg0K+4DoDI5p+/DfhOtII3Z8QUwTY9/2ceSHLy8e
YFdylUMBBild1pnq1+KkesFTat7D0mzqJilZoroHa/kIlLOXaNqMG6Rf5Gav0GIY
CF8uTevCGlhTAGurUTX+nliGkqnFBgcO/m9aWiB0eNjDCm2/ESu47ix6kd9RWERF
0TRFFvNVHL6e4DZW4uIz6t8zPs/6NC2ASoGpkR+a9M+SZE3SM2HDAZL8HxYmFSc7
PuYrta+A9mcSfgO6P2ODjB5/554lBBMLl7+Eef7qgsJqXJzTNTkKKsqo/DvK7IlX
LEAen7YhBNBC4+8+0ylxKJGIhJBbuNdpkay+p836O3ToBDGwExMf1KIpIr0EeRvQ
buACVQnhw8fIl3SYr7BjzjKIhVc2fTkJHs6ggSs86wdHooyepyTjwEnSKqHdA4C+
cU/On/BM3Ams+Fw99AF86H76BgAqvrRciNzQ+ju8uJQBwAoTTFhhl0LpEwbreOyA
B48tzLxIzXz1mIPoDCA/QCvOuFYGUgAyPdTAR9el/XsEgfeEOkgHXO+hz0Qr3wl8
XK7Y+ZpT+ddaFsuR6+V/Y1SECwgU0ZazLcfsBkKUjduOR/gxr+E591R8Ls1TGK2C
WTlW6nB+3jMefPXBuA0KTP7WbI5gZQxrf+ansBfwAHzHCc54aBzrDu0w9RE4UnI6
tmyxy6BkUWtLBS65ayFD5aBJXaxK6gd8haZA7IHON5v3u+3OPlgQ/UIWI6qyqrAB
VhgczgMw+YWatDkZrjg+J1Y05KoWxMZUQfG45RSBRy3rvxVTbREtSvNPGH2F+L3D
Y2E9eEijy9fYBVRyi7R+YjHdcngKa4Bb7b4cFXI5vEinrSBNK2JaK2FvWALGcdfA
DfJdMP55E7bvsCx5awhQGeQsM6b7ywdsLfQfsAEqkfWz1oFhw5RtNHYygb676f1c
lMVTG3TO10iElW8nvAW6H38AXElvLxoHyvgnjIReyGqWW7mifzvm/YuiaMYL2+4D
ErdvFL+rlK33/+UZpQvX9ryNRCnXFCx4nfJK4sKmOP4pPbHcuzkeiuNxYhX7IdnP
cBUiIcb+J0EkUYPHAVghME0Ib6MXX4Rwff6SEaTT4FriO9FWE86rbTUC9uIJBIWR
El9E6BzrbfZu6xExRcKuGkOklWDUMBJDdmdRDIbUkxtcmKIA/380Nkykh3u6ETzg
Qmvf2f8MI7SxhKFlqX6xBq4SQ3199pLKSrbUdG5msYGdAaDzidmQzLRp5ngUg4BP
B2qJ5wN3GyVeNkuRbHdiTbH4m61t06NRwtOZ2t0ACtyIBseQnL3QJ2L7Y6nyOphB
FIPo7Ne8ug86KR7Js+eps2jCD8NMVZE5C2C+6ap7h6VlzyRMH1jMIS0osy0uCaX3
4HSGIZtA584Rc+InUZlfc6cv4QEKXPSRxV+EAyevJs4oTzrjLPbFOqMQZSC667zU
M85yYMbCkOXGWofBz34EXZDGgoa45UGdExaPRQChKf5Oezw1/lVQf0iPaQiwdDuT
8Bh/M14MWfhbJpjKlSc040qTlVmbT7PQTXewCLUSnqpq09wpgmVghx2GbV9Yt2Vw
SnQy5u2bDA1KYZfolfDG2xZOS069uX4jldnN8fwIcmhTU0VUhztrQMOucyW0S5q3
N3hKoeFwMd3MNJeCtt/yLg==
`protect END_PROTECTED