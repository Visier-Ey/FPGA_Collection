-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "N-2017.12-SP2-4 -- Oct 23, 2018"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
FI1ik2Asst5T/aw+S81cYI616d3kodu7q+EaoP1JGt3M5wstNlMSS8DJh7IB59kH
24qMjBJUodnJzQGgJy5i5c3yv39rxK2bvr68xnLYveaQNWs5GOPgSxwmwqW3fMUw
fUqIhzeSZmi0KdPo4Io9P7zmE136d3oD2ZY9knb/Tpw=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 1680)
`protect data_block
lN1DUwpChfQSVyQH1KuY781MBGUakyJH5YbN66RkFSNrHCbUOF70cxaIgBvy8wWT
S/9xEMg4g6OfFJhAcCAl63SRktWlWKtydMsFlw5rBntpEiBVZQ9+52EJmNzhsqy4
CoCgxAdjs4ATpWnyh6dIQHkiovhOp3QlKCviMQB2f79BmYcdX5zfTrKSVSk5vEye
z4zIFmmY+ISc+GOuFrdJftnDMVKEDnJkU3e91QhcZ96PtdPdGipes61dPScL0ptr
Yf4k4L2tMRcpDdsB6soSPhpSJdhp+VbusiklhXNYWbeR62ES2BqaI5kwn8RGduiZ
AO7T3Na8MnoyTScxGF3w+3oI2xL2AAXw50QxmKZNUsYhn2YdrPcYc4qQSXIvuqG0
r/Y04+ZwMCL9FALjNA3ZztFGChymvVOwVYxp3YWnp8mEM/4HXuhEMtNVr/TXqgpY
KcfAQPj24CxbQ8sjbgEqdyMQlJ/Ry6RE/A8pKu7ejiSYr93ZHiwIPaYxfcgzdfMj
/F4MTAWVk3wvONbY/jNHkU31bfqV1L/P6xFVWwSMg7kPyGNvwoOrLdW7BZIGuhb5
fpN/S6HRM7GcOmZnI7d/rBCpOaK38CzEb12+ctDqvc8T9u7bz+1Y+7c0w61ezJfz
8rYH4NkK6012NZxr9MKxE80IiQY1QVrmRWDS3rM2dDwajmBAtDc9MNk34n8Vmoa3
byoFd6m7muSUjIdmHyc+Y1ByjowyFV26ZoM56j07jsz3Edm0pU/74a5Jjlfqgfgw
IGYCJlt7wMxZ4zspNMVVM7HTwn9ux5fpZEcDh6Gw7ZuWdLyCVftC78FpTUElMVsf
8TF7mClcrZMHdx4O8Njbq5Ppu0g+0FoR9x5/gypXeDovgb/loeHnFpfoNHLSXqMI
+KN1sguTGdO9dsf2j1nR/TBjomCwQ5yUBLZ9mfjmM/+2bjaysG4ZXxgUjEJdJBEy
wWS2M+J7bInZtwtDLPnYya1Pnc5K/PBh2WC2SQCeNcYYVAnmknXpdyURoAqSDrRU
TDivymEhO3QDP0XRpVgdGDHQb1T3Cl9+lW6Ln68TDBUTw667H4UqN6/3NbbugkYH
93ZLFrKpIJNCiWrk8jFA1SLdfqhsdWDC/dvMHbRhi5xCjdogAbFB3xR6zVq108tL
LzJr7dSrTdyB5U3yen9AQUk+Yh9yR5vyqjZu2zsBuKrvcl2TzMZh/FkvXLgArCCA
Df0QF1+sQAMsR+Fyihs/day9IKvh4WvtZWC51pInlvyFfqgU+i+PMMAxmoO47E+M
ZE20HuQ0ETdVCkPy9t1CoAq57Vceg+liNmUA4c0IJwKg+xwBpBxXBbg2duz+7V17
iMHuNY0YBe+HWbDWxnhudEjWl/jRSRAw14C02LYB2MFOcoYrsMCuxRnkzhw0f3UC
/Ae3A0oP9Mn0j1ZQwMHo8uI39CKEzpRZ7uMJOptUZYW8IKCWlPU37hhf+4Z57eyp
DDaKfUoeT26k4a1z7a2CunZMiQU40n+c6cuT8oFLSgxRAYwtnuRDOfydeUiyRrH5
0ZUVA26vXNgk0gkJZePzurKhIpKWq8eEiiR/ryodYPbYeEJ+iS6PEw/CSHezeng0
eFxSJt1ijumodUzlt3Bk4EBi5LYdaHrokJWXbBbq+TprRW/wpVSKs+zNN37A24x/
i57IlRZyVR0pkuyMsK9S0z1lNUR28a897NfvSLW3FO8hj8ePPaES0ehfk5qNiIca
NG/h+d7UQd4yhyezS5l3MqpTU1v+UjCSLc6K/7yJNfqw9ynZV0fEoU/de3jd44x1
nuCUQvzJ02zKD8Mad/kKHSu1nuTRaUJBXykwC4RtJ3vYcUTgGNS6JzmBBG/eZjpc
3mZVdf9okW7pIBkNs1+2ZzQETxFl73llmb2IFXIVMM4O3P3QZjHxuxkC72feK5Mb
NvruQosaB2uTOfGVO72kOUxyjnnZK638hkKK87/fjkPnkpfFYoi6Qul/icIkWU0z
3SCH1OflogAMU8mHze5uig2UX5sVEFQS3G72PfAEsRW2KsThDioNC+TIdJyY+ahe
e1r3UzbRoaaNiGfLk4jtTX1YhIfaNPNswvxEpFT1piB9Om8U4G+57RLElddsMOpO
Ljn/Co7ZzVLO4JlQbqyC8sv2VlWRUZizhrDr2Lz47qU7+/HJVcOT32QnBhGg9Tk8
ILaVur0/yw6ksEHPMSsnfMCX8pVhhhBg8zU0p/568ni+pugrd2fdgw8po1lIKa65
`protect end_protected
