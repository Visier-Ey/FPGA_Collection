// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ACefpqbaYroQD2cKh4RyHootXrlEKEpZA5w15c+NbijgMXawl1dOnrzgz8OHBm3ZYyH28Yfx7iiz
gZf4NeLnBtXS6W1P+KbFtqRCKZW9HjCMKX7Qtt/937rX2eFMIYVpUexujsZG2nWtSxtPXKP/EUix
qqvwRCnkhp0v79UFIRi6cmHCEMIltc+Cf7aoPlFLg6FQ7tcfsmeESJhlzxiuRHlHATmtgpdf5I7F
9VY4JUr9Bcn6QPDLjcReoy6lEpBixkpvrvlhMISdnFmE6OsTx/C+Og8MK8KZR/qyoLhPtROo2kyY
VXfgypmXQRsanzmOW684qQFipYviCvzl+WTVng==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10864)
TGHC47vvFp+p90NiF4D3voA5KcW9WOa5v6vucCzlREah8nfUjovdKXp2Oyup1oR0UkvWtrxJS1p/
f4s/RMLQGxELCwUzWd3jSmHpuomDJs3yyw4tL7FZokkUI6Q7RKraGmVf8omxiMOdvZH3sQgsxYSy
utTnJl5dzvgbUKNvmVOaqUmXTZwfWzLDhCkju/y9cKs3Qw7XDKGelChtlgieO8vtGghRttKJvjUe
i/gTIT0EINkAdsXVXuGWetDcaaH07NjEo6Cd0OGvWUoOfjPgGa0OALcwDnl1xBLOQRJyNS5qIUkz
krH0tJ4O3axSM6VICmVAl3BSTGuxqWQUbnO12XsRkLop4wgMRc33BKrNh4DhX/9859sVM8zlVvG9
w2l+k7XcxHW/XJFAtxFfO/u/HQTKon5mp/0CdqZ9QL2TSC5VQNwqpUEy8iBcUvlnjc4+oxySsPVP
fkV89wqIIUC2Phjpo4iX0IA87vFHiEGor3oP+tFUVEp3HJkjzm14cLiv6c6eo2YZG7r706oIC5gL
VK4pTADO8OIWMDIRAyHCvPjIxMQGpXTy85zIN5Qflm18iUVeT2GZPgie6P0AkYC3S5+CqIxciV0a
V0AwF2EdsVGTEUqACUxq41kXXWvNOsUizgjT/0YS5NdCXkmgZLRpu3H/tN8jFMtFu1424hAs4AzO
cT9LpOTLpQigt+WYib0cSmzj4cKUM9i3NgBUoNj1Q7PNqNuElgW/vhocY/LvIowk8ANpGn4433Dg
Svyn/kZlQ4M8npLUCrwOhCPauEd/IPUhh2s/nv6rlji0wXVde/yATr7SA6p8ZV/qFQZYwhw3NFdC
xJFeT+jKN9H9Fseofq8YUFLa6bovgh6vZDkD88KZYrfH5mgg6DJlqSq0sz+tEn5KkyO6gbbHxNOp
H2kXaPHEyPdFHmJ+0gd2SDITIUCspgwovcvn0iz65fxJRGLoWcPhnAM2Hha7Gn15dIlcExU3m5lH
+cx92NoCLabLJUtK387SVC/ogk+rTK076glE32KNrj9GQz/4UOCTAgAbfji2XOq6iwZO8NnEBzrt
kQvvgYp/mt21Ivk9rDZtQLqkkf7+SkMxNfAosyZUkIUX7UXQ1l2NxhZncDe4M73hBqIQGpnUVUmo
sWN8uajhWTFvSxjNqR7RfD5f6VMc6wJv6aSN6tH8gNhSRGNG2yOO5NzcNMjia8tVJT+16Q6XRPS3
8OhaS3wC5Je7kE5RA5WT+csNd6N9dUVbfcOS59NrDLQr1BretJ8SaqnpUMba+rOEmsSG17YlLr3d
PlcOc6mG98b6rOkDeBBDMqpQs4cusZNrMWeNcMIv/hr997IncqwIwOGjKuDprl4sId/gjqMxJixS
X0rXXy1BW9OeUk1qUenKuqu960as41BEF8/N2ahmCXGhupCQiCwnrYQY4Rz2so/enor3QlSKX7BD
FjkuOfYyimatDki21wYSFyUqC4g0bqnp07fqOGEEvr0+1qp0Sy6EidzmnL/PafYtbZib0nkEtELz
Qz5gosJTTxbplK6MlA1IHGp37bkDHuSKEQm+MdIXVNhOUhISL91gouD3gHgvuwDfop/OcewGRRn2
V8z5WmyHUEpaFAWIda86SPF1xTIPF+u/ncQTwpWVjclovDCfYeWj2hn285wzjGHZRCbgBeURrk+u
Y3I4Zz1HC6X/fulWyZhR5xLGcVTpCeFyL3DRp0uPi//aCkoTR+Z8Ne3R6/H3lpA/2ZwZUb7HHrhs
dbuI03SK2DYnfVWWaDQ2kerqcru2rtRTP5zB0qnFZbrigYd3fAbqLCaRsozKL+QlyepgoPnBCFu2
/bLesuvfXj5ioaae4q/K5x5+OpOtH3Zc4ekbnOPrn/YGV8jt71OiAT0NCRfG0UdFktK8JQxhx/fe
DFSGLe/9HcysCFvwWdcj5YDL+QZZNVLTYdqJCi65oC0E+GYOvpOnQ6zipGcvsf1MV79fFUrdfDVJ
57+laIGtNam4/KOYxNO6LYyVbeZhMjh9LjX20Xqmcyk+nj2k4qFmSUOCeac4NIHRZYzM848CiU64
EVF+d5OANnRHxUd69Y9sWMTpIc2nCwvjIUUdMZvEUHODn37TZIuNnr+bBOtHwIUiMxmoMRZpn57p
rSRIU1WT202brsJG7ztXGrG9vdXu65H71b9W9tfFPTahcAuQpjtoKGEGLq9tRDxEEJFXWAse61v6
DXDlZGHxMYAC5x/PJ04zhk5Y1GkWwT8uotloYlyWzXg+6yh71vz0CgaoJP2+BLHveBzs8ynQaKfo
NBbEegb3gTRuYonjyXsKbae4gisMLocoNh/GdDGtMczvj3CJQOlxelwuxxik+w/E7LrO1cAnTG7S
Li4xeMr4hGbSEQYQ6F78SYTiCYBj8dnRyul9EcvXstE5lHibOqtb1pQAUUaYqQ2q5id549FzrGIr
PwhCWve51fZ+WWQPOMU2XkKv8LY+y2qSAmQCOLYwGmvwns99Ipm888uRB2hVMSGQK3iZKqyTYTgI
Gb2k6QfZLNWh1c72kfYIjrkVb58HBQw5lA2H5NpG7e7N1cyksp57X/WCrYMN6aFvmVNLOkSasW/3
ulOYf1IItudgKej/+CQEHoeKeGyXOR4xaL7Aht7cvn4nsn0fh2gUsi62WFdHN6GK0Y3oXpmwnf9D
qEpflsmQ6F7MG2bMq2j3l6dd1qonGfQRxYYgqYxJ9c/q2RgYk/VcYbQW7fFpVF16Qpqo8FQVIe/l
cGosoWrsRmIibRMPNKDwPq2Var/3BSoagbufCyLpAHqlPlakce4Wwzh6szAtBAUV8CJbDdzUsVKB
LgNvIsnD6Qxw7NDmTojTskH0V8C3vIIF7f7uXpvV8Q64v442x7EPzySeV9/7m8QyYkJbJeTNtW+G
dNhv7VJ7vUWfqAGDcqTyroSKqf7RElYI020Sj4Y7a8jMB4xX8M9xu/M7jHuZFPni9tl48ntU3Epy
rYhhz0QD2I7ezfzZd1XcsGzh2vPd0Bw9nwhe8kPnKDE5Utay9QPBccF03tcw/Aa82pS05BRRih93
Yp2EkcKlaODeKW4Cbeg17/ChiZbJ/Lc2CxsrkCN6MznZ/pvgHnec8KT3paT40CLtwVMUlxy4Wnqb
npFjo65Bd8Pd3WzPLh1YZcHxNSuzsZmJGj+CLfFK5ZEpB6LM1dnyC+3dPhbR9Z0Wg0LdGBZHppsn
KpbF3eMzUKGS6Hg+VrAlaZkwvUomkBYHWiUTBqcCkXe9dciAGbBl1i2PXQOKOM8WvSozk3oyRoiP
3CTdhlVJbhRypg2H7Dko59nxpuff6LOtLkUv4cD/mqVDFj62glxLcIkfO4dP9CDawfF+aWMlTFHf
fn6wmL07nYZNCnKQlAKwYAAZFxXBpC2oebogN8JjFYi/2PiznRpg0lDHQ73+bVv8jc5rNBv7/cxo
DKb0BlOA7PBQRWvk4TM0mC8Y2upGe2ZHDJr2Dr1+wLOSyeh7pprbIn70c0+jvt9EnpxgFCSfvdnB
SWz9HktJ9ZziLtKFtzVEROH23OK3Yn9BUnREff/uk4YvCetWRrL7T9tMCBw6/7eOscRjAB3hcCsi
KdMMYBLA0yJcT7zEcZ7fSEbiinbpBFs3Cf7vQw/QUZ4ziKU1K68PE4nzcyUFTTxMLZ9/l3WEkdTt
7J5GT2exv4+FPMfor7EVi77pGtRSlO2KNziT9rUss+1mop6YKAl5/+grfka60p4ufm+qQ/l4kZen
mKc2QRckKEHPKmXEWdkAiEg7Jc/PT0YIz7IWO50uqce41UF5V1csREtSRQ760zZRZim4GvWRycPO
n4t3i7qZ497h+orFvNSQ6FUF1P+kk4D9xlhHJHJIaBHLUXn21MaHiK9jxq6MN83yDhpLwWEP92Hz
JlyjKj3KD+BH8kLnczwFj+zHXlRO5uHBNCSZxoVFk02vPIJiHJ8bw4YYHgWe+13ySjgBH3HX94k3
8C+q0AAutDnHxmr5WsbzT0ngfSBJzRb2/ZJFq6aXYLTTk93LgXTLkLEDD+VcCz7ejCmnFhea3+6a
o4EeJ7A4SYydsyDOifEpIYeQfzMDgcIqscWs8Sy2uLhm8dclAZryrFPfgUJZa5kJY4dH8ngVYQuP
s2JHoqQFHxIUrwc4DPOihDLGuf12oHV3qM455KmTxkJ6Unxf0YikVRX31HVyKbF57mcfmXssD/RP
/Ny2x3d1iFqfB5Qx97spHKWCBAzPPgaFQlqfs7xGAe9dNnmSxcfy0pPPl+uu5WqjIrU+EIvpDa6Y
en6oBu3uNqfmQ21NymjCFl2XWil8y9laQ9qJZfj7pq8UxIkxSLSTbxoXi4yz2pqly5kYbgoWghkr
u6PKfUTSQiz9zODiPKePIURbADWhD5UJJDsGIrRK6FJ6NMQg/Lzi8MtHCvIXWmz4b8X7O2Ty1Uhx
OzmL9anAhrO0nQWLxYH+Z4DgIK0g0q46o1cjmW3JKGerKsIppKeNWqx1c6veRigi5B2HgP8vXTNp
1gNiBIdU14FIuNm4RuIIl0rKrAhF094QMWI0zfVGCrPiH3NUoH9Ydim1o1CssLWj/ZZG2Kcy35Oc
IeSvrCeWvsh2Ld21/4qgHJobEikM/Zkt3Y4OpPq4ssMLLiKXOamctIWyogN1FaaBsewxAu7rFcfH
ERL8eqdpAH3HdQksVx6ikb5ugceqhQxyfVEJir4wOjRC7bWcyKnXi6JG+gMsyey6PXZN78nUmMbA
nkiukL1QBec/lNEYLNe67q7Rind47foFw4EThxJ2HVVpgSRrg488U+9bMBX+szmRNf6lmgxCNke5
bkAEdOZ5PXbmqN2cfH4FxInGd2ch9JnwelR7y1ngRXTf0Czbz936QQOZ3ZDrjekG3SIDDEMHTNco
WQplcVDZ0dfvhi+atWY5Aq+m5TrIY4wsBrGXU9KzZqy7lJwYX0aJDT166sGsjtFYLuH7miuyDJLu
6yHaBP97cq0rzgmFNkOXKZCBm+UtUdgwkmjJ7N8gQf14ahecX8bBgeFaMSmVqvApmcIAA7qMUDLW
WsfO9Y0kUbo0m4lhzlTjLoziXxaUDLtqWlNFmLjTmK2H+Fk4KHHUjQkIf7ipnNhy6PxsZoAH4YzP
8IhhOpy7n02wvWmsrM758KMrd7rWCrEvAGnSztv8rMTiFmQxnbjGkeZgaMr20c5i2upiVYE/taJv
yCx7ko9JfRVrPNd/MnTOOzWHJz4rYDEV6KDBhXPuI0xcJIa57HNKB2p7++CySshDG7OER2ZA5Egt
b8wQahIzit+6i3oa8JXp9XUDHsT1NYj+GGyCqTRKEh+jwmiOMmItx6pH7LtyBprAEPa0si2SRENJ
By6FrpY4K0mAVz3xdgiolfxd6VaTmcknu1qsoeNuObUbWfUMWeIlp7ozLU+581/4lr5XQ1it1xsL
rSRr9HDXudeL+2h6WWddMsPYF72X/wyeWY4/OrSHWFj6vprNEo1drgIPb2KfD1M8LaYGHHkVcNK8
5DmRqhyI/gPDgrjfhmCMABqHjpW7kLkALPawODu9Zzt/04oQ/BXYuzqExn4Z/h/qgiqyOrS2QpDz
1XbMqrZRVDPgJzDtdPcik1u6K/2k3Sl095o+MF0OqIMlYtnYP1NsiBbyVAquI/02Z3gE5nkcme4S
l/4TiQ5N3CCWGVqMSJkidprd1PUJMNmXuC4O9h/nN0pH+iv74dutjSl8IvfOnS738hx1ZIqBDGaq
/21aYWxTysYRWcG9RnPx36YBdAWvf3aj5nYh1njqA5jx5dQG5C9BgyxW1cuHUa8+Q0F2GTiEm3mW
Inp4jZ42ztio/tuDJl2t0bTIoju+cP7rAk0MHb885xlbdRUjWlTrEKfcECE0Frg4EPIGV59Oj++T
t40TBGHhITxptw666CTcRCI1bsYOajwV3W1lZws80gTwNMd/maJDyyOewo7RHEpd04gu9qpfV+bj
Z208dsHzJRl/6GX07OQZm4RJPDhMrfI03tI2PA9pezM69X+teO9Pn8azk4Pue4KS2r1nT1kjiYDY
MR5S2bw0A4VqaB7iCxsrbuSD0mfhOrO00Foq8dkNPv9p1uUMR7fyqJs3+a3/5GbtUQcAxdXXmi4m
uFCcxX8dWFe3F7wWCmtTO/39mQwLAx7mpp6eCNHyY6a5W/eDRL94W03fR1ABFa6qL/bClTpheqXz
wNDC3RB7oyR4bUXcWp++KvwUmtAJ9568N5Y6NFgN1d24BUPWnumLEoot5czP27sxobxxKvX/2evF
R4HEn6KpqDAT/l3xNvkV/51VX5swCv0bRfHdcz0ESxh5NTE562m1XbM4c7KOVFOjlO/VXvKEVuHI
8Ye3Kvkjct/o/gm/qB7MpCl4pUcHjEz/RdL2rsuTyWWuh7djWdFBS03LkK8wb8M+xf5a/TnItHOT
BWUc22ZdHnSTswUPmOfV9InMVVRvOoTKh6v0FLjYIBZ+SrcS5WTuW9Grfeo/Mbiin4h49nlS7UW4
4BjsapruOxUaSfmvbn0u5pDBBaP3ZFPOETXoQBIyYBpLPGE22+h/obvC4Pui0YPonETUiWbDkv0I
r8PWolaLTJNMe7KXKXlMDb6zy4Buxr/T/DzDZyaBbKXQi3OeIr55N5tDkc8GiAoNSyYB/QXCif+1
k1sNV6nBTXbirsLiGtL1L3e4PlZn/NcwMvbERB7RiIHAI7hZnuRC0Fbh+LkNzsiz5fS/Odkh3d14
UjwdvOC8dCYSY3gYY+h6v/gC5C2OoLhKyhfXJ0Q5PRM15lC5Qa1FS+nRBRDUHygJHsFS6JSRg5Yc
1781muMYxbrRZRGUsg+ADZYsg259DX56c+8ersNqnnWPDqlWX4XMH6Uq97RrOjs+17HBd8vmL2PH
Qn7+chGhpKgBd3nJvbqKi3shVeRMxo6KPWLU6JNsqyOGUMplK98g7zzmCkqPMpmOa7sqUnHbfAAk
d172T3vH73jx4ckOcKMAuANH3fBhwmBd8R2UETUJd/U0EWalNoPZwnglvlb5xbBI8yma3ZgL6L4k
7b5wSIigpORup1vwU8KhtnNl164lziGIFs9GysRHDfmJI1ubuhmnldwmSLgJn0pmurxQiAwA5wPJ
kqDJgULCxEbhIt1YAKM7HAPuzEgXDmrjNotxOy+Op8rQ0bAPtUxwv1PVuauw5Lohe6ReenLXyFYg
42Rqr/9oRqdOGyS6ymQDZ4FBwBLtYXfOCCmvV18P2teG7BVh6mfpW9Q9L/XlabkRzNKCNmnsLBVZ
fMIf8lEpp3PiXcWujINRWLonbSJDwifTBpZAi3tc9Ymgb7J7IeQ4UWkoV6MSf786TTE0K8Di9QtR
Wr4d29YSZdizQ8QudNCu6HneBzQjgZYD0Jy1q+pGSS3IrA1Zju8YpFBaSv1VovUQRFWgEmAxsVGF
IOo2ESh3F0bVnytsM43D6DUsarFNoKZYN9f9JVEEEaCHbxY/ewNcSyui5rZiBBGzXlPCLTN51+7T
fuSveB+MtHdDR+jugosju2otRVX2gT8ql47uA02Wlu0ua77fbdHja4s2M1RI1dwyYFW858Tv4Ts8
0uNpA6r+HpPcV9xQ5xqWbZj84gFtZKqkGpBexx0ELS2t4JiB/Uol8Pl3w9qWOFtkjcF9LlSEf9Sx
MaIPFqBJRua+obqm9FiQNP6PHoGeQri6ZVCNzpUjorqVBzR+ZPiHtNef0HQajuphE66RYBNbYOib
tunwpyTo6MzZBtEXem674enUmsW5wtP3BhqAjdjlPkL55mX1X9sztQmihc4sHdp4Q7AApFN7yGve
aHCbwM/rTqxAfhoSEfZr0ONKb8RR3qQ3WXFz1Cd37QX3TyPJGD2jZAyingIyCkyhl9sUJSXsKjPc
qaGfwzcF/DcfT5hjI3uKTIiP8kixFlrnqsEFmMFEQAXfWhKf0pG3KRYCTOkiuB3H9g+pw9Pj3t1X
VYLVBMPu9rOwF0W8HmySs1Hv7DWTGvVzlWZvRItPnCAcO3k6SsjcrOnFE+7qfRo27oV3p4rmfFW7
5/4bEBRQ1XV9PL230iuWvYrWn8rYPBfp3PmkC4VLMpqTtkXWDWfSvjlRZ4kT2huXpgNxOmYwAfiA
VT5uWvJmR4TDTXWWoJQwNx8yxR1MzR2YgP9n5aEpvbahPIqWwOlh2zlrcJNhy3u2o7SbrW3/ECfW
1sUf1tAcW1O/MlVSP53pqEUTdbx3qt6MoDnFyP5CldqQoRDgbkCrqVyMX/J4UTCe8aJiMvgl4syn
arI5cOQiMygYOJ85izss5EDWIeBBOv81uwoawT5DdPEcuooo61Qe/CqObi4RkKCSy68ff3XSqHnT
QLVDpZ8ahgSty0NAjPtjvG1qNxaHYnA0hb5l5YRPwgJZZE4W5RwJSuNoPKNi9JMdaSOzCCYeHE13
/m5ycyWqTzYiO6HSzc7TIyPZ2cyivycQpAJ1bvLhCnUyiQXwVsirmaD0+p1lGrMbMIuSkibmsciH
E5sn5OUb8V9wJ9CcP6Bve+e7+jvCT1X7TcrUGiJNVnr1I39NgBvt+3/QAIGKHJHPcYmsHTOCX923
Dc13K2ZjmugFFZeVY3cfNEtHpjMcFy87Ulbeg1mWk6FnLNOQae4A4FI3aHz9Yn8gIYUkZ5T+qp05
NxRsdCS2Ffam3uj3Crbc2KBmPXvF6GR6LGCyVJJ0ZHGSWHGZ0hfREizzcgMXKKNFiuGicWTd+QFq
0K7Wu/olt0D4LxyF8AmGHxh7zQJUXZJHYNSLmtsz9cyPYkjD4MCJFgfHpQOfUfc15meYjx7vWpXi
5k1oVEGzjEwUs04/nFJm7MIT6W+EDWRTHSl0kIQn8pgLiC7ICmwJwgLAXResuPgxid2uIFOMxU5P
YFP76LphjAmcInAwDvf9MtG+AKo/ykP8GIf7g3BAyR5KN0AQ3WVOEXag6OvSRhnnJ5X3lBTSIvNA
XlZsDhR0w6S5MLDqDLnRH0eEUNMjzGNFQa+QosznVOio0o9Ol0JMZ+Nvukh9sLFO5PxlH8Oxh0UL
Xsg0CI+jVge+gPmfD7Ey+tR8U57UU19qgsn9osyU58QNzqO5xRbbmZUMnlM5ZWYmRgCB1qf2v3C1
3EqwZR7ahjnMeE9kNSOHUMmXCuCbxD3XAlGELhSdGuFOMLBG4bvA4goL2bd4XPUyKvTJl+cIQ1bk
xq/uRI2+pu/cIYnDw3rNlLCvSPrYROdWsRuj/pyHGqgMrCKpw+upNu6hWgA1ocjE0xvQY6SO8sOx
LzDQaoLYB1EN2YM0+925G4fDJcRV36abldSGoEnotLqSBpII6HI5hJxgCxxolGHFVFM1Nm01JNqW
uDfSR/4WqXo6wO+BUtPsdFMU2BklmEarVy7Zox8H2HXdtlbd12JP+bcZKD21sQT4DPNduA7lhv5v
5mD0P07YZ49SFdxLdNLfOnk4fIIKZS5JqQnI/pkD7VO7lsR5G5Y1xGLi44HL6ev4ZuimsksnPBjv
uINmI6mwFQ7THETMkiDKIjxGt0SkMnj8Ks+PvVVYnUxOEhQiPy3JNPWYUtI9u6iWYg9aKq9D6VrW
zmop6COYZ1mpmVEVusvMgKGfXdLXFsQEMQlDQ10GEJYoAt18AHZmo7ROb1ZgIszJzmYsTL8C1Fn+
4O3Wtn2aszfYJ0jbz8Cwvt4EKcCNEB1dhtOJCOkIZi5pvqJInDr2FDL+K6/NUerQCIg8pkh8xhhb
krxuoUqJfUOu3DIYUOTjPi8R9F39mNdl2BQr4EI82HK3TwVZHbAFqPJkmeAAk1KNCsVevKugkVIl
QrWu0BundZsyTUfuWeMJayXByI4/row/EjEEJqAx2/tvnFnJzFJQLlRbjssatquStHggp9neJk9s
KfxcX4nx4ntr5Bk11Br19VS5UUTqKoz6BO6KlkwNZe59Y5ikEfbN0A9L7sh7bWGYrsuxBeNwI5RU
fP+k4B97sL60ahpjaPLAEflcDWclzYTTPq3HIl73BIrQbtQiEc3aJdQbrDczLnnx0DPq7b7FSCMq
B5NDjOTGSOiAv6SIpV8ieHBaKOmarjjurg/CuJUBqf/c3TYRIcJ3k/BS83mJXh6zYXdd5dpaaCNK
dGtIQn9cdAoptlZ2+yjzjerYgecY9M7ME9uwzImU1E/xJm/aSgB45b2Skui2I/LaZTPrXBo0SBKQ
2HqmaCpZ5WTgs04wlFEtast/Xt4TCrUQvGlLsdBp6HqiYgM1QmlBLdqwb9Kqi6JyulcnOMI+nGIs
Jv7OnTiKph73urvKuGd/TinyohjO6Z+fHd7hybt5v+2WOZRVrFkNGkpAdKlVuWuGz/RhGwKiqRm/
DfFSx0+y6sJmBHfDYAbnbavsUdmSBLJdxm/FD0pf0b61f7HMlTxFEoIXniRWmzUXNgmTQYXzS6bX
KFPpz+KrO41jExwuV2j6Mbx1NwdRVE9gsG0t9gLKqgo9fN+1xiKNKTdiL1VCPDaxnHG1bgtZdc9D
seB2S2/cY/MvhNFZbq8TPxvcAD/k7G7dr0XMyAc6auJcmCEAlkmWRys/LEy/jnvaZ9z6Homcd4P+
o8mwgo2KMgzoXIXHXm9sFkFLRYLB+CY1W1rdlpm3pdE7n/Mr+SBL9E42jRzUWp4fsKlC7IzEzcaJ
SOA2gr4fEKbF4gQouOJZNfLRaB7B3HDaDUTh3WQhpnP/ttNWuNyh6/hwp+W3LkviDRX9oEH9sGmH
XU0Va/TMa2aUQCdlIvlNnLFktANJuf+feJKefdxcgS/g74+8V98ui+r/Q72Gubbk3z82yDNNPdm8
Q7jBVoEkaKE67ngKzBB34f14F/RAqcQujUj2Bk2YIKKpzSwwX1O7MA5p+IdLWpokvd2lNngNmvi/
Kn/oqxZa568kQyJbD0Cpq3NcDK7EWuJZXT6wBU0ReBoOT5aMue5TfYgBIbeOXlsrkoog6qLfw4Vf
tfUSSi3KfWrmIva82IyqPbkg0qTpGYl9sdr38BYp+Oh2oN1jB2w+Vw/ZBuuyN5NI7OVgJQvM8dPw
BA2MqjpPszehv+YTKYd9kpYcxTU8KXaFbSxX3JtLlvvvf4R/6sUfYGffo0CtDFjx1wbhNZKGoXk7
D2BUvDN/jqn4UJYidcOIdD5ZOz+oZJrTpolpbQFdssjutQVQw/8D4dBr19ZyGP4OImMiq2pY+u9U
moeWu/5g7CHR608WXrlBj4yOeLjbusCAb9C4uKnMJHXShloBSW7XuNghUCzURJsZz61/ZNHPsci6
thx0pZexJSatkM7uHUIGyTzBgXWHdmSF8vNmYbsip3l7ulpihlaLamwPLY5TuFddZvuD9/Ev0jfU
S3VLkiOUraemXecu/BbyEyjPRBOntpDODb4hLmZxREg0QcdLPJgwKbE2jqGD7q4sIOld5Zn0wBFz
UB2jxUkvSRsVkaaVtBI1QvCO4pjhKo75pZcrPuEmdVxhyKzztpufNNrjImzfykbQsS82oe5WPAis
9NG4LQ6d0nwyv+1pZmytkjrc7eFn4R0xTKi+SgF4V+qv1d6wJzNnqhzb/PWyXPAKrdSzndrRA2FJ
OGj5M1X65UdzaXcb1NFAsqVS5fmIEkzAXyfa0sgUFeZUQ3jAs0lDBgx2+TiWHysIvXaP9+05TQe5
ptYPpGRxHjXbChlOnGUQO1QZqwqwJx9rg5jFsFGYw8go19lsLFm4L8wKRRp+acC9UCahT713uL50
CscCORPerO6l7kVi5bdSdUr30eFl/91vQY+xjqwqudhgvugpnbRfRM425qZHbFruNTqmG4uz+6oi
UQhi1hW4/xMDWR8MasC9BEmEtSTMhKCgmrQFHVgdTX8b/rHw+d/CABz4r5F/OU6uXNrSoejXgHYZ
JSnjhJ9OfdPXrGIV19s4ERcgRG6MD7Mv3QHnKPl0A8YjrUdj8UX+ZqG8GxBO5uq9THzNPbE8Hk+Q
pSbibb8tOLHdkpoNd1b0JcrkQfkZUxeAowzgw68DjSfJ1OygIQ9vwBcvntpUBs5BDvj4bRmeZ5Gt
wEhyvbuoKf/dfU3aVDhBFARX5uuVNVUChgIdBWhMHToA0j9pvz+Tf61fEhlT5ZPv2Hmb7Bn7tFsV
ebmDLOgQ44mnEPDxEvie2OfstfwUxJB+Mmq6+U9FiAeDgD5etEtEuJEd1VBgbOTS6CL78b1Aa36o
pPCXdIGvhrETPCQ+IG3Ftaj/w75fwuh4FEvZw7dZpkFmqJoIbZYav5/DrBF+rYE2G9Un8gVh0a2F
w2jy3DMApojheiclgbfCL/1Y9ao3Q+//SM942bHjG7eJzP2Iu5ctfQc3NBhXEEFtRQbSnU9z+iSp
feuyVIVZs43keoePa6ahRceUIM9jI1lM9cPmxdAHT1FDVf5Bor9uCr8hRfHy4bedCLAgOy/+rKao
OJpiqn/ZD+6hUvbyqiJULywCUrW/vySHsgZgd96sYIMluMDhvhs/hb58Yz2GB9J8gr1hmCPmId7a
Tbi6mwgEBjD0k3vFUxZb+NlmJNymT8r1mOPu7TVzY2me9jpHEJbdiHDoXFuu/O7sZn/ALwpL7ctB
YR52jigHpGL0tkwmAEAyd7nmGMml9iis4tvRevi2Ha4+2I35qf6jO2pCg5SFgEwM7ouwcwlMG95B
cxSASbiVpa0bmv1sBmw5BiXmvccl6pCoZnhB8VNCsCXjLq07ddOH0QV+MPaM8oB02T9R6bFuR/v7
n7aGP8FWQmETleG/7ZOb4T/uiKjzHz9Z+i0H6Qp/2t75ehQ3i/bzA6zYY2inoAY56YeqYrj8e4xW
HkyI8GmqPExfKwVNfsQ+LR+IA4iSYTkvRpW2KcR1QyUncIrAjo67DitIbFXHUVFY+fZaVB+xWNt7
+iwFF6Pan3eiORpQquNNYe9nsuB9J7KhpMpD/rulbDrYqL30+zCLfUSmXUMWyznPEP0IF8r8JJ7F
wjgx92LP1hBToRt5XkwVqo0JxcpRuAiKxh94oV9j1IcWr2WMc5m7CE/qXxr3XUc9IN/kLQrHGAmc
JJZRV9gngGydCe/7nBG7u2gP3QVFS/LXuc1SHBOQMoBr6vSXNXei/Z4bn2bp5mmpjhKchHEN6ycB
+dwTr2+1sIY2Djm7ATJssjaB4tKtXW+nEDb9wdcdrBeufLfBaGdqOgbX2uHqjgzgT3qYn2JKGotA
C5B5UDBQuwsfvKps/vqrx9zSZkWpnULfYvBaNHc5imXv2+6GiKgwkKqn6q2zlIeOK+uUBMS/EhoX
9pGvvBSG+NRhqrvD1SZWNCtvkRNeeF3w6qOJSEq3Ty/KjUxFUZCsPGeYIdQIWwWZKujoJOKj0HNu
ggv/BXNiWrfrWTjBhT1WuzzAnYpXLLAn3hSmETJkNaMzxTkd02oNwlc/PVbdZedZVRoiffURpra9
2DxhWci22+uZleBYkCMK1hipuSqmBgD+JsEXP5N7H6PzPx3rED7uIvA/PFnQmbYp56sQS7FcVhIb
0SLApUvWZqkaxLDkv/3yJ96Be9phwzK4bZq8h0Tq7eL50mmQGqV8VdS9aZba6GQyXOpWiWq+TXls
nEit3okn5VIlCvTqUUs2jSxHMPRceOE8NMisqSkIxCiTuJvyY/v3shPkC9nYlWt67hfCxE4lq1k4
CsOgOJiZlDKepjJ7xX/jJjTEIPTVYEMftPQBEH7/2ZSpM2ssBenIoy8IRYKbTLhbzxS+NRss4neV
x8J+MDcSUT67JhvwK1jllmE1/uJ8RvXYpLGkshM3awOZ5E3O3blC99SBkQxK8SpopG8328aXFh/k
Zra5uELGVLQzVs8/2humN9oXujtnhRFPLbcwVAC0etXY53WjUTlSE/tOk64JPkD2W8Xm2uSQlnmB
yzK9vqWh49Ctm1ngGwWcqvihkNBYF5syd7VgcjPclB6CZwVniaDId2a1M6qpzUMStuHUL3SiTMm7
FKcr1t/75k0eXE/O4sF6fk0JXk/xpFoyJvwtfsDcGAbhyefJuVu4I5tTBiwxwNoa4apUnXKbK7Bk
3/nJAQolgtYb3cfhFfddA4teCXps9fWF/+dq4w+W6nElVH2UA92DyC8O5q1BJmWLkd/jm88YE3QR
Rjg/TrDBgQMp0ssQlmqiFdJ+7GhEzsXPmtZsTg8cG7Uu8J91qqPa1GC47SAP2GdJOdkE687dPglt
xkS8ESKocZtbEix1KKyz5lVseLowBThA/QERKEc61aI/XkKxLfHeUREfnA+JlfttOxfAkAHwsQ3o
FAGKXQdiB23BZAIIWRHIEQkQH8fTzNyZokcY1bALav7ZT7zwpLT+zyF5YEURVe4LNbtIU6lqvGqm
LII4YgbnFFqaoH7XAQYz02MdCFWzJhsQsBfuQ39SF8W36//vXPUoVuI6H0IvqCsug26Gx0SoIOig
ON2WLMd94X3QiMR+iIJqFCxisn3c9l6iQUCJZrVLrKFv4lJuTVkGsOnV0HU0gBn96bFFdk793BXB
FapmxTeuh2hf//XXtAtQMImy6CQ69V/zJUA8Pp/rncfFJiKP5yumwc6Fg05yWBEx5Jg9EUr/8TOa
A0cuZsw0Gs+Fppr3ImcdWcXH1ZBV15+wbnbxDv5PzPFh6A==
`pragma protect end_protected
