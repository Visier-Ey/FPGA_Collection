��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F��������n�BJ�F���U�FW9d����T�+�wt3��^��r�q;\��af�י,��9NL���ٴ�[�Z��^��Jy���0�T����l|�x�5#B�o* ��J/�CO������|�)6b,P;����t��ew�u��5�v�u�E�8����R�oIk�����Wb�A1���5��r�5Hڜ �r�n+��MS5��n��þ�|R1��������E�%��0E���;%�6�׸ۈ�6��:�!�#��L�jT�a�S�N�LS�[�&Ϫ���]/��nm� 8K� 7�H�be��
@��1>��?���X�U��&��P4
��J��tz�6�^�O�A��S�������EjS�V�6�$�g)�H!�uA�����.����c:k���:J�G�y�*aio������6M�pʫ��QZkw5~��ΰ <�z���i����Y�T�w-�q$��k�d�V�5i��[�r6t�`?�.�^�v�
��l�;�y/��y6�]*T�۔"N��d�V۬����/S[�B�U��7 a��p~q������~�5�LPؐ�V�T��?*�ؓ�C�r�����	�].o������߽o8+\i+�`K��+darwEi�JI��4?�}͍�<<�,�j��'��u��K�C���=a�X̉��37�Z?�(ȣ�$��Yl\e���=~�Xa��s	 -~����w�N���,v-�xa��$a2��hA$]��g���[\�7�x���{�MO|���1Wc���C��e,m�"��$�O��
	��M_O�~���jCL�"����V��P�h�Jm�_E��HaT0CS��&�L1<LJ�ګg 9Tp���N�Hm�}r�NBa<��9����-L��s�/�ap6@^߇T��!�3��`�[�� [ݭ��O�>F��� ���&�	��A�A��.V�Sk^�%�M������P ���v׮���w��]���B��(�	�r>���a������{8��Q5��}�;�9k�Ԣ�BK^��J��'�.�����Z�B�y�"��_"brMV��" T^�J��b�{86�orWf����)����0Y%���I-��3Z����K�����N`
�ui�^ͱ��fJ�������)�zYf�Y�"�0ɟ���q�W1���h`>ֲ-�wo��a1�n}���\�'��a��k&�����#�-�'��7]��=��o��a��x��H�ӛ
h�X" �_n����2V�#�*S\yԔ,�e��F�]%2�ƒ����Y��W�L�P�bӴ�=�� ";��HS�zf%�vK�c��-�����_aq��E[�tj¸�@�����pҌ�q���:�1x�$riʑ�����l���M`��9����1���>�~fh8(�P"S""������f�D�F����>��P��l�z�5ඖx�U������
�p?|X|M�m>6��ܵP�x��,�q��M%HQ��tE\����R�c����o����Xm�a�:=�>�Mej�t%E�j4���=>������)s��πr��CMq?�3�=�ݍ�o�#p��aZ0�3l`�?KHՎ=ǂ���Pǌ���A�������3A��/��ա�7x_�٠ƚ8�Թ��
���\(BtvC@	�Y��	�?���L�^u��]�u|b�.����3����rδԂ�<�pھ%�s��,���*]�Q�*N�ٍ�鈼/{�)���=�0u�7h���E��2p��i�'�A���̀��9`��.�'���#9�3��i�#vD�ɳq1�X6gZC��@�]��O:��/�{�H�ZH2ډ'�� =��cp�!�$`G�@Qp�1��d��4r'�F�F��=0�K�.�;=�� �hh�z/�'׀�Q7���q�Dԑ/1x�G��lJ�[1�"����J�jb�>Z�=:�!�+�W��D�Jp�-ox3��X���:�3h��h�m�&r�=!E��:�����+W ,��}��б+��9#��f��L���=�����ٷyl,7���6H�MF���&/?.-���jP'����]rlQUO���%���A�,�u'��jU�`��̇��u��s���Vo��`?��~ׇ�~W&�7?g���H���,L���~��Nf ���y�,/�>;��h�+v�6'�?Z�F�:�ʊ���2>�Ã�)e'w���3w����}y/�9Q��a����q*`ʀG��;63��ꐛ+�az�1�ʩ��İG��e[V&���rv�~K1�Lo��oc=��!��X0��QPa[>7yi�/��q�>��W<G麸��A%��a�	���u��.��)��ٺ��<Dt��g��jZ�~���qG�A3/�Q]+�y����JS_>I��	|XR�Tl���9�?1(��q��/M����!_6�tRt��������+|��pǟ`�HR򋦍ɩ �����q��
 ����v��Ē*j��.�fp����"����(���P�om%�%�\.Z�/�p�KVY)���%����4q0��%���!������l㥱߼7z��M�1�-#�\��L+zC�~��$a3;\�2	%���d?]kE�]���Kc��@M�A� 8%�:wQw��#���X2�~��N�$
�d����;2�w���G�D�[u����}�f��6��"��ʌ]�]$Mre��a��Tm"���������ԍ��:�\����ṭyz�X+���V<9�#���jd�2C]z����V(0�0���-���"ǒ~��% kEk�Z�=ḻ�xKgg2�峠Tr�\����1����9\L�æ��%��� �5�x�aǳ�1���]O�p�g�SX�E��i�o�GR�l��=����#�j�q��c����>�������$����ɩ���>0�����ȅ�F�s�����*Pt���&�xx�Ӛ3��J�o��wN�n���Z~����V���}��|��~�dc��LM@�@^�:OZڙS�ˇ����}�_��c~� �V}!�]x�K��'q�<,B��;�7�Hp�<D�L�>z�����d���%(kA<��n�.o�S�>.g�8`-t��*B�#~('�2J��3c��++�'����Z�el���mz>=�H ������ڠ�>%�k~?����)8���S�`>o������/�ǅ�I;�<�6��1�e���0�����c�����\>7�3@�G�K2� L��Dt:jHv��웫-����bA���y24���x�6k�����