-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
Dd55OFjPh1eVAENTejZrD7/Phk2936G27FOg50a8vyG4PNL/T9OYDTmhiXwCQ/fG
xow41CIdeW+noYX6R4TPMe30j5owk16/4I/9x18XnfQ33+uZzOEt/5VVLuYAvy1w
V0sicf1lZaWJYzxhPMbYmP6gtONWTlkK39JCuT0cjp0=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 1651)

`protect DATA_BLOCK
5CrfJAIVnDbW/bzwu4fGritcIWaEYqzoYLYy+SPzpozd9BOjYnypRJWITYTC1xuc
qjEKVHjFtARqmPW9nP3gwpVh5qor9d/290meH/qgqjQyc8xS/atUM4HYrLuyN/+2
dbTEYHugc8iBLOsTQpgZ0yFRl+YysqmJjBLvpsNFL3qJHgUAmG9QljtdDByccoBM
RhAXm7cDJvkcP5v2A8ukvQ2hZw52dP7J+MoYIggoV1d3ynI9ni87so+OMjDGQzv/
jttjES8iLTUEbw8OjavizeLsbqECPX21a4mOrbv5fxypRXmdynPQ6X73qM1jlSgw
oo82E5cWhK183Q+n/umyRZifFvdL5sD0O9RkbW+22+w19ULuD93y+y5eMy3ULWkJ
TFXv4LLe5qHh4oD++Us/qm3UzzR0gh8kcp+6MAJ+QZVyb9drMQrvmvFMyQ0YumfS
/rK3VmcnthIBiJjT0jZkVUihF4V3xyS8gbO+10uOmjn0d3kjQl/UtmG643ReBxNw
APTObQxQFwfPF7FmXc2jH4NlfAN0ZsnpnY8IolDtQfyN9hpIx69i1Zea0ksUXxgi
p/8fYGcUks+Nr6SWgWTs7cRhBBP4pyMjstsBM+5gfNOiKdC1yEuQi/YbeLXR1Ghi
Z1mWioDfdu+qR2CiwOl0YFU+wWc1D8530L2cYTFNZdB1XAe5rR8FgETq/JaRm4Fz
iinOl6YABb4O1G6lAZhJvYlsJNfC6P4SkNU68sv7e4kpWaEaOlwDXm3EKR6cNHwl
lLwQPWpggzUC6FgWqICvEDMEkpmZyPxA8TbgdhSt4SoHHqBAMc/KLBspOTF0TCVN
E3VsPRaogMTF+qB+0Xm24CSuAzXBD7HuQFvt6DB7rXDew+HbjLWwGbjmu+TdCGAg
ucep4MYl+JVs/1JmfGqoyuq5jBP6CMg3q3zPiT3k7MUkiLxHb0O+XMA8WUBoX6Mu
O2Yu+wDLdaUHsR7Kzn0beaxzUOKp8cnC+nyPqe99QJkSHzUqOvL7MAOBIu2Nq453
FyMd7HB7jzJlVwxn2XJAlqUJOSyHXg6Lam21MoKBcGxcHgepeNB+XeGQjKh0+FWj
eU8GXN89BQiw1Jfc/wgu0ZpfxQXbl0tBDNohOGPiKcqQfit7vk3ER/MryQbJC0Yj
M9NtwtPhA4m7TTq8ysguTqcjcCtJMPreRjkCSvinX5U/Ql69TxRH1iw/WLWEhggZ
7G+dfKnwWds8PpFO97Np+v+6FfX0zbTSRsQK/xqQLCvPFxlwl3T214hGFKOw1vf3
n3dIRsvEmfQIA61UgXFreUdf53Flj9hPyZgqvtfZGh9kVhULdhAlKW+PkT01Rya2
63utPe8w32GtkNhzp0kUf8nJ3jJaUMMuh8W9V7LjscLyyXqx0F7ijO18bOpdwkPC
e+UeDvZlSkOf4ykC9tG7so941UlWo5iicMFM9E0dc5qEvCwgOCfafTZdttBM+qxE
jg74nt71IUwdZK6EkAAZLIuHuTgMZY8XSJK/6AJmG3sEafZktaSH86jdwWNYaxyE
Dbbi17uYBtMl1R8yCaMRSsJ0kmEEyQmHn5T5utlZ1d/xhr6TtRgK0oJI0/m9jmwi
VEiqGyi2+w4xHM7LXdJmkWhOogoKXyyD9GDrVH4ynzcZuPiWiRt2C/U+VeyFBf9N
mj9XbG7HdP2JsUKsOQS+qDTGl1JHBlhXacR8a62JPc0eYRJg7ZnhlMY2b//Gl1xP
RsI5IjtWXZ+OLCVSu39zj9/Vt2T4FIDOEeD3s5mHK85Q6eANQMJ/2Y6/SAVj3tNe
jPSJNYLzO0+SWA+IVZxk0FVqLpgz/2f3o+tQ4YJj1AyRjL+ufGNoYFWSHsZJ6Aay
EM01p7coJ7rab85WL/JL9NI1wbO3dvqozWKQ+vRdPCnzsuwAKgcM2PSKyDFy7VDi
zYmcF89LJo2cy5GUfs46Vs8z2xGCBJrEuBfi0ItsRRTA7bgxD6BN4Mv4W/v80MZl
4InchIv0CXEm32jEVWy+AYDJp2fzGFs3DDwYDfgCUwydaV7DSVoImnLHbSp2SLgg
LWwHEJbInFJ0U/MJ2KO8VppgYiaOFGNfjU0hvipuJBwVGcrPeCge754wnXB8KwrS
xq6T8WPlbwgTy9kzC3KIHzjbmn6s6Ory5wDii1sjwNdfeYA3KGF4ziyk3V/NDjN4
nddvzWndaIhYjbt8hCrbSry41JDojSGKTmm7hN7pPEMUWkyoxmM+bto8q593q9YP
`protect END_PROTECTED