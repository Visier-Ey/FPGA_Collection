-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
--pragma protect begin_protected
--pragma protect encrypt_agent="NCPROTECT"
--pragma protect encrypt_agent_info="Encrypted using API"
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
--pragma protect key_method=RSA
--pragma protect key_block
lLd2v4tRXpNcfRAtI0sAGRC2h0jePpWIRwt0edZlITBfpQeS2doGmqmal3wp9Yeu
hn0VF18WVhsxvpKzENKu7U2VBRQq4TVFPraIjcDIYlcsKCLJSjOmmuZlL1983UMR
4x7xKldHEHVp9ArHPxC9qiLpcc3Rl7cZvjFM8iUL2ppybSdRYebAPfEhVikyk7R6
P4XnLXRfatUfB7N6Z2b+PMuJozGavQm2waNkibqIxUC9eCWsfSosOMeMyx4A5wex
vkMc/rGY3aqnVaVdaA+7q0JcAHBGkUcP0rTG4wXAcXCpfaGKRCAd2psgeQd2vhhl
1tFuSkZDaHkAkr24xmMx8w==
--pragma protect end_key_block
--pragma protect digest_block
lRPZVa3D/rno9wQ3yM1Q58tcIf4=
--pragma protect end_digest_block
--pragma protect data_block
UXIeMmPJcjpniwafL6N3BYYNubcurzza8Vh18tWNkq2LX3iLFXqrJZ/MX875Ovwm
R12GQFN7LwvUaMat8+AykPRwIO0LyEV4bfj3YXvXn8obtAQpokkwKexOEYR3HsO6
4ZeDlw5zIRMl763fJ0deumge+1eCaI6LeCSlXdYVo8fqFlB7szuXFNx0t/qr6xBk
8p3bMI6O+DBWl1VKOxv4AW7ihn6+t4JzCUq+1Kuc8oDPIBmDSTZwqEZukaQ/lsBN
9uw7cEWnMntD+fnDi4IDmOEbS7TRekA4kRXskUjkZU7u/ddCJKtNgw+U8buciSt2
cGI3baReqMOpKMOvPFgkxvMhWWLM6dqtk/R2mTyKA8ItXP/t1/HnwGbdiJ8epw6K
BmI4/oX3vngWt2gD89ILqgEQSkJ1aH4nctEJcYrNPL+4TJml8d3nv3OCxpxrVcBQ
1Nt6pqf20pQJEWGIQm0ArURu+9v8NxYc/ohrLEUYBjt+ASWlHKblmvkDZc7LMKJV
2trlId18dNiXc5hBPKj10MbGpSbkLro4/4f8orByUQBWAO/uCkK2fnEt87rZarNo
WPQk0TVmk6JeSHZyf9Avx6fQv9QrTMDrHa0vGB0J8MBhqrtSC4ZVVw8ab/zBESk/
CnVad5Bue9zuLMFUG/LmiL5OJ7cOJgn4zyQ9f/8w5quus/+ijv499ZlaJGESeZPu
f3AC+q58rNhjj1tlcfvPvgvVrceEwRrRjxBw7UjCbEW8dPPmKFt84TQPdJXaAhV+
cWHCTMRsXb0VGY+igivZHv3/f0wkOuWebB449YXh0Fu2Dn2804AwGnhglJFR/G27
0dmMe0pj86kmLGQU7nZ7BTHkvLMkpD3hacq2WoVP9IGlT8lwO48wi/faBCRZ2ozb
BHeiPzgQ361462UVsVFXyTmqj5dt/9jwHo+/x+EeQ/VGpAZ4A65ws/dH4fDQE78u
/oEWnw5Xf9OeZWlPnHynAt3dvhMrrWbh/4IbKufmBVBNrmVDyZ7Fs2SGE1qM2QGS
QXA5sKAcamuKO10HgW0Sjkgclz2rYim8F7U6NXpQ2s2ahJPGb/EjE2010PGTkYQ4
DhyGxVhEFOT5qIfSO46u1Xnm1aaVIh+vTEbqr8FMfgk6Xnc6fN36CxczLNCNrkbe
ADQ4+UnUApy9FlbSo80BuGrDO6zSnhxT7aA7uexlSBROg1N2UuUvONFa/51kERyr
9SygqxYQ7KbbgDOni/CpKjf/rqcO5rRSeuVWk05uaQyOsQ5phTA0bI6jIuNOplWa
M0PF+bLbaw7dUdmTbIiYhHWqwEnNPwfAudUyFtV6FK6yqWg1jl4/urdhRFOn+2I/
G9ZhYOPsY/DJKRUDD5QT1ittIC7u8R1JbzInI5K/NZNscbvrTRr1q1dU3y96lYI3
G+sxfz8lw1V1uCFCk5lIOkw2AfoKXCF4yPpG4UqzOfWBX49lHOyMN5t8Z2TqQ6Td
ehn2LQ5BljwSZ7IGV1U0CgcAhVL8oUfHlIUQwMZu00N61Nwj2bq7/nkKM9+/1P4s
rquS7xF0nrJ/XjKEFtfa4koNYvqsNIHNWaOJu3ifAvb7cEMl3tKUlQc5djAMLy33
YN2ClO7lO6QSS+tocythADxSjGWmlPKVWlaIcy8HNE1F8wlGJcy9EVbSOFLKc/s5
cW6sBhGExEx8UNrqysZP1dlaqmuXuboufsBEEmaGswpWKLabZf7XoAjfJjaq0+/t
2mxbIvaABTn0hpeSDVD8ynjf92j76bcizxxIgY+BU7tJGGh8h+RyRvh/bOUaUgKd
rVMiOpUMxwSSpnxXanvyESS5Tz7iu8WRqnviIw7Lf+ONiKvKrHFfT4Na2zzEegSI
BUIahWUpulLe/pG2HIqTH8ILYKLDb+yU6xuTplgKcFOka8bz3WyStcr/9GO11KLN
msoUl2iJI5VbRyS88bRJ2sHq1G6vXLdLWGeamWUBSzXT+fDrq9cw0yNAh9txjHCQ
Egv7/SKEeh3fub4EgyGLYfqSPLYeEZKZ9YmpRBentSqBpEVV29eJyat7JSBmeiuB
iA77/s1eqWZDDtX08FQ4M3oW3eY+SA9CXVs011KhfORYLPgl7baSnW2TAvdrPhuh
CPRd8eLvk2zMuM/yeMtu1Dq0zE0dUgqgqq/4Il4DyF+B4e3doXzhs7HMPWNpPkV5
oyhyLay3TcM+9fTgK2gmqVSjThA7PvgDHITNQ91LIhCzEJIrtt62kQ3cevatfKAJ
tLrG+eXTYCZ6RvatBuaaSsEg6VSV25nS7OYnvIKb+ABHhOCQmZlS4UB0HVIhRnHG
WOXvgdSWRFM7hp9cBMk7qtHoTJwsdEtUTzKv4/h/HgYOpdD2dQ5BkSs6+wcY0UmM
wJAW/uYzPY6Q1hT0lqNoYk7W6kQOl8Z5QuhWDAQXGn0AEm+dDqBXTX50UvIHBWlu
1h7dv+326T9lZhWlw9Qm1SMXrK4p9KgpvC6PxFnxd7nSi88+kJjyV48qOiPIYxyL
k00JMKFNjjErP+tMWNUsPa7Qa14QpcqTr/1QoglR5OmHdNE0SF0GcG8LG6xiMYJV
CcdC/a5/T17PYYKVI2d2jYzVvbADxFtrUU0VHkhqmL+BuI3LAKIZmIiQJGQtbJmV
KC999zrRWcYCnPsHFO47rNFROVfjR5E18uTvUbxWiVFqk853X8AN8fFofP3I1QcC
y2Kage84dNsfPMgTfBn72lACJ3D4nJFkdxoJBs6zyStnBLMpIpL+n97dN/pi/m/n
6FSAeJTVCnNNbpQCiktJBudYhLyfHv3xa9m1Tm0MKA3m/EkbAQVBGIbQRG59VvUf
sOsvWhfNrexAsgfabKH6XxfjzqbSdJAg7+RvZdFrzOt0BSmZUArgH9TT5MxfyMyJ
2LD8dXWQ7hUOsOvu8/3YRmRap+DgICD1EkAbjO9I6C4EIehCwWLZ9PHFQ1G7uiL+
MkASzAuAo7xgUYmwagI2omm996i1rxozA1Ug76IX5UXcctLj9c9px+j51HpL3r1P
boLoKCtz6ziyrlqPeYgVdEnHmEs4FQfsczuZvUL/tYb7JtUD5tUqbHRcqboqmlwX
MuhJkae0TLA0KdgccY6pzZRUS/A1d8yfKApt6bbujbnB5Xyj/Ma1aYVQyIj+bvZE
/2AfxUPEmJ2ltuLRmII7Ts1QWTYWXb/SYToyx3stK73X37/5TE98Q6ABrOZXch9f
XSnxUZch0Ua8KbF/oPP/mlDpohturwIAxApaB8wzap50BHicvZ/1NEm4odVPhzC5
Ixz4huNVX60nOz2aDI3x+ableCft2Gg3itIbZq9JXxp1RBXQkqIyPq/MA/v5TPeM
QeNxJods5PFWRgVPB5+eu/Z6aU1raIsMpvwHZheY+UEV7TMqIc1/ON+bzTgzoMOI
uCmFdI0vFuVIOQyK32/WLrpa1UNxNnTDOw8s/mReXDrVv/J5KR0YVlQR9RuzoTJn
7VaaVQufzh9xfArT68TCZE2gAU9ilHiTIABt+EHyhaeV5g2ts1tdj20SFeAISC7s
62S61xuYhCCcThabSzqIqO25XANlQNpD99loO0TobSd914sVzW8xblL3G+Uo494M
LiVp2N6TFKUZ/WUVwPzbz3BD4KttJ3XcLsMe5l45Av4vBC4u8QNu67tB4Fh/VzAM
bIrjdGFhRaPI5AmVGek117M0WDLXvbdt3HTV2Jzmj0M7MSj9fUPVK97FOdgL+BjN
7s7Fy46dws0/r/ovyv1vl+IF9/spqG3BFgmE0FzRF1Qfyj7SRMsLpVac0+a1tzER
PIB6/Es3pzsdg5mWKaXxUDYOqRwMv8R9BFMfsTPaVmUGOQrKwk6hLIWYLcc3qb5J
Gja3S3HHjG2v9oBM0+lIqBpDqUrBOGAShEtVKzbB1y45PMVomyMX9mCI5Kou8LaP
ufKmwfvYhXYzNukfrTq+bsZZe5CoBqQ12YrHwFLzZARvckfcF+sPof74TV0UKXQs
3h7vV8ojt6N5onGAFgFei2wkB0ZH8zgJzeVw4PvzyFtucXTUmhtbq9DYJKI69k7y
iuUxMAC/mMVQvGLWgkTsJLGiz4Gc6PoDD1V5uE1mHulAMc473bZutv/V7HqOpFyR
QCT9oZwek1qz349GGwGdcUBMwysp3iQuJ6/B5dSwDYmizY7QgH8t5bZIpRW4Gy4j
amexEUErdRFSevJ+EvaJ9qXs9Ipw7bNjYmeXdSDqNngsSpM6JjsCAjqaz2A2ParN
ubxELvr/NDlLOT9SGUQC0E69xl9T546CXjKcTzFRIgZgBxTJ/PUkYnPmuZrhc0Tq
vZaYnjd6RSFHMsStmhjOYB7asXiwMpfu6tmlwkg9eA8YcyARCEUsTtkej2Yo5hQ8
tMDkuoG5k3b+tZ1uly2wd5yWaPN/fYJqwM/hhK5FfBqIeOjoQKhiKXcIA7KXT9mq
NYm75QoeiuqNTRnJ8KSQ/VIjpJOgVWMOUrqfCM1FdmJsu30UD5jcSovS59gQrOoE
wwMzqtxBS5Xowv5GSU0KfEReg92qvlv8LIpICZFf+qdT77Qx8QMXyL4o/0Ox1cBG
kFbYwtnhZKV2GgtLingT7yQFuAWmsTiig4UWtESTwuplqrXdNaR84mLt8umFwFDV
/UFjIS1SwVa1iYrny64y2eL5YH0S+3tq8SMtegLv5ua3o9Oaie5o9+EPkw/sv7Mx
oKSLuovyB014vISNJV1tMLy6ahAg2ExdYx2YU+SqdJf9z+ITsmVBbV5CGZ0eeiuV
KqFLa/N/pXQ31Uh8BPZY8iSQNDQXeIK3R4XUtAzSd0GRZ9fwHvygezvEfiHoFAXU
LiYrUegc99W4ye4zK+GLH6PGVnX6YqTeGBZWg85fie77QA9R5Hz7S7mfhaykiAJr
wVibKwNIRGh3DObAu1IQxvK1yKGFAF4/aNSIeT+AN3vILNgWVqL16YUJOe9z5PTV
Mg6W6i8gJ045OX+x3/FaYYeWy5Zxo7/kSzj+u502h6Oc+qHgUfoBFxYNJEkWy7ZP
/21lPXipC5Qhl5A2s8n2ipOjd5eLrBG6brhr3POH1C7Bdkk4TGOq+fdv4EZBKkG9
cMOBCO+/uYORzgeiTWEa/BEgzczI/fO4XQtnqX+7hWODnkWGFWiFZnNCEDprfSJP
5sA6M4VdZC/8M5TD77J2iSreSGSTkZAsyzIAq8uXeOeXGSbfyd5Qfzj5eEO021eh
oa9xdikbWyu6C8rc5GuvybK12Hfb+n6zZYjPrj3CnmLR0tOd5q4oVllixtYRTK6I
Js+U8ubURO8NjsBXiF9AgLzjZehqjrXC73DwuI/d90TFTXhxCIcATo2i56bEYyIC
eleT3ZZjsPzugE+GPvBydjC+f1oG9uG7Jm3MGHuuD/+1yJs/Qcn08ruhudQGM5AS
h0b73l/iJ91opUEWwK5/ZMIALlqO1ExAvx3xDwi0CKV11iHatlXnmBFxZRyADEGa
GX3nwljaF0vBsePWc3EeK4sMEMMfIPgrZQM7NtiHNoPe363p1XCYOWMj0AUqafCC
xxPKsHUUtRYfok3zj/iXuiBvr1v4TVyOeDz+aRyiuCOpsAtRFUtuIzcENG5ayUBu
xFMxv1NNzLywtx+6ONfe/P5iA16euWdOQ+5Hxx3L4YSTOdO+In4ZMJJWpSTWWev/
bAOegHEyp/V/+CfDhu8MrnvG92E8+wzS14ttoDQe53zMqve2MFuCsQXTZBCSMc4V
/h/50D+1T8hlwac+cNHLj5D623juCgPW117Esn5KpOsjFq6Lx7HuGXUvmZcYz2Lq
iEXthS7LiTC+SoxsLYUMY7Lu/r5b0Px4eOqsvnr/4laCEZ23Nn8ZdQ+H07HSco1J
pzAwKeqFvCdHRva29MGC5jN7INsPg3ZltzuwT5eEvWx5bJYbyYh0TOYYJ9TrQbJF
w0fufSxMQzGpC2lu0swXVwjwyQuQKNn1P37ZORjIz5fyz7S5hy7Jg9lWrzGvtQvx
k/7X6M4IO3qHEzoNMkAxzVMHqt3edZl8upk6Uv13HNJd8/hOpirmeykw3BtE4fZV
EtjPbZUdazbtKfoOgSFEryAjJ0k5b29nVYMzPuZNCoWt1yqwrfBdCHZjPL6ST4GM
MX8v3V2/baEWmk7IZtmyQMvpyO9qc6Mif4sEWB+WWUsjdIRQqg6RtkMRsPxXhPOc
hBmUFaDiepd7+NE7qqmVx7/+m+fGYKPwCXsd+QwJeMIsT+fZBR3lgcJyqsZ0wqi7
DhNd2co7Wzox8QGa+o3Ep7jWgMFbSAjiDBzAFHfoYnz8T1M7ryJTMb2yj8z9aaWW
zi9p9JPdRSL/s8xaagsBKRzdPd12Z5/DpwEefKaePkpVJGndQinXITqUNkXF6Skl
Ybc2UF3FVzvxSedhqdBNHb4Uhpdm3chgMkQfu1LKP5GwtoqRaqrCntrU/Bg00Hpa
hkP8I6PYQowzYUnhPNV5N+oHUxoYM630WLwCO+e/k1rb6r6i16nLHH9HgL6Pp1Xm
Oc7fvTp/r6Q7HCVKqMeDVX/RIcGO+/Bqgnpor55kVNc2wDrgt1Y9c9bXjcsMQQVS
6fNC5aCM7e+El3qpR/WtyrxL0Fvn7b8gmHmvE7SDKqKOCCroTZy65yC8KZ1c/+nK
aWCJgu0QL85c6hLdPXhXhe/g0sxk8Zwmx1rPdNEk6EEna6FAklgnn+vFOe3cpo/N
XeFXgUNYN9yGlnl+tFFC0vEmDJ7JAsU7D8+qwpQmLPwoBA7rYhTfVojfy7+5gskC
7XDFLj2a/T8IhQ7yhZmD6aUGsWxmjbyS8eR+tXCLDIuDdkQec71h0gpMWmEO9gyo
C2SYPDxslzckebALPEGzFcp1PoAJG3l/NSwf6YPPUbMAGOQEI+qBGN62wTgRlH3U
OYaCk5epLv+qV0FaojA5r/6btdeoBzEfeERUS+Mu+SUrpNC4LvFe7wMdAieFAsx+
ApDJUIFGveq6CvfEFmooACgPMyZBMhbY98f0rEVCPZKR1CjW+lhctnSQla0HAI7l
b862Er7urO/YiCtFNBTXDFGI88ssHkWcvF4WPcVs8lr6w+bz+UKM5J2114cG2zJD
dC/3GWGOU1e1y33qzghn5HXzJaxTrbcx/noPhmG6n896t2MyCBUDtQmlv84TEp08
+TIY/GEhqPdhGFmPSCU/dQtfPRQgHzrxPxwzBUtEd4dQ8Z7qTZPULqKXffAS2+/c
JTVpysc99CAJqpYRetFa8FWFoLIRDMMI28G9odefMZ4A+taavgU2oEC7hIORauZL
PK+udddNCHnDYCKurfop+VIsnEPB5hxGfcCFtqKFKgz8z1mNg1gyJeO0+sy9ALb1
ch6oxL639+UXGMd5SfNZ1sanvCKro6kHO4I5FW9NTxj6BPyZ1nccmRPOJb/oLt8b
ZHqdm6y53FghZt/gsThAca0Ne+ZMGUqJABBWJWrX529JoRE9/ggXNWAHtAHaHgBa
w8FN3F7zMWKZUy+0xNrho1UyCPlgpSF1ry7g2Ug89qG8SrafjzDIIuvwKLRUgxmN
57RQYU6QgGByPlpSUabmvcivPQZm1eZzBtAVLkRqEt0yoDP1Ny4DCjNlAF04tqRN
MlUPKaHrjDZJrBLbyUOzRbqSvdylEHWh24w+gqFJllHz1x3voGkW9tWf9zZKI4p4
CEw9kO9Y58c2twSaMQOocBxXTcX10x3bOHikiul0J+kF3aZFCtTn5cBpPP3F9zFv
KvTel6D5h7DDQeGLd5hDKS7WBU0/8rM0n0xuY9x/it/DoqwETE9C8A+LnA3MbcWD
Qzwkw4ODHvlQVyRwAn4fbrxnq2D4/oap/pC2jQ5W/qJuSHNpbOcvm75n3Psa+gX0
97OWeh/iKSM/sR1vxaCrbfIMxoQ9ds724lkqcP59Wu8yJqGx+atG4gnKWzmrVN7C
1S6M0vE5ObwfcPrwtG5dnTC31ndqktfWBB8HvnP0YRkHzoCDL4WJgieqfbVxu6Hh
aBnvCP7tTWaiqIfiO4+yRbt8EQ79ALGfXQGU0x5/69hTa7jFUa76IxfWy6/VKdYi
QvdMkQx8nbq/SnAMZB982FrMiY0jElGWrAQ3iELHRGyIub/Xd8pwjdCCwyNwHivw
90rDejVkrz8zS0DjskJsvAIySW0R+CgTiI99fxVkb/ufTqleoq54NLQv8nutixtm
m4I1lV7YgaDU1kmjO/xlqaaggj0yVUGkg8fTHOjcZxK5gxV+g+o3KGU9XySA879o
BVAl1SrHKIkWpWuikfFxiuz0NjvjtYk7YUrsLae+rNH99Chlxr+KTD65c2G1Nu0M
Yc4OM4sSDncfsoIxbtpp2vvPoWOhEQ+5YN1bVQSJV0AujFuaFL030sJWcDM7OtYV
uBq/66oAZBxWJH4Xjf+rmS+rq28lS6gJO3naCZl7EEUHZnveO1w1Fgco2eQuLWrI
dHtnyX2Vo5uFZBGXxW7weymGs98Zl3VS708HFaeWAAnlKjw9p9WrEKj8OMov3UrO
dbjsUYUA2M8z+ktTW/8m1x+xInbmVi3ZeqeNBEhB+yplkMkdafTHBA3W+UTi0QV9
qwBu/jftWFAfniDnEoBkVBifg77TINJXj2aR4J6sW/2xK8mU4kvOJbbbHBLJ8CLd
TRbIJqfA/v2a+aXB8TkSIhvzVAvYbuUIPgOIpLf1VEg6aMIOF6RlBYmleq7KUHw3
WT0NKlkcTqZ/69GEPlNYX/rp/LCNxoEYQjGB0d55CJ9cNje0B9Ma1cQOYy4RRrUh
HLjDxXxc32Dn42NjwheKZLvhNxVUf97YWhGZ92mqQaD0f6soLqaK5JHSb+lhSQs4
CrI9VN2uvOR84yrH+e0oiQ2LCHeqAQgg+0W8sLsWH3dUq6h5Q0oB+6QTnLpAK2i5
Y834Og228DLwQ8+Hv0wW6k2kUn0hrqs5xH6Ny0eGcaPonKL8Bmn19oqKLFcIA20S
5jsh3t9/APV3umUtFUIQd37NsOHl105mYCnL8GMYzZFP/iLiiB5PMO+5CWCqbLhu
do5fAh0bgcJtyNxfIOM4KDzy44P9xVdmXrF95eyIRjx6LvpObqsThtuRdPo692yk
/x7MW0vwjkxK5Es7AHhzT7ntZPv9BCFuUqll/k51LAvRibuedyvxtopT+iQufXwh
RRgs2SqSndkN1Aa64lK/jFw56zOFRbjmvSup7UjV0ZObgwXCWJsBmRpBo14aM+vM
W3WUBLO9d9Z66mh3rwVnU/lzV0HyT/SrRfQVR/kpuDmsZT9uPPeFFX/rqzt4115L
vkyNSZEVBfAnJzdytPnFmLXVCCpg2URHLJ3v+gKSrKtg171i5tAO5+HFmRog4nID
9fDlcvhkM8swTvYjOFvWog79Y6heF1ZvBgPPXAl2FZRNbirFiIfZq5ciZNocuwSi
IuoYXKbr0e7Wn9LG+yFhK09JQmJ+HFRsvuDWvI018gpVVSFPrDlrlpHkUrqHLjoa
2AT98CRBBGeEECVSPVeOPkKxvOA5NaeAgFUKNJu3AbI+VUm4uu5BrU9fdn8S8bSJ
61FoOrv5+DLQXVGkOscADURo8nlP5l8kTj6gu3ay2J1VvrN7Dz+Sa4FuGqLxJAKC
4UyOkHo3CXdIMpSD/h58NaEpiKveO9IQ7H7PQgaeP0y11gny+N8XfwdwPXT4LqNk
tgHU2T+kkZg0QjL4WjomCenDPn8x4E7dk8YgqeP0HMiBvg48G0SdmuIWzHKVttiG
d5AnRw96/QzZqLpgpysYhTM3PxScywIHUvEpqAKwNh3zdJj+ukaghUDsZA/4I8sA
5k6db6TZasGTVPLvLJarcMt0UQrVFyu0e5MGr5n5TJIFw9/M2nUewA6AzgW4Wrfl
ZnudjLq8PITjB9SIau2pxO6EEGPxhXEDFMNNMswtVVNTzrMTl5oGPn9uQzFhDpP5
saDkmDAebJoASiHPsrhnB+rp3N4WqhMQKarICsgTW+2sh19PldaTGsw3gj7fjx+z
OUnTpPziNw9ZCsAb5bwqGYXXr2VmFm8yNWO3lQwp0VAZxFE/XB48qtLT+4yg4M9g
ap8HRCMm57KilZ9HPafN5PduVer7uJDb2w2ci/mLfdpAf1+EXRF29R08jE2r0Goy
jGE5daBYUxOw3OSyE5dxSjd+NQLAR5CZyhXxEAZyIISIZG0He7pZTfHXZdTVujTV
fUkmaf17f7yc1hbnGnUvV127CjMNTBzEGOqvKF+mKQa1xCnXvbw+9xxKhScYT140
nE8bC1Fh9abyosSS5LHRZQLnUqtJMiC9Bnqu3RhqHyuoqwhoSPI8z7XHc7tHCSR3
hHtYHzfFmR8LPjL01+NIWeL5cAKotRkqMY5/MH5GRWJnmKU64l4k0YOVtwrahn1y
We6jkkAWh4IiFpbZeWdwDYSijbDp/3ISpUNvM/N4JeKA3M/nEmgrqrdQvuuKDyO8
Um4GJfQE/PO0N9tnB3wxeQC8xC1AQW5qOQu1O3YsPmOPHH7V+IsqhfA2K8V2vQlO
7CUb+YIaZu/A2SK2MWS2d0iUxyCkTXTdFQOfvpMcZ694ANLJ5IdP4wmKEA52dZ+H
/1moT3RsTdcrbN0hlo4j1lIAEV29gcR9dJwgisg8nauHHas9h4eteYcuNnZQTwqY
NAmMZ5Xety1evKmu2atM0GmUeN0w+K4QR3ikSimOgbv2OdcX3ZabAvulr6ViNGO2
AT2Nl5qn+tEKsUeAPeIOz0tRs+oGiPIoizY89SQaRqxQdTSZFTfGaFQNPCI0UJ5u
74GgsoIGu1yzofzgYenNKZpjxDUQu+IkQtTxNNtgqHg0wOEHJkgpBP/r8ddSXmuF
lrM/SjoxEesVWTYxLpLsAR7zmGtKcRn+SSByF9eGvIAk9TR7gREmfNuTTaj2/BhX
s4U+OmgkoFCrRbnUjcriy4yxjJNA8eiiVAgUxgyMagMDZkkhuJpiPWsrKesRxGqE
ufnuDHXw3XFYojStU5RMyngcB3HJtZr+RQlcF/1ls+i2KqPRX6oYNfdmk1+GZgws
wMS0Dhy1TgytPBN66UahhwTFot8a9Sz6X5bfsgoqolciDd2pQf4Y9NmKdXErlI82
utovvfsANDBNNzxdPswOQFUCQMXHkBkPGpQEzDmZYqaXIJN9TWxEXeb8c9rCUcuS
D5ZpwZGwHdxO3f8hEZYtf0jjnv0TMLpuqKf9+TV6v6cfm7hYaBoWU4yJNiWa2Drj
3Rmvmsx74Xnjn3aoMupTrLHkCzZjfBxj9s8nJvTp6vXIk3T7abSD9SCzKPHzi2li
KDKe42CCpXgQ6yHp5IjFgwF/ACtRoonLRH56IhFVCcmVRi1zp7D1aqiL64IU7JkH
tXm6AKRVJG87vXHiB0opVKRj3ka1GVl7a8Vad9NBtTgUI8jywyPoo/rAyW09eWsk
rdFvP2Txx6JqakEukrREgCJ1/n4CVEoJsHb2oQbgSWEFB19Hng9zh3AKxaf3VKCQ
w6ekDWEaJ96avk6SUucF8N7zVCq+duPgO9QHemt6f8guFGyDBol/3KkKFXkjY2Pq
YeZcdzfKJuShM4aE2snK+OVlAfzaT2bJVGPxYEtDjV+uVB8Ab3u5aV5Z0NCQG22I
pAbzkGSvzoMdW4Rx9Z8Mx5CeWXk+EEUdur3YivTCabwnVSz2f61dNcP0ezkSUNw2
k2cPA6ySZ3Uwcez2I/7cUWquqKFzBQm+/ivUOjqfIvW4BXNjAJGIhfIxtjz5Nnmq
qaXV7L56L1SX/8BqalX0y0L9lokk7yQFFnVmbDA+ZkGSnVrfdJxgfB9GUt321UAc
Dehm75BZNfWtxfuzIWv3jnjM06bIMsm+O/tG9gTQbn2yCZQhuieYhcR8DbgNDAsb
YA1ERhcrOQ2IDcu/VrNoOEq6gnGCd5NZKYC1h/k0MKChKiwQoB/oQu4g5t9kLgQj
b+xDyTcwZ65DBKBN5hGwfg/JWFcBwObQEbM77SdLCE/TuyhlJ6SGYpcvZ1RWqVHj
J9c+5zLnbCx1foso8t79UjvXTzYGBxW+nRI/Bl9w+3oOIXDPlvIrOEhE705Ia8Er
GkBf4N34XyySVk6LP0LoAoe2PRUKMeIMTKchAZu7HYCx29vm8USqE+cd+OFNIXyt
Pu9J2c1pwNpvsMLSxL/jW6zd+ZBhqdQoKTL3yI80wrAM+zAdCuYuUtpMT0SD63Bm
WAi+yS/3IxDnSI9A5Iy89zYKb9dNEVOWtUiJdYibGLr0wdsQIdQjaWFRCpMT2Iia
6o5KASSj9FuvTcPLnGPtyYMfUR0iCIwGqjq8o3go3K+pC9n38RfwaBv30cDezLfq
6MDiWJX1C8le3RS2pOM3Mve5wE9XdRVrqqm7V2yz/CasoEPDBefckuMW8v4TA6b5
cGRxrmDWW2437Pf5CTcabIz8BDTgrsmBLad4ZqpmjVX/Evh8zPbNax7dZjzOZN4K
WkyePa+ti9X3TxC6JMjQTBWwgONYp8DlmcGqSJG23GP3gg/bR4N+KLYiJNIpmGSf
Ir9LU0ax80h1bUuXaEZv69MWOboBfexX9L4XbZT3WIycACjtKFsWg6IZAE2OFf6o
sStAuar5cXgW2YbPj/mnHojCIrQeVGSB/MtyAui43jvxYW3+j5xSOmnK/AV0T8oq
q3fAqIloXFxHgTQzjFsqQdRwaHiZs2z5q0iyAvRXF+CI6ReB6vQojYVR7uhF4NpE
d5gKLqaq+rfJ5lxRCD6IaLtNygl0/RR692ZejBiORZwZTQXu/BYNX4heeP3ACEFU
6Nuh2U5IXMGBC7DtsMG7SS44Pa/CQRA8hQ3ZkAZynCdhm2kQ1hElse6iwBLe6G5a
8b8aLLbzVKLPpHPmpfIe2IhpHPWQkUVxfFljpG9UYp1FZbyAf1tVSTv51avBERB/
9nWFHQZ3XvRd08eq/6k996a5f9nWXHgpPmHPXabwl3cmPMwiV5SZdjA6lWmbXpPT
WhRU4XZKlluHededC/uWRsUGaCAtwMqXlZIwrW1rJ6AadP8gV2h7D3pFDFkpgRLI
QMKZ+vhupZ/8pwr27DzTgCfka/Ns2KhK6Iv4p/w5VCQ6UoZ9+6tFRU5RTcfxk9kA
HUX8hV7VigkW6NRLdchT6+stBXOiic8DN7ib/FJir46hcTQ9xT4yJK+ZRgr2d5fP
GL2chBNPf0JaF0kcxZB0EHtlpjfuxoUlZ+hGGVGSj6PAOyMSdvwAeVfCuJ4r0t1y
dB8y9C4Bipfal/WUhF3q9msarx4ARcjmjmfkJ8wgiKtACIfcIFYTUPxxXananGHt
VfoptWg8yoQsWVLv7MHs2O0mLDsznch2n/Tv8M5y4oXQAcJbCM87TogUtMP+m3/8
1f9MnBuOa1OaXxSsa0Rw07e2qFleHshqEIbz8MaEUCQUntATJ3kC4Nk69N+jYO24
pBWpxjSm6Bqx4fWoSD1nBlCSu2r4k5r2aE3YMr48lp0sJ0LxQrQNotISMO+7BO0v
BHu0SwNPXuR5z4Z/ZiCWp/AQTLAi7KbDuD2YtVUCiSAm7sLMwZmftxG31UIrsKj+
pXbW23KZhzuq5lVNnXf2YReC8ymMZomgO9bTq7NaVLPudDDKwHdjk+39IN7HhcNw
S7L3TiLjMT2m9kxkSpVTwv0hjVuBtNgLfJzuehSxxTCuXskB3OdmFvqDUurU0Juf
q/smqHtbxnIg9XOmBFZmHub8g1pkmaIEVffEZLHEnh2J5BjlCB3JlDvreaeGVksX
HguW0oHXAdEHXafeUDgjBUpPXK+O4qR1C5X5U/Qr7VsgmA0EtdoaovmkIx343owx
--pragma protect end_data_block
--pragma protect digest_block
+2uMTb6hUZ0iFopZ+zC+7i15y2k=
--pragma protect end_digest_block
--pragma protect end_protected
