-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
SUeZ4WL9sKrvzf3CtFBQM78OAh3KuQExumTOTaD+fXesdZrWrEvVpK5j1dbZitCW
p3kWOg2vyF/9Fe2GczzrGz6i9kMkyIhotSXD8Z6rFVAvVaps+SuCTPp7rKb3DHEl
WaYceUWtxrkJlRnyNVv4HQnDf7ZBgAgrEIPQUSQ29Bc=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 10018)

`protect DATA_BLOCK
s2PDJZkp7HZZeAujWXQNIxP0rNsfkvwJicsjsUXaB3kHsQTNMwsQktQiD0g+y52v
DafYAK89Rq6mHAnQ9flfeJViMO5k2AygoqcIn0XkwrAddTecJz4sym5kPHWH8drc
cTqfK2wJo+yfXqnGIHFQXR09fkPM+51e1lcW1HqZ6+B5M4KTXAIjqqZwzwYwUBo5
RdKeYoOsU/WJU/355lRHbR+Sq2PVGEyIs0NHnvRVzrgTtTzrtOw5x4S/VKJD9mCO
nRrUX8FjnX0HwJxE1KTlla1ICmLgUUrY4oe1SCMsr0iy9p4UhUxHq9LbZzxMvnT8
A6r257Iton4AUjNDVMXEGjKAfB2vKSfzz6YLxrwY98cKvuE0q/XGJ61UfPVey1aO
KXIkiIgledgTlULJGheV97hawpN5IheF0llTxS2qD1+n03yAkPzb1kQaG2Mg5zM5
bZ0QDeW79bbnwA39wchUNVK/7BHtgdIC6V8WeVuo1VOdnrc7yHfYj+4UMomOHdkg
qTU3F8NxfeUjvDlKq+bxC/JOIlqzCVwsWt5ZzvQWJGS5L2n3TAjv3tXSaPk0FtgG
pfI4yssZfCFDwnPd5G0G7MAGTl9PWK90GrB9EZL2qxk4GJPnvt7l8091EK1KdMyb
FHjhQGpU1GARMFdPExRGWoPHmWFPe5L1iyZr8c9zjpTJAzWHTd0OahmJ7aYN2HiQ
WVTMc8ZGXM/R1+EnqiE5ylpm7EpXU1D/snQm1CpHDHkTkqvG/EXzPN0UEIAgY5mp
IkC7ic1zc32dngT8nH69YfQYFvMdMj2YFwszScUFfnNLc2jONUfzjBV8IgKZTvCM
O0R8NvKKBrIX4KlMwGtcQOGody1CFA22j6ARDlL1ErfD/I7wSjd03tI4aeilclt+
OYOEdaulR+tbUk7uWpdrWf92cnKn+Gd7DwaxRGr+G8brpcu9zef4gtWTyxPYU/XL
uxWbT3e41sakMjY1bmy+2xuNw49iCW2DKhTVB0cffg+a1bI2Q0jCd0Zdt6E7i4Ur
QPptZUhnHpqtayyuSWfccVIQx4puGjs6R3JqibfVBqE/67aGX8nX28HAn7gYrTg8
b3aJNhBcqv4VfJq0BF1v8f+VlUcYUSHsiflziiC7kU2Yv/XMLZoYljdcdL2ZzZDf
71zZbd2XVF9uvgxGZYywpg1zlzda5nh5RfnzL8T0BmRN7sfntohrhoo9a6w1xkWK
8Ic1SHyx8W2S7KsM+8gnwBO71jjKT3AsaZlvtdr7SMcCQmHofYHTrOWkVYYuJGh4
NTukXvsBHozlNe1gQ0sPCxECEGj3wKtYP60E0gVNDCHylU0emuudHhn/Bghl/8X6
XEQvG82+5pk0A8SNVszvaSOBtztqiNeCdXLNCyi4oYOJKYTlTQtX+9gZDU/sy+j8
pEs1rJqZXI2lSTG+LX5WvyfeofFCwimrV4C/WzpjAc81ge5h5kQl+Ydb2tN2djc8
5NdHsFG3tw3gT2QgQ1jmuNEtuedDd5xqvbBfB8iugTbmD/BP/1RgCJormrQ6QjjN
F7qQxbxapryyUltFnIBEPbEG3gW3xowFROZ4MjS34G6d0iI5ZKQjpQPZbE3B+PWS
+8Rzl7vTm++OVDBxICg3fTXUTVDsHe9Y6ArBaVVfCqxnDiNvEYjlu2Ubn1DWwnzK
X2b5rk0PSi8vuf5YjvpEv1KSQ4veaI8V+DDMk7FO0WTP9j2MhsqCJLjrLpVDAxFY
ipACpiVhq7rG8/nV1PHvd/H90GT2i8VLQWxpdtqwHOL2lue+gJXgVK1zTYdflCVD
SvcMO/GrUNeym8LA6rPGEWkBSyJAWpJ+2yfFrTsR3OtiHQisy3pBCugykLJ7WS3K
p7vkGqYbtDzFIynLJKvzSs0H00/R5Pi/KGrTHaSL2sHvqDQ2BUZZeVgyiuK4pPeG
ICgm4LK44Qz/KC8T8ve4dvzfpPG6NPTSCoxShG48RHMFKe0iLpfPRlfdJR81mjKv
O4ptGAl59vTgyirQYjU8yBiDCCV6i+JcBKyA9+w3eAafvvgHSw3RddWROEwlUi7D
l2RAe/1N4ijqciGkk45McGCnZWCpefyUpnRDhM5hG0+TgO32H0sbls99buxB8iLV
lTEZcCrjDIE904qWVVJGgUNC8tBoSn16A5Klzq4/4f/WbygkS3iaG1kWHcyrKiTP
Wudbz0WshTxBYVlKhHhM/zIOXf7YGLA7T9g0vNuGyNqDqyFbfcj6pJdMhWywNM3V
pVvknHa6VdnasVkPboERHYPqzthfioOfGIEARPOduiS+Y9UEquMT2Hg/UcSI+ITm
u2l+9jRrdDvKY+hfKzXXmnbWc7hmRE51ApZsFf3NiveOpF8ibYY39vJzaz/AaK7j
CfakKUs8cPLl+AJeiwvboS/3ryrh/FDNHO+CLUd8ynW7rIbreI0fOuJbVbofyEeM
HZays2qQw29SgOg8gfw6hClpaV0uk5gW1tW9rWQ2bkSJoc/7Jr36ajCi9+TWkZEX
eiLkLSsJiVBL/6R/0vE9CO4LQN/J6g2O6n8P368PrX+XM0VPu5fgs1ZyhdXCWSF2
LnRezEuxnd5dnp5TzBHYjBDJGaTZOFfcLc+q1nLLbXLkl7hVQffLoda+bk1iN7SQ
fT+ALiapxrCYtTKXy+zzOteepGPqEoGnfdF05SaSkg1i/tW8lp407mprTGbdOCXW
cOvn3JnPoblvVmz3ixhhbFiNRZQx7SZxveopX1tO3peye9e8AIGGxYDFoJI3abEy
hgmoG+A/YnirzFwRgP5LZDyMIES6F6whDs3QZbDspVjLeYAlpFPUm+lXjwzfQBak
TCR+w/pzjxcBErMgrjgBsrls0bxWmNPt+ngmf0MhnyBCRGxzgTryloj5XyiHVHyd
ZjgM4OBUUzOP/cNYrx9pHqa3FDFugZNP6jwAt/XxC3416PxcLjYImvFUkFtWumfl
hy9WGGj89isEmJLhYolTmVK+ZCsjIs1kVs6oHRCPXa4iKFjKjLWU424ypZTeaTBh
udbRKOkicJ7Obidy9OH4RZtzdY6swb9lZukclh+JmxqC6dLA6bDgDT4HqKd/NB9K
feq42r1BCzS01oOXO7xk2VRKMSMGTW95v9qnRTEgMDjQdAo7ASqvWPDmfEXRjEwp
R0KxXsRnX9yjieKSZWP/vU9lwH0JSZdnVXxovHjBXqcbd+GbY1mMLNssKus+rvpe
xUrWI8ASqDv65YLRQu6F/eJzRWtc6alcP77uIOLc9vlT+Te5hCeVf4J7woojOfWH
UuokQ1uhChtL+F8Ha43zBxcSbeChQJYJBxODn6edWYyqSe6h+hA2cq49kK+93frn
oZ3MrQFUb6aSk1g+C9Q5Nt1aueBIBDqpCpJvS0/MPGKXwadz6n/6ClYBxQo0WlOR
SQXCyj2tvwl5RioueYBaMAmrQorpBFjTqHIQYRUsX3LGaQzcVUis+Nr/fSKx+0NR
NFMH3rtiHbtlAbCWnyWwEjR3TlmPjYpwLPO07w6LOnuyUJMtVtqrKeX/InZsRnua
9ym7Y89FiDxqM8i0rmI5he1Hzo55+cYBNSnwbAQFDTB2dwVG9bQb/9FCjO+uLrNu
Jeb+zwfZBSLF/n7FMfuHYQkfrrx5qmDv+aqQPSPdd8srSCfmYG+CrEjwnJOgDrvK
YQLrgx+3qQwyyGVuWgbOZFWYqX2HoCtUDxE1jpJlJtnzsUgzwypfzGFwK4jrgtlO
JG7PrB4KkVN9iMKJJ1Exk03s03w9zCFlbTLm3tgeZxDr1X6xop0kYta0sLqz4ibI
Yx95Ty2kkaYg4awiz7ExIiBQr51zC9ouPeCzPkThtjn+0a61yuy9I3ox+2ke78Gb
uO41Be/CJmlZzs1sc6Vj6lUr2UtoOtJpAcgm9Ky9qL9T5Y4Gb+bPEWHWIUiCiqhP
ertN/cnsqintLTAgDJEjVFCZCt0oBTFwtAg5KrjQVBHhD+fK1ir2wZoqGplOKcuF
rwFiZM67nibuTPbLEPpOow08affcdL/baQ4bdTd5weojdiHK1+Url+PRKGbkLlMJ
ajLe1477giKJbgkMDFq/PfFkQ7q8hB1Pe8qyWO8su7oNQ5wu6KHfuEGFw/y+75zr
3xz2R/dgbjW8HxHnul8fGoygKEKXn2l4IwnnHuFmLWYXYe9lSpu5GLpB6AgPQL/u
+zBNn0YIgKLPbOzL6kzYcNsqb/2+lE+2Lv3VzjtHaRUtZo/pFRbfsE5y7IXjw2pt
mjFwJmXgeRGdVbvvF1oWXC5GiGdXkStJbpCw+C86OcCAZN61f2PnxSfr48ffUTha
CpUSr7q+s+EQGB3DDABipO2mzivC25vApdF8QHhQITmJPmc6j7T8dw0+3DsrF25X
77SRLrgDuYTdWnymuJVjPcCBBTayT+d6WfO54W9QvXSIUU6dEYCO+b9v28FKNG75
MzNDKPvcj/yWaAy8cZaz4S+2Il5oLNlNYurnQS0J8EBO4rrwgZ6bfB9MtET8tUiG
lqz114hj+cCAeaXmp74brI5lwt76JHkpxmOVm7wEM7DTsPngeV6CC8D/tafLIQdA
XRwgwaUT9ygX6OR7/ZlD99/l6ykpZyjk8kRlZat43IP1UQSFhqV17Evgyy3c2Cd7
d9/Ch9aPqXnySKR0l4ZCpV/cWndKEWXWgRkgWXlZGQtFB0GQ6ZeA6cL3d1R16ZwK
x+lhxJMY1qE02fekGbkD/Ai86AkL6uWHfdZ43y5XDDOj7WVqURudxw8AbSozATj7
sARfxiOSrqeQNhbXHwYnB2u8t/Y4gIAIstuLSW9VLS37H6+HkWhmxlKGW09ygS/Z
R4OPOmS3l3so4aWMRHPK+TmcB9ky6ZjGX9CFs15nLC4AbTXDBHcCMmHoUVz4X+JX
TOJrP2ej/J6DSm5GYh/gcGirXZOvvwUwiLUSTEAcgqHk1xrrhDoc75JNFO8vOR9l
1BLE4JY3o/6A4NiH5ir/qbLGVNzF9VrYyABJoItj3tqT5bFKHn/gN/fSWJHIhjXP
Esl5+7IUDrSnycLkMrzr83Qglotw1eXL3r0YNt4g9lk1tlcga/D0BPpmr49HoWHE
MZqSR2N1i79stWA80XoPZSmXjqWw5Br1USvOKCOdvqkZhy2xCGrhpL+eNINCs6tJ
nYml0/vW1Xv5iewoscB96/nhLgtOx+WCKjyycEpHbUYLjeIBOypQQBm0b6bdzcB4
+OWO/cHaAirvKM5iirFX7NEBJ0hfHJj4i3Vgr3KdgPo66/tbHzfzuy0X3cRikMR/
EdZ+xSZGgizRmBmauJN2CYSAj4L43Wyzlcub7BqavbU4/HeUPT3LNqeLfObQhEet
ZQs/EYHmHb14/uTWYEPtHqaVRxgnXqyuDTyPg9tH6TBxC5cn9WHPtNpiFE3G0Bvy
fhFwsoc8C7YlcyyNRD79MsekY9NFX1ahAZ09FVG8Heo7g2MLRFMbH+dZiDDws1GP
XNK2XnYPe6h32/StvIiMdNoeGYAMedsYqtMih3kbs8PHiu3ksHOlNyj1T6S4DCsH
v8+99jV2FS594O3zwaBdyzuSWWBr0CgMo68+UiTcgj7+zOM1RQdULEPBR3RoP6GV
s6NlFp4Jr+68xvbioLlhqz8U2Iq6nLrzGVLRY97mloLmTehK+j2xlJWgce/IdMQs
YfFa3Wa5AUoMiLrqJWionDC2lnBbSvZSDLGBzv0IR0yCEdJKDilXF9+prGywbBIe
WHrmgwjRQg7gTlB1AHE+LWmu9jTfk7NxV7wFoYedtB2L/+hd0YPj4rLXYd4uXUdh
Q3vBiC2ybtwW3LNpVLbGJ25BkrAFKFTlATiexrAs0eeV+mjSuRchzCY1lQbb1LEf
KoaTikYjuuIEHVu38gNZW0XeMgCU1Lbs2jrPRe6ZJRN8EpK7YY7qrWnaDyLuBiNT
lsZ5Mzh1ZLof5yE2vSCeopXWwZ1k7QgUCW8CgE3hlq9wArEVbfxGHKgzwWtTrgA3
aIN06DaMHDd5rEMLz1UsM6/KY6HXq1xJFsduTKzu9nTWVG3itlnxBEfi8o524rAA
+wcf/+QtcSA/8tLvAQfs8Ok+Dq9biQ7lfAtHqXF+yUfEFxNnOROoiXrILlIyb8Li
MzTSFG+yMGwiDbrtAV0n6fyy97IKdyHkNW1Tk7Y9y7eCAEYnb2tVa6FgGJbRtMes
3OolUwV3qXUtfNWDhKPydO/qtExsGRxE92+3WhrkWZhTG4qtwBn2J/HJdfO9Fnuj
J/cllg2lHWAJle2n+gZkUxjHdCn885+RRw+uvEgyvw/KI7pDAFWbbRrSbBeLoFAD
gHwI38oLk5cSfETSaJyFSN+TgHKBByKIXgSlofTh1C17/TjZvTZVLjF29VNaSIR1
L6JzE+nqBznVAOEACyu2plVbdgL1kk02nvyii1Op4IvTvSumfCNdd2gZyF5FD6y7
SEbM/ZLTV25JReIeNLX8Yma6AQe3wNGzmaYuavyRXoyHJYqi0r98qG4T4SjxOxiT
mSQ4cQYMtVWuIhC/7sS0Se92z8B5047e+gwJpe4vTU4kDG7Ml1hm/MtkQXCPQIfi
DSzMLZ88t5YjocL3QmYb3LvS03RdcqElV3rs2OkypTwwMhzW/ZhDvT1QLcze4Mdx
gXatQmd42rMrSKdWjifATVJzVgzM7XyU4R2VZln19Iu8HVVJzplaUtofu9YF+rJB
yMnC7cKpRTMFWxOarBm5jqUypUStUu/gCzvowH+R4IvFMPzp2G6OTD7nND22Bd3P
lrGMMMuekEy30SLguIti00cQc83muitYNj0caOothSBjDq5+Hj2ogNQ3aL1uLlQw
4YVMw0UJjsV32joTABSNWgSXYz+yYXHCAK1uopAkqNhKeHAuO8vBnq1M8pH07j+w
lAeFVBxmzU7Fjt+KSlHf6c3fd2JGX6tIYHi/M8DZAQn+QFNSXEFH6WJbFljG7tBX
wjjdrk155hGpvxu/ubtoTE9ayn58DQCV6kFQLwl5GYmieznOrMQIgXK72WECpAse
rA2lO+Mx+d4Dn+vWFBPJyPASAPmRb3A99fR77MNe2bLIDFKQtUY+mCRWZXrIihL/
k5DQbT5mJWaSbCf96mu1+nuegx5aADQxybBZ8MzC5OBSJSuBNDtvTo0NBgwel49B
0eImSWZTsqXmxSAeGpK+vuAVwSCGU7Y2mQjOfdwjO3q/SArt06MMF5U/A8yCS5QG
XiCLbmw650B4bXOyvnNuGiv+oWQNfGA5WQf/F2+9zkyHWhhss9j7x4zZ5wf2u36T
y7vjHKmk0YfUjPkHOdCD6u15UwE9EWw7UQqH0FOtmSaN+yyRt0/EtWMWTp93zZnw
Y3EKf+GrYIKzEz8p9o4rZhhSgqLlxqTthS8doNfRTUqHc46A5eufJRQyo8RIpV95
SfPw0MR1Rx7ZgriDm5QEYjytN0Ce3NzZM9y5PEfL35dCi9K1wkYZGgBMkqYXOSkB
hkWTJ6gHg+nEF18K3SFgq/dXDM7iuigAgWd8hORd7eDKOYtkAk2FLAslN2rgnk+s
UOdobiQ511rmWBdweK7gZRbnGVb45gv0IrBzgegjCdMP5wLDealN0EesLPPEmd3l
Pfo5Iul4eMCxhfZ3h3OCbTVeqHrrVcP6fSev64aZKto8v/CNegQQttnAQwH6Xog+
VpC3GuhATM2BeqVfQpNV3bMdOZh7YqLPPaRx9FqS0J7Skc+R72YrTzMDjL8HXONe
cD1jz15HyW4kdDIHzeXFBTpMzC4TDeXlOqVB14Sl1cqkNdKMxwDVd/0r6YpHWnWs
7cXFyMNHSKBi3XVvsCi6eFaS8B7VOmtbCZPMAZ6KhUU6pK1snoPfgr8PR20Tltw0
ETgL6Pk8Q0IHzxKnXmYW7xMDA2xBGuJ4GIJlnq+PuwhzyHW6xmBSXfwdwuBHZGxL
0inYwzrN/FSXX51L3EIu3eIk57pEyuw0T0hulGXmkpdyk263ErbtA4Q4qlIFRIxi
4/bVSjMCxJGPf+VG72kTfH42WM8ArPlIH8IvedChfmsqS5yIwvN9l7kmtC+QctOE
qLI1HpVbIiDcmufB338V8ph0KDGBDzFXNZZ/+BDgT3BtBCrBrcFUR/XEiVMLqh8W
M2VjNM9pRjhpoyJ0SwtcGKItd7zywc8UIXfPQ9iC8wPF03dWcP8ZjJE0hsnTaHMv
3adCIFYoeffFLkfxMSWu8OcFe/la/YkomOfbE43sSRFdU9/92n2plIVHaEsu67hQ
wyJ+OJS7BK1Hn1Fj8gLi10+Y6AGdtrv2h+eVNDcUE5hbU5FepUhDb3UoKc7Mb/E0
ngYgcRxDT353YA9/uglvtdbzd1JXMNAwpD2Oz4YP5fr5gjtMb8pTHRFUNWNuo4Vf
jxKwRqcE1LAUVc9A1OZ8dVCyBboenmwS55Cv8vba9c81Gqb8AbKDLo2pvuKVt+8S
gLBb8dWIrIFPedJ6vIgUlA/0mXkCfU4TQwwbWIyS1eZ6VwYiDR3ZQw5Y6X4pQZ/f
5mZ9XGyFGCsPbN2lVxKIoVfwV6HuTHMWGZUR2MOzGfzO4+hY/tE4YiTwtz6y6D4I
eEBJcMeBJEqTju/r4kuAXn385apg7IALM++vDBkEoVds4Qbme7saOOkRpCt3s9W/
ISIBWrnig6y0Llzt8MAdSVf6RQkJFiCdvA/93oeBUJVEeOTN80HyJu2ARyg8EmBE
0QJaN/5uj7LY01LsN+0zrm/TPfYVlvI2H6keB+osdO/pfaIvrgzsamy2P+RvPPXI
tueZ4MHYZ/ZFKpnKoR04fSJHJCsxJ0/4C0/5vqnUnXCVT8fsj7Isy66o0aflEdGO
PEOZaKXnxHmLMpBPssLD+OUZch0PJb+3ZSyuqT1IBOC9NVRPLzkShMMChJXHrXcR
xJVw9JXkjhp8AnbmEPn2pjwUWwhbDNXIIARmCZbQN9yCkGF+onQAKDcJlG6+nU90
vm9C8bA2x9SeYWU3wW08KCuukqhjxVWqndcvpN7/qDICmOHWSiQBBMcHwEU0xaAI
GjaCzvhGVbccPLayd1u0W6t8uHyzkW147zey+W1KSr/+UYw8JvXz81wZHBqNZRoO
sKjmrdUmiMprdB+JKwqR9U93R/KYYHiZa+TZkmiMdFefLp9aT+ficr/0aePo3ENb
7qzDuPgyHMAKi1xSufOv+KL3Gs8VDVCgfJSds1xNzjOCdwuQ9wSREYf9O5nzTpA1
/UisMmFCSLj6ivzzaho/ncehcjAu8lfx1GYwK57Xpj67GiGFqSZsLjbpUfMtY1nH
a+Jna/O3bMX54fPaIXOaGdnG6p89ycPZQ14YNrQL4xs9AHw3/nT7EVeQX0+9WJGB
cy6AW1voJRVJ6xlFG6DTcQZQWYQBBDwguabgQUoHFhBk5utWSKrQxQ57HmpQLjrB
euHZsuToHp4l6HYkzD2HaOEPuM1KyT95dJnrlPSfrbiHtIwVAkNBVjd5AntZqlu2
3E+Sb4w8vfQeyVRANB/twG5qRjoilTmr67LbqxWq3oXfME4TibzgWKSKwGn89D4M
Nyh16XszI2HyQYIHeFtH+VchJDWPfSvJ9AWN40sQOYNtUQHf9YSDjfAH6fl2THZ0
xznRqG42qJwJsQFtu4X6CMWN6uIPoZSeoom3ugkdJYLC5VsSiGT1hGTTguLG+/Oq
FmY5QxDayy5SUkW+6hzzse5xWIIAlBsKcR0vPSVqwg63MTm5Ee7YG2VpaEQk7A7z
JmifGEV3dZil0ohflhAAzUFImKiU8Vh3MLIc/OpCGMAz2HYc1vtlpgwmnsEN/aaB
WKRMB6gfjILm8wPwCFgtkaW9ifVnISSPmdQ3Q2FxnMHXYgtT+vkKu9MPAuLOwUIQ
Nx1Ap4UUDJASYsJbt1Vjry9bDW4wsr5LTNwMyYwA6PQCzRJIIkKYAJvqx7UsEoa0
FRriSDsk8aBovU5OQvhBduJ0hxpQKV2MMMWXTQ2FUFglzqrJmGizD+hjGGO2Sja+
A4Mj7jAbAeYREHJaKXzOdAU/MuJqZdiIL/AO9e0XfMuG5EdcMYbfgZO4qlCLaN+K
r4ybElxk+Axr2xOA/tfszUI8bgfGRsqPb5tM00QgRBEAblM57lJJ+N8IXvLfpSpA
LXcLt71nwiCgtHZKBzYdGJR7LJE5QKUiUtu5NMZZfskH9JrAezOfvYORv9b+3/k3
nAQFl7lonzp2g8zi1hf4sIoKlErmMvfEVW+mVog3YOSoAnpLkX4zjFFrOukweVH6
dKEHCur1T2P5AaMAQvJYcsXqGIJ0BTvkNrhgptxI/9xJLTpUt4L0XWEX1JD219G8
ta0NJ4/C5mKO7RCzSgzhVyOGKie5vuPeqz+7f3DHT0TvXZq3pHsfKTODXOkjeYmh
ODRgcp55wJYgTPkCEOAGWhSegz+P458lT+lyI0AJBGBs3TDsWhNZRtASKXRmdn0M
gLcUw4ugZnRKZ6ajC3NONiG3ApWGj6HtEa+1OC8u55dNOfIZ4y1fAI9UAApVAS1j
Tma0rfZXOKnHYy8N3HBVsNUKbJ0hLFDsELF7dGIrr1FL/finaj2dq26iKigY8wF2
36TVRN3KE0F64JPVaDJxmK8qRQumPpNAgoFwlGlar1gy/pggnIZXtt1/LdufZjCV
Px4xkZzSkGDcSd5CFt2IJlvQkZWLsrBv68T1cIKsZtVU2th84A1GyjLQp3LOPy14
XNFiAQhY0yldvXUTYp2d0vEPBBjG641aTni+9GfC5VBg9Zl1bHH75XQAqXxnVpRI
m9iO4wM7Afl25atAvRJMMp5OLx19ZnjToR5g7w/cXp+MKffE2IK5OXzHmsnnOxBD
dmWEZpgOzzdEkoBugh82Mxk+czeo48nXY0fB5T70r9G13yjqlAOk/k1k03uDxA5T
u5XZNPmbXErwycRKTkAlCT3T9JbQ5luYNR7OB3WuciuEH/gxmZ8PnLNOA1ptnVle
xiuDkkMB2DpRKClvM6CMfasxWyF2z5rVkSA8/g/tXn6NZW7sml2o+56TReLKQDQg
RlkL9bg3fQ/Ln7kFdBQ2b2WQrApHoK9PwaysXAN9GLfBQj7rRR7DfUj210CvnMsv
56GHjWfwFI4gdnInWc/T7Mp/SrTEsMd/7vdkE7nqL5lBjdwgpEk0A6dchtmY+NbS
BPg18dr2XqVXiwFiz1e9BBdty99HI6G1Pu9BA3Eo0vPBozO4r+xJ3d6pajziTgKs
MNJUP6UpXSLWrf5azivhCb534oxS71b0DRFcRimmKhyKWD9fmlA0smlQPUoG5Ks/
KS5UKgxKERDepbzguz2MTVlEVEXZS8DmzzffdMae8EjVHDMmTX1Vftf6PST8S5fz
KwhWjBUcEnePjs9dZusNu0gq1eacPIT54XUZEgc8xCemyJLptudlWEzielIkww2T
oTk2v6d2rAqMsyyZFpJrGvjSEM7gawFKpUprJzwnRx/gvGum0+v6QFWg9UqSNvHx
wv5IxAzUEYpC4S7uPRvj8MFXClXpuAuHmYGLmiVMT/ir1/41N6tub/koI+5M0y5S
nhd/Bxl5DcAMbXPFVd70KDbT7MvZvVTweJ6tDr8Gq7X1TDfc5OJZvoVWRtBFDhlQ
x6CqVrO27DyZK9UjiYwZUP7C3NftAU9DR+E2AGGzfJpIRmZ2BnH/6dHvDWCgZfNc
gbIs6Z7QHuW8mEA98o1Oo3J5+TZH1l0GruaK3XEFx0TVGEhrNzAR/7nckOuLxE3n
naDW1KgIUt3pHr+ePF46BS3GEA0i62mKFZt/uYiLWOUFCOA/a0VDC6RAt8+i1eV/
ukbrnuP1LBq5VuYr+Xa4iQJhE1rD334qh0L+5NbRY1/i/24IZLX+23FBOn+N8H+n
5Cle/6UUV494JCBaOAartBMiO7Tu9QiX9+w7x6yBUYLLC5T8dt8eWSjvCWVB+g0y
0xmVmQ6TiMuurj9S/GiVdedeXzuCGrPbzqKxlaLdTJHDc3EhRrHFmIc48tJDbo/a
d0Y8O5gnWrG9LsP+VtzMZhcFgjxApLqGIO898bjvpHe7/CoNLT9cdKwgIIvZSLVc
jhbiEjJ9UP4CTX+D0IAhIm05UliKVKuhMHZc4H8PkF6zVHqAYEt1i3EG5vj0GcVB
GbCpwFsArci7G5RRzp+hxrWOk3VBWYheKDg4tl9Accw5qFX9ljrMgEmWI0o9WLbI
vRM0BkrU7x6/J8uchJhuK6DmT2UgW1LI0hvjKLTqp05614deHokEgZn3Q+TlsPrk
DvT+GlPGNyBu1+hzGEeeym7mjKnbPqVXtwqVLrv0zHj6vKgcBBLYNQOByc+baRPa
wnTWsk01GpW82S3IRfOeTvVcY8o7CF/65Q1LKtpreboifkud1oeypEZooJ9ysSub
gdwFFbvmo3T3F7iIUM1vJlnBPZU0clLlQGaUA4/MgzmBdFUEdnMX5QtnPECdtsRf
EEPGdqQcOl5Aw2+kWL9aP6PAjAhnZPoFUIdfD+nLD3PCAEColDlHaAxdAZEwAEz8
cDI1JE+zu69C56WJXBevrvYK+0N6KNe7EZv7l4t7afvK/9RNoVvVzZD3Q4lAX5qh
ZA21aX9W5LeyTEJCbZ5yOzaKNgJ8tRyLNUpafQebt/3KOJOTKITady9vFnF+wse8
Ri/Z1JYf41QMzk315hZFy1wB7BgR/Qea/jCXTy4krqEbF0vChhoVQSnsxjHYueQx
Zthq2vlKyauRCr1EeudkTnRhjhebe6udLTJmzuQZPmgR+DfNiYn5T5lH32EXkb+R
0oDONATTQ802MktVMxovLHCdCLwQDCyr3uD9Ij2lmGrCpGbqAJSPmYDeww57lajj
zCbVntPi6owG7Mjbt2UTuQlWV+5geVlvfTNjoQVyc2++QH1n56ahWyjngfrJ7D1N
v1A8ctmOAS1kdfmiFIT47hlwn3YiQrAdyVHTAxDs2Gpo6XEzpiI2XVnVnBvPa/xg
CRXs4PcEP1Z/2h7ktytGlaa9xlhb0TBUvkCvN0X6+qw1MRXqIlxhwAxLPkZVnjWu
C0zZSO2LTZQh0BbG0+J41rs/loBeOvOtoTUBSeNs+fGLm2MZjKS+RKOWRLV4LmAM
UOxPCMcumxgMhVe3mjqvffyTGJ8TbSscSKdnQfcL3hhPmX3Lx0YQZBIc86mV5XtY
2sBbj8iNAhyTr+L0/IjBKGKTZU7t4tjanf1Q7ziyVxX6DpBNfuXIzp380pQxIJYF
Fui/gV3PabJ6RzQaRqTslCpY/69vA03oB+dHvaSng9tuDIsKoge99gxNMUrI53CK
jas/eyqmOnSTbHjD2JAH4pl3rLxi1GvVW471Fece0rHU0t46ntcgzo78PjLi49LJ
cqO7w9Xtbsy62fZsMRorqJvXMHtMVMyvFkuHED6gyaOijoh7MYmUA8BFeZBQNH9q
aONBAiSfSg13OVyad9L7uCoXL2UbimyyQRJyI8tYsm2Y9bX/DFwsbV0wT4TkxUUB
I9nUcOLMu3qQG/Mo4hbrYQ==
`protect END_PROTECTED