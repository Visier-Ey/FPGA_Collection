��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���d�v����0�i�=\��A��?��� (��1_B�f�	�Ѻ+|n��y��Q4�]�aY�����*2�y%����>��������K������ �
�D��z�z��C�y�B����
_�U��hkF<�~x�ܕ�c�g`�vQ��0!mC _�e�� �ý�j�
(��6��N�����V��iv�y��a�2@����<�}*dw�4:Fd443���f�[����*��g�!�`f�ޚyP�/5L�6T]��4�*uj1�PS�U�n�T�m{_��Q�#�M6�6a�H^}`_�&�?�_�m°�P��9s�wܲ���DcJZhh9��[���+xF��$�x�63s�I4~��W�%�2f�E���Iq+���J0�a�K�^��
r2���{x�{��h��+�����%�^o�?h��F�O�����N�*̆�6����Isz�m�HC���)ά,�\ ;,��2�!�#5R	�YҒ4	|�f�7��ٽ�[t9~mDB�_�9+1�a�!N؅z[ŝ�Nut�d�P/�p���e���t�0������j{ݣ���S.�^f���0Ms�-�bx��C��z��=�F���~��š�y���XxBc�X;�%���_h^��+��`.T���^;x�U%ev�¸��'��=ݜ%���� f,�XS�5��w1��ӣ�O�MML�欧�רk惕��>We��/Nvf_���P� � ��\%:�v?�ɣ��$M��=:iK������M��K {E�UXvmt�j���`"�BuH/V�:ᨑO.H
4"�)ת�֙`����0��&j���ϣ��*"���K�`K�@+�=��.�E��N��J����%�#�����f�=������ϵy��e��Ψe%L�ֺg�3T�J�)��R���b��> =~�	�1s�kE�b�T1~�ڃ�{s^P,�A�Nǵ�2~w~-Y����q6�O�: &���3����*�Z�y#�����
�j�澂��'1�SV��:��(���d"���F�;�2V^a�;�*t)��+g--�9���Lwt�3�4I�"��q|���x�p Eݱ� 2սc�0j{cƄ}6�$$Ą	������i^t0_�<��R�ihsքdr���@�F(&F�$��tj,�!*jӏ��<o8�Wi? �bl"���4�$ܡ�����N�k�:[0�	G
��Y�"IѾ�1��d}��.b��<K�W{��nB��pޜ��ˆZA���.{sN'۴H0Θ��}�5� m��Q��F�_U�	����:�s�֦��(vs���K6C#�	���GV�2Ȅ,}����ǙMj���N
3���&Hq|��<�|�L0�&%G;#B7tX�en�����̆���W�&l�&��2t��~�^�x��¯��R���\eLoV�q��n{�<J����ef�9X�lK�N�bďǯ��5Ϡ1A�y��w*��3~�#Җ�.�M��
��QuJ'Ϧ����޸{���'vƈM���F���L�T�גv
b�o�[�M<\�� �+�����C̖�����/�ͥô�u�e����1i�'��$���ñ��I2�_846��0�ۢ�����v���U�T�Q��LzU&C����]�Շl��d#З�x#]=S�y���.���,"J�l[���f��ƵQ)��"Xzh#�c�Zݤ������M���K:��a2Z� ������B'�}v!l;��N�_\X�Q84f4Ehh�|ow+=�����^ �s�#si��f;�^�KӚi,iR��u�w0�p�N=_
g�a���I��q�"]��?ND,|��ַq�N���2a[��v7��M��,O�e�6S��z�9@�e;+\�d!�S�mO�fL�"�i�+���˂<���EYE�F8��<#��'�o}�&�.���Qj�!^%��%�B���.�88�̬Z
>\��iiߙ_r\��%�����/�)+F��"G(���5D�����O{"3� If�\���j�Z\!�s)L��P��?�;���u����dr�1����v^~�VW5ʟ۰��4z�n�hh�;��~\$V.X�Y�P��i���>;1�Qn9�[�2\�?z�W� 7�M���֝L�Dmrq�V����CMk~�����H|��/^�h�������O�L��P_�lA�;XM�.8!i�mYb�C"�Z.SK���S
7S@��M�6k2q��s}g/�?C=r⤧��J �]�h~p���)��ZWq#NKG��K���`AP\_k4CL�pY�Lq/��ꉭvnٮN*o��ʹ�4r�a*����M����M�R=.Qx\�tZ�Օ���f]O�c���fD9� �y1�!�?]�x����ߙ��؍eb�58n�����t˚0���~����'�f�i�7�.���
ܳ�"��P�7���s�[vZOW�l9��!���q>	�S����e`�����N�����3�7�~����Q_@yi�n�p�;SW�E�?��T'��������jc>�	F��W�Y��(	�4!1�*�)[�h�㜰:�rլ��<�������ng�������'�`g�K�&�@^6����.G��(��S p>�u�o?�c ��*��t0����H�3մ�:�	�%�
>�HP� ���;w�f$�Ê���d�R�&��:����)d��<qKs�dl#5k���t́����q�^4V���'��S�������)6:�3E�U�RS��J-u��l��^Wc�7���哦��0xR��2ݜ �~B���(��ONވכo�����m
�^�G�u���摱��	��6z6V�z�o/BZ���B��=C�F���[����##q:Y�;d���/L�������	�59!�������}�&�5��y~� |��4
�2n�Lކ���V�^�l� Oi�8�x�N�^�&^�&9<٢�d�w%?�F���j��+X��\�L�k��7�����0o������6O�G	������\H}��Uᢪ��� Nm������S��r��������k�6�bF�H˷��Ǹ�i���)�Y� �����d�O�8-�% <���"A���n6�L��
�dX}%���=thw9��E#y;���Ӭ�XJ���Ve��\u�s��j,w�2Tb���b��R��v{�,R�w� �T8 �Ҭ'�_;}%�\X��w�,�{U)P�%'tBP��9C;�O�|4�>^Ta�OX����Ê�c_���l�PB����E�ؓ6gw����.;S��D����ݍQ�{�Ϩ�� e@�l�w�6ʥKX�����$�&|��	���\2���#D� �wa�;T<u"��IM��x��m�2�'�/����b#�mp�ͫ'"�^���vd����)�{���GS�aOD'�/bߖ.j�֧���r-!�.��cv ��nJc�i�vRxy��kڒ̏Xcx�J�.�_̯Wl���%+D��^K& �D�55�"��.��"�o�'Z�޸�Gbs�"4߆���--��ʠ"�W�2����{gg]Ϋ���Ih�������]�������l+�}���.�mk��.Z�A�ٺ�W1�\)sk��gG0Bm���=ǫ��SZ�K��锶��sh��?d-R9�=mg��GP������;��ŏ�e����[����(_O'P^�U�;�L���'���p�ѵ6��5qdD����ь0��s P.̠*���Y�\��~��oyF�fk�#��T-}�%�pu�v��O�������.�=������io�`�0[|1h*�t����	l�WBm��歕�С1�R@�W�Ĺ���|��h]�M��+U���b�?�@u8�)�~g�|��F����}|X��@��P-4���Bz'��1ݼ���{ �q`���>wZ6W��^�l���5���G{��Di(זh�t�����K���#pC0V?5`X��o�c3�?�:B�ǵ�(>I����Rv�]�~դ��܍m8���Xe�H�L��� �R�~����0a���gF�q��%1o��(K+����Ԯ���g�N���"b��t<�5����̌�B}�D����%G�ًa��'�'@�0	���_3b��~o�����!��c�E_: �Ib�K��K���)�����͎��=���։�
��	n�&	zVž��̲)Н	�����k�r��ej���	R�t��Y}r]�LE}׉}�5���S9�.4����KЍYw"�>��M�l2�,
s�zQp_ox��;7H=纊c'�}� ͯ�W���"��L�%�����Q�G��M-3���P��|�>ou/��*�@.����|�HG�z6G�~�:殱&�ʌ������z��`j�"�2��+��ٺ�$���3=/�|�f44�[9�LcU��cA����#��0A�<C�z ߺyKxb�ix�A�<S��Z�r��'��`	)=2L��,�fƳ����9qv�>�������oQ�YT�����:���������.�w�͗�n�+ �7ڜ���2��a�U�E��a�N5�����K#�'Hd�4i�t�/l^|��+�NP- P�؆h~<�5u�y1���(�Ǜ͡��Ls��T��Kp}Z�LQ�-��:�	c=��p�}�F	�FQ���Y1B�:�qO}Yj��k�g$8q�ϴ"�J6����Џ_iܘ}�ճ�Ch��i8�ar炠Α�_����]݆�r����Xפ����./Yt���K��ͽze���d�n���1�ȝ\�g^7rY���l�hE�6�;�6��5� P���R��+&T6���U��.q�HLR��ec2)�8��.��UR��0�D�z�;�]hm�lPr��4k��.��@_"�b17h�,(|G���|�����=�{�Y�
$�"�p_ѩeJ��}�5~�MT�Nġ ;n!'�zΠ�t|�#���O3fc6���A�(5�\�8/!1��R\���zb�5�J��������
�~�[��+���2e�ܔ�^h���������L�5�-�� �_v��3p���o.����:}�}�]�>��:�˳����矀�d�\f�pr�?W��Ⱥq��1�M��W��v\|�Vbm�VS��n�]݉�/���"Y��k#i"/M���)q�)�Gʱy���Ŭ�8�H���΃�-����5m�cx��q�u�,��߱�R���H�MW%���PT�Oa�:�H�Bws�-���z�*.E�=)��oN$�d�knO����#
!��nHp�8�͍��$�Y�+��Er\P�OлHrb�w�~F�D0��!-%�N!�F�`�N�tS"XNb��o�Ԉ�V�Q��	YN�AM��2k��JE��i W�\����q�cw$��B�̄��:��;�j�VW�F?GAO)��^(Rћ��
!D�#д"�.���|`�4:�x8��䞦!:!�Ga�e�xD�U�/���<9��4(&B�/eFyF��l�*I�����v��O43��V�u�j��;Q�.0�� �g�fehSz�38Wp(�S�2ݔ�@�s��h�u��SɗL�}���ZρF;��wa��1���^}�@������9��R#��A��|�=x�c+L~i>��x�˿�a
UM���^��W���=���f��L�Ea��9я��ĩw���[5��+�ʳ���#Y+��p��Y�" �&�"���5��I�����D��}q���/tb��fWoSzXx�ő���T@H�Y��Ju>@����x�@��P�$����� ΛF��L�аv�4k� '2��ځΜd$;fHHx~*����q�3Ȗ�v�M�J�o!W|Jpb�P�N���y�8~��S��ޥ�Dd�x��Nr��e�?���}�fY\V���?`�^���`cb�4j�(x\'ϔ�5̰x]f�*��!K)�K;��ϔ��/o��	����ɣ���(yJ�Xm�9��M�w�#R��9Ư��0&�#1�`M׬�͇ �Y_��#NR��_��qf��b��|��?q������F��2���AO��Vɣ��y���6��I�/�%A8d�9&�&%����asC��q�~3ʂ_�#@f��3d�.n�ս�(!
��y�6�Q��h%^��D\�zH��6�հ��m
������P:&��&��V��L�����xt��?���E:��ޛ=;����`�������i�_��r�3�����R	�A{�����u��4G���X��˖E������)�ï����Zd�
�q4I5S/�X(�0]�����t~ϵ�e����b�Qh������Z�v�!��	�9�~D�m8���$1hs������"e��^�'Hr�+��]�G�3;A,����S�r�����{����>˦Y����֗.���}�g�ʣ8�6l���v����r,^�~jԨ�@�6P `�H}�[������ �Q��p\��Q�f��<�<�a�CGx3�=����]� �Oˎ��M�]#
�48�O��7/'���9�w�*^M������?m�Q���s�+8��Zɲ��6��:��#��(��x�r��R&5����୿���\�t�_��q����ݐ���+/��5VէI+x�|�[�����V��6�L��_���i�5[����ž��!������c�qZ8H�P�%tTN����n�0�� ��̉�� �Ug\�`e�v�0�?�d���X�6p�+H�^�����5��E5tnSW(��wCF�Tw
ٲ����e�h�Sp���G@E��v�W<��Y�6�L�F�4�<�:��� �Q�����\z�"-���D� ������\Bq����|�3�:9 =�2ef�S�Z^d[Oϒ���mktr/�{�z愉�?���@��u��,�0;����� R"�f�c�R�H��(���_���N�O�M�<�ܧ��r��y�"�H*��|X</ɨS>zH���Jd�v��ux>d[܀��
%a;z�*'p
h�3���;�IS��
��F_Kz�c�L�wI��&I�,�pQ�L��-c�4�q��bV�M�H��JXG����h���yQ:�%���L�5+��v����0�=3���9r-�1&JN��CK� KѸ&_����P�ҡ�vm�J؍SavwI����Z��Y\��! ���=�+��;�MJ�M$�?�A����5��4�6�4����3�<l�P&����v���
gw���4#]BZ{NmM��Ӌ��X<����{32��;G.?�ݱ��_u�<j�s@k&\��g���1	`๐����2��M �Y�5i&ԫ9`{9��i���"��n�i��Ӡ�r��:��B>�w�������d�R<Q�L��}���&`f��q����)�(���aH {�?��at'�rS��!9d�6��:"�T�?�T��!���G�o�L��.#�H�/��Oݰ�84�\'u�N�0��&��=���׉�~�W�	K7�@�ߓ��������Ou�!x�ɂ��d��
���Z�X�9
�3>^�d'�vY}�cxg�pUԂ��jg�n�D~�״���XcQKR�^ͷ���E����w=6�ekd�̣��@{+Ǵc�q��W2��*�w��#s��h��a�f���=	o�H"Ld.�
�H}[%ÛK_�T
h��j�H�k@��0�/*������K�իN�󞺄���N�7���յ��u���j�d�ə���Y���47�(�f�π�ц/��B�.{,TM ��x�.�Q�<���^��� #WI9�זtϡ:T�,��!9B;Mc�{K��5W'�QU��B�n(��m�׫�k+�T��>"4����xys�-U���0su�9$Ιrܳ@�tI35
��[b�دm�9M)��|�'�M�g�mPA���dޒ�Q�7?Z`\��Sf���&ۭt0��[���:�K��#;*C`9�&��È�M�1�T^�6k�
[1�5�V��|�Db_��]�O"�k�	�w�J�&X%P,��9M�+X�	|�v��A��.��n����i��p1���Y�U-�Ӣ�1�i�m�u� ,��Rn�(n]��W��y����m[X��v�y����Ǹ֠�� r�T.e�?	'�h�γ ��Oȶ%��#�cP�Z��x��1D��ЇY$����R*p����4��]��=�Xcv��"�L�uB�y͚
�enЃy���_��_�F�vY-��U�0d1�pg�f� ���
s�j>&c���^��JB� �B�"T�(W#&i����Z/i�$�ˏ��.���ā��2�����-tC��L�xn���v%5�xKԤ���Ea�d�/@�2J�Y���2�=i�i��'�&xz����=ʋq�'eG����l���&,��!�
3�3�y?I���Y"�WB>a�
AWǱ��W��4��/m�����>\k,QP���גb��ےo䔖�o2O��p4�\����e�z���'~ ��1\ќ����;�
|����F]����0Q`�^�w�7ҮA;�nXp�Ԝ��h���,��JU�}�T�Ar�rKj�*��띲�6�����$�UU)���7���Q�R��n��m��CmAӻ�l��H{���=n%�[H���O	����E���q��U� �D��1Q.DY��h=�8BY)�72���	�C�2�Q�@B̗&|/s��@������Vr���'��Fk4�b��B�l��a.��Ө���"�mܬ��Q0uK��N�w�Q���c�bѼ&X�MD�yAg�ѱ^!g:�W�H�(�C�-��)��LJ���p�W���}���Ga�����4c8fa�Xb@�o���#�5���])�L�%Z͗J_��G*���IvZmc��!�ޗ�-���,�qq������lx����'�?���S����[oa��Q�!��6'�"�b�,�Aqݪ�>�S�����2Ғ�	#Q�0aݲ�GinZ#ώ,��1�Œī��[ka��v.墒�n@rse�d�����[l��� Mp}�ɘT���bitSxwX��'
ݲ<sSAм6,Dľ�Y'<Kԋ��tZ�|�4��3$��/?��1:���B+o�����U�grɷ�������Μ��T�Y���J�7��pxIc��§��܀�4T��\ �D��1����b_�X.M��~��ח��1<.�_P>@ߕ�1Z:kZ���x�m�o�ַ-�Ͳ4m�!�ߩ��}a\؝.:���@�r�Im�Z�y��g��CJz�]���F�F������mR�[8��BF�Ԇ{2��u��b�~�Q�]���\u1dՏ�V��TU%��o �$�L�+r�Ȥ+D�"ʔ������Qv�}߭����87ݯ�ml�5�O�9qo�U��g��u�(�cڗ��=m�����],�<6����R����:���r7w��e�s=�/�*L[�t�.aTm<��V�-	��qh�q�¢10D��(!M�B�������h
�`��S
�:����/����X�"y2���1<l����D���g�:�j���N=P��6ql�s�q�9.|<P��̴oI��`�N�vN�m*�V"�����Ԥ��gw.d�^�|4����W��)��P�Oؚ&���þ�P)HL��J�7��wOe�+3��>�_�c)�)�"��%��b�����\�I���o��S���\�&527]z%c/= �q�g�=��7B��,Bt��}qK�m����A�.�}��s��WPz��$�R �t��m���j��րb�D��x4Y];����g��`������ ��pP���+L�7��kɰ�5�~l����5�1rĠ�������D�W�h�Γ�Fm�^X�\_�sR	�G�D�P?�4���Le��ܭ|��D�
�x�)Ҟ�������Oϯ����^�%�f����Gs	��tE�(N$O�ewÛp�ܠ�x��YҾ�1�_��p��.i$�K"�=�l2��d���,z �g��t�t\�i/���3���B�����
q�i�ډI4�7��X�/eܙ�λo�?��\?$A��Y}D�¬VeL���V��??e�+�y8�k�ۻ�#��c��H�|�U�<K� �#�T] �њ~Z��J�mMA������Q��.��)�(��[�lD�\+x����R^��V]]��,����ٗ�,�|���L�.k�(��$��"�o��S:��	ȝ����S^eW�l �j����-sۻ��T�� |���Z��U�#T���l����y(�7~PF�C-|�I����
1�Ay�<�$� KǨ�Yy~��'Y��^/�Q���Nұ��wZ����Z�b��D4���K,�(��/�@�������� ��ݜK��.�V��2,�c� ��R���M7��6���?�_͍%-�p�9O�,��T8$� c��gJ�'�dxv9
"j��4�3E ��ߍ��J4Y��S��I��9_P�Zޣ��Je��������!>��^B���ŋ��a??]�}ٛ��,�����pM�}���MP7	�Y�f04��}�v����<k��0t�Q��s�z�yI��K %�B���z�읇��`b�3b�}��!3�0@aLt�>�y�2���xqұ5W��3@F���]�����;}b����eX�k�J y�$�����d�(|��%�� ;���c_�ʺM$�ȼ�VO�y��J��t{
�J2�Xr���,�%L`S4s糾�ez".y�P��E��`�q5�ʋ�gx�L�����7��s�}��'t����oS$�w^�hw�]��:!=�����Gi�p+r�N^D�g��Mm�Ӝ_sJ��9ΡVza�����\�� 7������q5�UZ�Yy�[0ɍӺ7��ϔ��3�ď��J��<��b��V����|��Ϻ'�&=��GlJx<Ċ�P�< wW|m�I�j�G�%�"�����*Sg�"�T���'z�0�.�J�����],�O��Q�Q��n�:�<�UT���cC�N��Q`��O06+\��Ie�7.T$��{B�N��7nHn �=�v�]����$���~YP��[�;��^N�.2&�P���3�,}�~^�?�k�d�TdCsu�j�4�����$W�{do0]�(���i#\���CڜFc�VV�$����\E�<,�D��^ݥ�5D���r��G��c��O�<�5��GPW2�}�HU�ݫe0�3ܕ�RR=�h<������د�x�#����&@���lޒ�b��C��]j
����"�=	L�R�<�OB�w
*dH����hCk^ ���v(G��@��ѻE��T��K8�� N���������x{���촌�ꏉD_o���<���_UӇ���3I�Ƀo��X������o�=HR��^6a�?:���e�
D�<,G|��~�^tj$�
��_̺�@�	!����Qrӵ�N�ˣ�>Dr��
Kn����Z#Ý�웿��%�)��I����5NW��KQ�{�~x)ٗB�挒cP�[$k(K��0���
�%h�4եm =�]�>����!QQ���n���k�s�V�'�VQ��\y����!q���R~�^�⒚�?M�ʈ��tQ�e��u�sl���y�̈'��C�Q�`sU^&�jp;g@��<bb8��DO����7����j�#�2f{�߸q��k��A��-X��i�j}����EU�#c��.-?\��N7���j$@��MG> �-��}�$�E�w���.�y��E=΀+K��Y^ .�����b�k��Wsz����Z'r��>�݌b2=N�K��t
`��V��8��	"�H�*T��@\,{,ISq�ε�bq�N ,w���D
\8֒�=t�"Z�"�<����tP�	�� ����H��?�\0��_�@��n=�e�T�������|�~O.�X�}��h�^ P,} ;di�B�3'>��-aۻP#��N��4�KC�$�eV���Xv��zM�$-��ɶj���G���O:��8�>T4um(�̍R�:U�j")!`�����a0��Ĕ)���Ո�1�R�s�n��� 82u�7�w�<K�ބ�VIx!x.,XsI�߹�rI_�����`�姃��|a�^�E�Η%$�N����'�4�C�!�u����a���S1n��/��9�_z/wR�
�M�=���S#�Op!���T�nw��dXf�w���bdn7��;�D��G����{q������O�3�k}V��.~�S��n�f��Jh�kς�x%SII�>jmɠ�jt�U��M�B���}'xG`�	-wx�y�?:���0��_�Eq��ʗ`����g�e�7
��!�N�廔/lJ�R×����,mK\��w�@jw/ʯ&�P���2||ĩ��U3�m�^�N
p��� q?&m�U�#vQ.SCӢ��y'NL��5A�,.��5a{r\�0O��y����`	�������_��_*��_�=�(���ً�
�G$��q�YM�X�tA��X�{�/�䋈��0��΃��9|�\!��|D�D��5��#P��:�֐SL�6�[��8g��%H��sX�($e��1�4p�i���x���Rjg��k(e�)PH�f����ͥ����H`��zS�^�x��ң�n����>
�||�z"I�+B(j?���ԭ#z�-5\�&qoX����ּ@��A��C�02Y��Z�뉃ߊ#)�KX��)F�e
����+6����e��e1Ć��PR��4�MN{�,W~dԿ���'����=�F��=b�+���s��-�Y����%��l�P��u�ejh0?�Б�$z�M��s�%X?���L[q�Jۭq׍6��'+8n���3�;��[�!m���K)J�FlTX������6�m��i�?㧷aBi��~l�&ˣHΩƇ�[w��G޷^�j��S�pf�����͑�͞�by!�����=��S%��Nj%��Յ�(�:�$0�T)����F��|��Ս�$�����Q9+�
F��O力�Y�mXT&��u���`�����E�2R�BT���*79�6�zζ �Z5Cztc��|7�zQ���#D�Q�)�X����u#}���D�G���upˈ2Ap�%\V�g+�D�f��V*"Ԫ[z.�֤TKy���zMѸ�k@>�4�F�C��؋�1�W��0�:ծk���������O筄!��>��^����J�P�/D�/����8L�1Ģm�7�#�������XU#m��r���0��R�x�a�TR����� �E�1�JM!�XW�`✧ڿ NP��.�I4_*�J)my@��WF�.� �T��L�dv�S�b9v2o*�*JlH�"�Z�k�^�����CN�U�V]�;Mr��U������((�+���$�_�j%h���/��h��(9�W�+�a#Z����-�S���#��b~�k;�o��Y>�7�6_�W��%��ã��B߄�+�HA�z(�E���۾	��6��!dFJ��@vx(a�;b<�T�m+�*ϛ�"�D����P�u���%<����S2�s�>��ɑ��-���H�ܳ�|1���|5�׋N�;�1]�g����K�� Z�SG�b;y��АV)~j�t�a�A�l�%��/��Z��m��B�D��=��]�1xtr$�B�֌��~��Ô�wI:��`D~Vq��8=��q��#OL��K1*��2�0�av� �~��t���6�Ӣ��:��>H�|�{wDc�O#��l�]���=U�T��Ä���m�t��6�;�H&�����V̖Iyּ�
v�"��J�N	ؒt i��ڀ�&����+�?�n��l��P�*�;���J�Nq��.�'��EZ���i{�Α���[�'^����
e�hء���GiӊO0�n�Ys3M{VS���sJQ
��l5����F���k���E��$-#�ׯߎ������W�b��!�36S�	����]ɑϙ��R?�ʫ9�f ��������=8�>6B�������OF���__�~|��Q�t�kо�QO�\qIT��C����K[�Ar:�TB�^�/8�_����_$z���"�ٸ+t���\�=#e�tIz9�SZ�y�&���<���:���&�(�xd��q!�<���CU�q㾺�M�p�%�n����RB�c?�k��0�= -	�~q�b;�g,�
Y@cV��dw�p�կy]h����=C͡�s�9��SQ�-?�p�7	[ŷ����=}�o�����ͬ��X�Vb\3�G���Ku�����M�ݻ'/�}K�?`�,O"�R�*�s6��8��l1�#k�yϕT��1��@R��Y���)0#�ݶ����	��#�H�i���J��[����v�o��֮�s
���q�VK��q�X6��J�>Y�\	���?k+u{ځ5����s��Aw :63Cx0	�o��dh��a���SLX�8��u�%Us�v�9����E���R͇ry�\8 �#<'��*	-�9���%��:�C��@�B�E`��5��E�ѿiܚ ���{�։p��m��{$�4;>˖0?:J���G��.����F�F��i;��	��샆���z�$?�9�N�7�7��ҪL/�0�`��/�<� `��z� �}�Y�GZ�#+�G��^��d�G~�e��q���	kmg��R���C-ƞ(y�4��a|^D �	]�"����?�{H�S������.�7����XG��)?�v�1-8��Z�	G����[y�ц)X��Nm�a��7bq� ���A$����.4�Q���/5�G[HE�=��&�q��u��p��ɂ�IV��5ÑSh�]��活�fY����0�W�x;%�k�S&��R���|R}^JWg���~/�W���2�8La7͛
'�!Ӵk�ѯ�[9i����,����7���US�'x'i�U�Ȕ�?m���WQ�{ �pk=Af,��,ЪQ&�Z�h���>�X�d)�[��1t�2��T�?�k��$yw�ط�F��*����$`���U���w�[��6�F��܅]K����N���[	/;p��G��|g;��556]{Q���
區�q�Ŗ�q+�&��^n,O0A|k] �����w�@��H�|M�S�d�b�✜��3�U�hU 3��"�8�!f��U*}[+qٻ�x"�~o%F���U=tQD�+�Fh�a�kp>���BzDTFc_�$B%WX���2��x?�Мs)װ�$C*�[!_��j,ڣ�tXV*��T;R1A���g[Ƀxv�߷���>7�ǅnp�U�x�5��Ӕz.
,���p�g%��6h�K�{3����`�(ͼ���ډK� 5z�;��j&�9c �꒎&��	
�$�>��!p,���4��_��{�����/VnL��ݭ�1���pʎ��*s0V	�|�gWƼ�������QLT���%fŻJ�պ�_���_��F��}2���.+�׿�"ڰo����o��$����-+�$P>��c�1�wL��h���:��3	�,2tŴ�m<�M) �[��`t�5�L>=2��ۡ�秛~uQ�A��%wDX�w��V�8R}&l��_�ޢ�<�� {�\�W�T�־ݫ�Q��o+j�l�����6.�&+E�<ȑ��vQǍxW[#�}[�SȨ$�P8e��������5�n5G�'�k�:�N�7�QA+ �Aw��D��x(
�����M���­
4�+�x��Z�+�a6i��~�",�r|$F�M���ZN�K�~�-jci����E.�V3�$.9�[�rS-0?��?ؼ\6,��\ى;b�)������� җ����D�Hqt���;ݛD�&��(�J2Yr���8��n�OW�,{;�kw�A_p<�&p{^�7�>�J��x��Tz��e2�l)�dv��Nk��䮙��2:OD.h����/сk�jr�D�s�댁���٠y��J$��IH˫��\��%��CƝ�/~j�ca�/3
C��Q��ɱ�!�K�:,7�G���`���<�,0��3��Л��I�����}�'μw��az)ԉS�2����
��nt�w�Oy}�q���������Ղ0��~���r��q�/����s_3}z�ŞA�����GC���v�����v�,y��9c(�59�?�Q��Uk�y�4J5u.�6��zdF,����)��t������k��	�	��$��m?���������u���*`�0rТMF]I\\1o��3jZ{����4á�{�,`B�y�����U#����^ �l(s��>�Rڙe�R�F +�.���w����d�8�S�0��q;޳��۟ʡ���?��#��v��$�u�+X�[�vE^�P2��;L�(j{KN�0��[�ܢ�e��r7}YS������B����)�:L��$"6u"�=���9��bv�]���S�x�aR-�/���a!���cD3���d��ʜ���(�;`	�[�m���6 K�`V7E0��zW����>�<����=D��RX�O����\�������I!��/���h�0���'�0G$+�T �5�	@K�W�ے�(�V�㐧��6%ߞE��%]	��ꕶwԔ��)�C��`��f��öM����E6���k{,5/�4=Y�d����_.������\�!rU�iZ�FJ������bN�{���}��f���[Փؐ�Fu\Kб�9�PJ|p5���Kf�n`���3�З��p������>�'�Ҳ俣��	z�m����D{�1��0�K��K��`@0� e����]q��79�L'̠�%�.7��=�$z!�QӁ��Y��3��%�� �M��4n2'�|�j��i��?�R������Y��s��f, ~�@��p��.pQra>�����m�@��(m�����I?�Pl���՟��o���Ɛ�'��m<- �;s�Ku5�~;5��f�2���u�i���C�
�'{��,�;߬m��s���I���؜II��V��^�Ye�E��ݻ��>Me�
%]��Gn3�V��9�o�ctz��z�݋P��3���o^O�L��U^ -����>D�^�q*������@�(�O��Q.�5Peb����um*
�Q����Ʊ�Yl1�@����VRa͓h�w��� �snLP'��� ����� �~9ʘF����vїn��һ[�r���ʄ�0bWB�z2ɐ��ޤ��z_��68T(��06�.*�|�H�-k
��&����"0hfY2�Bd�^_�vQ13�b��{�L��^�%4�*4��ʔ-�0�ʼ�m�<�#/+�u�� �gv�K��:a�^������ᓟ@���'��r�[��ќ7�o�U�#���[O|�;x��-���
�&8�wӔ�!}�w=���ⷓ�8����c0��!5�S�R�{e(�����8�A�Z`��$IhqGϗ*���{��!�)��o^�cA��]��}6���6�|BN�*��wQ�%Y�} (�h��{�YbJ�>�_l#j[Q��JO�	z�0�O�R	��J&LUX�F��a: a��7ur���<�K��!�3v8�l�}o���+Zx懕��r|�hE	���M�W<h�����r)>�
*�}f1(H��Ƕp2�`ba�^��|��rLL{`�o?UE0mq�����Ix������¥sN�D����f����B+_O�������o_�3�D���NQ�WJ�rށ��Wݶ��e��~��_,���'b�Ux��
���SՓ-�NھY�u	+�nN�!:kx<	�X�)v!�"���0�	SV�%
F�)G���pHJ��u��wd&���W�\�Q�2��ɤ�Dͭ��v���;2W�v��2r��ֱQ�^�� +E��3@E#,B�[l�+i-�q,����b����5����Ҝ�p��(Y��6a	(��ڡ�@�	��		]g���V��=���(L1���k�sr�Z�{'M�5��|)`$�m��R-`d)��H�N.5ݟ�r�$V1A�	���!b�
�z���,vȷ9q]֙`�A�@���.��8|�}dD�`�M�b���{�������5p �j��j*g��L��-Z�M�Z��:3�Dx^�6JE4���SgJ ���`��.-�浖�`���C�IP����6���=�F�Gn3�녥鍦�4Nnk+�1�����e�6�?/*W�v�����m�"%�dȎ�@C0K;�] ~{�7}B"����1��:���e�����v�iG�� ז�P��(�O���jɻ �8G�_���o�;!�_���V���Q��^��[����	�Y��#��)�o�WSq_y
�@�HÐ�6�:��-"=^S��&�h���NOrwqh�&��AJ,%6�d;���,�`t��f3�e���g;(�V4�'c���~����ⴥ�+!ڿvcI(��*~zI��.�u߮�ź�d�Ϙ��|�46-O�kq�>7Ab$�(-��Md��#�;0Sb�C��d��|�+Ro��<�߄J�B@j��AWNH9VtA�MD:uR����y"�n�
��'bn��L��,���
8�]��C�}Ɖ�u�*��<o�2$ߐll�2��?%sj^@�����<��i^a�h��(�����1I�<[@ڀXacC��@>�Ea����*�B�ܣi�q��~d0�P)NPa`l��6����y	�?�ܚ�eq�ڸ��j���ɽ�V]����m��5&@�};��"	�:Ab��MƇ	k	�E��i"*�d>U�kZ*��t6v�	LDm2nG�d�KϑkSɗY����vr<��2�H�ֆ���7�{P<�th��t~�wG��/���c�`� ��x����`M϶��I��]q��Go� 8�$
�0�ɬTH��AUqb�뽲����X��@���"�"�4�[���A�d[����It1?��X�T�?X	$0c&��J\PM�Բ7��T,���:΀lV�����F(^C�y_�fߏ �L�3�H��Ϫ�fu�Z�q��?�&K�%���:��XG���0l����Q�}��\�{y���i����7�B���w�Z�erVc�_�<����:��"��S?\��;=� �PFח��h�C,������(��j�˚��)Y�@���Ym���u�rw��
�FΕˏ��������
���%%���3�o��A��Ht�#b/h���BT�%���)�h�R�Y��}���eU�]D�QI�BZx4Y��J�`�ӯ�$w�_��ؚT����'����_��%�3�R���W2◺��;��k��$�ۢ�uzڴ�A�e�@q� ���a��aEZ����������eX�G�����c$l{��-��T]�%כ?yPW����@���eO�m�	��	���*G��Ά�aG�i��c+��Qr�u��vҝ���v5�����=�YۄE�PZ�H�%ʌ*�~qT�������MT�:.�[(��H�^#B���>��D���{yX�j� TN�k]���=k�b&\
�0i Y�E���b?;�|Up��'�TDh�v��FXc�����FⲶ�J|���J?*Տa����;8ZL`��dE��$����>�~h:ցvCK*���)���o�֟�i�����c6�NNdbd�ټ�Gp�Y'u��)W�4���X����Ff,j�$ɚ�v��T�<(�V�|��%��k:�M�]w�B���[���
q*� &��P��{�Uue��=�`��]�$��h�7��iز�/�'�I��n�Z���N��J��,)\��4�Jb�U�F��CAal��b�R��є0v�s�j��W�� I�L8�
�h���m6�v��A>w��'ꊐ���p�{7��$�]��#�c�l��#�XޯH�E%J���}o��b�Png�_E�
r?n��YaD��{)�Ȗ�א�`0��i�Tĥ��	�S�Qu�З�F��f-��U�ʀZI�g�([OHS[����yC��M彛���U��`�J��~;��9- ֛A�$���k/�D+�3���=����L���gVΣr�+�7���7��4�G�nO� �H�vER���9zt��o oFiT�=㺊����y��Ƃ�k����d�6^�A����c�7y(���w��u��uo���i^T�3����}$�$Q�"�Į,��f,դ�� ��D«Jy,�%ݯȓ��~�N�X��j����B&��������/�RS"�l���Aj_$@�Y�V�)k�j�<Sx�w?�P{�QO:����.�LC�d��e�w4Y0z%NX��#��G����������?v�H��/�X�k��I�+o���jbx���a�K�7�
k�g�J��]ՉJb7���V��Iޘ�
�|�E���%e�[���'(��G�Ն�oBo���~���7F?�LV'�$<���D�* �G���ā �*���4\�L����X�L5�B��>w)twb���p����1Mh5$��I��%���rqа7c��+
 o|�A�U�f�I�j��:+�ʺ�f�_�4�/�2}��w�H���c�Pѭ�s����x��z��.��M�M�O�'��|.w�[֤^.9m����.]�"���EӣIE�L| �'�	y�������h6K�zc ����L�c~�/\�V	��ms=:͋"�͵��
J�Gq��q�!y�8:4mS�Q\�&���l�����R�Ɲ�e�R�F�擉g�\I�ǳN����e`�]�����$F�5'��;Xm��5�J�Wk�"�K���$����/�o��a���7{�jIǺ���,$HHI:)�z�f�MUm�م�?�+��)E���<��}C6�/4 h����i���a�.}�U��8�z�.Vk5�0����	���V���a�d�j�؞��;t������8PT?�P������Y��Z�ي�K��#6߯W�ͳYv�Y
T�}���=�=-x�yǶ'���%9���$k;��a��H�C����㼝 �6�O9 �٩d���:��N�7����DN���ZτT�����\ ����n�U�D�&�8���]�Yݫ�ַ9��G����m%�?��\��\ c�x�,���O����������۔�i�%Q��|��d�T�^[����eY���o��Ș�ф2�����z1!��k�_*�
`��3�/��3x�9�?Pavw;]`[�-YN\��x�X�&���� �R�vLdu�p�n���$�F�8�3�L³���=&0����XĴE� ѧ��o����n�Dl������:ݩ����	ӎ^��>�8*E�s;�O�����S�ԫ̶ɨ7�y�3QȘ>��]���%��(���?Y o��<�Cɫx�|$���HE(t����T$�A��c[��$��p�Ӟ�bbӉ}�;"����De L#�&��5�E١)��O]Tԉ(*�g�j-�ע%��5�hB����=��v|����	3$���kߢ�_��Q�Z�l�a`�y��nG���_�[�P���*�N��ʂ&�a|��%��6�op��W����� ��kR��n٤=�<J'�!4�ny��@W�h�#�E�Ff{��B����Nu�sGskn�s��"�&^R	J8��O0�!�TiU�s�rU2����׃d�f���Ӏ�W6�&L(b��N[������}N@@W�n�*B�u`�y��L�|�тV���lX��`Bf&�Dz�j�l�:���6dԮ�u�cϴ�
�j�W6�L�u�#Sj�M��Z�I%I��mx��_�j$\'��ogmV��S�=)h��n΁pc�=�����=�y	U��z����M����? el�>mj"�q��&Kn��m;�^r�4���{��i2��W�� ~�>�k�ҹ(kE������6:0$��o��/]�8�|U�ʾ�f�Ԡ�ǖB)~���s`�#����¨�}�hs����+�d�0jCj�*cdC�^�����	���\ʠ�7V�d�> oA������S?H_K�L�2���<<�d�V�m����h<%~�7M��(��l�O��ڊy����=�Rm��n�WT�|Ȑk�Ӏ�'��N����@���^]G$U),?����G�����������"�ٔQ�Z&hR��[.�A27O�����!�n�X,����ه	��,�#����JX\��Ol���9O�"�B�b��"k���_e���P�����o� �W�}�T
��{'\޴�}"�Ե7{4ðM�6Iu����Px���qR�#��S�+6���r�z�-��y6�K��Z�A|m��p�����?���v�(��{�R`�k�ACT�C�j�`��9���$&aG���W�O\E2���=�#jA�c/L�ORh⳴������&���{�|H d���C$OHs��lt%�7K�����m�Z�`���aì���z����I�ܒ��f@��y|�{�9�h{��,z�����v D�=Ԃ�9~�\|��QD�s��I��p?�;��7�lơŉ�F
&�֞Zw��a<�6�,�I�����L[�F�u��-��w��uIl���Q!�&���P[�^W�����:�0��;��{�DǳI$(��������������l�?��d5�{�-6��y�]�L��Ê[V�!gY$��V�׶���Av�\ō���ՙz��8'Sl`!���Å�n��4�Q�3��9�_�4��n^ו���S����3S�������1ć��jA�A�('9r�?�E�42��lf���L���Г�ЖNz��m�Ӟ:�H�O�a݋k���3��%,��6��m��p0#+��F>���π�T,�.b�V��]��^'�f��_5����]%)��d�/2������|�`%eʸYt�����%6ְKl��{lΊ�s��� ��-s�����TY�̭"�1�6BQ=�v�R*��[��$$��f"��v~��$7U�����HHX���bA��RUK�^�&�\q <��6�3	!�e�	ں�n>z
ԔH�i�.3���kQ��@�ظD�-~�I�!$Oɻ�Bd��E��7ms�5)�w�t���1�������}�g�&��pc�$�I;����X�^�R�{��a`|A��Su3��u6z;�.	���!��t.�x��A<pC�)�)4�
g��7���R�#���E�U�9٠M4=k�-Q�~�Q&��¦��B���كN`�'F�\0����kT�^����s*�H��R�G�E]>Yª�N�9)l���x����rڨ�3�.1J����PˎZ�s�������8R]�m�CrP���܃��~���i:v�/�Q7��X�w�_�GF�f�Q�:��x�H�b��P<��o�R~IR�K̅�A^
�������7�i��H'щ�X�Txw��m���B����ύ�B��W=Q<�l1�]��������-�����`8�m������y�L���m�y�PzxE�� �_�����m7J[R�	v��쭄
r����K���X"/�v�� �䊒�{H��4��cRZI+���'J�gH�M�vzk>�bHI�b+�}�d�����UO����-x����}Mؑk���$\,�T�VT|�e��!Y�;z7��u�eQ7�#qZGl`����d��tK���P�*�,����%;-�)�D݉�+�?~�T���'�7Sr�[����FdE��^�F��h��,��<��>ˈv�0&xH�0���{�D�y�$��m�\+�<^<���h�:�հq��N�%�5�-��2'vsQ
~��M�K��~�'�J2-��Tj�v���R)$U�=�n��0�+8Y��T��� yҪlzo���b��UȲA�����{~i��t��e/�?5�l%�J�M��ٹ_n
�4�З (N���W0�aP��Ǜf\�[��t������{Fp���	/z��`��M{�%���������`ĥ��i�f>�2�66/ԖiI������E�ء��RK�͕�w�l��)�$��ʪ��9ά��������@��z��7x*5�^I�&����@��1d+���|�a_��;ߑ�u��U8$��YEK�lP����]p'��l��������]��ؤ�fa+ �i�\=�WM $�����N:�(�����d�2�|BB����U�;��l�'^�M���Q��9P�]�#����c ���޶����\�0��.�Uu����_�LR]o�>e�d��6��l���E�0�d�eno�/R�b���"�f4��`��3lT �#`�|�>��l�$ݨ>�,%���G�;+�⃃��C!�ʢ��=  5����Ӈ>+�o��B�����rˬ�fk��C���0up�Oy�o�i�L �����u�=W����a6n'J(��Q�)L�*.6b&R�52H�r�?� '��Ǧ��nF��9*ѳ��bH�,����l*��H)#׬ ��������d�:�z�!�_��wHC
�7*)mr��*ph�0-}����������dY�u���4��=�wy�#� d;�"/���:g�O�J�=���/�bC����Z���ٸ!���ZiX�O���e0���.�'!��d�Z���.�$Bm��|ѽ\�2I�-��%x�����^�׃+s����}M:�뿻N!�G�{9�aQڷŔE�U��2���R%��W^[�����j�)I�k�"~.����p����3� C����	=���WN�-�U�'	�ܭ�>v����mE�E8�qPI$�/��S����8��{��ܢ�>�iK �L$G/ٻ�c�	l�1��3@M��n���rsf��S\ �P��~Vd����t���_�U\#���ȳ�`�K�C�X��ϑ��]�$����3���e'N�HXe�G�ys&jm��od8r�PX�w��HG]�a����1�z�e����Mmb'2~7eY��M����Od_���&�\MT�"T�Me�)W�����\N�B��â���rU'ϑ���>��0��D=/��u�\=DY�����L���R�g�(��.�;�����LPc=�@@r�2�>�+n�J'v)������U):繇I����9�J��$�Z|�%�弚Y��������@�Ǯ_Yp�KS�Ę�5ȡ*Zb^_O��o����] �IԳQ�jO���f ��Z_.s���r�?<����}�����jXw��G����[]}g������#[���F���o�@@0��F���Jd޸Wӹt(3�e��˳K��sy�o�2�|f�EZ~�A�����+�	���~���� ��?)������[N����m�b;���iz�!z
e�r뭮�����%�<�wL݌/q�atc����]���U��a"ey���-��+��p���h#a�����Cە7��+N���:{�;��]��e%/N�x3b`�%�:���6�$�E�>�e����wg:D�z4�=y�����i������鰢������^��u�<^�7-1��3ֻa`�(-�m>�%���+�Ĳ���G�^,�,O�Ⱦ#�K��P���E�I����Qi�%��[�t��
�t��<+����G�� W3࿥*�-Pk׷p��j����rZ(�]%G�V�i'��F;���{j6o�9�h#ٶ���.Zԧ��r+�  �u ����X@�g���ݵ�<H���Z�AM����	Թ��+�E��!���-���� �[г�t�Q�8�;�m������lF��<�fl�^�ٌL6��c�H,�e�!y������ʨu;��W��}l��A�[HL��|�c%:'���a�&s9H�l��ha3z쵤Oa̤�ٝ|Oq7$g��F����9'Z�Z�5�9#�R��b�Bѡ�$�$5w���-,J-���9�Pg��טD���2v�;�z����\��f?�h;ӊV�����{�\@:* W�<�Ү���Cxv��
ũ���	��|��,\'C?j_����#�-)g:d�D}������U��4�6:"M]>l��i�;Ak���v"/\)NيwQ�S*�*�w��?ge0⅕읤 �\��.i��a_��f�B���d�k$���mI<U�-/�y�	����e�E� �]��g�7ǒ���{��Z�T'�Ӌ1� ��s�|��
�J��	�̌�BS�z���/ٓ��h\��E	d8��<�^�n7� )42�Y`�R�.�<%D���30g����L�Ё��qq/�F��ޓ�7~S���K[��TO�M�]����6z_�-�1)u�SG��ǒ�<�J�˸|M d�o��(����:�"J��u >���/e��!�7ҹ�Bׄ�\�'^�f�)�g���ʘC�[4<�9)����HUW��aі:m�j�G.�J�b�\j��h(�.�ͯ��4�@u���k>B
�2ݓ�3V���L�01���`5<��7����� 1i����l1�	��C�Ä���d�g�b��x��^F�ա(G#U8���XN���3�Ɋ���؟�.��,E�#'��)kb�7���_Ġj-�.&���{VK�ҹ����h�������^>c���q�e��>���(Jq�n�f6�4�1}.��vՄ�n���=�-�j
�a�1��;�}�{�� ����DT��\�_H�R�rv����`���@�n	]4�AЗ║��?�%�o�r�{\ԍ�(;)��u��q,��q �z���՞��T�&���2��M����cr��'�o�Y���r������Cp"����+����?eݝ �3p�i������i�[ǯ��+�J{{��}�^���k�(�fJ< �"gt��ʀ�����ܖ�s�5N�z~�����G�z�L9��*Z:쾈�XR2��tx����8x  l��甬ƀ�6�#?�,BP��'d��v��oki�V�9�b���f@y����@�;Oh���.<���H�٬�����.�-5Z��w�\���4VW+C��4��mo:>D�7Kr���d��K��f��r��kh�3u��������W�L+�E�#�D*sR��)�P�L���i��٤��ǖ+�!��Έ'�`{4�T�s��ym>��S�8O��Y8�r�B�ddÝ�M�L����d�0�j��+�
�2���/�X*����ΗF��/��:����2G  # ̮����2�!�y�ֈW��;��_G�5ucX{�N��о�Ӊ�/��uU�k��g���n{Έ�W��O>>|0 4����v�{KU��4��#����a*9���K7��e��l��+�\�0!�*Y ߧ1�i[�b������k���}�k2K�.��,��@OF)4-K��hl��zU �Q�H���P�Ov8�H�?��ُ�63A����&b��^������	�h[VF��h�*
Q��r�43���I��c
�-^�Za�^+&�[�P�hN��U(j�t��i@\x}i9nŐ����*}�� �JQ+D`��uIL�;o�	ӣ�Z�%��/�ZCI��Z�k�񷬴�(��rS�X�5�~3�fvN}�`X�@ي�Ƒ�.Y43��N��:a�t���"�����+�t =�O,<�t��@_�2 ��E��3� 	�)*���++��ŅK��Û�[�[d\���!\�=���׸9FmY�>��*�.{��b���rf46w�n�'g��`����ڬ:F���2�
7�8�_~����w���9���~z������l9��}3��abQ��V3c3�<��B"�ݧ2oo�2QvUq���"]n��}�̂[��v�q���R$��P�<��𴇄f�ҶO�VP0R�2P��U>)�j,�7���l��Ⴐ�AK�[Tp�f�{3&=����p��
���A��y4}d��P��y���0JH�I����y���'�7�=��Q@�.��2(~����I�L}�<.��簰�p�r�}�$�Ri� ̀�I���;ǥ,!�~oc{�}����WH ~�/�޸�T���i��Q5��ٜ)�ѡlN~3p*4�*#�]c`�[������]ȃuN��b7�a��_��8�k�=���p�g2�o�xF�%��H��B]�h�|��9�d7���L0����?�o
l\� �M`����^w~5R�{==&ƺ�&2�↶���ONH[P�R��8Ag:��՟�Ѽ�5(�R����[�r:�����QƩD5�/-��o3N��0'B�8�~cGQ���PHHS*;5�6�q��vE���jgKN�9��f��(�=s'i�z�t,�4�E 9Zg��ڱTZ�o�m��q�Q�.�^����|x;��g��!|4�hhr��oz����Ij�~�&e����Ȫ�)U��V��sS����!�J�^�����d>�F'��'��F��!+����T��M�� "���u:x�Y���B+�����ʒ�����M9<��1�T�y�"�?���0@^�%1Z���
ĠCx9�|������&RoP>Z���,^���:�m�3"ܢ�a�%sf��� �<���*�|s�iF;;�����נ�j��d�,�w���j�$͗��D�<BA�����=<�����Z�9�(��)�k��#����4OE}x�^N��x�0W���I}~��w&�6S�+ol�����$���s9�݉)�W7����?ɐOb����I^@|Z�>l7L+�>T!?����.�Ė�(��I:�l]Æ�wa�钱��	�v��Ч+|`�a�o0N��z�>0��DQ,��\���״��@�@�,?���E__@���!�;;`Q��9f^"���*�����%��9�`��BD+/@+�{9�`)�MC0�vr!�1HQ�I0.,}��c�#Ne�țp5���Ӽ����"a��=P�����!����>d��,iO�����;��<�kaC����ODb�Z	>}��#�Q���ՕD��	�,���W���f�A �Gf�v�����i$�C����ⵄ���  ��Eݸ;�� �g�u+j��w�lae�6'��vǁ��L���rcx����=���&<$�JX���޴%4=QU��=�����LP59 ���44)��M
ߺl�^UCk��C&�X��d�t&O�̌�p�t�!��'��CMj�Sm߽����"�}�>|�5="�W.JOc���6sp	)q�װtd��N�������}�@l�w�����4���`�itz�鶏�zw�����IOh�u��|��P��.��^VZ�8�P*+M��9��|�UD�e� �sO�zk��O�f�e�*y!H�Y;��ݎ�8f�����<���nǫZ��e�Z�F1��K��5i�����m�*�1�k���/�'vH=E�i2�3:�&�
����B�@)�ǡ%�{n�#r�>.���K����R%�1����d�{��6B��rzjd������:�~*[�f�}��>)[u�P:���)e�9������G?yE���e�����S��ݦT[�}�p��-n��>3�~�ex��~U�.<�/�tM�.ɂ�צ)�3��Ζ����ԟ~�d��R�����K���:�c�a��-��Ǝ'IC�a��b$94���~��pOvHa�^W���c��7�>����*/���7���%6�w��'e���B	``�>Zɯ��d�<���/�}��*J�&�i��g6�,=a�1o���2)�5I
�E<E���3����ʤq���J����w������~f8�/qk�^�b�M?�3��J:i�찴J�i��ZI�-��G���ߨ�1� ��l�R%a��|���F�=$�̙1)lC�Ⳟ�Ivwp�˸�仩T,����9,r��Kg�c�8!B�n�E��?��Z��j����A!�ݕ�&l���w:���_�E�� V�
;Sa�Z�~+�+�ڻ�6B�Eʹ�2�R�o�4�Q��䁓��S��9�(��.�==�����s�>R�����XU�e@R�Kn�`�
6[E�������&}g��	 u���ʪ���I��n����<����6�#j���F�L_�������w6$y�7� +y˶���(��e0r��'C6	C7;�=��{�b��?NԷ
[�6�l�F0u紲�F��g�>�e�_��ԩ"t@�k�l	jR;i����	�@����!0��n�Q� �l7\�hv������Ӂ)��H�+B�"���%�Թ��E�ÛV�rM�'mä� }๿�؊���եO*j�4YI��lS��(}8��b�E_")ӷ��'�\���c�^��׭a'���n�O�z��,B��c8z�F�� Ȟ� RGL�-�č�s|n���G5<|c���e�}_�����l>��;!_��ۚ�����s�s�V:��L)�G�iǗ�Պ�&OQ�l�i�vk6^� FX�։k�oR�d]T��~�
��C�+Z(�u�s�˿,aWs��D��A�_�M���/�:��޷��Xv�|J)�7�a��W���<��PDƕ���x�RB�\NW�.�ja�>\,�G���+����Mu���f��g����ŌyE�װ��q��3����j2J��� 5�d�'3���4M�g���ě����>���A<�/�S/��?�^;�|���z��i�4���3k�:dM��Y�g�8�g,�xɧ�Sj���9GRo��e�a�`ԉ�nF���fc�hg~���as�M&�З���?��6^mAD1�-�z���hc3�YX�t��KB���̶k������^~�i�k\�p �̱	��d$��I
T���2�.7_OڦGUSN`�Z`BуX�]�nU���$�X��r=ٞ�+��:p��L	��R���4�7T��Eb�\GΓ
ܳЁS���1q�Pm{����$�6>��
tU}A2Qh����Q�*�[F�!\�|�wGn��F�86`����S��F��&1��꺩�� d�EW���C��1��c�K%��XUfS�3�}����֍�����e�䒕�JOf�L��M�����i���e"}x����@!��UWq���(���v�D:�<DA�;i�=��F�4�
�lƫ��$w�DG���[s(tәd�"��{T}��+H���QB�#�r�׋[j����ɰ�Y������E��Л0�DY�ї�*	�r��sǔ�=Ed�Q�u!W��&�����)����+uzђ����<������Bj���^C�Ą"�%G����Ʃ� /��`����i�b�9��$���Xox��^�g�hhl�!J��0��ʴ���������1��ɶIPqf{{����~�α���=�CAw�T�t�>��(ȇ�&{��pE:.w�E���g$�þ�iY��F�wr$��,��N��{�c{�Ƙ�-�����RT|j��4�G�\*����8�Q'�N��E7-��͑(���.���]���Tw	�t�E����{D�J�ӸE�0/�;b`Q��s����Z��W�~0�����Gf�F��B�O������+-�uDy���k�M�)��m@a>S���}ilG�����v����sI�'+��gk	+QQ\�w��j�q�{$��2e�'�e#dwї�v%�\mxgAd�I�,y�0w�Q��w `�[M��T9U �Z��P%p����`�D�����j����Ƽ�#�:n{�W����v��i�)�ś��r�O�n��s5�Cܭ��,����1�T���J���;�fj�6�rS�1K맓��x��{��7����HB\ʇ>�A3c��p8�c�����*������@p�>�߁� =*��N��X'q�++SX�F,	om G�=�'&<Y %��q� ��;�k�`�e�M�-K=o)~jf���8�B3�^��/�Ԟ-����t��*s0�{QQ�O��<l�/[�a���ߝh��C�CH�RP�X'�=�*7p�,�g�\̨��.�=�:˄�n��W���(p���O^�n�S�eJ�m��;G���:U��-����*P_ѣ��:���>�lg���Y�E ��A��Z7�Yi��T���Qظ|�L�����T+-��0-1�p�L(1�L]~�[!36�����I��P9��ᛳPe���ʘU��m+��Z:�F߷7����Y�v�ؑg�e*NF%�T���p儀�(#O�����?��f�M���b	����>>>j�"�W�� h���Ļ(����|lh���n�t�o��[+%�j��+��}����E�q)p�����G��%Cb1;���Xr�녽-|qQ鋱���D'3<�ݾW�|I�t�8�T��Nb�2�Σg�Z<x���8�	�~Ά��0���Ýc�&��<<b�9̽������"��eh���9��O��Яl�9"b:��.�E���T�)�/��g�ǀ,H��h�bMt˚����Q	��e@���0���bоU�B"�Š[!-����`z�6�2�%Hg�$@���E�,0�����ϱ	KG���鲧����Md�A�S6�@m�g�^�ˍ��H�E�%~��4�tȘ����~���>���(
Y��wIsG��Da"�����r��JBXX���Wǈk4��V=�'!�����Wp�?�Շ���\�yW�����,�{�耻}�)dFԼ��}���e�xf�`G�װǨ�����:"ha�b�ϧ:�����C�/1���Է�մd?p칮�����
t`�n��� #R8.��<i^�d�8���!_::�>RJv�t�;����Es�nռ�QxB��^9L��A���70�gi�'=�=\�9�(�/ޗ�I���Ǿ�"�Rb���0MK��$E}OE��\�O�[vg����R ێj��Ǐ�`0�pa[�n��o���$|g<�)Ir'	����[?\ֈ���RS���֩!/��<iN��p�1����tM�4����8�BS��_@	{�;��w���9.�$r$/$��a9cg�n�Q)�td���fR'訠m�&�1B�n��_rOj��3n�i��to��Чf����"R�i��4�3"�^�r�Ĉ��w&L�3%7]��EZ�B�0E�
ڇ�w��[�݌���Y��,�y'N�,%?P�|�x�����j�tz|�d��2�u�xUF�;��x.��m�ؓж�8�#�[*����,��ƭ��3S�.��D���Ĕ�N�����(�6u.���!��+4�J&��D�����)}Om��������
�k�Ms��F�V vQ���'ǎ6�J&V<����?��cf��®�>�F�ǻ� �Re�k �_9D�%vT�v3[�欝��H�'^�E׋/<pZ.��k�x�L�tDG�S�L��L�=���R��B��,��V�J���D��K���|� !F	�p���CH�iiR'�f���kc��A(IcφC�Y�d��/O!7;Ã���Hen�rd5{�ɖƯ�xD��@w�$�����:��u�����[��%����,q����\���-��t����8ߋ�/H�^_��AH�$��ׇ`Q�c�pv��D<(��x�j��v�d����
�I3��H�Z(�4tv���Ira<0`�����w��Ja�t_�q)�նG���}4�	u ��{��C��3L�hMR�n�C#��t��@o1�Eh ��e(�q�O�����ȟ˘g�ٞ���p/����;A�t��՚��i��Di��d��.�xH���]��(��I��(�m�����'rĖ��4S�H1C�7���Y3��g�-��9�%v�ղKC�]΃*-��8��6�����F��HHp �^ދ�d7q��i���0"�=�Qne�$dT�o���J6c�
���"؞�n�R���s��*���Zl5��l2M�B,	�6_��G�ꎩ1����Z
03�wJ�$Hq����u[3��O���7z�F�p�g��,�y�?b�*�&2өw��<D��ym�T'� _Q�'��+a��X\a'M{G7w���o���3CN�I����P 2�[Pڛ<�њ�P#u��?��b	-Ri�.�����mK^�;T�S��F�E� N'�ZXF�B�����a\H#�+�ٓ��rq�ű3��	���KӉr�u{D̒e�-�@��p�|}�l!/�ќ5�O��u��LE�sr�*��1��n����(-a���9��tf0gMm�.��T��0�2��BXIW=��]a`��f(���<x`_w��C�F���D�r)�1��A@�ߥ/ハ5�7O���B$b�|��z�S��<�iX�	������¦WV	�������٫�U>���nC�̝��v�A���d�ic
n������&�c�e��k�?噒r�l�qh�Yz����6,e�2����ikR�1�"�Ⅽ��v�j$�q�UP1��%IQT|8���u5D`R�s>��Ve��Qr��iH�p�E��7�!����������A�D���%5ߛ�%(0�Y�_���V��y�/Ī�+s"��0飯�T��*�"�s��G��B� �qs��8����.?��$�Y��(�7���	iJ�8�
4�&-�j`A�駺�U�D��}�ڟ�?�Wx4?�s�*P�4�@rJ�{�2�QA��}$�J��sh�V�%��H�	�3S}J"��SU��tj�5��6Q��ر��=LM6j�{#0����&�RU���"s%N�7p�ãTX���kz�\�&%�F����c��{�qTE���6�ɨ�D�+������6���)}�N�J+o�����ւ9�T��!�job��!P�[���^��R���:�sV@�)ҕ�0��4ٗ�J�2"W�b�Z���#�� �L,%�e�9s~�e��)k�OHl<-{m�G�.`4��V�αGS>̦�T���{m�m�b٢lvIE_�x�����^�"���׋-m���q�)�\`�/D���9G��?�B�)��=C���$����.�#��>���!��W��'����o.�{��h�Ȋ��R^���Pvi�������zW#�֮���
�)�$3�I2%�[n?�ܼv2�l�\bYH�Ers�Z�Ӭ�&¯�����DA�܉�����=�`���h-<��&�'��v��d>���a�Nw"�#UAZ�o嗅�		
�8�XV�����5c?�V&q���`U6�1���l"��������U	O�K8"���GVsF#�t�V�q��它��#7��-\q��0xr�=�a�~A��f�(q�Q{�f�|�{��k;ZB���2��i��'INVĸj��b�S��r8�$J)Ȧ�D�F��~C�Z�5,��$l.����]7�@�d^%��˺�������\QM���0�H�����Ɗ6�Γ.Tm-����f.ʷ��cE/*�w�~�dd�?ى�v�&J�V���3�a��ٶ�����`�Ö�F�����i騸���3(C��B����q_�Jle��%����U{�����ȅ�)�B�j;��0� ֳ�9k����Q����@�F�X�uay;��R��"��oC�^炅�v����.3�\s縣ߺL�:��*z�~N���9���Mq��nJ���,t4��o�5a.s����2ٱ^�[���<򾈏8''7�!��o�5�zߧ�b��/�P�o�d!�Q��?��2o�BI���q�	��v�W�N�����Y3���%^��N@��aLt|W��Fڀ	�r�|��\_�n��U����Y���W�S!��Fl��6PrBƭ[Hw���W��̩[�����E�t��y�_��tY̓�\,��o�7�Zݽk̍ză{�{��]�X���ȨK���i9/��aj�#1L��I���?:�5��n{��f���wN7(���ӽ�wi+У �D�G�R ����c4���݌�����p�$�q�쌠�qP�"���X{t7@9oN���Is�}��6L<����}�$�$!R��|7��F�q.67֡2���w7!�g����@V߶|�g��"���JC�僕6��iٲ�.�5��8	����[2n���䫀�weQ����6��u�q�m;?�/AbK��F�ҷ�o؏a(��v�,������:�;X}N�q�0�����&>����:�����׵W�H�+�+3>���F�C�zM+q���ߕe����}0� �Qʸq3PY�D��a���j��k=���S�;<�j�(�܈��MG�P�����i��o���� ��#�Nh�%��f_��t]&aY,*���)��m���lg}]|��'�\�ۜ�����-�I� �k����u�#c��5�ƨ=m��I@k�}V�(���t�;��S�-/^�-����j�?V �|m�K�֮��*z36L��c�eBT����R+[n-h�JJ�R^�Z���MA�R�B�����a���es���1!ZikUUU3n���F}kb���������B��_�Zj25Iw��g
Wʕxr�jR�
�6^�]�����)�K�jF��I�9��b����x;w����� d#��6J����B�杻��[��pW��ơ��)-k״��z�el|V�&�TḥEe��o���]��ZH���nm�s�/����2��@|N���ps1�?���&ɕ�g���p�����tZ��#D�l$*�k� ��-U!�Z�Mťp�a|Sx��͒K�aE���mq�`��-@�
�YR�YF5��8�'h�(�Ԭ T�
Ti*��E#��D�Gx/�9�i���H)ݳ��i����Т�|:�F��
�h���t����,�#��_r@X?��m�Ԡ�cm��$`� e�7�H�?D��#7���ÕZ:�ee)���ܞ4s����=�I�����$\9�~�$e�"C�\<���"�7o_�{����'��^���_p�ɮ�n��f�=1=+�
%�l<�E��X��z#֎���~�ۘ���i���øI��;-���oV��qǊ�����o���D�r%��@���,��y�+!;!��~G�u�!����O����|�J?�O�͔�Vx,��l�Q�0飩����jEDN��C���G�����J9��=�{�h�v��\q��p8>������&���'.�=�Vfe�BAv�@��� g�g׫��e���9K̦S��Re���_.��C�yS��仴ӹ�c������Es���^o��������� *.!��-L�B1��N�ӇpR��j�N�\Ə}!�	�?4+p(�IQ�_	�5�qm�������~h��l	d�fU���>	O4)o/���7o�a�ɒ��5I:�&X9r�Rm�@��O�c@�����a�jYe"�ǜ�[,���-�_��
e%�ݔ-P�{�� Ф��۵���Mc�]ֿG
�����a[��xVG4>H݀�7��ص�����K�[���|]�	*Ud�+E��7#3�G<�2�/q����Ɛ�tG�4�7(�8�Hh���d�I���s���z�� FYLD�(�h��'d�T.���p B�3�&=�ߎ���:م]`�X���a��n�z�F5�Fd:�^����b��}��?L��vz��V����������^���%��Ծa�^�x�,��/��S��
�Lsgφt<���5:6���';�����f�@��f����o�J�o	�����4t�vR�Y��p�p斲�G��m��c��X;���`���Я�h1�G�o�ΑiOƊH�`?׈��RG�
ܵ���� �.H�K����&��]���ƨ�Ro'��&�1��_�Qb��H��/��{d�Dh/�@JJl��F.zÉ���?*����iv+�����2'Fe�Ls�q���i|X~��G�Lv"�{ap����P���ң�e�9͇,�� ��.C7�o�+��Z�1�8���ǅ��Ε��<�Ʊ��#%���j��q�����H?I{5�H�I(�)�{��L����"���o>��,~�g�%���]a���R��G'�ptK����i��~����>_�\u H���=��WZ�=E���V�G�E[ߠ~��jV彮��G!����絹n�7�2O�o�j�cd�;��NKO����ۛ�S#���PvH��Qj�A	c<'��xi�,!4�����B�ߠ7�H���~O�S2�zi-.�����{�5�$�mC�b �[�#'K�Y>$M@�{��lU>?M)ȑ��i�{�!*�!��.���%��X8���y�q}�?����7n1q�U�:t9Q�LOn�^�����t*ei�0�lä���.�*1b�3b��m�s�ҿ��,4�RE{��D��>�Dgm8ڷTE��������1�Cխ��o�GSW�@�V2D��*2��+�x:����S�u�����8��+oL��s"��-��5E	$�њ�o���Ņ��x��P����AK��	+MWՇG���<�p" ]�(�jv�bPP�M���L���e�&���+�X)M�������RTA�J:ܶ̕�=d�&3�Bz��J�.k���H�|m����KkD���r��!�[�KN�Y�(���#UI�.�j8D�n��q7e�,����$�B�us,_����r*����W�cG���k��
Uox��	�3u���##�(٫���f`��`H��;�x9ujj*w�Y�w�3���!�91�%t�pi�S�m��nP�dF�O�DYh5J{�tZ�UA��}���CB�B���9t7��U7����A~���(�ls�4���3�@V�3?�H��Jqg ]�d$��(sa��N�Q�kB=����9!��Cy<p�p��R�[��j0�iV�w�ܶ���	��d/;]�q��Υ+�IW�7'�]
�Zs�q�l�?�����H�gh�.����7=��)���+����~ۯDe��$�D��N�wc�����M>8Ɗ���6�Ž�����Ը�V
Z�s9i���*Z���4�B+�c�
D'����$�0ש+?�4���	A�jHt9�]�t����o��|u{H�Ȇ�e�aa��j&�~��w���4:������Pp��u�P�*[�ϩ����BP�D�t��Wk��ݙ���p��g�H#=rnG��j�eM$=��n2�o~v[��܂�޷d���s�hݿo�v�Ք���Bd}	�O5d(E���<��ք�ŗ:龴k�A�K}Tf��fנ����/xD~�/����;AP�,�w��.�l�͎���,�<"��ԅ��:	۫�(΀TĞ�"�D��A���KE���Vh�O��f�NG8
ۦ��C�v¸��6^�Z� [���H7���^M&���Ηe�ggO�l
��EI�Y��5u@�P��甕�2��B'p�?�x���T�V�����c�O\=A�r�Q�d���C)
��(bT��w���/��f��B���VD)Hl�ZB�92�wє�`�0���"n�C��ǵ����;�,_ :���Z�?�r�J�����&Q}Up;���?�fmC�?[�[��=��,ߍN+Օ2��:�O�4�8~�]Ij@	��S���l�]���Q�E��z�D�~���UFY��B7����j�n�p�/��ŷ&���Tu�K��o[�&нY�ԝ�|�q��~�*�MKG�Vp>�@<�]� L���@���ב�/
"�w����&[��z4���A��s����f1�ck��#0�Բo9\_��|8Q0������⃒e�$���S��;ClX�'������æY�5�ka�,�@d'�һ�'u�Z{/�):p 09�2r�SUa�lda7�� �g�\GJ2Z=��.�-0�N�r��*��o[��*^;���CqHv��go�sA]�ʗQ7�M
�o'�#KU3/��!��^]}��a?`���Z�~�[N�iE�^Mt�:��t�&���9�����-�'����c�uP���w+��a��F�m<�d�(����ɇ�
��Oᨂ{��8�D�"�$�������sH,F�Ig@�M[Ǹ~
��H(K���_�Iq�kIǰL���K]L�}V�b��t�0��4w$�Z��G���.W�Mu{PK��xEt��X��Tꃌ]��y��R�Ws��N��  q�NO0�&�}�{�d�^CY�ӵ`J"��H�s3�fi2X�L�e`f#�ܢ}�Ϣ�v��$M���;�rJ/��WJ�V�O��c�{\u.+;oXu�t�
�Z�C���oKT.���G��@Uݡ��8�M������6S�"h�?�pX'w�:kڼwʹ�a1�QY��
S7����"e�j(������ \US�V���ݩ-N����ۀ]O��o���R7�[�\��5���`���^��5'.Ph��	�ڦ;tPz�X��%���Q�F;�Q-m���x/
j�D3�!�ÙgpdWB��g���v�m7N6�:���}�h��[ /�XnO�Es�*1È3�	�ִ��B%�z�m��N��b-_iq21��{�BD���>��˶�۪(C�������V|�-�l�fh�7DWR�-�,���x�W�+�ެ��EG�gy����sK4��FN~a4k�����p`?��b9X�.eZ�Fd��R����m����o��z���k3@4k�s���p��^�x�^/�K�?�mj��	4wv�Hc�^/���*�S�eAV*�j|��N������R�4��$u��b�A�G�������<������X�u��t�L<������U�+�mВd�XB��b�X��$E�.�1�%ɩUn)e�#2�0��ic���D}X(�����*��ȕ4�kN��n�k�Bwi��O+%ܴ��n�1�|^����"`t8��%��;�W�u�Ѣ�h��v���׋��p�?.F���K�ՅҺ��vӎl� ��+kN������#�v{����"��K��/���j��w����F�u��]an�2��+)t�����A\��ѣ;��P���*�ơޔ�I�����<H����	�%լ�H~K1�R���������&͛X����W+����d�=��o&�e,��:�~�5��d�� �&Zhs�Z�"֧�Y��ӫXb-4��\�X��"�$.�z���R�~*��wU�i{�~��[p���
��PL�zbz,���\��Q���k��u9��l��*Y�8� ���D����<�B],���5`NC�%zeMS��&	"_o�Bƅ�oZ�2X
*�a���������#J�~=r@o1��5U���~�<肞#L�#Izu'���>��5���1i;a3�F�cdk��A��{I*�_�����9�M���׿ԳX���;U50��C�>��UFc5�f.�x\ˁ�M��KF�;���gJ�]g�����f/���z�S����qT����Ð5⊇�@��A�at���*ú�ք���}��fN�*�������������A%�8ծ��#�0jx/Dg��'�A�N�sYFp�9��{��kj+~�*n���ޔ-]"�;��桎ij��YDֲ|i�*dz�����#AI`��8�X@��R��a�n��=�
+���2Y�R�K	"Ir�HN��Kh_SN�Ȱ�}��[F��!�_x�1���%��:>.��SJ
B��S�ﭴ�YD9��jH�2����PŊ�ʋ��ə�_̥A��k[r}����fB�x�8nA��"��@�*�H�,�":���;�xulwzX7��`j׭пK���s�� aKl)t/Jĉ>����T�`ʼ�/�* �"����Nj�H�t��4��<�?Y�|�<�b��l�B` �̈��-�K\DB{�*:��k�ÕDh49�\h�W#䩢��Fčo&����.�MJ�g��&�B���VQ=�70����,wq0�J�b�̖«�o�)�\�I@���-�2��}3�^[
@���>�T�:����x��`������@�x�{�'��Rz�(,��3K0����@��^���F�` C�H���eS��l���������X���EZMn�jv���i��ƞ?�8�6�!�N��@h����C�J�!��	�'�pT�{��5k��%/���V��Ĥ��3��с�b��k�dh��*K��z�8�CF�1�Y�M�6��<��A�3��>(Ұ$9<zw��7|	��܋4e�/� *�WS��= �������6d2oa�+��I��S�'�,L����J�Q�-C[L0�E� S�d7b
R�Y�/�IQ��o4gН$�<�`��4%�$x�F����[� ��$`J����L�����3R�zȮOV�����{(9H��(��,������#��>Dˆ�q<n�����qݛ
�)��{O���hk��N��b5,c+���}~�@ϰmBvE�-!�%5��`a!����O'��'4���@r'�Mߍ�m��s{[4L�T^8v�m~�d�ꕯ�:�څ���P���>����Ķ�?Kk%7�p�2��7D�b0�p�Tn����"��S�ڪU�b���ߓ֨c�@�1��ˁC�Z`0^�X �J���\R����wLY %k:���8yȼI�u{�^��s���lg^�yI� >@W��_H�7yJ�j<$Dg�%}��ҍ��;s�]X]r�^}�/�U�Б����K2�X��Z@����;b*g��_p��٫:�!0nf�+�8�Q���1t�N��_7��O�J��>�����rM� U>��_���{�pGc5�)u��/汶28b�˚���S+Q�����y����P7@�B��Z(ڗ�v����ͭ��-eG�s�s���ޱ�6;�mMO�@��� ֗���Y�{} 2׉�M-��)s:�Lm���@��L�I�0M:���.���]By��FvLf^�V����W��
IB�7UI�����N�]"ϼ�#&F<�/�٪�]q!Ok}8[ T�,<�j5����M��m�������x�����s˝��6����%�'��Q@�*�}���%�p�۝$�f�g�V��"_U�}�r&�l���DO�	}�����H'�9z��X0�����<��6��N�k>�ti�'�8ƍ�5>���h��mq�ݿ�ZEa�n,�:��'�xW�u�����ꄞ)��)g�' BTSq<�����u�4i���������t��p�.m�I�M���k�fǚGg�C����N�����y����?Fp�{ ����J�����n��P�H��o%�d6y�}ܙQ��b��%���C� �����KŅ��n���T�½�w�?;���:HUe�ɮiJt��/�z��b/��cx�󖠮#AT-��u͚�"�/��U�R��2*�����X�{Z�@��d��"	�����<����u�c�J84��̐�.5�_ȯ[e�ob�e�Be4�Ґ��6�����׏�G���/�/�nx��˞�h����VR�B�i�(�ĳ����7���[��#ls�R�	"$�qŦL4gJ,P�=����/��#�|N��6�MԱ�+&���H8y��߀F�:�;:�_n��9Pq�03S�9�5,������{��3g�!�.���z���%���X�����1�BL/,O�Sj`�6:�c����ό="}���f�-������x�E�@ T�{�~ҟ$�q�'���ݱ�<Z���>}�>��WP���
B���Y��q��;����v�C�.͌����A"6x�&YT�g!*o��U*��&���3���i�$�;�Ҡ�*om[ț�[.�|&��X w@ؓ��ڳ���
����h{i=L{�n�;r�,�|z����V��w��G3MQʳJT&G�vʾ���}o�0��)�f�V�M�<�-tqX3i(R,�����Y�Y[~a*ʭ���R��O��፬���m�FpaXP9�Bh	���Et*��u0tw�p���{d�6D��(|P��9.��,�8�aK��f��AH�}�]Y��@���W�C/x�v��w@���N"�&M|1Dmͯ'���k�\ˍ��U�_!�.���S�`�6L�M��g*�c#	2���!�	'&i$q8���;P��VA{gx�q��~C~�!�]dS9m�o��à"4/��hd&�h�F���s�X��Yv�X�Zx�:UG��B
u_�\��'#�)JG�'cOR���B̆Ƣ:��CӃ�jy^��F��A�@P�VMM�ѧ_V���ݙ�h�_�֤���gK�ה- N�$4zzۼ�~�>,I�D� �J����]�q/t��.���fv�E��%��923"wb󆼗�|}ƥ��'�!b�| �����^��@i"��g3n3��ɑ�6�۾����v��l`AL�;I��n�� �S��S%�~?@2�Ev����-k�n1��	�eI_�YVE���V;=�#�Z���mI�,ع���x����xN'Wogl�RK�FD5D���TrN�6ƿ�i�h!��)�'����~+˽�2�:9���B����5�K����S���)A���HH��e��}��4�Mf��E���u�S��W��y�'�S���;�'�$�>��k�ZX�j���!�p� �^z{ff�G壢&0Н���o��|�-¶	�6�%,����1�X�v�KúhU�fBIx?rR�l��	��t8�3�^��Զ9�%ܴ�s�{�{Á����ss�2Аa���a�)����8����{k��)v�~p𒙹��� m��ǔt��q1�m�ȣ8ݙ���i���q�!��C�6җ�ET	�3�M����V��a`����m���[���-t:b�U��/�7x8q!_W���Nu�`���@Q���[�+�:���-��td�i�`o~>P���,�����+n3Q]���^A�<E��p�����om����4��J5��'���~�`4=0hڂ}p�ԙ���2�
D��u��lx���En�ζ��LIѸ��V���uo����!�~zu} !P�z��б�U�^6wDP\+i���E�a�؄$1�{���_��6u1(�&����DӷNm�-���Ë�m�?��ɸ 1Z��7��Z�
q�4k����'9O��6�ק�T-12n]VKB�p|��_b��B7�p�L�f)���_��]�ʕx4���� ��T^�T�^%&{��
`j%b�������Ԧ偐�k��P�\F�2�R������.T Ũ�2�e����%���eT���:���E�������.��'S��o(������YW[	>;T����|E�����x6F��ء$D��h&����:yj+ֿGv���mɽS���7� �ڹ_��ձ	�s��Jj�tG�$�����G�!�g�^��d�A���Q�RYk��3�lp5�����J�+�P��Mn-��&y��h�c?J�L�d��)�左�Ya�B:�O.�S��p=����e)jn��I�������A@܀�(��	e2U3��eUE��4@z9��ǒU���̟9y�B:̖�VV��� �]��g^l�X�cݱy�L�T�?�"�X���/H�	"QP�9DdߨV�7���㖥'9��`)���~3n��X!���M6u��b�=��Y�U_įD�sYAҊ!�N�^nƗ<ޜ����=�Å}�G�*�6�������w����<>�Oh*���*�'�g�Z%V��i�i�)w��&�!G��u>��WV��ڶ�ċ9Ԏ�T��^�;T��nj{}R�TBx��Y�
�Mo"A�d�<�x[$Z' }���<�X��s���L��|����&:t]'#���&��ep�	�Z��v�B����N���7�U��Id}pW�`�i 6�M��R�Ek/2P�&]�F�Skψ�n�#$�|>v��3�Ʒ6�rw�Ly�q���"���k7�!7L��n!*���O\D^Nդ���fm�6���$W�wÈꕩ��af��,���?W4�:0���Y]I�`�������z!�L���~j�n��v��]�s���?�q��C���ac��}�_`l����ݼ?C�W���Yf��,.,�J��	[ �Cݳ�*o7k`�M7��p�S9՛`��_�?�*��Jp:��13s��K����SW�|�{������2zW��^+����k��!���P��m�>���}�����E%�ڬ��q����u�}f�c�k����Yc�oh����� �ƞ�"��8-+�����{�ۛ>ZM/Q�7�
}S�G#3Ƥ��[$  �
��{5�����TÅl�S�A��Β=ˍ�N ��NA���D	�P~&$�7X��Rgt�y���r�E�H��dA�E?�p�G�!��|
�(�q~'ˊ�5r�h@�N�4n��/OxOh��A���f�]8���g�8m`޹rͅ�Nvjt�ms�ʡ����o3����އFj�u@�q��
�|.���$��Dpvge!�ā[�/�N�/�׭��|�%�S]VS�䔕X\��@� h9��-�h����K���)����,�o��6�;#�#��/(�cU�&j�H)�oç%W��8<@B���cu����>�h�c�j}B�D�l2�ÖٞQ�x�{�ɨ�6�+���_�A�-�(���lS�Y���:�r�dB+��y�H����G
��� ��M�	U�f�h@�N����v��Ig������_ ih �(�M����76����r=N��E2�c��Z�Q]���B검Z�%~�c��x5���eկ��>�٫����f��m}j�l�ć���
(���M�P����3N� ?���8��C���Z�
n��B��<�W&ˢ��eb߁P��Vp�H�yc!X�XO3<{UWV_$z�e��g���0^$L��"dk���Ht\���J]֨�su��p��>���\�^)o��Ql���ֶ�N�c'l��[��8���ԉQ�3��� A�����ܞ�����F�\��=A�ƀҞ�@�R;9��L9J<�z���t_�D��!4ٯљ��d��Nؓ�l�NΠ�&\���% � 3��I�C&�uً��^�X�|۸�V�ӭ��-�Pj��Ґ�����N��8Qi���߂��'��o�R΁ϸv(���x� �?E̫� %�W�i�lH�?���"�DS����aw�o� $�zsベхŷX���-��
�}s���@ڷ�qq �r>�C�Ӕ@N4�^��X�S`��L�>��3B߲U�)��ܛ�6����~��	^�xσ�,f�,��N�M3Z=plrM�������¬íݞ@�.� C��FIb���"��utOT�q�'prw|��g����r��}_^����s+iNx���f�d����͟N�=�^\�Y��@��ݙ�Gm���)�}���0��N&�>u���\[M�(������%���M�������l8��ha"��(s&�þ������Z��Ϣ����a�PI�*��oi�����7YK��=�:ız��"
��s�&�~���u e�쨦�)Nͱ9��G�42SG r�T����I�͂�3v=�����9g�^������H/���{D������g�tˤy��R���@� ��K:��z��5��'!�^n�0�2O��|p����Ou���^Hǳ���Y�E|��I��E�d�_-'���q���I��ː<��bI�%��b��Z.�<�L~��_vmd_V�$ڢ�
�L���6q��Ov�?UkPCh��u��x��.�!�q�0Vu��uϿ�Mjd�9k��H�������k��m����H�������1�,����*�����k�$N���T㇇`���<����:�]{��g6dZ��!
���Lʥ
�i�gm�ǔ���x]d��b��f[7�5n��F�9H������w����N왙�&g�F�H��$?~�����P�Z.��Sc������+ ��b�ߥ܆�J���<rb<Ar�︪�3~bOT�D�Al5��3���J~r�@���9����[��m�JsM��g}@O�D�-<k��|By�d���ѐ�i�� ���;9�����2[<\�H�2��K��:z�P6�_2}<b����A�]�-[b��yw�n�J�o�Oze��K40�����Ǿ�s���F���aM���\��yj�q'1;��m�@�6�;?S�x�8�Bl�-.�m�,��=����_׎�%�)6_\so�K<㎸a!uO��C�e��_�!"��-�Yl�!��j�rl�ʤ���r��d��6- ���ٷ90�@!����4�5����1���׉@�Q�:�D�QB�sD^��N�yʔ��l-5�Ms-~���ڰs�8�cɬ/GZ\a���8�W�ÿ�=�
�fY\uhY[��n��j�����,�ɣ�3���J�?ё�H���10����[�~�R/�0h����n�.B9C��@���+�o�i�.�+�N�@ON���>bҠ�H�j��'����yW���ٵ7��|�0�Bq��o6��5)�\�&�FvďZ���B�d��CT<����~|�?�@���|}��(�m|��L�p��!�yi=�.�^����74��o<\Z�0xmT����N��$R�i��@�-נT/��-qBz����ͬn�,>l��`��_~fS�+헇�v�N�*I��o9����($K�@��{�X2d����3���� ��pL̈8��@8�6~�ofe�>�x���#�m��i����\Lp
��}��+V4���Q$!���w�3<�I>#X]���g,nz{�R��+J�q־�GU@׻q<dSn����,���Khn+!+��7�6�{�@5�;�,M\�O��4�"��pH�ū6��K�_����>���C3�پg
�����
�f�e�E :8j�	�7rS�R�b����v��t8A}��h,�0up�h�H�_����>����d"�����֢m�Q�F?(�I͢����k��vW��&��|���O��7��B�>��5/0��6�&�Dt�T/A���n$��GO�e��}EZ�]ܷ�e�?ye�i�����v��T	>^��*eҿ������J�����e�����_��<�C���/.��6�nd{KMa���;0��`��R�=T�mө˖	����s4�P%PU-r�&H��}�,������ө�p��Y�+�QN-�����_4i�r�c�}Ԭ5�Y�����_Dj�t�&�q�U��5�W��|���:	�Q��u��'�/�AI-פU��7��Nˏz=�Q��4Y�N(҈�ܖ��ϠCW�>4M0��&Ȝ���s-�<���Y��f�
�SaٰlV&Cx�FX0)q�c���]�I&�� =�&�G:T�z[�{��ޅ� ��+~^|��ZVQҫ�e!G:�˖J/2̌��EF���1����Ыa�3s�m%�naE��P�Z�\��ȵ��\����I�,��:�
w�$�̍8^�"��+4b��	�7zy��v�B�;�l�M���'��	�f|G�m��ZO�V�� ���<���Jʀ�j�2��DΘ��O}�> aI�V"��d��T�֚J���܌i]#t��;F��՚�@t����y�	H��xX�����iG[(��­��XlI$�?��aJ_���j�+@c�6nGV��ϩ���@��B�!��D�$Sk�;�Ǜ���i*!z+e2�ʢ�ب������5��{/}��$����c�T���sԤ��pmt�@{��𺦟@�o�X��E|��(#��H����9P2�;�VYF&.�BJ`y��u��t���tü�\P{���W]u�<F6�E�$�����te�Z�BI��X_w��g��%���p��TZ%|�����ZY�V;�{b���N�:����IC3]l�R7�4��	��N����W���g�uXr�g�g�o��Mm��p�|��3H����G����(&V�ۇ�CH���4�`��vm�K]�j�8��"��ǒ�C�y�v	j�&P���8�9��'�̤%�W��X ����3���}�ٴ�\��}�-Ԡ0+dY9�J��r�e�0�i%>T��#��BHR>������O�,�#�li;�'P?��_{�u
b��9i H�$��ն����!��zk\��.J2�E>I/1���M�8j���_�/���L��や��k�˞�ڒ�r� �ul��j.˂���ݕ�Nˠ�_���|/�9rj�[!c�X=ȒQw+� ��p�J`�Ӄ�����E�������ͤ����t�N{��M^�c�.���i��Q� �ڲ�̥\����{T��0o�n�G���%G��3��t�� ُ5��������s$孢�k)V*c��(NS�"��m0|��(����Uq������8��@�x
H��)�!a`�E�rBX,@耥Y±(���}������:V�$1���Q��Ӱ�TC��h��55Ab�	rEqp}�r�z����W���;�SOv�y���]�݆fa�X���_&�����YS��~�qJ`4A:����{G��.�c���OjeV�H�mw}��vK�sqH8Mڊ�W��6�Cc�vI3D�p�(��^s+�"--JX0�>��/p��^�ӎV�G�z������7��p������O���`+�~��Q���P��˞����VN}:��ӃW���$�Ą̊��?Og�&�#S7ſ��)%��4e�^�"��\xP9X-�f�w��Z����(u/3A�j����r3w�X�7ѓ����, ���P��I�>�>��IY�sCp��>n|�)q_=���ݙ�
GA��L����wL�4�`T�
���ȟN��cV�N:;@n�A�@&"$�@�	k7X�.	�d~�p��:)%�
��X�
��-N>F���9�ɘ�m�>[e%j���{��P
�Q������&�>#�O'B�=�
��P�{fHurw�$�.
��?QN�`�Op[^�@_&�n�c���̭c,oɺ�L���P	n�!�I:��8y��7�D8`o�M�hb@�,A��7ǖͯ A�4J$��$���|8]�-KR��Y�b�� 
B@z���'�0M�Rp�g��q#
Y�$�Wg�aa9oS��������� ����c<3�\����$��.����&�)���Y���Ƕh�q���"u�J&;7R=QQ��s��r���e�"\�ty(x��4�4|r�^Ve��)��0��ր0��=���s�췪��$Gm�c��>��n�q�	�VT� u�ns6�M�	ևpJ�K����q
r �e.�>Vr��e�:7��<��88C���`��p2c��d9���Q��#.O��Tq.i�������N{��7<E(��C��[�#���_t��Ϧ�xC�4� �B����J���j�] @�Bq�Xn���S���n�yB6Dq�Lg�-\���D�l��/hL�����o�
���F�B�FV���rł��q���U����'~t��G��	 ��T��\PϽ.Ã!Ċ�e>m�n�Q�.���]�������$�t����v��Rz�\���w��;�ݤ�}	��� o���ҥ!�&E8!�t�I�5�ٲ�<p�c]0��pӵ�Ys'Ш�9��D�#�g1k)��d�پ����*�a�L�����
�
�Kc>o��y��t+G~K��2���A �W�J�}�ɥĬ��� Q��WNv"�U5��ә�A'æ�Ҝ��K�xFɨg���{��,�%� ����%�"���"[kx{��f��ޱ�(��M7q�fp^�r�=�S���s<���HJ��S��V�F���&��Gl�9e��j��GYC��t�HW=��#ô=^u�D46���"�&��!b����٩˴ؑ8��խ���&ʯ�E8���+�4Lw��cR�D%u�N����R��/�_Թ�_g�-ĂS�$�60�=>;eC&Х����Ӗe�<�gf1Dk�^ߪe�����k�w#��ʼ#yv"+���4[����B`o�7���d�Ҙ*���6����D�	�V�����U�~�N�� Z�_|�A�Ev��8��Y}/D����6���hB��@�"Tx�屼\\�2i
���R�}�C����H~��<�K8!`��m6���|H�Pl�� �5z�ｬ�JK_�W��R�w����#[Q�Xwh')I�obnl����g5����0r��8l?vI�������~V�V���=	WJEy�`F�2ڢ.�e�E}��U��u�ʒs2t�8<�Ě7�}��<���<�X�M���T�bp�ai#��m(*Jz�����2����VqWi�Z���ɉ�A��*�J!"���veʞ�x�9E?�����"a1��0�̓�h� �0Ӥ8�O
����� ��Z]�X4�DJ�|�Ӎɻ�6J8U��v�X�H��NZ<��U��b2m���*HH5�[`�vԟ!�7y4��["��VJ��8�^b�;6?JKy��S#��� �Dg}Z@�c~�))����|&��BۯҠ���A�ZYV�f.b:?��KE6� ����<��_r�s0bA���FþHM�uq]߾�3A�̧�|�0V��)�m
��#?nԶ�����V�5N?��*��LDj9ʪ]g��~bA�Z��wN��-i>��:C�.�4�l����v��[V���~R�}R����E��{��4�:��:�|+O�#rG���}���5�����4�AMww��Lc`�����lB+��o�HP����Ϯ3ם�;����!b�q9[z	\" +���K��B������ΰ�wT�����C�'���2�+3Q����"�=-��	0��vh�v���G�H��]#�:����/LH�����w3��<��L�I�u�5��G�@q�������J���y�Ҿ�v'�'�+$�w����8o�4P-4�TW�
=�@N.�[]�d����#ڗcT�����{�a	U��'���1.-�a�6�[�PөM��cG�>Ӗ�jX�ʫ"N��.�ΎYB;����$yt�O7f_���x�R�@�0��������YOu�"�F�9T�t`t���3�Q��K#��M��ͱ�H!�� ��އ����vʟY��}�	��K[�g��u6\�"��f�m�d����Ko����s%C|�%���\�c���
b��b[{ֿ^P�EE��ҙ1f;3<!w�b�I��n��4"�'�e$�"�7����4�|��ݪ��8䪃��~��8���	e66��K�Hx���K��qDU^;7�r�I��{*>�.5���X�T�:.�ח�7���mu�}
�//T�����W�Ɵ,�7`�I�ۈ<<T�5ٗ�-G�$��"�Cٖ޷�𱨋���1��E���M!%|W��m,�v��^�q'�:ؓ)�_۽���Z�W`h%�0V��Knz��(E)���ߩ�%��SwZTY����Q7J?P��8����9]�X�W�y�q��5S��*N��w�ܬ1�YLB@����B��.�\I� жVf����}z�&�v⏜�pn��9��Bh�����k���y��������BR�
Y�m�/�I�w^[��V}p�K�����|��v��0�:K'L7����n!U{Y���g�mN�v�װ�� ��f#�>�}"��nˮ�5U�wȠ�`^�&�*�pT6���������|8c�X����'�#+�q	�KA�C�#��Tퟄ�)���/v��{� �Np;��^6�^�����ܟօH*�x��0�A� ��c.���X�y]L�E;��¡�[�m��3z� oK�xP?�s��c]� ��t��l�Uz�i�5�q���3��§[����
H�!�U�e��[����T���1	֊j���K�`#-��ِ�K̉�W��L�"�M��<�������d�5A4�2�¶�ll
�cќ����RG���ԣ��bv2h3�߾�e��B�[~!��I�Ř�#�
��V��$��i��"�Hyƙ��֝��DM��h�T2�(&�{�1S�[�&�ں�����1� �H����~�=�����n��ٔ�l{���ۋ|�6؃��� �;"|��~��a�|�7�θTQ�X��J��$�����CP���w�mtSy�f�N�-�鯛I�!�͹�5�1E/nE�����$�C^�x^��H3�@I�$gV���<ʞ��R�NԀKc#SHՌܫ�f��
v��Y��j$$�2��M��n�8H�������wH�a}��o��;Y�`ǀ��`
�I�I%u���8Z��g��J�^.���u�u�_t��8���>ԯ�E8W�X��u��vM��Qg�!���R�.~9ا��˼��e*l7��=	еo��C���,!�z�Q	�͒]o.vQ�Ĭo�C�tztd�giX��"s�0a<#̔�������CW`�
$��O�/�����,c���Dҫ���;Gi����i�E��;x�O��qݽ��{�+�Y�#@���,�Sb�,M�֙�N*L�U>`��L��`=����06gj%�ϟ�:��%��u ^��?�ڈG�tm"O�	b� ���N_�$~rR���:yk���$^�=���Tv��@<_ ���M!0�F���8��{J��F[�D�n��k���w�����2g�(�6��
����j�7���x"Qߠc�fW����H����F�/��={2Z!�Xs�g	[B�w���ó!��>��lv� �&�ݹ�2�l�GWu��Pc�p�_�)�֐��b�߃0�Ѽ�D���J�ĸ�5�f�fB�,�J����W�ٮ(4�L�P�ӥ`�
CB��'Q���k����་��"��e�������f��*SQh����ꄊ��#O<�m���n+K�4�u��c[�B�ެ�a̎�F��]��E�er�������p�ڂ�y����w�f2�Q8������~�����0�2< �H)k.��<u�7I�;:wI_������g�����:�%�t܍��dH.^>Xbm_+_�jB_�c�IN���U�Dޛ��ü�]:��7aS�3��lm�k��yZB�m:��4i�����S1�3�c'��<�3&�b,��WK��������3� �����;{P�d�,�b+2T�p���U0:��[���j��i��{����B�C�"�[�T�0ώ�rQ_qYԄ�����:v�_w1�X�?F���g�D����O���8=���.e
1>��sD�Syԓ`s(��"
;���ԩR�2�����aT��6I����9^��t��82ܳﶀ	�<_�H&Q�L V�ܞ��1�������
��K{k���2z����1�c�Ҳף((�Gz]=jB�#�$m������o:��ZΊ{A-A�~��v�t��]-�=��=8A���hN�媉�J4�6�� �'J�W[bt���\�}�/�/V/y��A`�V��n�)'mĻ�[SA�(�L����TC�|F�X�ݍ�ph��I���!�S|5z҄(�qѪk��`��G���|���8l"�-A	���0���}�$� ����ϑ�&ޤ�YѴ����h��2Χ?����?����(�m�Y��%��07Z�(�}%z+}�#��<�޹�+۽��Z��x�(/Ϥ`&�gj��簡˞B!f��عJ�F��.����2�w���8B��vkg��k9�	�^*�G�-o�������v�a�;�hp�D��y��$V(��
G�٩>B
������$M�}ZvB����y�@RM�2u�O��7��������O�{R���|�r�44���;�"8jo�<�EvX�	/��ՁU���1��޶�L�*Q��F�J("�����k�*�7�=�i�����o�u/�b���Й�O����vF�Y�mf�!1�Jn�?p)d��KƵ���1v晇
�Z�������)�v3q�C�	������k�ES��g�;�Fj�s��`����]h,ds�Z���xȩG�'��/�Q�q$��e�-���Qµ���a+;'��郬�k��+p	1mL�]��� ���e�Kɔ��~]�|�k��ZՄ�iL�-�aT�O!�eG�h��*j�]��6���^�S&����-o�X��"'�K9����G�&	\˱�Vc��j�����c7~iZ1Y�QI���� �X�2��e�Ą����`�8���~���,�Z3�!����x�g��ӻ������B߁����dF���Ֆ�zBy���h�5�?"�ZsL���fK�1��݀����c��8羥�g����濩:o)R|׆���}�+_a<C���W"�b������uv��p꓀��w!jQ�B��X�<�r�4�K^���S&�c~��<@���b���q $8��m���sp��wE\v݌����)'�B���X9'Kp����Pc�('D!n>�3��CV�CE�iA��������w;#w��'�����J�OtMGTk8�
R�=�o��{$r|�(R�@����|f�v%�ь�[�Ɛ"V%r��=�i�
� ͛"��J!Yc1�[�nq�'CS�G��;3@]�Ȏc����?L�e"0�x6�A����?�0��48���Z �K8����|?�p1�F)��������nz`�ֹ<J9�
`�b��P�'6�ɠ.I_�5�:�J,+�5:r�=,$3�L��CEȿ7`�q�I��1���}���+�u��M	'���^���*��j��2����H�d�剒4�b!��= `mo� ������<�Pʰg�DP���J�TEY��Ie���ɣ]��ԳL��Nד� t��&7nN���]�̖w-����J��!,[�~����*�"4�qA3� �����"L��RQ����8:�Ԟ��Ok�7��c�����:���!��`)a��t�o[P���PTu�4�Aiy�5�_�49��=.��]Z+s�A~�������F��D��d8�.�m���~������u_cOH�}1
�?�(�]r���"��=~H��-���L�H���
�]�z�-��(��r�]-�%���^�n{y��gLL���� 6а\6)��|������E3�Bg��3o�u��[v�!��_���v%�z^�r�J	���\@��
2�}/��/��N�y�}����s����Q��r��Ӧ��
z�'�����xb�����(����?��n|<��x�Y����W������U g>�u�$yg ҟ��Ys'�;[�� �\��&gje�L��T[�ST�X���sR�54n[������m��LJVR]���P�,r�,�ե_������K4����i�8���ZH��9ّ�4m���r�ʙ��ڴ<�a�^�t,}���Jҝ|3z���w�1���Q�[߲܂��wm��sr('�����'_�zXg-b��5L{��:�c�u�t��F0g�x��0�.8[��������t�I�5��zՓ��F�^l�h|�-��Z��[�S�f9��%����x����'�����Z�q��ǁ/�ww�I���a��R��!���K����%GD����3�c�<*�h���@$��H�(����9���d�E��6��;�`+�M�aж`c��Ľ��W�Nē�oZ,�6�[���0���FP��!�Y�c�N�/b/���+�q��x�aF�fW�?͡�VrY��R�C�(匊(IZ��W�K�\/�� ��#X��4�d��\��3����|Z�}���=���5An�H\��
.l���@��#H��a�a�4p`1��{�;5e�Þe�i�y�͍vb�0��H��`}?�R�PW��k��n���c��������j� X� w,e�r0<��i�
jh*8�'���}�`��4�HF���BTKib���(� Mw�f���dV!�n���7`I��ǹ�
��4��K��-��e1��� '�@�A*���顬�]'�W.���֝sf�<G�m�] �p�t�0���D3V2p3L`�f�g �\��ϐ�M��>1���1Xn�O.s��G�Ě����Ko@x�bZ���#kg��Zz�Q�>Q� Fi���_-�P��颪4@��\[G��CbR�9�wm9Y�*�O�:��	�)e֞�]�F[��;g����������i�q��xtu>aW�J�,��Оv�����,�n`�+����3^v�j��T�W���ߵ�6����(���#|4Tu���x
blm*�ŗW�^2��mqN7B�l�W����I;���y�?�#C�a�"2��Ř�#N40h(�U����r�M��04I�&J�ݝ�sm�1�4�q	zEC�8zm���"_����Y`����~�����k�Z�_X�������qT�	{�40wPZ��ј�,iʅX�x4��
E��aW�o��Q���q��~�ڷW�����7u|z�x�S؎/�K�/�i1¥���NDsY�ů��l.���1M6���7[sD�'��3|3�YG�}7���Վ����Pl A��C�*�m.���R��/� >[\ �T����2�����ibb*�A�K�qh�)��-����Ś�,ZM�~��K?|J2��oUଜ~�<�Ip�$$uA��g�N��S��i6��C���|o�Ҷ�zW��RRfRI�ڒ��$ E�[X�	��W4������s���p�^ζZqνfs\�P��&ρ�Mb�~�u�w�Ls��(V�R{lj{���;d@�����d��[��-MYTI,ib���à�%��L�f�ж����`�f刏ȸ�RT��~����6� �;,�U���>S����	�9>÷��^rĝXx҄�R����n��\���>
;�|@�'@�b���%A7��=s'
�,��p����=l�(\�0caI�SB֣1�^H���u�'TTeۺ�J%	4f�mj�� ��L����Kg�a��N7!i%�&]Ԋ���zZ��[�5�9�>O|Y��z�`*�%w����4r����5��VwU�Ě�a3��)/�5t1�ˢ�W�@
]pԑ���ZO�]m]���K�4䙉�|��D���!귁���(x�����Ю|u�Ky{,�<���xF��ȓ}ں�W��,�.���4��4����z5��H��7�[$��@B|.Qk���{E�)�D�[���>[=Z"Fߟf+���I�}��$[��n�P�JsBp/B���FA��/�	��9�K�9=S�M+"��D��m4��*`�$�/�0h4S�MTF:j.P��	���6)�����2�kxg��kB�ʤ(Mun���3)z��c��$�4�@B��ɭ�y}(�~F=�g�.�-pK+'��N^
t⨖s�% 
�Q�އOs�@�_�n���S�2��Q���Ravh�ê�j|`ǚ &�:�z��K�s���6��(�0C %߼R�����Vj�DH�������ɡ3O�o�m�偩�$�A�����R++FD����s��HF*�}��)��`�>����34C����u��]|�]������țD���ѐ�]�_E����N.�xX�ƞ ., {�d�ڀP@�O��PvRgbf��|�b@�|���-Z��O��y/T��L[�S@�\����jKf|����%������؅x�)$��j�:�����9��[tK=7��"yk8��2M�x��aq�;�:�M�ܒ�`@�����9Z(�@t>g��_�]*�܅����ܴ	d����J�a�]�U|B�K�(~ nj@�<>]h�H{RAZ�
U�,� r{��@s$^�b����ا��A�of$l� \�U�]yV�|;�"д��Npd5�� /D�B��E�]8��.�z�3۸���f�s�!����"���N�v���1���TxQ��1���SP�@��$�_�ah �׍���⾨���_�^��+�V%$���]V�γ6uz�]N�6}@8�{(b����&����/"�
�����D�܌�� lp�3��;$S�d��M�0�g��˹r�B�)��f3���v���cg���1ߡy�F�|���̬��'��B�944q��������|U���ln�Az�&��3)�qg<à��j
yxS�q&B/RV'>��j��)A���c�������C&p��n/�������(�c���@� �z�>��g��Ky���
@<�+�Ϝ� �<ծ��/aW�;�w[�Qt����j<��pIl��": 9�I#VVE)���ĥ�,(���JL���j*y딑W�ӭ��q[��䙵c7�u��`�툖ؓ��K��M2S|��1�i�����K������uB�ӏ��tſ�l�LM�!����(��i�s�f�q��Cta	f���Ga��H�c��|v$D>5�/���^�8��^� [x��64��ρ?��T\��h��P�1+[������&��[�d��ǭgz�C��_��kf�㳐�m�af�R�����d�}��2��xbD��#���I�\����ZԨ�Q2�do����Fk�Xv�#D�¡.$#���b&�C�#�����>���B�Y�1ضN�ʽx!��7��y���#��R�g"�i#�( ��-
㰡��f�Q9��l܀9�"�+��^�;�R��D����D��l殫~^���������k7Y�f�Sz����+n­��1ʿ���/��CW��ӓՒ��9��kH+��܎����r�9�$���a#f�)����̧�Y.�Vr��&`�f�w2(2�&2%�Ɲ��9��'#�E��\3mV�	��E,F�,R�Ea`�s�;ϑ,_/���Uj,�2G5>�[����(�d�����]�iV�m�Cb+��1��<:�X��QK���:,���	�7�A���h���GL]��`|/�<>��\eg����<t?E��ӑ���^��Yݟ�?��	1~oY

�r��YxǢA$o�a��c׾bI�k`�'Q`7?k���P�}nK�l�0M���q�7�U^�3���FvG�'�[l�B�����*y��.�9u8���6ŗ���_��p
��5#�q���ĭ,f�x�����˻�A�<?n����n�WIjPтɷ�ctή���U`��'��Q��㒭���2h���
�ѿ/�'Q�Ix|�*�p5��*:W������\q�;(�R����V�V���h��e���,QtlC>o1L��wE��D��2������H�	���:(R��UfTUvV�y0�l��I'F�g2��n�5Q:�S��^4�p�ϒ��j���{��ε-Q�.�h��Պ��8��j��m���P>�&N�m�w�V�ٺj��2���?>�}¶6A3۵J{ pn���r=���%��XG�.�[4:��4r��#k��3�(�݄Ǯ�7F}6�F`/W����Gi)��i=�룻�������������(���.++����j���;Su���?�ɜOQ��u]�Ks�^QP(K��YɥLR�2��I�۩0@�r�9E"l��1C��Z1à�����G#T���.�Y�[�^@���:9*K��Ll)��*	3�?*&m�,��(��L�y�:ŧ�r����pG@�do:F����WiU��[%	M}�y��0�h����_xr�/��k�d�c5�q(��9 �"wF`���q$��p��1t�������5h`'��+�Dk����L\����T���`|�_!���*R�ٗ���z~OkDvE[��	���-`�54�y�)z��XmrM*�{L�L�b���� ؜�����������ʾ.�kzq��<*��0�Pg���s�@��O�&��a1��p&�Q %�U�/V��O|B#0�g��r�)�|��̜�
&:��;����5������~�*�n o8�^�F���'�Us��w]�>�G`T���8�Y��,�_�P�C7�#�$]�fv7e�H�ܐq�IPї �V������� �#�v��q��v?q`�TB6ݲӽ�>���fp�;�l�󬧒��.� 5q�n/��}��~��N� �.F�{�d�Ϣ���?n�)���� �~��i�bQ���u-s�]<��_�xص>9V�^�?~����I��C!ƴ���p����sJވ��b̋� $GUׄ�P]Lժ��%�+��EȀ����Aߊ8�n��}����eaO�Q��7~A���g���义"�.��1(lmq�S�ԑ�Q�B�!M08
�_����&���M"������Z��Ij��e�2CGRޛp��V�����k �_7��``ې��%���0U�Z� =|��m<��V�u�^ ���G�QN���%�vڅ����,V�H.]'#{/+=��5ɿ���}ˠ3�s({������� �j�J�	Z�`@[?f\�,K���:�`fV�euܽ��\�Z6,�i��2K�3��ET�K<�֤Y��q�0�ޠ�}w('���f�)�N�2?s!������i|JI2�t6t<$.�χBs˂Xm��mh{)\��k�״(���E�/�G��ٷ��2}�=�o��o�V<��jV�䔆�p�ke.s��a��>Mх:v�z���+wD}��z��]� s�X��N���#B���(�TU^blm�
�����y)c��o���r3�Қ��NB�U��gjb9;6?�Pk�vq��q�)�<�����k'������U�̰�E?��x�S&�>�^?�h�F�{�{v�d������YLM�]z�� ��\h�]�F�RI��xr{�ܓ��wj�j���Btw���L(:	P��h��OB�I�\�Ǖj,{�թR�@�E��k\����	C
k>���d`�З{�5�N5l�������i--��z�Bb���hT��M���PtDE����}N��=��ɲe��a����/Nnt��nff&X��.:���r�nn�/{2��0B�O���"9is�iIe,�}��C0�X��Q��c_O�v��+�����`)���Ф_��A^�����yS�tr,�/��IS��4Ut���w|_��ɋ%6R�[��Ed6E'yJ�K);�3��Qz�D|�٠m�O �H��8m��H��z�U�l��Qc���	��=(0��n��$B���d�5[��7��ިZ��(�a2 u�z]�>0"o���3�R���_�ó#!����vyp�K1���[�1���4ۑ�Gꃦ��d��'ݠ��~^�ƌ�<�Oe�b�����(�ٗ�,�1hG�ުE�}Gf���޹
X=c���NL���,|�|g�.�zj�$���
n�&X@E���}y�\{�����3KU����VD�^s#��,��(����h&B9Sq
�t�c�+�P� �1��+Ԗ��P\u;��x�C�O��U��DC�+'�	b��KLE�x�9ZS���\���wR�Y���m\�o��Tv�8q���w�g�"��H����7��N�{H�1�!=wQ��7-�EW���� "��N��?SVY��������:g�=)h5��o�����m�|	�^�~��=��Z0��?>��H�ʛ<�n6Ib(�v6�xP�\�L�ј7X/���Du�2Xj��o��1�$�[�/�f.B�?m@�-渉jd�y(� tY:�j ����⇯��Qd�L��(�ems�*�z�����z�j`1@	�#�zq��/��|Z ꏕ�qY92S9�-p*� hjt�d%���<-��
n(a���nK#y�%l��5J{�Z%ۿƑ+�G�8���4�$�*<���.�:P i�Sk|�j��ɞZ�$@UR����M��f�=�{;S]�I�@lu�^�=랥k��Z�\��ٴ}����o����m���Px�Y��nX@����r���i���#/�a�	a�5[��,�v62���4w�!�gVo���뮐b7>�̀v?:�S-�@��@�>04!����F��L�&�|�A�,V$�W�K&G0���9}��S�/�?)��'�l����:^?��v���:u��|J���~2o�Aㇿ�N�t�4Gt|�ӗ�8��p�{�se��ݯ���nc6(��z?ǌ��%��-���9N>H���u�Fh��.��O�^������{��EO)H��ӎ��ɺ��qH�� �S��]?���x��T�ډV�Ii�m�$G��h�kܤr��,Sa6���B)p,+���_��
j½�p#�oM���kͮ�Poy�g�@����L�hG~��=
P#�A�{��}���{� b�dI�K�n>�Ī���<-����yY.�<�� ����ѥ��v�� ۦ�cGd�����v0/�,���͚i��&����]�@)����B8p����E8�`��i��I�)Nb�8��ۮ��>,�h�uj�8R&X�tr��\eu��7���e�~�`�m>D����Hj����w��^��<�����?ꊧ��Mx��*���@Hy���N
 �Oj,���=�M"6M�:��,��e�k���<���|�_h6jv�V���~�i����mjd�6hE��z��e/4�n��t���bYX0���Ƽ��H�K��9x��ϵ��7�dN͊�iD�K7��Db���!Y|���K;�D�u?�Ӻeo�@<��r
���O3��f����Y�\��?*��{ǉBU���_��`p�6���^�"s7Ny�/�3tn[iB:���W��t�*`�'�6�T���>jhv1�4�JGv�^14��$�2�,'���8[B�b��"ԡԄ�V�e>��? c�&  ��2˱��%8��a���_�u8��fUz�'�m���E
�O�Cy�$n�n���[�X�P?�Ή:qlN��C\
:��^nx�Ł�/�M@x��Y*'���V�	�(��?���ݲ�Qj���ͣ4Ә�\�~�A�\ɶ{��To*Aǡ�����N"xd0�~�ӻ���*�i�(U;Ot���ʂ�M���x�d�Puh
���(��gnL�c�E�$�6�ى��x�_�����q��3a�˼�.|8[s`�5dQ"
u���������P{oJG�ĸ9p|x�_�21B1�	�J4���î-�T��=�ʋW��]�5���%�NwXLBǆ#��+����y#t6�[ql������/��|��H8�D��GkXxC�u|�����<�HPsi!
A��6��G��g�v���W�P�m��"��j�r52kr6���b��\[F�����h7��#vCA��o9+z� �+�ΌU���2�D�\�r ��]:�!rƞ�$k��]0:�'����z�;l�y�&l�Q!�4I�vD��h�?m��"����[=a�^y�{��'4�nx�лi�=����q��u4#�d䇅۠`	�a	v���~�G�!��������f~�a�l��r]���-�~��\y�v��#z������bj�E$�Uя�c
&Őc�+��0�q]�F�.���Ԋ~p� �<���%�G[�dA"�dy�:��R�yM�opu���]��� x���1|�|M4�̟\Eupr�6^o �� ��lkuٹ��?�����,؎Q���kݑȶ��%ia2���D��y��x
�L�w��eukͲ�WgJ;G�c�Ұ��Ў��^D�8`��'5G���O��g�=y;d�Ԗ�i
^'b5����6L�,��W�a���uT�v0�f��%ie@�h�%`�=��̹��fm\ ��p�,q�x��f��4�n�@�l��A�`�4{
Y�X��MW����
���社��:2�G��a�Y��h�ֆ	
.2~���yۺP���,,��8�dw�i��N����a���|�p�#�Q��o�[��a?�V��$b�J��ļ��[���;�ye�ܣ�����)4����o�(���A5��Zb�);Gc�{dF�� )��X��I��ʧ�
M�˖���^�������z1")�;v� :�l���J�pn�T�K$#^�Ʌ7��Y���'k���"^/�Jt0T�D#�H_�ٻ=D����zD��&"֏���
��}���p�><\�3�|��Ёlȧ�*����TFV���(�.�+u��ID���N��Nɢ{g�X8bg'��&`.l;�n?T�?q�L�ۙ�.��o�Jb���E~�S;W)�ɻ|oN��l��(M�?�ϊx@��2�3o!����O!��Ъ8����b��/��o熾���ܷ\�QB�8 Qq6�Kv(��J7� @�\���#ѽ��b�e�I��bG;
�zsgA��<pt{���6�H�du�Z��jBA���X�A�N�|~-K}����w��tOT�!��cg�Hz��ᄷ�r�,^7�E��w�W~�+e���)�źwP�f?����Ɖ�eG��M�*\�D���Z	��(�&~�۫�H�@4��L%͐�i���t�#=��k��=b6��:��th���<t�3��j�&I�d�����2��&��nNպ���?`�Ѕ�z��;�.�N���֨���Q5h;��H�¾g����'$+��p^ ����7� �m�P2���o�W�ÕS/@^n'�a����L����1ܲ 3���(XHϬI$Q�QZ�vf����,L7x�z��4#᥅����8��b����c1�ng%�Ĺ���̦YhZy�:5���2萐�5���� �Pش�5��is��V��6Wh��aq��,���Rb,����q�S�T�������ֺ�PK�J~� >�7Mc=�&�h5�3}�����\����cl���c�����(�2$��MO+ m��D�H�f�Ѻ��s�BZz��6�p�$�v����T
�'��[�8��R�E��-�ۤ��N�<��/D5��<=ɘ:���6K+Ā}*Й���x(�a���⷏�~+ݤr��\m a�OT��� �/=2��n�D%$�؂�Zz�>y�z�Դ��Y3t�/՗��2���m��F1~)3�˕}U*�~�p�� �fw��z 3r�Y�kc7�bk�gl�u���7�ٜl%c[�b�?�1�e�%�o�X���u"8ܾ�����nBy�Ԇ-��Rv֙����~��0�0l�Y�귯:'�;�xà���f[-?�`<SB�Cq]�C�_V��Zɤ�͛��Ϛ�Í��S����e� O::�xh��G�Xh�2��Ȍӵ�1	ٞ!"N�Cx�G���z��+QX�}"#PElP ���X��2��5jw I�{g�:���UٹI?#8�(y�p�uZњF�C�d�x��W�|�����xu��C���c�>���2�����v���������_��������YHq�|3��Ʈ5���9k��A�C芲���׳�_C�f�{at���vm=�V�X��;��S��!�2/�Y�H�k��b=W�m��\���6.�;����n�mi2��<R�h��>�=��D���Ğ�����3w�;km�>RiݽR+�8�x$�Ս&�����-�q�]�vU7x=���@N����nH�
ꁈu�)L���(Ok��TCϥ&9�Q-,�a�ho=L��h�O�
�8嗹�\(���^�j0�%UQ`v^�U�b��Zj>sE��5A��.�5Ҁ�|"����҈ϙ	1F9���X߭l��GO��K7g(���S �~�$wgW@�-E��,��Q�p�{�G���֞}~)���{%���ȉ�ȟ	��d>>�뽲����Vx�GVMi���g�������~���ţ�Vf=+��lg���/6�.@���l�=��RQPc�0�%,�/ުW�����6ĭt��$�L��c3�y�D��)�j����t����0�[w�ͨq��AN'�u��/�k�t�Nǋz�Q���	&k��w�c$�g���5Β8�A�m��}܆:\�ä�z�(>��n��]�ͳ��,IH�,6��B(Z��l�����R)�k����}>�x�'�p�?5�w'?~d+a�����C�+"61��R�J��p������}�ã���������8�؋���ޯR?���љh�/�R���(�a~F��w�gm����U��I�|�Tb�郐���~�n�g&�)�X�����O��)��9Q��*S�&^�	�.*�}�:�.�x�Lj��-�����v����/1\і����L��ƙm��ϟ�&!r`�4��A;9��-$����&����l����h�㪿�Q�Y�2�嵺]�+��Pr�q����c�'a;�֏����i<���t�����3�����+��<��I�tY����%�)v�N�.0�Q* �Y��w��U?��'gk��	��~�(���sx���z$�o�q��:�$������9�S�����)07�D��))���U:��`���h�*G%���uB�Ɔ�t��x?�X��._�r���
Hs� ����V#����g��u��j�lВ�r6�h���!sw�/ɲ�(�@:�����>?��}�t�V��H�ޥ�����-P�&5mX%$z�D^Z9�@�R���z�� �?�'����|����'۞5)@�h/����<Oj&iIUj?,{��Gê\���u����iK��]7����#��>]���"�[��Q��Ӈ�����GD���kE�FM���g��K{YBy�2pk�_4Ib�Bҥ,e��#�F1�tD6^�|�%k��V�\��y/*���:���(�Aͫcb�rE�\�U��ؚx��c*r��}k#,[�h���>X�S)Ir���Qj���I'w�bK��8u��f�.���B���Ja���^��'T��z�A<�}���"CP�\k�Lox�
Í�Jzӽ��9������F���hG~��ӗ�����{>0��]���!/��hp%��A�7CNm^�0e���[ǵˌM�"�q��;�ۑ,*	����Qu_n9��^�<��KY�j#��?�u�;rNU��Eg�T,�Ze�,ͻV�%Ӳ6Q�ݮ��{�`�n&%Jb�5�9#�o��{��t6�|
���8��y'���7�&§��8��f(���G����Q�bz�Ǯ{]���Fk���l#�R��/������I�̒m��OCFa�3ט���n1+���G�ט'���R�Q�����ꛗߖ�'��O�G��RiD"�����c�x�=�8T3�����-)#E��
���P朾{C�S�yv�@4]{��IβA�䓻C���x������E&��I��C-�eb���G^Jk�vʞ�͍�Sf,��M�o~���T��KG�M��J?�Zk�$�J�]N�zO��mf�Y���满�"���{�Y>����\}qA��� oG(�W��n�{�r M�GϤ��6�ư��K����&T�m01���,qd����l�X�@c\���|<h�0�@�M�>�gA�>j�������=@T'����Rx8>&����F�� rW��
v%�I�Q�����!J�:��9D�T��$�����1���^^��5��P�T�q��*���{�e)q�7Q����{1&���B1�p�R����^d�lx�L�t�lb�����K;S��v��c��;���u̝�D�� 2�uY��VJwR	i�*~�F�Y��}��ز?O�[��J����/�5��%���"D�Z�GaG�NFx]�x ���M���̛�`�֘
����e
��]PP�&��O�h���pw�g���9�@\�	�m$��U�=�&(_F��"�:�I `�"�t��H[������s��DE�f�3�݉��@p�g�O��$�9)2��^w袰:�ʛx-�V� @�]q2����Q����ӔH�ô�!�ʢ-ٖ���	2Cs�xe֯M�ټK�ݺ3�׌:��D/|�%�N#PI=����$�1���3����pfPD=��W��t�JX�����L�n;�h���	>����\�0E�(���s��ֈc8I���O��`�O��?�>_� �_���ݿg֤��|LF+��v��I'�A�D�9B�Gx۱��m��%v���ߦz2�
7�:�N�'��]�ao��>��8z�[ek��a��>"����^�Q�?V�Ny���a�
��!�=Vj��W5f��}���=r`nI��i���������o0۬�1�r�dJ���-X˱\(��-�
鄋lm��0K��^s~�Fp����"O���U� ��"Z�([�uf������Ed�l��_X��.?�g�����:1eѝW�UM�2f7��-��L���Z�L��T�YxR��Cs l��ߗ��}ju�ѡejV8y�_V�h�Pr�2:
�)u�V�Y�V�i��Kэ����x7~R�&�0�����Z��'l�v	f�5~�G!M��`B�O[�k����ڄ���j����sS�!����z
�>�>��{7k�J��If�mQՕ�Q<5ҕ�Pl���!�HW�v���]xw���V}ћ%������R}#�� Qa�(��}���'���9�[�%��4�3,�ꀨ��m��l�v��q8�V���t8LG�a��˓K#7B�$Z�����--�s��*�{Ӑc���NI~n��=�}QO�b�R�B�]trZ�����~��n�AB]X� ��}W��f"�`��[�{	¬,���%�W􃕁Y��ư�I� ��)x��,^���w���֏6��YuKd�Ȁ�X|�m798LDP�]��/y�6q�wv��$��O2$-��T8#ci��^����F��V]�ڝ��(�0ԥ��C�Q/��)��?c�U q)ɚ��v ;�>�m��jN���o+_��uA�J���g aN�0��c�ݒ��v�����KG�j@ܦ���z�~*�c@��V�q�]�K/��	�s]%�P//��hm0�|�$&i��n��'�e�C3����7�m���Q��Z���V&��C ���yx�y����OC�w�n\J#�#_XDq�E.���8{���/����D��Eb1�^�SQ6t�(��+Jb��%���������8���'w�?�@z
�^&�����,����r����1�M�8EY����� ���W��d5r�ƒA�21%��+Pw��*��D���
W�;��~j�
�}p�R����;����Y��!���NjR�
�f��{���(���{��!ͮtոd�T��0��>Y$-OY!�`E�i�@��k��S&��(2�R���Q�W���U�@l���=H��L2S�r�����Ex.���/<�z�L#F���ʱ�ԗ�>&:HI�TE&�eB����wj12�^���e���g$}Q'�����c�n;���*	
���<��o�&�Ƌ��FY��%g�1��R���x��������E�t�1��:���`�y��x��P�ǥH���}~f�X���sC�9����y�T�������r~}9�=v��ه���oLb�j�)�?��2�����'�=.�I�ڜ	v�<[�GÎo�F��O����M?6���s�Z�;�'�z�ַ+,Now^���\'�h1��w�< �U�h�U��&��a���?��%�[��w��Q;����o�<�0�LT s� Q�j�/�S��1䦡!wBqm�-TIe��'!d*�!y%Zݗ)��[2�2�|!��؂R��3ő*U^���޸뷆��C}sf����s:�sC0R��Ĝ*��]<f{�����f"C&�UA$�#Xn�2l-@r��jG��,���l���Z�H���r`�!$��5k��;�B��U�1��]���H�8XRC�/:��QbÑ��)�G�q=��[�8�j�VQ#�:���kd�n��^��bۛ�� ,t'ZN��m>�<�C����ڟI϶����~���TM�͇�Чɬ16���o�p�g{��^ǽKF �f4���������<�:mT�0L���J���r����	N@a��]p��ƛ��e�:']5��ù����)WM��=�fk3��c�L�ق*Wo���F3����&|�q���A�D��H���%�),����TTz��HCh�=[ѽEܓ�R��_� ��+�9i18��=��
�	�qC�$d�����n�sc��(��4�D��³�pD���*G�/�?����o*�B�ܽ��1+�ܢsA9��;�#�jDI-w��Zv�q�S0������
��?��}���ζ����?$ނ�OAj�qSlر�H��u�6��g��;�9��S/��X$G&/��>�r�\�c��!�4%��`�&,���4=��[�SCM�`ܦB)�DP%!g��a����h����-p�H������ȫ�{� ���ˆu����D2T,��H+:6��S�9N����fn���,
����:L%�K��22����ܷf�V[��k��V��-r��xG����X{"B�t��u���^Boa��1��dc����*�V�%y.�A����T?g~�G:��� _��fY�D��$h��~@k-�H���
j��]�������r�hy6����PY}���Xb�R�g�B�?<�>O��!(��ז.��c�t��/e������}$��M�M�r�<ޣI#�v,�_��1��=��.�,bl`BV�v�������!(�*9q���)�s�F�p�� �J�dp��E!��6=2��p�F���QR-Z�p% ��X� ���7wFי3�e��I�ʃ���.�LN
4��J�  [}�ۊ�k��s�TkO�S2@o@���n��������0��H��6!(>l���3���z��Q�������n��z��u5�i��f"qxle�2�0��GC8e�go��@���0u(Fq��,GJ�EZ]��u�	O���fXO3�g�|G����b�F�I��E�iE���yC�mn��o���� ������� GB�yۓV�b h��"h�l�8B�KUk�v6"vEPwF`�,׫��5:�/���ֺ�0�F�"��!xP��	�}1]��sgiV�������|���x&�Yq�y�;�`�@�:�,��s˒��A��=��";�*1�`���"��ߔB�V=�|o$���dDQZe�%��H��`�a�3�_��5+�b
�K��&_�;)x�;�G&�	�%@��z�ٴX�j�G����b�	Y�;�P�̅��=T�~kO%�,��.��8��ɹ�ț؞����ݜ�QA�g[�Ŝ��3R�Q�0D�Y*��)�oP�/ϫJK�x�m'��e�⍶�IJw)�X%f�`J���+z_Шe�5p�dC��]���1di۩FĶ2��'�ۺ;�����U]�O�$଒�^��e4!SUQ��`�mz��Cԕ
��"�<�z�=B�w�[��;��י�&���c����<���	�����e`8 s
���rz����7S��@9�Z�U��͆j�p�9:k�꼊�� ���bY� �+g(r]dٕg��L��aAz�+s�)�f�ësZ��5�`�oBk�T#�^�<#q��%���{4D|CE�aj�㄃+��9Q?�Z�5l����P]m@�o��U6#�ɵ�e��۪��l3�N�>�4�rY��}u���>����+�]�mH���jc"ā*���U�i���Q�M��ߡ�(f2L�e�PЉ���=W���(�hܒE|\"�����*G	~e�<v��L�]���zócoG-I��:_R��"�WgK
���P28��-~�����Ur!Ǚ_���'Z����=I�M�?!������nۉ�<te��إy�.��`Ƅ-v­�<�e���}X2f���9�+D�1��B3-GI�w�˳�+�w��G�p��|�XL�o`��5w� ��UQ�+Ȯ�����>��f�{�$+��Ȼ��<��:���ˆ*�b=aV��̽�'Ha��Jn���!���$b�&���:���2Ɇ����at�R�~l = ��7$�)�� �_��K!�ɆD�|��M8]��&�#I����W��ҝĂ�-"5�0��Q�������������&ril`0���x����=�R����� Y�Xf�-\v�TWxm�\�.��*/y�!n��m�b3Y~�2�� �-po�l�7�G�����$���e�@0%�CQHN��h8zzu�=�ξ���R'|�
��-�ot�9�����1��æ�9OX�$�i�1�>ದ�_2�0=��d�F�A�iz�%���C��.�a��Y�H��Az���zjT���F��2�1�4���:�{*�hr6W~�˾$��Zs�RD}�����5�c�р褗�ˋ�=�O��ߜY�o_^�h�0��ù|7b_a��t?o�+<�Á�U���jh���@\�*�b�گ֦B�%-�DD�X��m��=��z�;z�$.����s:h����g��ކn]+�/=�#�Z�~�H�-m��W�:�X�[��BZ�a�s�0v����W������M��r�0
��i��LtHu �7#��;qH)-��I-�l������bP�mR�>����Vd���~��#�5m���us�+���6�����eb\4�yf?Z�)R�t<���[���k��Q�e>�=�RP!��$�7S2�ۡ�	woz�|v��E
�p���1#���j� �OΨ\������
��mSP'�c�U�V��=;G�G������~W���L]Մw\��|� X�O�?O�l��w�7'���ĝ�s���]Fv�?�"����v�~��;EM�����ӱ�W�)!3�cd��&HN������W���Q`�F���b�d�F����[����%Q���e:��@���F�}�/8���9��֛�+bũ
CD
ۼh M���7>x��=���]�'8n'S�/_�ų[p����7`�<Iiy����L�(��Sw�L�n�!�4��}\G�j�>��8�������O,~秾�5^ψ:hc�2\��Ja'�-T�r?����%��G���S=cc/>�T�c��'���wY��\F}��e~���+������Ω&��	�Gs�2x�(�c�����h��l�0�g��6�%��7E���A��׶�{�=h�b:Z�&���b<|5�D�����>���'��iX�Y���`�2F�cr�]i�wʝ�zb�5ʚ
�kv�{�+i��j8��4�o�]Q�X��%;q*���t�ds1�w�#rʎ�w"�ᩮ5�p ������⊠Z��U��(�+���t�S �O�~�,�M,���;W��:͸��/4"���KfA_��/:�nlbP|D��wD�W$*K`�<�۟�,��p$g���UC�\+T�鳡ް��� ?���̬VO��SAO�>�0��>���e�<G �p�?����^���׼ߺ����/t9��J��\\��)&DZFG��v(��)7%�Բ�A�U�A݇�9zG��x�����6~$gM6�
��@���HWw�Ͼb��.�@����.ɨ��Xz�~�KL�Q�,����>"�p;�I�-% j�	(�}QN�'�1��hB9�W��U����b���ZvL�P��"��y�� hY{!�`T_CN$l��D��mN�(ڲ?��OO�('�{�1��26�D���n�.����I��;��<)|T-�>vl\�>܉�}I�y�t��t��8��A�:�%��aO�+�-TT�P �ѓz]�jMFqt�@;���]�����^�Qa+~�H��s�E�i�����[`,�����N(�M���3Sa�^KFm�����&�h>R�R��"�e�1eJHB���Ù���o�H�;%�(��$at9>_1�:~��gB�>�� ΂f��q��j���<o�\�����S����@fCi�棯�p�Mޏ�O������9�T���S<ߋ�@+��Y~���#���@le��7[_>�_�5^휃��i]�v>�	�O*�W���C��u4��ۘ�h�J#&�xZOm��[�ߣ��H��O<���x��W�����"vw�0���̓�ds�J�P�-J���|��e�||}E;d���Y.���i��l=馊�D���U���� �ódV�
�$$O�[�,ޟh?���'4�42z
��2��HI�=���U:�������RA�x�N�@��=	���G��y5�L�2H�<dМ=�/��q�0^j:���$	3�rY~��n�F�U��l�W���G`�k�r�U�>L�)��:�;� 5�}EG��QC�A��,�Î.ƾ����V.{њ{x��'�OxAn)�W\XeI[���:I�� D�N�ҭPc���(��$Ԙ��Y�U��=����۸H 	l�賫����5P���\�OG��Vk!��5g���������5�\z'���蓝����eZyh�/�*��j�( ��ۜ�}����=��`��FXUtޅ_�Q!=� � wSA�M- �U�=1ܻ�N{����+�ճ�4b�q�e�Q�p%�_,sLA��=1���M�s��X�j�����؟A�p���龐��Q[J���C`��=���F��1��T��S*�'1�d�*��z�JН.[E��o��2z��arj[�YL\I���8u�u�ݯzϿݽ����~���ܟ�'=�u��L�'���r�kJyٌ#��Um��#���c.G�ϕΎ��b]�#)tQ�#nI��V&��:>J���z�2�T�L�KJ�*T� Wj�>0~�K����6�2��w趇�X�@N��Z����Z�d�e�/��<����CpJ�0�e��3�_���ŧ�̎y��)-8[���;)֞%��l$��&<�e�6Q@}z
u�Л�{�"��T'�j��΍_�����X2��S�+s>"ƟA��vӫ+��Yc�^0
���ؾz\Q11ۣ��7_�������+-	*�@�vl�Gk�Geam5��^�u����.�Ɗ�"�1�c��[L=,OH��H�
QFw���?L�>?����%R� �n�M����\���K�۠��fl.N֖ň)�����f�*O����Š�O�;�rەn �)~M]�_߀k�x�r5�6�` ��.��>�r-�5���p��x�*������^�,j�����t�j\�_A㯳�T� 	Z��!�T?�	�puU�!� �Q"�hB��J�P(���1����c�E-�x�jx��M`̀:���94�vD�CTy&�o���G���n�L����Ы}���z)���+���~A/e�����a�q�b=}�jF.�^�q�T�׌�iI/���B&;�eP3&�n��ܲW��R'B��l�W)񟖯25����$g�� w>��'${:{!Mh�J:�׉�t`��(�Ի�h�ϕ�`Ճ.�u~���u��5�Έ���`�Q��/�]ݥ[V�;X��<n��lF��r�)���^��N�dR>���e��J'�w���2&�Zv��iN�� Ij���HU� Xr+Ր�X�A��mJ��� �Ts}�/B�x1�rDO��9�c���K�]�v���؊�M��U��fnc�%�0�����*�UZ������>MP-�?*�� >�=0	Fz�s��˲����vO4�I�%=�Ǥ��Hۡ�1��;� �kZ:}��}t����$Z��n�j���Շ"�,״�-mh1������Я1��~:�Bh'M��s�����@k�ܶ0^(2�ɦ�O� Uh ^q��aLT�pL��Z(�+qN����-��f_ᕜ�x���=�&A��}��8��VĽ}9����4���yw��P�a1>OHc�H/�ʰ�+F�h=����|掎_<jg$�;�v\1�0K��yAj��\�8�<������A2ce���]ǆi�'a�;��"�����%�a�����8�=eF��Xb�G��fKn����$d2eRn�bSg��C���Zg94�}qQ ��R�Z�z�;E���.��������\���(�:��)�c��v����K[��};�W�����}�Www8�ܼ6��E����G���q�>D�D�,�������y�,/��i��e�
�/�N'����ƍv+�0��?��1PU?R�W�M�~��]��$mD�v �j���lP �M�x.|%nɡ�1=��[� h� ����f�u���ި����f
qY����yj�&⚷;�����楪����	�|v�f-��qF�G��T�Âfqg�"�»)i�%����ѓ���pY����`Q�IY7��QSo��}�!2��E�}�I�(c͛*\U;lF6��}�T6���\k��� F�����ء^���$���Q1�$�QsN���O���Bgpb<�&|���K�����H)��M3����:2ZP���i�|]�'"��n�H&��,[��NA�-8BTYK�C�Bn���1��� �m����LWLA1�d�4>!�A�K= �L��''-��`}L�+�ӻ@KaFl��%��L"�G��>��E���O���Y��[%��o�=�m�66L�[��?�:�-
 q��F�Z�,&�r�����'(b����N�P�XlU��o|UE7*�_Y{,Ud��ةx����X7n�H�c"8���ϙ����� k� �l�-�]�Wޑ x�=���f?���M^<�������z6��*�̨w3_<?����ͮ�)و�y���+S�.$���Z��6BB�'҂w�]�N1�C]�`|��P8�,�e�43�%��1˓�R���1��s��`:��]\�SX[1@���ǋ��kW~��D��d�n�n�jqc�T@dBR#��E��e�\ߣ��#}����S�pLb��z[��D�����?%r�*�P6�c��Y���0V�xGݝ��@�ٓ|�1;�Zv&�r��~��;!��@���9�Ѕ=�|5|D�	�J�5
\�>dFR�&_
|j5��S���w]��j��IG �N��33H�������ю�j�(���Jx��)q������bu9fGȐ�<%�����˿�q����|y�����d~ѫ�	��2\"�*��i'Z�i��?��pH ���iE��n������t���*��<L��+�
�co)	�j~�K��>���y��o��`�62�tG����R*�E��P� d��e9%�oq�%��"#C�8���b��a��Q�����.���Ag��y�,(/3ɜX7�|}v�R��,e��.;&
��eHK/b"�b�f�l�����vИLbl9�,�mǸW�^m�)oK\?E% zu�Œ6���N��2�R⥧9nu�:�M�t�?.���� N���y_���l.�����5���Y	��Bh�Y��/��"5qØ*w ��2��x�Fᄓgt蛓ͶH�1��^0���آ�x�L5A�p;s�%�s�Ӆ�w������i����̩Ip���=�I�yq����x{�7*OA�Mk��7� �Fԝf3�3_b���7��wm�N:�-���9;x��r3�M����t]'�9����|ji��>R������|��76[�>�QzY���� ^S��0�WFO��x hχ�Wpa�+kt0+�ջ�|8�@�<��\|��=� J�N95BQ�fm�^�N :��C�$�����8�߾z��ǈ[�<�E��Xi���NfF���w��#�z ?%Y��#ܺq�S	��P5B-v�ґw�������I�Y�g[p>��)��H�i��f�M:G����� ^�+|���pm*��ʰ�)�Bo����Ϡ*"��k����Vp�� @�R~�F�	1����t����4���8Y1q\��)s�@N�C�t47�����,�M+8v��;�a�ܽ[Tb듐S�G��-�[�3վ�A�/��7D,EF귮����4w�;m�F��04�JD�D�&$_+Ki�/()�7���?3�D����4��|<��;(m�_Ƨ�s�QT��b	�(d���B����"�} �1|��Ӛ�`��ϟPT���"Y���U�u1eq�^z�V}E�
�t䨴�s�n�Ç��M2#�G��JL�K�̧�Z{� � ����Lܡ�;�f��r����]��*ߏ����e��ZV/U�OYV����9�qȂy��?Z9ï'�u��P�R��\��¾5�
!�3�)��F ��<w�F��*�g�܁S�ɼ�Y� �E�f���Q�!��v�j����YV�d`{�V]#i���4�x������v�t�rfYC���,+0i��ؚp~�E��#�X'H�
�EO���R�&pR�-�T��\������j֬3�C�]�B��W!��ޯ��a=��pZ��$"01û��z|�Nl���� NMed�>�.:+D�U�S�g�'��Q ���	?j��k�
܊�!�|s���h@i���un��O.!�XC
"��>�N/�v�v�Ӓ�{�չ��,yT*�{�3���}13#�b)w�OKh�����
)��Ѱ��SO}#�o�.؇�b�2�D�d\��ꦝoP/*I�� ���f�Ĳ�Z�=�Cͯ�̓Mz_��أ`���
� \�w��]��Ӎ.�P�eu�C�HR��(a���<؃��1��ߵS��ggؗ�)f.x��5O�������H�}ڍ}1����d6:�����D�li�>�6��Gr�U��H�|1��9r{I_�Ur�s��O�=��W�,8�.l������CL�w-N��ů���SqB*y��dH������&
6z�~�\9<�48��<�()��āf�z�踜vfWT�v���\oު�<��z���f��7�! ����RR�c���	��;�	P��>(�����OX<����:W��K�I��>���'�V?��U���Y4���Wj dn"q#	��t1#|� 3���̵�gt���s43͂���O�Ͳ�eB�S�_��\s9x])�zz�~:Tv����\��j1����mnL��f�܌|�Cq�%���H%����D�䊡}�O���h�\ʮ��q�X�$|�Y��v5����z��e����!S���%L��2n��D�ܤV���O7����:X稡�b�eO;~�V�1��4����M�'�M������u�:��r1A5�o�ͷ��|��ǁ��$�(s��f����W� �5o\�����Q_�o��5ۮb�<zT/�z��0�M�A��c�m-���z���ʸ7˦��R���too�!h� ��0գ5�Yl)x�&�*���o`��7\`ا}y���@~f��)�J*�a���1qO����Q�2u�]�-�"~��0�=W�tb��d{�\8u�:��)#rx��u r ��7`�7�.�}u���s2T���e��+-_�s���;�K�.s�Y8b�L�Qk�(V�������&��[v`!.:��r0�г������X�[��,|M�.�U�����NӐ�����7�\[���[5Ӝ1��T0޹�Ltkr�Y߾O��t�#�}n]<�:��B���vgbP���#�6�t
��	�d��0i��P��	�%����\��'���	�l��!�C��J���A����kO9pM�:�2�T(_Z.���
Q!���(n\�]��JuR;[�6A\I���a�[��8�C5������ʦ�(XO�e�_��*7���0�leԦ�K8~z��:-�}�k� dE��Zs*���Q�>I��UHHN�&e˒0��sȞU9_�k�ʜ��~�� ��T}���̓z�ܳ�_?�*�|�W��b�%�%�ӫυ�� ��ìO�؋�vLQ���?"u��Ł��Ae5l:���d����%��G�x~���-+��+,�G�Q�%�{�)o�*�6�3�<���j~B	�N�%�=SPW(`���:�([����h�H1����C��y�|�W4�O�n��oߡE-�з�T����2�/�������^�Բi�b��RĖF�]�2�($��C$���V6n��IA��{�V+���zE�3�ťY9�Xy�9���q����M��w9���<=)�W�����Q(��6r��2 ����F�NUP�(�(��8,$�N��5ˤ[�$n~��� P�믾O�+�ߵb��kH���=�Ӡ0�'��UBNly���t@��&�y��`5��;RW��zP4�xNi7}r���^"м���_����a�8�m��nĸG:y=��D�����G9
��Z�p�������?�2S��G�Τ>�������;�!�����9��)\��G��	���k�1ʑE<z,�y�h��wU woe��v3���,"�z�@7Ⱦ���cf��`��#�Y��P������H��� �R�T�p�yD'�M[5����n�[�����ŪL�ipϭ�wrE�d�]��$X�\,7�۳�({��<�r�5��Y7y���S���ս�E_v+�n���|���v{��0����+ ��y���S�3��b��v��%�P&�\���/D����"d��5f,ԇVY�p�,��������t���"��gr5)N[a&�sf4|C�&բ݋����e�`8�^�U�&p�w�Dz6/o-V�M&��}F>K�iʩ����Wa_�S�mB����m�k��s���@Dxm��ڲ+����ɉ��=�����h�U���yGۊ��;����ޭؼ-��R��F /&"@�:I�<���Q��'�e2	�Ÿ+X�������9N8�i �5���́g�����gE�`�$�3>�(i�Z�K	��S��� ��ah�a7���������p[A�i��L��Cd��t@����!�s;�<�w��Rh�tEH*1���[��v��Y=wDâb�TB�QvH���a9�2n��l�U��������;��̱���LY����.M��ZxYdLl��Y�� �e����p��f\�-5ʃ;�I_�ls���|��ugm��,���&�!O����Ru�����th�x�
�Vٶ��M$K(�ƞ��'��ؾ�S{���iES�=[q�fq�
}�����]i�ЊEx\�^�Ã��>���3 Nw�ݳ�{�8.*��w����\�;/��u~r��߅|�v�EkRZ7K�G��y�Af|.�<�ׅ vF����?vT$�ȇ�B)c㒙w�W�(�8/˴f��eU>�[�M���Y��ݹ�Ⱦǌw�/�A��� Hb�.�O�^QA��'�^�}�[s��J������U�~S���N� �`�5lvj��[�H��ۖa�D�.%�.���<T�C|o���l�������a�?�b�<�I=Q򁗝q،\h�*PP<�{�=��*1�G��L�7TL���ם�ض��|4�N�*�lbG���|�"�gi�tP��V���>'$yQ��M?���M�?*�-� �_����H{z�����@w�g?�[�4ŭ���ͭ\w�MИ��7>�:Ҧ�I[�Xf3��_A��4�;���[����N)�����c]��~�[�j;{��"�G�x�B�9�Rl��xZfB��� �-���%'o�����YoKU��-���&,V�	% �8g"d�V��ɺG� ��W��{��b"NF�(�}V:���)F�PD u}f#Rm0%6�B��@��:7����9UA]��(��P	B�렾
�Sƚ\ի�H��v�K�<ُ��M�GKX��DoX�K��C�CuLL�+оV�R�D]0�	?GZ����C`�̙V��Iع寫¸uς2������l|ҋaC�X(���%gki���~�^S�L;}��6�4�ϋ�0l&'OYj4}�g��T�Z�$OI?����n�t��9��ӶSJ9Lck壮f�h�k��w��M�/�N+6�m���ֺ��@*�:�[�L-�җI.Q-���ʀ5R�����pqc�`��o�@{�����"��8 U!�ho����s��Tz��i�z�E������7��6
IĔVZ탍��و���Ì{�چY.\�������j�?8u��r?{4���p�}!���H'���C�G1��G�T�o��f"wP���=繦08$G�j"�	�A��ʍ��$�SFi��t��S)�m�#��20�ӾB��#�==���>��az�AW�ڂ�i����b&&��/���r��҆�z�H��'�U�:+��鱇� ���8Ǟ���>�?a��:��r����Y��?Y�W'6:;g��C��ܪrk�}�;[T
�7i��)>M�߳�3T̄l�(��o�+�~am%/
����4����ؑ�ي�QJ1��:
��DB��[�����T����*���o�=�?�uGUZ��8J�s�H���v��TSa4��aM�[��~9KbܞG�>-�k�?�#���B�+���NǮ9��M�q	� �ƃ�n{~䶦N���E��?�v���q�t�&p\��Gy�L�{��[a���`��������!S)RN;''M{�Y�)
C�������O�����Ah����E#%L�j�w�y��_�p��zM,)Qчj���I_6�t�$�)ߴ�o��
�0H�꺖�Ï*��fd�ZN�!�%r,���Fb��'
���;:��$� j�M���v ��'Y��;ȮS"�F_��58��)ױB�,�!�sU��������Wkk�
["���+6�U*�.r���W�ku��A���`���:,�fMH[���s��2�Р��S����[!��?���[H�k�2�`N�\��<$P�?<Z�m������A��66��0��J�`=��/±��)M�\#���}$5�t3�bg�ķ��C�D��?!�gH�L�(X��Qn���=;����AW���x������e�����Of����
4��Z��P[�V����L7"�@� B|��fqR M��`�(?^n�V K�ԉ����.�6�o�&N���6oh=�ʫq�H	����9�v������$[XɎ��$�<��W#=��-�+>(�$mٴ������L2��}�1*MDF�1��؉��f��>6�s�h����qa3~s3	W�<�y8I������"�w��h�B�P����[�Jm�sG��9�l��'���;�i��.�F
o�ɣ���u\݅�I�`W�Lm�(��}e�T�,�v@MZ��/��r�#���<����ᅚB��sS�!|([f޶�*'C�Ҁ;��5��Q>����v�׉aV�����;X����n"�j�����m��uh���5�?zn��&w�F���,�3`s*���19�7��Q�J|�B���&��^!<���=��(��`�����B�6����|^��B�u� ��_&p>;�Ӫ_��^R�b;	F�>�)j6�71J��0]Z��,kı�Iޯ)�0`{�ocz���z�R+�
�\�L����(ƚ����Q�~��F��F�@ЧlQK/��k;Z�x�g?�Q
y� �s+��VR� #�M 8*,B��q9~i�����=J��L��k.g���F�X�IV�Hؕ�#
K�����e]������P47�w2-j���Jg�����iꐨs[]�,��ct�Jξ{�,�b48B��G�"/K����	��5�ǣ�Nk�D�c���>:~����)���&� ��J1T�����F�ђ�i4�^]g�����]'&��0?�Gz�TI�!,��ޮ��E"z����p�K�8�[�iBw�G'� :�S!�X�R�O�Z�XW���IgYN�AAI�q�юE!ɕh�ib���l��׹����XY�`���`�^��WK=�zmn9{�Y���f��7��M)R"�+&��(��5��?�Ƈ"�s����C�g �@7.ܠ#������6���5n
7i�G,�D�����ݲ���
��3&h�x+���Z�9��~��aF�k�;���<A�������ä.��?qx�ۖ���e�z^��������c�f���UnHlgh۟�� (ݏ�*��2�.Ѹ��w�&�J���p�����(�΢�疣��#�� R���%���Y?F��މ���X��.##�^�����Y��?*�ˠ9��E Ӭ�f��*{.���$��V�b�zKÐh�?}�+>��#�+�Λ[E�D�����6/��B��(��(7g.�ޤI{�?G^ɞ�ȫ�{G���������8⼄�vB,:˪�V�軤y�[?����!jfJ� cS�@���\���ƫ��H�����@���X�69���ԥq�|�y�k�>���A C�v���~����S8]�����uq�wS���#7V_<T?YKV_|��]��	rs�os�94Z�G�S���"Te֧(��_7�A`U$$-����Ϣ�3�'\UNW�bj5w��v�e�p�������W�+�Y)������r����8��?joL��ڲ!	� RE0u��Xb�u�2�a�jK��[����⿵��vX�b�d!��]?�] �;α1G<�vp�5�X�p���/*,ʍ�?�S6�F֮ժtN�G��,�)��^�w�)�<�^ �I��n_Y0ҿ����
2Gu5�6��i؏�~�Wa��030�@;�:�>W^��<k6K�M����<>TH@ktk��WZ,s�.��q%��C��R%��{������S.��j�5o�8��<+�j��c�/��{T�=#�ywXa��Ac�ͧ�҉sU��q�5��x4\��s}.um``�� ���D��k��"x��tQ���ү���?`6̻*Yhu�ZZ��[�Id�^us�Z�v�� 5FM�{���7�t/RV>-�٧�u��%w8���/ }�<�՟�_0�@�cwG,�A�.��4[�^���X�yL]sY� ����
�e`������uv[V�~�r�:��>�=���_���U��0��>���YY��8��xJ�c�����x��c���{Hj���w���ꙸ� �j�K!�$����l���%-�����f�Dc�Q0o�Gu27%�n�Ϛ�[���l�Ŗ2�{��'��8�G6��Rh��a3gŲR�a��{�ۉ#=��T{��({ H���鮮��|+�Y-�;���G&]T�!Ov�ώ���v�K�|'�V��G,��*
�0H0M���h����z��]`�J�Q���[e���хY���:\��t����y1��6 A��o?O�*w^�4y�&ԛ�Z�g�<�)6[<�f�V�AL�f;H�B*\�I�o��޾��#ϓT��Z����C��y��!3c�G��҂פLq���Q��{�b���EgV`��q��Q�i��46�K��1-����jz�)�$���,c���'K��U��K82t��������j�+_���J/����cQ�0�KuvT >B�.e�c�kLy��E!q�a#+Qw�"&��'r�Lh.�N���ѠN���|.�1����6�\E��󭾦9�~�j�#\�3����C�}�K����C5��'k�{�f�WO��e�����ͷ��N��T\l�2�<�R���s�W�h�P����o @��=�>}y�����B�۰լ
;=m�awY.'��f�.m��q���aQ~�����Z����-�T
貕6���C�) `�i}'xŨnJ'��	2��a<T�hdI2���Gf"$
.̤����3��	}���C&�U*B�y���(W��.�A�'ccצ����t:h�Ѕ˖p�����ݔ`o-#g`�v��x��L8b�˄~+$.k�A���z�X]FU1
e�i"f���#�o���w̒��_�w������2�~6�S�\|��0:G���RK+�Ay@��kײ&4h��Z�b���������+��#�g�F�� i$��~�/#�;"�+'x7����	�G�_ÔP��i���L{��ʠe���o�����Զ�Շ�S�Rė{�v�������t|&�8ΝN��0cp�,X��eU7���V�ͭ|��DHSo�5�F+���Ԃ��Sq��5����~)o�O�O��9lj)(F}q��^��Rw��w�R��դZ�*{�qo��R��>� 5r'�v��/�%��H9�2�
UiIp�+��cyf�җ7��/����kNm��^�=A&�	e���{��D�< 4�e�։�c%&�b�+�t�av��!4/\<��|�lK�F��G����DAM����VZ�˨_�����u�������.����x���q�rcO��r�<�-�2���C#�fm��k�9NϹ�ҕ��0����T�P�+0�K�PnA�ٲA�G6r�����:=�,��U�5>s���n�̳P��9�1xӁ4h�g֑?��a=غ�淌v ����&�/��M�Po���=��,�(���q��lh^$mh�PZ���Z*su"�R�jɪ�Q<�eS��f��sl�夹�
��i�Oe�0e��<���,�z `]�K'3���=H��2Y*��+���:�6SI^��lZ��r&%����Lu8��/:
a��/���Eh�G��(R.۴t��u,u��U�H����>n{�&����˯��2f�m�����H��Ġ����o�������*��7r��|����}�#}Z�@~���48qdန48�X��d��Py�(F8��K��g�?;k�y ���l�d̻f��a����/�O�;���y������5e�Bm�ۥ����J�+�c�;^zڛ���*���<Gb8��ϡ�WT5�8�X|ffJ&�*o������9\p=����ƢA���lR�?~��U��$��P��
	}�6�SX�N��V�Ī;:�\9��%�r��"w��|)bV���a��ܚ�T ��S��*I����'�cEu�W�R���9a5��TIr�[}C+����Z����f���YХ���Wy=MZ�ً�\�  ̉rM���Q"���.Fl�x���ч��UCu��'8鮦M�vs����}��>��9��K�)}bL¥߿��c4k3����%~�*-�����;K���?�aD`��F�����%��DW��Rg![���{FbH4J*�t�>�4Z˱#��z�6+��z���y˙6�eb�L�؁�榐"����U��X�p���F&�o�=��]�%����Ye��Ct��o5~�98~f�~}��=���`��,�?�U��h[�D�;�\��m�bo�"�U����F�1���PY���A ܚ@�a7T�X ���i��"��)T����T��$"���%za�-���H���G�& �MG��p��j[�T※2�f�� ������}�$�W�]پ�J�W���3X2����V���9�0�XG�^���2B�:�*��|�ݷ��Dt��r
aO�&Ӥ����7
	�Ib`<W��u���V��q�!8v&�(݀�Ju�ͽ�%V�~C��u����B��HB�)
?��Ry+��P�s[�n��e���Zl����@�/p�����+o���f�,p	�����!���X�CT��H#�df�A�b9m?�zh��6���n 1��\������ȧBd���/���=�M��R�fXd�����(���A�54@��Pi��%a��o1�v�1�H�1GT��E�zj=3�D�^�����4B~�G�F���W׈��z���՚�%���Ң�Q���NdY�IxS�⁫�Z���l��7����vډ�~An��Z�S ��?	_7C�~JҲ&�!.S=�إ��b��%�T�}g񊘾�e���K���uk��7�%�Vq���FƝ�Zd�����b�q�^>�&wSծ�	�U- Hp�E�/�;uw�a�w"�=ɏ����_Iy�ԫ���$�\�j���MX`�"���↎](1h�wڄ�ғ���Ex�65��tSN�xdI��*�T+��wL>brB9��7�ݼ|&����ٱ6r�'N��4��jXF�ZF�I��٩��o���`�u�������2�/�X5U-��rV|YO�|/4�
i=�؞�L��o�+ː8�@qP��U�>$�<�[�\@��	7�m\"�t�5�k�
qy��&2b��S�!�I����D~}��ť�>��m��#s�����nL ��!d����uI��o��~d>�I(`��I�P�Ƃ�%���Y����q�f������q���`�)¦�%�U���@a=��|�t��ʒc��M[�]�l�>L���s	��D721w�J+���ӓ�EŸ�K�����=D|���O�e�=����o?Ub]j���2�`�Kob7F�`�bq��j&�_�0�>� �`��G'�п��/��s0r~��BM4׊Sl?t�(�qSj^�{��v<LL����K�˺Ca+��O���U�&�y�\Lj8����!"�6��L���`��*2���'�|���ӮBl
<�uu���v�ILp�i6�{����
:}	�崏�R�Ԝ�nE�4�(fT3��M�� ��0�"�c�!���q����{�CjP�X�(ɗ�2���~�K�	g5$M����b[��9�l��ɩ-�H�r5*�:G�H�\��x�~�D���x�8�U�3/O��P/x���V��g���ľ`}h�����4l�Շ��O��ZD�~���;Y�j��Q)~D�h\�H���0l����B���k��W��H�:5��k�TY�ѣ�03�LM�7�($d�V�Q���!���@,�?)�T���ĝ:g,���C��Vk���禶�u���>��Q�޼�
��**�"��(U�6�
�M��5�:����A�e���zǔB��'��
����0�^�{��e���u�7����z?�fq�گb�A���$n�Q|�;�U����fŮȷ|�@{+݅z�<���WW�r�:w�[B����d���f�_o�_zߠ�ċ�NwB�\;T/�炉�5��N�
r0�V��hؔ8Յk�B�a� �9C���^�2���I��^�7����&�aa�B��K�0}lUp��'�"�4�};W+2��jN>����B�������2I[ݚ��^�h!Y
��As��f�b�:�zJ,�2{�ň�����YZ@��o���U�ܼU��fz��"I�ٞ�#݃-f�T�KI)A��Fx�x+�yZ��5���s��2���Ɠ�cȂ�����Ӱ�|�����cѥ�'�\�5�n�j
2�9X=ƨ�-7Ay	ŏ�����rs�]�ȵ��w��[
^(K�
+p��&��f�4�.9��w�����V����#d��j�`\*pcF
����f�J27�i���d���)��
aY�^�K��`��'~X��T�v&��V�`Z+TFUp~��6�\Ő�?�%U=:R�P���/jl�Ѻ硣�1�d�x�T�-"[oh��`}7(j��֔�0|�"��h �	F�O��+Er�hg'I]L��8��L	[��ܡǔ_�7�B��|o[$���W�1QO��\�{����փ�Ow7ar"��O��B�m��R�4K���9��.>2=�L�y����OQ4ܮfCƉ�'�ʩ]jFbS���68�B�k�Zt�f�m���O��НQ�Ԧ��Blk|�'���9Avf�@8�^`��Gas��C�J��6�*Ǐ��LX�ܵYot���<��q��&S�Rʇ�믫���3H�1ؐ�ٮ�9�q]�Mi"��~<�����H�ؿ��Lg�5�����a�4��"����@�1`d��J}y�{g�8���`WD�}�Uન>%ź��ۥ����Ko��4	/ch��E��2O�]>�4-\���'�ʔWBqn�Q��#zz������i��<�X
��ba�X e���2�ϼ�N��V��C�NLkjN��ht��!�*�2��8�]ӷ�Ǐ|�Y`�5��L�g��:&n��|�7~�ɩ-4N�}���f	�HtE��9��e�) 2;�%��ڼ-s�����<A�1�^~��]�JhQ�ugS�p&(K��2�/�K�.צ:	����x���(�l7 [�d�2v�R�Ԓb2f��8ʹ��/�ȯ�^�Ɛ��u�־u@��<�W��uN�� ���/�5��q�L�ÒM�E�o����x?�������Q�Pq������7K�k[ܹ�:��W��.%Իkb=�m�yG�1-��MA�K~�$jϘ���+���j-;]���&>�c�9�9l�Tc=��T������)��=a?j�� �O��#�g��, J�z3��;����u�)���9�[W��!��F˲��R0�揶CW�d�3lAG�)�*t�p%�lN�0c�Sڢo��i+����.ݷ���h���/�_ÄH��m�Gg�#�+~�~����B��~��!��)E�[*)�. �E]r$�O?���F�Ƭ�/h��0r�������f_����Kvd�#򑰷�&L��&UHq�W��ͮ.��;���Y�:�ތ��_R���w�}.	ҫ3�� �X�!4��(�K�8��Q�MIl �*f`��c��]AZ�@9Q�ǻQ����i�0�D��q[+������NzFq�"�}��b��U�h*,�	�Lͷ޾���8�3P�c�y 3|>sU��$�:�C0s�Q������<? ��BV���l)�r?3����Űk�v���>����t�@ô˰A�uf/� �o�����\DZ�Ŭm���'��%,{���G�n;8P�J)��R�_�'��M�ٷ굫��W�����0E\�'��B�E(C��k֍O���X��#���!��]id|օ=�h��cu��Rܧ)����ƶτ�d�$�]��sQ�Ć9e�a��E�1v�����(��)kse+Rױ}5��ڗ4��*�����"�W�������$G��������3�7�k���4�9��Z�#O�N�R�cu�F���(��A����(�IS�	��6�?CH�������ɱ�6�
_�|�KA��)��xuC��fc%�l2�cc�6�5��0��U�����ބ�غ�VSK�H�O�K�춬�n�~o�����QH�$�l>e���B�ϥ	zm��u���W}�wS�0Q����0��nT����kኂ����]���y�}���E�p�::�wς` F��IvYq���ah4�dm��f;;{弎2Р��^�st7����l#.�ˏ���Zj���]�;�y��|S?,O3�!��\��N�e~��۹�|��t�0�yȆ�r�G���I��»���x=�b���?��Մ�ikDE
q���G`8m��~��ᓣ���&�opJ=�I ��آ���WԮ/|ԃ���Q��W�kNL�o�Ua�7�K�Cn��cL! �gщj�mJ�r7ԅ5L�NԠ{EM`�h�KY�-�_��m��5T,y�9�)���%�����c����e9ފ�]�	'�^&�%�9�L��tDd�u���X��u�cj��"����C���vr���oy�wgR��6i���ڂ'���hTS��K��������%�ź�o�?@̩t>\��j���х�����.���a)��5D��Lp; ��J�O�^���b9�De�`��O�ur�|��tڥL�e�Ô���>%��F�8M��Q�q�{G���ąfB�_^�&�U�?'���S2$�g��CK]�!]�N�G���P�lo�ߥ��5'����q!��@O.q^��P�����z�w����hA�[T�x�j2�oK�e��:��z��,�.c����+�!��X��9���Xw1�e����{
r>?g�K�,=�G!�����y�e�98Z&��2� m������u�=�������W��(;�d���'� �yT5�~0�=g�2�	,c��Ț�zy7S��9�њ/��&�)�U\
�Rap�ri�#���4�,�=/���� q)_���]x@Y}!���cW�ԯ�o��7a�:7��7���Xn�m�'�ۢ�H`����>��o`?ʼ���)�q� ��VYwa�z�D������r~�P,�e���v�Z�{T����� qI3�u:��)�ӥ�4���^����ԣz��_W�\^���:tS?r`��9�@����`*�z.�o�K`�ῥ��J	�Jt����L�uS"��o�쓉ZD*��� ٤��p]߭;L+%�*�T����Hm6����>�(��79ńh��U�~�N.���p�<޳(;V�N�M����K;�I���r��>�����d�:�����5��{�Su�x_9����84P�_��Ц��LL�{(���A�Q<[9Y��<:��/��ڕAGyxe����T��V����ҚLo�3��b�g�ߨN1)VH6e:�?�cۏn�O~�ވ)mw���X�s��~�sSH��h[�6ߠ��;�O�zb�����B�x�|�J*����U��ֲ&��A[�A_,D)�<���7��v�jqJV��j�82x�
q�m"��b�~�v���1�k�e�6	�Yv���Z�)�:id��van�!}�*������!υ�т@7� *�k����h�4�5�!���uoַ��2����(��f$�	�<�5<x~��w	|w�I	��b��'F-�И��� ���(w3�𩑔HZ�t��+d�=���z$:�TܪY��^a�2����-{�w�Cn��  N�q�(C�}DpW�p��j����G��	gl1��,m�	%�Cx�aJPq�_��&_��9ŝ���fa"����I[���H�QY���(N@C$�bFж$�Ӵ�f��h��[7;+��D=�j�!�l[�كJ�U�����2P� k~�e_���4y� 찠�_�[�Z�dް��*��������y�؉S�D�bVw+O1����j6�BS�6���ܺ ��z3�1�<��iC����?.�d�$�l�F6���>��ė=��se{�݉��}T�:�aU��f�Z�������Ha��Hx��ǿ��ujJ����d
bE��:�!�V��N^�U�|$ml�+ű�VNqA�r�Y��[Ns*���9��S���䬪�M=9Q�c��'���{���)9��3�Nu��c�o٭��7/\E��<�}L%2U;�qΊ�<�;Bg.�Gu�T�����	��[���}D��q�3�lg�:mr�^���J�S��m��Pss�.��J���ъ]��,%���|	�ime�D���f����Oꈉא�z��
wGY8(9�{{�<�%�*�ʦb%�aN���;ߖ��&�0=��A�	��.��fC;^���?_|BFv{>ɕ��(� �l.�h7��B3ݷOҒ��;���(x'��%�{�,�{�2���!p�pӗczf�L�lDCT�q����X�b^� ���&�N���N;�d��E'�fŒ���EZ,4���,f_�]$(�溳aiP�DJU<���c��_�l�br�{"����TⰍ�	:bq��	��)��s�R�/���d�n��%W��Y��+��:At�"����)�y4С�1�FQ��3�*~,�� �Ď�qea(��ݖ@9ܷ�6%��%��6��t_�H��>�)�@|���2Ee|������㑇�9��Cv����[�M ʯ{���h4���ک��S+�jFc��ڀ�����
�;<B5�&@D7�+j2�H?��d��_:yjj� kAE1�J#��L�7�-���رo�K{�#8��ER�]��P|�����
xv�c���<.C���"�m,����v���&�qzN�_[�Y�0a7^Wu��F�7�S��7.���[/
2�J���IE!C���Q0Yeo����?��B�����קH�1���b6.�}6�te��"�tp]8l��4�m�sfc���
i�^���c�ȑ�8�r�/�|X��pA7���+ӂ0�!՘�}\a�)Es�J�� �T�1�p�}�,O4?���6�R0iHfg�d�W���˴ �zR%!��3����`�P�R���7v�����Ջ�l~���'����! /oSfNȒ5XZ.\X�z�N͍���_G�Ū ��i���%��_��9u��n��W�w�M^���I;>�/~f�б���Ҡ��(k�8�.��׿T,�,�gI�s�0�Y��-�7�y�e?��R�gA�n��sG���}����Ϟ	�,��O��5YE�V8'�c<���(��B�{q:{N��L����*�
sC1����� ��
Y���A��7��d��Ŗ�M�ݼRi����u�٭��Mz�Z#G��ώB�s۪��'�g��F�rx�M�v��O��+ ��(�K	o����"{%�eH�3��ylt����F��nf4q)d�_��m0I�=��Q�����m(�������f,���v�f����ֆX�bʉ��m��	󯂡�D��RLJ�Y��!��Ql�ྣEٖ+�l��g�.Y�L�˶h����SM|�=�MCP�5�e�U�z�G��:�>&�혐%<�ng�O͏�96�z�S�b�}ncqY_^�;$r6�墂�4�'/_��9^cP[r:fh�_�GR�iVA�/B�͉�\,~�/�	~҆3�oH���U|,2�=���T;ԣz��*L1��ě}��O":�A�u�h�r{1� ,�*�C�c��&��E�����v�A�k-�!*�,��ɢP��0:��B���a���Zj� �.����gb�q_^��,F��z
��$>|Ҟjz�ë��e�7t�N?���hD�K�����JNt*1Ns�8�*�7,�A�����
�
��ӌe�U�~]����[���A������g� ����T���0n@t� ��~*
k�ң�!�In����Y�m� ۣd�tƠ:��o�dL����nP3k����Q
z�^p�%M�ګ�k�P��~��IC����h]n��o���!v�J�v��e���-b���������S��}\!J��6�.Ѐ��~���0L���w�	�7'���hU�B*k�UϵV���jP�&�>�U���i��5ó�ZX�цX�\s��)�g�Z��i����/�RB�����O�}3eR���#+��{Hܓ)&N�*��C�z�(�����u�a1�3
������[t�s��T��~�୅��{;
{���@��JJ�S;��pp�6;��W74U���x$U��� ������j�Ȅ������)��
Z�~T��� 7�j�[�Ǉ�dǄ�,��z���x؉��ꃲSC.q�OjOȅ����ȠI[vm��Oq�*�ސ��F�Z���,��%0w��,����z$x#u�� ׬�ӂ1��d���3��Y@�<�0�ɼP�ب% ���S�W��abb�c�.��������zF�cZYro6�j��5��X����Mh5��
��j����~�����r��s�#��{���d���+*h��聰~0�[,H~�z&I#��� a<�����P�*�ɪ>� �:<t��3���e�K%��%C')-Թά�^�y�s�1��~?}Cd�P�>�}� ���'�\�.y��m3�"����Uol�1,a҅ ��ӧK&�P|cx(�k���8��%eH��2�����@��IBR}M��)3���c-x{ӄ�yP���/)��Hi��tp6���>ϣ���.�.�u�gcvIU]��9���Z�+Tm��dvʧK��x8��Em��f��>�)i��S|O�0�.���$҂a�o�:qZ\�B��q,6[P�D�[�)�H�%΃�Ƶ��z\ER+��KeY7z�����G6��j����X?���?S�/�C~`����VN\5cL����
3E��XK�c	�6�@h.�%�.y$��R��<�}��K�{����(üZvR��������Tf$�x��?����uգ�m�"��vQ�~���qG�S@�d�V��u����2H�-4W+���,o�6p$��Ά�UH�� �4�HC��m�E5��wh�"� Z��Y2đ��ҁ=�j��MGc�2��[s>8ޣh��a_G�q��������e��.��7A\����:*�f���%%��/��X���=�C{���DS%�Z�`ͪ�RW�:D?���[	>cJ��DF�������M�ֿ@���l�`N_.Y?��>Ċ:p�0�waj�z�( ���ov����h��P(j{2�˴��+\2��4]�g���:E����v�7�F�m��Z���p��q�
���7��rBxC�"4H�-�cH5��ݗ�M.��H���Cx�v�'w��_L��tR���[�ۂ�`F�����d�U�(���� GӴQ8V���"��W*!ۼ�;�hۺv3t�}�߾UF���+n@r�!9|��� ��zXM���E3�[�����d8�j,) �9W�ă$����|�� vW��q�K��ijrJ���b�x�$-�A�#�4�����y�i��=x�����|��[Ʋ��N���ڞ=����]i�l8rUˏ���F":�[�ᣒ�F��d��D�0qt鮪Q��Cʈݟ.馚��AJ��- >cc�>?����Xۖ� r��k&�\ߠ�S�t��~9m�����l��aX��S�k6�ΆA��:���W��d���3����V���t↘\`����q�+��P_de ��=��E��v� j�9�V�ѷ.X�}̟I���w�-WZT;^�~�Ka��-��_O�,0�Yۢ���~|Q�}Q��`Y��SH�ur����l%K��Ͼ����J��j�)��gpMH{�3����s?�B�ԫ4$i�A)Oُ����!'��������M��~JhE�|���nӇ���$�#*�B;,�x\�����[�	&�t��gy�Y(�	 ��g:p�Ǝa�r5qӥ��U��ɵ�̛����^��?�}](e����u/���>�|j�G����,���D��0.��7���	Q0D�Ѯp��.qA����uY��7~!�UiH�%�M�i��P9٧�R���eY��be��F]��	�7�lAy��`5�߾����SL��� ��f�Ѵ�v��O��n�Mؼ�a[!� $�Bq1�t���c^��]�n/�-��n9`'�c1qb#�Ȭ�J�� {���A�䥧��W0��t�2��$!LM���P)���P�_c���d�_6�*��F�#ب�R{Pɋ���㓢�#��~2�ޕ�X0f�}%`/5F����ԏ��m�U�s�׷V���j�w�C�6��0�VK1��X��SI�"�(o\�ї�ȶ��.@�F����*]�����G��0P��[r�/�����;;[O	nV<)�Icwn[(v�Xߧ$�5���VT+"�)z'�����%Ph"!|�i�����c!��_L�v��
�>ñ�'���Oz r�(�[n� ��i6]t�i���l��ڟ��s�wq3�]� ��t��c���CQfpYo�ܺ ��dR�� U	�N~Q݉�S�C@��b6�~h������&H)"��±L8�#� M�Xe�hNc��i"^= ��L�:
D�P�������@�gq�U�X�yUL[C�/&&�ް;2�L,���7x�*�"1��j��
�^=�`����S�Pp��?���ɞX�$�C�)Vp�Z������h'��&�CW'5�ꍤ���ؚ����'���y=UL΋,o�9 k�L�Р{B�_�g��Tq����o녧�N����K}�?��"�.3���o���
������V�IB!G��5`
�R�5��]d91��j徴�r�h�dMf�����
J�;.�Z���4�'j2��cΣƔn �y�^[���թ��@e�V[U��$1Yl}̆�
�M���td�vMּ�C�@V���sm��Ep&�j<�	Ț\2��}M>���b���Ī����!�jCp9�V0�kR;*��3�29��0������0/E��5�͝���ow1�L�z�P�w��Ӌ�)�`"37�_-Я&N@B>��s�#���o�=�+�Θ�Z��R��$�u��du�!U�gc�q��X6�Ϋ��ū}p��H�+�� މu�?�b�	ؠ)�t?��?X�I].]�6j!�o��\���RP�rL���G�'@CR���,�k�E�e��@�סF:�	|���P�ع�B�M����j�@]Ou�r-�,�J���.���"I��(�X�a�����-��uc�%%;����wj��J�E�����1��)�~t7�.�ٖ��釋Rs\E��\���K��Tr�^J�����\n��!wN!�&Ȑ��Z-W��ǵ�L���˶��'¡(r٬\)*�@�x���!�/����� OI�n����r��ȹl�PN��o�&�H��IS���iN�����/6v�}
� i��G0<K��Z,Ƞ����B립)�8<�>����etV=��� ���G���IJJq���\7�Yݱ�>����N�|�������_��NT�^5���z�C;��u;B0�B����;��ɹ&��(�6������-�͓��-v2�=t����P(O�<�����ZJ�o���#Z����tYU�����^�3�O�!$�s�3\S���t�;�դ�7P����:y��@�q��R-N�h7��hlI��]<��Qe@G��-�Ryt{����#�P��P�.��rC��?���t�n��O"���[�@ϳm#LT�Pi7 �,�1��5�Z���{l�|�XЗ7f�nqP�e���wL
��XG������m����L=������՟�dY-I=�&S�(�f^���c���Ei��4��!H����^��<�I�a���Jl�F����L2Fg�Ԅ�%	h6c�r��&���{<Q�i�I=U���|k����Xp��a.Di�}Yd�ӊT^����p:��^�0������u���-�ñ��8�!��X�I�lS�YS�8.�뭁[��.�.
:�(Y�tD�k[� �\-�xO��_`^M��̅jP�Ĵ3-��T���y�L��{�!",�I)KX| �D��A��7|��?F�����t�e!�Oǹ���`��*�o��~u��O8�l<����7=�6���)�q�&xr�ܒFT�wP�.gJ�D�A��+��|�����_� �4��j\��X0"e%��H���	vp����R��PR�u~Afw@_z8�lXs��F�9~���,�v+��H���c��I�[���6+,�z'�O9&Γ��rR�r�׫%���Ie��_� �q�+�8���T�SB�jl��1AB\j��f	9� ���feɴ��7�B�ܘ���R�f��B�Qb����d������:W����k�)�n_��D�{��=���z��r_?#�j����W��M�k��Uy;���+��9��pP�����O���� �AF�o.i��"��ya%��w_�@o��*~��x�H��5�G��T��@�{����`��Q�BdD[�y`󢀗 i���+u�!u|�G��Ȱ�v�iF�����0��Bܾg���↧Ƭ�/x*��ҼX�9�>R�dB�ve62�-��F�>b��L�w�IQ|�3%����uLz��0N�WAy���5�ҭ�.~M	U0��mS'��M	-�&�Oy\b�}���|&ǓH��g#��GO~����&�E�T�0�e.9T�|�}�?�{+��0��N��m�o֤��}�E'��*ͮ���=,aۻm[���'Zt�K���C�~�����]�Aj(1Ɲ��$Y;���/z�7e3�0q�䮵�bBT%еY�-ODWb�s֘��CI#�h�~U�b�������~����-Ȟ�=�L�<����o�x����E���-�#N�3ԡ�4 �>�E�q���=a�?�\ք���oXu��ד��ֈ�{��	�G�`�L:�y�ޠep�5+��ǲ[�!BӜ�0���d.�Q�M����: ��[ �����d;�,���n`�O�)����@���� �8��B��?&cy�T;s�i��8F��!�����&�t#i!�e�P"�'I�}��xrZ1���?ai_��$��	�!&���޳E�b�p/=�7|ntx�?��_`"m󩨧�cf
D�4۾��oF�w$��}����Ŏ@��J�ΓhI��sC���l��H��K�� �&Z���_l����[jM��ҡ�*ňI[,Y%��с'�r�;mLP��"w. �"ɣʰi�SG����`���x�\��q��w�$t	��A� ���j�y���ŭW�f�f]0���4~�==ϹOD����f�Yݺ�=���n�[ᘝFFc`O�$���҃�oR�ի�
���&�5�M�G���p�G4x��n{X;����d�G��I�q7oI/x�+�g��7���dGp����-?M����B���z��d��T"�b9�:y-�^�e6�߀t�-�f�7`Zn�ۭ�����%�y�J��|Y�|[���,b�c�}O҂|S(]��-h#��tA�6o��Ȥ��I\���� �bdD���ѭ�6o���m�z�1I�0N!��$"6S��)H���ٵ���WFr{�A_s{qF�&�AV0K��䱯s�۟��¸O��a�ݑ4uBe{�_�8b�v@\���W��3�G#�BH]�Q�K`BI��A̮>ٺ���G��i+�R�����-_Wܓ�Ez�N����u�	��}��y�fMX�F)LRBK�e�\8�'�Y�M�Gt��>�6d^��o	�!�-�{���P_7d�_�dD������ר�+�;O6�9�J�6z=b/���Zxѿ�c�A�@nq�}>)�j������sR���Ia!�%\�^������2�'M#�[@X��
�K����Z��me=��^�'Ұ�Fr�Nɭ��G�rYQ6�.?<43Vg�����0�e�].j�*2G�Qs�&�W��v(v��Qy� ��� ��~���[F+],t�讨(̈́�9~��,L�塱���pȑ���X6��f�m6z@M��s/�m+�Hې��VNKף���v�_�o�Dd���sf<0+���ˢҝiT�x���=�t�p�K)w-�2�P{,�o>.�S�1r��Y��%1,ͪ�)n��#�Z(Ӳ�{��4������o�}i\ԡ����u�[���nW�R8�	`e����(�ڊ?{=�����2�������p��q�.]��b���'���$�'�A�kl��3 �w�iVY;�%����
L`��� )���y�|@��{V������P����N�`���!�ƍhV��GmBT��{�f@"~뼞p�+1����H
3X�HZD^�+\qw.����
K����V>�r
����e�M�.��'OP����򠎅�����3a����OB���M�������<aJ�e;;�n�ſqVY�?۷CS�9��f�5?�rS��6Vd�RF��K�����,q��Ԁ��G����޳�ݥ�����,������ۂ�1��BV��Uwm2hl~��V�[��@fC��G��`�y��
�{m�����l�_�gc鉒,&}���v.������������
�䬐�y���^��0$�׹�a7���-`1=���� �[��6q+'��S`��}��+t6��)���XR�kUb$@�d�E�S� ��͌�Z[�4���f_�-� �c����yG����k� ⽤γ�*��F�ݱ�	��y~�w�7���� ���پס[���E�)����%��m<�j}�T%7yΗ�\�,}�M�����pp���F47_��-�#F�C��v�[ 9|����2�
��n�R�n�������F��I?�]Ϧ��0��ӣ�D��o��W���9�*d�����*��d�%�>�D�"no�Z��^7��_��ͤ�T�qX[j.w�3��ڪ�Dr(׿#��H�0�S���d�zִd�>�v���q�!3��.M�5�
=�j��.བྷ9�F�ʳX��j:�@a�a�M��M��q��i�O,�#|�$q�Y�)ѽ��~���:5�)R%�����F$�u���zԫ�oo��	����қ
�ۏ����;�?�������a���Xl0�]0;&�[�*Jߛel����w�{��TT��NEfO�-V�n�
D)k	�8 !צ�U��?N���eu�'���3�9�
���_K>����w�]JVl�ܙt3A~�������'��;j��"�.[���(,��f����c�(du�&�c�-��Il�]AFa4T��U��}�@~��2�+IO��nP�^V��и��|����}��z��o������HM���f�ӘySiE�Q.�)�8�"�2S�=�N���2Oȏ��L8?�lJ0�RpT�f���m~Y�_]%~aC����9�"��,�|�� ��� ����i��7�ӂR%^Ɨ�vw±���m�S(��Bw�Q���@��"t�����d]���ù_�[*?�/-�1��;,N=�f5G�¥�z��d.	
�X��T������g��i"�膋X�(��gx2����E������"�vX^"���5i7�'���驖�b3���:)�4�]�c�R���J��m�\B�x� ���"���ܡ.���k���>c�Q�֊��n�1Zuz�)�r���pTx��)���
u��Mk�C��G׹�{������%W]Obd�µ
2Ѽ&�F@R����DC�w1:J J�6�ۖcSW��GBz�P}�q���y��`tn��`5t/�jl��+�y�O���J�|
 B��ۀ�ʬ��)_�Z��r���G֥,7�`���s��J�T��-NКH�\��H��"L*�M�$U�k�*���UM�������xm�&j�ڔTߛ�=�~���� y�F�}<����U���m���)�9u��ڭ����s��QK��'p�B��XɃ�=�Cs��hJ԰"Z�O.Wb�G�+3��oԌ��u����~�ݒ����4�a�Ӽ�ѭ]�I�..^�����|�W���&^u�b'���I�9�ƅ,͌�O~)�,��n��-�#�\s����a��v �:M�#�<��Kci���dS5��S��E}zR��N'�'�D��+)���/{h�n�}[��� ,U�wA�o���K��{6�S�z恚����>������s��(�9�kS֣��V9�Em�%�W|�P��!&-�\�Ů>�e�
pڱ:f���Z(����4x��g�?���M�՜n%���K�=5�@�m͖�Hu�2�'D�=��G���3ql?�Q�څ���M�v|�f��5�����<��.� D�;�Y0$ņ$~�6�c��{
�N(T�a1�:�G}=E��VZI\pV��ܱAgO!�w4��)x.W��V��=ٽ���؈��JR9!nv�V�;0���������.�k�	�<�D���T��<�E�)�Y>Tc���������B䁄)�Q/_@�G@A�Ks.��\G"���h#��H���I٤��f�݋�`pm:�Ǜ@�\�������~����Ğ�!�V�����vaH(�� V6/������P@e�^Ո��3�:��y�O��>?<�������=������2��Ri�i�m���*\۳*v����,�Z� ��d��!�ǝ���eΖ��6w�I��w2��ƙ��T:#權�DPbGQ���c�K�`xRqi��O<j����Tǜ������x1����d�(���1<D�]�؆���`�����,���Q�{����;Mc���ལG'8�����M�♻}�a��l��j<������eCƋ����;EnXJ;Q���?ZYQ���̢lV�B2�׎��=���}؛Ydb	�L'��{�O_�W�T�:üq�(���?��j/���z9%�����4y�Nň�V��Z<.�]L���w��1V~8�	�C��H�6+^�z�S\ ����WP`Y�:�Htl, Jc2��8r9�t�p����1�����^�Ĳ�";-F�%> �6� 2vA�V7j9����z�\`�)rc��KQG{g%��v]:Q����Uq�/$P7�-�v����ksF�SσnC#?Ԁ�>��ڠ�W���)���KT�W��+F�F��j_���h��!�<H���h��l���]c�h`�������0^�4�!�|�b�#Q�n��k���7��S8�IÏP�e����������=�k�ɘ�-p��ˉBt�1�=DHթ���;v�EX��}��r�.�jZW���\7�����u�*	��j�~�J}��=��9�*�&��Ddl��|�*���y�Vt�ʲ������Jޣ�Pw��p�2��-��s5h�g}_�)�̎����y9��ń��g1�}-�:��{h�1	��@(�$��G�������͛5�}0'�[f�5��?��������l2��u1�������r$���{����-�M���x��X�!���I�{������j��T��"9Eљ�	UQ�_ʜ����5~�"��Z��d��ϔ�>{s�d�̏b�O
�>��^�_1�	-٨;���%w�X?�bValA���Ʋ���H{���Z�ǧCnv�[խ�x��=�a��"����{���2�/��B.�q�����ks��}��'�@�I?���o)��}�ԡZ���9@�3�����-v(��E���Xѫ+j�5JQ�]f����Y+�����=�� F�{|�5��ݘSY q�����y�T���En�g�1Yb �/��T���$�6E$�t���j�h��|㼩ZO�f~�t��	ã�M�?3lW�JjMO�p8�r���^�.�u�oC~�%��WQEAh�*��2m&�G�_���,u@������]���|�Jŗ�R���$U�e~RD������������M������~�0bNE� {G�R�����C�҆Ms�p������+�} �E��60>��|��7/��5,T�$�����c��UY�i?��q�$8�.0]&Y��c�oo�ϻm؆�|3[��n��2��_�"z���r�N��MËm�$h/Ԁ���j��UM�j���A����1m��1���4�f�&�E"h�ʥC���n�7g��$'+�i�;��Λ̘?a2#Po?E�s�Z��}0_12�9nպ�b/��r^���<�h�/\�ֿؐ���?_K] ������M �������Xs���0кc����L�K�V����<�[o���d¼��mh�w�틧��J��|��a���@qA��v�F�E�{w4%5�DLZ�[�������Qe��h��=`z(I�%Ն�[�W�]��O�d��2l)���:�LQ�u�u n��N^��2R̮�������R �YS։�Xf��%��p����D^��_��/�7�ON�Oc ��w���0u�Q��������!U�� ��t�kNl�w-̆�.Lۏ�h��}_�~�Lӥ��U�c8�6�Foa����=-=̭�~]ED��E�9��I��2W�����.F1� �����7a/���i�\>7�;�[��N�L���rP^2`N �U �aZK����)�?Vv�2��,�nJ����Ǒ!��-GZx�5�q�~�)SX�3q�rs|_����6���j�%��L�9�o_5��S��}����^��z���FJ4�l^'KP������W�@���(ӗdyL��ZU:)F� (�-�|���-��+r�Ѧ��	�	�VRsX�n�|�n���C+��]-);7�j#/'�R�6�iJ�������w����,|�F�|�}L��L�����Xu����6G��
���
���<�)rY$�S�2�;ǎ֕f��!|"k�8� 1GZ1��=bR��ܻ�~�6ܗ���U����=�����J����5�5�I��홫� j�h#.����U!%6_���ӬЮ��bD#kY�*�7�e:t��6[�@p��0�Q�6�{�h��(
f��Ȱ
8�U�R�]���xU���lQ恙�y��=��6�)>�(���4���g����X��·9�n2��+�Ѧ��m�mN�촚��IM��n:��ox������݉k��=@]�6G��ѧ"�Z\J|� ��9��]]���6�;�5���~�ozs�ɩ�b������t�W�>��:f�ֽ��͂Arܝ�8�`���]D�q�b����+,�ֺ���-����E���w�<'����>y���t��р
��^z/�o�g�D�.�M�]ڨ��eb�5�������l�1��q��|��z�rU��ԧ/UA����< �Ru�e��NX���υT��:���(���_7�VLQrG���&I_&��3���8U� �b50[x�&] @�x�=���9�p!�������1��W����Ǭ���x)|�A_4����˷JI�n���		)/�t��� L<�⯘(^*�d�\_��n��T.�z<��Pc!�����Y5��M��WG�Qp�Tu��ë�U�F�떎��U:hʢs���Z顎��?m�v��^���Gw�6�N�w���7�<kڬ�`4�,f���*]a��}���j�p+��n)?��KV�l���e���s�⃷��Ő�ǏJ�-�?/������ކ�-�-d�{�����}�ٟ��~8�R���+����8�N��U���N�z���.�������%��I͂Z���=�^E�љ<�o�6G!��˕�H�#scɫ�����,I��3�����[�a�u������0�2�l�
���<�У� ���M��>o�w��a�{���{�H��K9�XTQƯ�ÞTؐZj�N�DR�F�o8)i(�+����V)���!�@(_�|����j���90��Z�Z�X;�O��o
k��b��ғ�GCT,�ג���_��E� '�C�����7 ~�zz�+�VV�Œ#g��U��ʉ\\�ע43��)8>x�aG��<P��Q�٤�7 ��\VB� �!�ؼc9֢�K%''�LZ��7��xѐ��o�R�O{>�~�Si��g.6����Ƿ���t倆��wIr�\C�q0�5"�?���a4U�Iz:��ӹ ��e��]��	��R!��g�����
�}47�P���Ў��Ml�q��w�~��������J*�̷o`�F�MF&�g�K�缥R�88��`�1@�f� ������Y�=�t ��aQ����Fx�M�;u7����)����l+���e�`8,Pԋ��va�mk�M�&֫��#WJ��"N��	�TA<��I�v��n�~�.�%����ld�]T-�-� �
2�h�������֐r[D����\i;!��P��mO�p��G�0�r�