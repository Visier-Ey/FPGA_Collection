��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���d�v����0�i�=\��A��?��� (��1_B�f�	�Ѻ+|n��y��Q4�]�aY�����*2�y%����>��������K������ �
�D��z�z��C�y�B����
_�U��hkF<�~x�ܕ�c���bǳW�}N��g:��-�~9�R]�K���&6��q�
�d�d��a*���}�GPk"��uA����u��NzII�9�$�%��Ҿ��e���J�_��){I���Ґ����m�S@<�����v!�b��hA�]���L���SR;!8����$ܫ��{S/�>mU*����v�1C\�5��|�n��..�K�D��\�Y7��it�n��~g�gb�aC1�+M�-��-o��޼����7����ה�׉T��B*��#u�'�zi�_��m����l�g�ȗ�ޖ��#�L�C�=���B�Pah�4$~�yB4y�Roq�Fr��ln�]�cD�Mot�k�G_G~�h��}�ͫ����q��=!�-P�yy�,3��q�9�F�c/�0S��M_|�L��2,	'd.C��ˢ]�a��V�����5���x�JHJc����A	�B6DC�~Epj�r�lI'G�Oǋ��W�C���yh�iL �T���U���X���Et���8� dWnP�#z~����.q�ͻ���+��|ٮӲ^�h$��LV��QF�!���D��}tv8{��j�$���Y�d:�C1|BD�B:��]�.G1*�����aX�{,=UN�O����:� ;�3a\t]���艪�Ž�&��9x�pN?G�<�nǶ\]���͢�	��������E��?�Q���� `�<�X�����bՇ�k( ?-�f%ɦM�S빻�w���7ؓ�j=,C��l�����������_���x�6�	��T��Nr:=�x\Pa��#D{ػ|�V���1���'1{F]�5�v��ӻ��*bq���̳�%�~%(MǓ�;�s⮾�Hg��c��^H�vG�y��V�9�2��!�휁+vT���@|�/��q��|?�t����gAݓL��G���_X��SP��(���k��4w}��3��L);��N2i��}	�K KfCJ1к<�،�JP� +T�A���VF^�d0nP��T?����L(*0b@6㼜!�ٴHȼ��po;T�3ܹ���O��}��JE����^�l��X`]��ĕ���B�.��㐵�w{l��XԢ���s��2���훚���$�O�F�s/=Cc��k���P��r-Ek��?��+�z��(��e44���M�6�FY��{ZV ���3Ꜯ�W�|J40�⦧tK4��G�6F�Vi��dcBy>	��~���z�
����=����S��w���W|�Ǡ�s�H�l�+�F����#f�:Q��V1��M�o�Gђ��
A�j�j|˦�9З!��֨T���5�tUY�v%�-S��?<a3����8�������6�vH������auR����pW�u�ˉ��DB�s��/k��Q�9O��og�	��j�}Ɍ_��/��-^c�
W�.ͼ�YI��9��M��E���piy�C�R2�i�F��ZM'��|/���JB�ƞ��d�@+��"�q���~Ș�Au\��-~�[9�Lh!Vq$�@�o�)�G�(\#7�{�]KSg9�5C3M���ٟI'!l�r�D-#,���1G�*]��G���L\S�
�����\�
�Z����%���@|��QR��b��@+ndx�d���A4�8F-v�H@�2,�q�yYyj�R��F$Y|�J,mD���zT�m�ܤ���j��뮰<�9�����>�*!Ǐ��t����9��"�	3aW��7�j��O����#|�~'?��k�(9�E���E�܍Dc7TItļ�o�Y����y�d��d�
�;6�nNw��=�$)_aז�����]�������%��&ؾj���
���9<@O5Nk�_��}� �c�Q������-@p�A�����s���!ͩ�T��$܁�1VOtN�m�M#@�����[HnR2ޯ���P� &j�����ߩ=q	H�[4�{�RƂ�����D�]E��T)�9�q�Pp�h�~�ĺ��a���JaH�D�}�4�v��{�#n'��7
@*>�3F�T��F�Gf��M����DX�hy�N�7�&��7,��w8��7)�vr��(@ExF���"}#(�z���l�ϻ'͎oO���;�[y�&\��S):63[G�e���NP���|�[ͽ�1c6xKEΒ�JX���|��"L�f�@�U� oZ�f ����*�+g!�& ����|h*��r�}�Z���6"!��%2�]='�go���NQ��D�W�.��S��B��b)ѓ,�6�A]0�+�zA&�<���6 �O�mƑ��	�"q�C��f���6Q��r�VV����>��B둜���A@0HWĽJ	m�!�v�̟]�����0<��v�F���f*}Fh�YG6,�� ���&�0垓})T�#t�G���A�#f��c*IKI~I<L�#@�d[����-��S41��@��9pʫ��=a�Qq��M���
֑;KK�n�$1�iy�)w���#(J�����a��=y�4��C3�s經��<��������{ ޹�C_(�7W�y������R��m���hfy�����u�G+x�S�,J��L������l����©�×B�В�pUm�^a@�7�]�:c��2��L��?���d��a@�=/�Q��N�F��
ڷ�5�b�ng6�d|�~^E T�[����4��V��8C�]Z����\b�5�Ռ]:�3�V�H��@��I8��, ���e�,U��Q�xzMؐ�H����=gʣ��K�)�>�	'M��0����1�3���b���F+������g}��oacK7�M�s_ǷԒ2é��-���u	��:�Ezv�XuTJ#���� �θ��d��S�g!����}?���[oNt��k�d�#;U�َ7�y����]qljw��-�EK
��tz_��N��=wWǃ�y@����SJi�5�P���_���m�g��d_y�`>'�P2�h/����M3� R�6,ج��l���l��*Ŵ�N��H+>�I�/��0�ʹ*ሓ+�X�� ���YH�]E�L|R,�r}qw��\fgO����7i����תn�p����ۀ\$]A]�%L`c,��~ߎj?��u�e��W�Ά;qfJ��M���y��l��4���^�_dm�hs�&�w�*~1j����3�%��V*zA-��$A�����Zv1��$��l�4�����6�R�oX#^�l�)=��Hz�W�>�2!�Q�Am�g������a�..�k�v���K�~7�!��fi��B��NG���*�<hvl@������
G���wc�  ����