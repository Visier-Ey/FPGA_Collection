-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
IdRkKZe3nxHdkZcdU2KesHajmwHrJJ3BOvMjb1byTRqvAKCnSYPe/Vs6z8BZgyZp
SbETAA0xfImPu7GpMhvd/azJYOMmqLj6bvF5FHaVmlb1hVo5WoUQ1EYE/XIUYBng
8FDVJNG/E4PRrD3udng7qJQJfUAxSCN+S9eSq+SLe/E=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 6315)

`protect DATA_BLOCK
JRqTwIB+6Zr5hXosDWCULYUN/+wqQ3tFB40Dplr8qnZktbgz+CQMBhjOi6+/f/4w
dFYYATwJcaVe4oZmPhMpXnmOve23nuXsmOwtR91rkF/7830NI3ZUeoYrUnn8WZ1C
EH3pBwi57UcS+iruHt1eFLCYHeRl7HshXfQ4jKTg9C7zyD4oR/G6qrSxPPNX7v9t
8a6EHXBl9gyGMx+6GA/fxK4cw3nWtL0DxhnMA311IMg+UDiQm9cUMA62Ovp1MAgb
PNjcPa1icHGqbML8cm/qfpG8tm/gUKZ7lnYS0tV0DvPc5VM+zJArxU57wWmypF5x
tor4sN48ppYUplEw1XtKU3fcMu9LwuSYsF/SoHipxB3i+NqZ9MxZ/vGNPmu0ufaS
uOUuI8Z49xx+2KEpvDVtOg41mjep82eNEzkHvkb8cVHAwOJtMt1LA+w+0bAaybNw
pMofxWVWCta31RmLZ/gxHoUPteMvtGCpZ0pxNyiUrRVeua7kiSXofEtfJ2I0lTe2
N1GuI1ndfau04U+VgAqO63AK/JAgu8x/Ym3Ms8qhKU++v5q+SSPt66wdt0c2OO/u
7zlGt2GKaXwmmHOHSl77sRbQd1TppDdanGv4skJ4qkEWaH7pyGVNy6ehJ7It1gUH
jQ32Y8emOrVuym5XinTod8AVSlgrb4KCAhsS6zqCjSAppE3zqqmiCNAC4m0mKYdl
Eu/acSMH2kMDCAmoVUOCNlwikdHCcFONR5WHUWLdUyjlDLzhowa/oFmnnMCjLO3P
UYHSuvS1+pru+liMc7GSaANOar9u/5JCSW3rQJJ0KfGT0MvDSpiAvBrKVpy5onL8
RQWw53l6rHfAkG/7yewQjLzONlpyzbsuYpCVj7m4YNVebFokGg56HBS7JWAEoCEO
d3OQUbA5FrRK8K2HDFRQOPvgZLkWgyDpOnHHkIShYiSfvDeiCLIFtXVJD98FTzzc
ftv60dD2gM/qOMzH449mXEL6CtG/A2CQLfuxzDA4CElU728+wZ/GZsMjRPXzXUTR
Tkt95ZvvWtEn/wTR7Rt02IuNuj1E3OIwwyIKQEjM8ub8qxgKE5F27p1WUgpJJ3oS
GIE45Rd9a0f3Tt7cOQJ+94c3qJcrhaoHiO85PLDEMIIHvDp1Xjs+MyDguImSI6y7
rflGQrZEaNZCUU+2+s1gt9FpM/EkUqFZ6jHceAjOYilRt3uHYCrG5iwGbLYEVJ8a
e0t9lSWu3R+r55FP6/PRJGA25SC4KBMgzu6nF+sZjiC5Zlx+r4bDGkjGedty9pq7
lXLBE5T56cDXZvxJKmNpZdEPn6j/TVse4G9b7vRGq2cDGBQ5l1uKBAaJBO8e0ziq
aw1JGi7YMAZkSbTqvTBXYPc5CLPRqfbFadUfrpLLg8dsiAYAPfna0u90UTRylH9d
uND3kjJhwB5/MStYd7Ab8q0oGjAawX33bRIQ9NCKc4TwfXGm34df9swDXvXsh9j+
IW3MEKjwrgp6Dci4gUxuGK24+BPibBwfNKXlzUJzcI0N0+ppfMjs6UQLR7+JA7dH
blosC4kqOjewe4GtpeyITagqHx4M3VGo0JKv75045Z8q0l5jQsdm19nQ7MQMKIZr
1ExoBg/ZiZpG+gfifQCsedIJ9IoZYbaHCi1adXeAFNEtqKRJZZHt14Ogr0Drv3PX
Wi11x4SosLc9c7d+gnRa1RUlzeAeTSeKLRUw17KJbsWafl4SjmutHZFs8zjtjYCN
GupCrJi7b7R83H8Wm496J24E576ebgomn+92NS/5yl3AhgPra9nItqMJRE9KqV/U
vCmFckbHHdk7gpTYfT0rVKYRBasVTQ/pUJha/5t5AiLsM06TbxwZsBiMSmGXiPai
WSUIDIWPFSE6q8j/N7+PcFAq6JSRoV+MhZ+FEO0h96WXfVhMQUjYfa8YZehRNy/y
uXJU4q0VgDKu25Bh0xDaQT8IaERBsUxDMdixPV/3c8rxr4ObNhefVkybnDR9g9Sp
Fx+JY0xhNAq7Z6dLznbgDHuYKrg9xoYyYv2DurOXZkKXnMrauNUmk0l+V8c2iPjc
7XoFxOLsBlyererVR1/t32d61KZ65gQ7O3KuX+JkSlh8hVqqwKEp6drT/TWsvQz4
w6jhL5zeJdst2oBOd8rPgaciye5mhYnp0H+wScZexRUcL5j1JiKNyfC9BkknNepR
M3XVEEbEdAXAx0fJyA7ZuI+PPWfpIRtxiC3Ut7b5YlANn58uS0XV6m1wfA3ATh0E
edI/NdXnYYjv72bJBWBtFdMrUbFSKO9PY8nQ+5heW/pTn2ZJi5RfCxoI/hoO95LS
dCuO4dgJDBrtqUDFCVc6hyxUDP4np8Gd2ID445+5Lve9W5dreXa/XjKcXODAtPNU
cS83qip8EZP/ytBbq0GuB5p4u9ocKnflN5wYuUs3Om6t9cXHkOpwconCUQS/k23U
NwaAVBgGg1XGooJDoevdnhgOgezvmvwOhmQtR8lc8CRYyXnlzU8t/MUGa1L/ttD3
+3uU82XJUL9gJMfzTdleNDjXASNFm5xgf1MWNJkyR/7r438pF3znm31ol3DnS6+f
oX1RmmAWExrPW/I5N45Ks3IIXx7xKYVcSUzImnCW1M2ShxyMttheVhac4e3zXja5
MJQCDEXog+/uc+28UVpUaEDINFHgNI5i9zCB4iSpe+DOEtCvs7hRXafApKSCBYNS
/rry+BGloUhvgIrKRhAZH+CKwfNnpxC0VUeCm2EUouDL5MzVxRVweP6cF2BgKKGM
XUs2g6ztQ712k4oCrD8wLWxqFLPUagD06siDVzc8RI+U/mHi5MmBRRhxiP9OgXoP
pUIjZyeVLZzDSqXmj6mqTwbjjU2zhTOYSGjXiv9Bui4MVNz0FBMhtLbMHb8ZJzc7
Vou7zxZPGudbj5YvZywziUXjkuziLmyTgfu8/8DdEquttIwjUVrDtT8ITL9qovQC
izmj0oX9G9RLVAWTAKlJaJ9fIR3gn5TzaEVaxzy7V6Xm8J+LNcQReW7nxbMqjiXV
6Edt0RolFzv/KmZ3X3/cOiLb0Vp/7zl0KqGfQ4IKzqaiP1uWBlLP3GxayLDzHr/a
j317mMjduiJpJ/Lv7u+5uQJfp9yTwUpU0kIs5KriYUnS6ICrGPdk/r/r81qBy1mn
LSlydvZKaSNI/xdB0F7b7szYTTu86wvP8qoKF8MXXfu2LM2tXRZknB3SDx9wqyNb
os5dX2fTy7BhNHNdOxikWnEu4S6p9xqpNWawK0vW+927evpSxtNPSFTY0bmA55/V
pu7mihFH08l+xHU0qGQgJQmd+tnitgZBUg1Fg6QM3OUw+bknmel1F7umSTa5Saxx
/OhUErQQCHgPeurVPnwvTzBKMYnF8SIa0QvLaf5C4bWp0cNxNNDlA60EyZfcig+B
+mcnoNwTAyQXdqnq0Qqpb4k+Qobt062+E3+ZiDAYpxj/gyO1VZ3rFq4ZhTDWKfO0
vtQLgJeneZxqDxKKkylb2mtk4E6ZK/8yhUZb748miducq7yjt+NcBxnigeqa+EWb
g4qSQ1s24o90Td4h2PO0pwY6IXpGMioCyWzGRCNBBNfzjpQ8RnJV6X4+r4JBpcZ+
PLwabM+neUF4ehdjLFj0VF+imvS1zHLo/4G9RqyRVDWCAsL4c0CqimdtanRNqeVH
0lxE8yMNGt0zTZTDTaqZHdaabcuTt76LpCipvTrd2VC/LLVmEpWIvUDR3qIEjqk4
ZNetaheHnmJ/qFhNW0rC+yPA+EBGmemu7GmWUpsIQKtU5RAyWEuxlmGh38hMsTgV
aOV+v0S3xU/CN4kU2ysNJ+/DDm/5LHWE9+nvHVEOhirFOepXNTAxzC2HhwpBvTXS
l9DAebpa1nX4DRFi1lCLYtmqcbEXoCNGM0onog4PFK2rLKxxzWBPT9pvhhEAp7xf
2eqLTF8/mKKIFSd+EUjZeq/WBvNvVZeEXkWQ7U7EGIHmBPvVFNSQdyYtACsYh0i2
la/wKJGXTJt4Aqa5GqPauk/b1XnD52IQoS2/m+M3v1hO/4E2lBw9HaiYgokPwZl4
JRoOqjEdAQ2Ky8T2M+xDjrZpAabtE98zaNZO8Ll92/2nSZiafsMA7iz3/seM3CtJ
o2Tu608ij+ie6HyV7dsmVBursVljbITl1d05lFebTHfXELX7Gn3RTxeW6z4pVsn1
5uM86FSZuht8baxzf0owUQON+BzDl46azlxK+NmozcaCUBmR58dvrWZsgIAVv31+
HIU10jEsc0YGmiYyLNnvHFnLAJvJ5vzbj2JKHfQMwuQzCNE+UK0iMM0dke0FzLLQ
krlcm9hxLsRjshdbpTuDfZsPO80EH0g4k6GbzAG+Bc1bX3OCJvCZaLmeMRbzo1Lu
roKnefRKfSzyUvJM7AKOxrhQn2qv1cls+DjFQ1KgakS8nJ8O3OE7PyeUeQI39txj
KMW4nlXmuzvZu9m9G41M07q+AvwXoR0hPOhR/8y+vBK/SgPzD2iJCRW17RQrpzew
0uIl6O6BaRyz/Ra00FG+njr59QRd6P2x+8mJ03F7Yr7UXg3yj4+AcVC4Le+el+CJ
oXrE45nI68H9osJlkRHrE+a9w27JKVk/56Nfmwsn2NUOQHbhZk9o/t3xPKDsqtuh
k/Urlp19FOEGmPED9yod9s5rgM/6TUPAXM7RVFdRfeW3dCh73Sxhv5b3qsz+f8mp
Jg6gTePxlvxXkyUMiLAwgPZA2SjndZ+p9inDJ6Z8wOcVvEtQi75j9BRckSmPlMcW
w/zvRWHWEQdsBcnUyqyRcReKD1zQ4RL3Z6vKwQatGiqS5UiJq5F4Ffz6uFFhhXuz
qeHRNA1xY2zBLaWoks0Jk0T0MibJyl5VYaGOh/kAw3FIjRBo6CfLrkueigtl+eHH
oFFWIQ3oOhAiQ9uIHCCmDpspPnA1cm/Sa+bnpNwZuIZvMQvPRAD7tP33kzgkOB9K
03OPD4enR6tGxW34r5vw8R3MDycL56rdBy02pYM+hGX4tO4HcaGV8OGsL7ufYxMR
WIeUa6yQOsU65tLFoYkPE97GJwPs1EK0j9pFsmYKHkFTsPdd41Mm49BsyfpMCMUh
QueDsJa3u5u9MPGHDThfNQk1Rq7SSfhg6m+nVrj4ef/mfqh3uHO5N3uaCw8YuuQi
1MRzBnfA7KjpJ+T7yfvXDlntv/rVTfuC0lc5WZhHVRmHLVwDjMbboryEvJDJcDwk
RcKRHB7083F8TvpFtiPl6fT6W6FpKZjAsIikwer6i0GpACBgGqOjemU71/xbGd5I
L6B+9hlbZgpSPs+S5k/2veW3ZinlywQniwkwJCiPzgG9JGKMUc0lhkM6l3VFb6UE
FXYJZpdsbNz0r6iPcfJvHeUbWSAIECEm4ja54jOi0WL1RJipoG8GYyWpGbKohmJG
QjFjjNLVrv5MntQ+flJmY1RwK3253ZhuDRA1rJnCxQEJE5Nt/4Qgzh/kWNhsumbo
kSqVRKSHEzr5CZTMUe6F/Ran4XqJXXAVSNfOtesfzk63UDgFxZi26UvL8lZG7oOs
TzvFaTIRiHdDFr9aNE2DSQoxe66GVZrO3qqjh75zsAUTS1d8jvLVO9LrRIq706nc
C6F4/U0Y6dPF4VrxM9Oul7baZ9Bkxj2wNKfUUcic6BQji4oY3BAKy0hmVxKX+hpe
3LZYNqI8ZfsUdgKFyumgCDP24eSbw/gl1uRNXZiXKnAbn/gh2b2g4ytk9kkaefbc
L4e/6kDE2McWNhEzil3vRaj1fDEfXNcnVmdViJZy/DihiYBvl1cHgIImE3klfNKL
1TNEwpmJlBa2PrEquj7in+T/fQ9roatyJcOXdKoXQZNDPtHXqFvGKeZL71GpJNjH
ZYIMwZxVBl0k+SsaZMADgDGgjWat7omvCBlbLO+0OUYbq+kuJY+NIQeLRRLnfBHT
8uP4KoSe1xP1vCDcjNJdpSIZH/FKlyJxHf9NwIzlJu9yTDnPMxqhdaXgYeksezgo
TT4ORG5OuGl5o/hEWWp0z/egkNnUNyVIupIov8RmQH2hhmADoUIFc320TU+IrFdL
akzjD39MQhn2n59/9OSBLe3M4E+xMweDhM23b+El3b6JOwY4ALv+3PpxovttUgLP
39gewrwH27qPrqNtLjNPj00NtBB9OkSNT/TUn8LbPC0o1AriOc85MS26CvfVFAUw
Cpan70j4+YpzAn2F09gGht5ZQrB5BIcjdU7Wj7xOygD5YevGzxaFzv4Z0U+P7DDz
WmV+pxDeGY+chgNViBVnCbCALB4iB+oYet8nA7wUTjn7a6E3vYFEBxugk9VKgqvG
imZXZkqr1ARlW0i6WhtIgDAEcw+PvdS1jVTTfG3UtDACQMBe9bVPdyLJwUQ3+D14
0T7CzilKvyGBixt6i+H6iHX+K5bZqST9ZlZa1lAYFQfeldt6NqgGF4FzjjnDA7BE
8JiYog0GUWXpOXt1FZjnxr9wd1fr/0VFxw2PgKsu3pnDGC8dQb3VtEcQAHNr5sND
WGGGHja+zL2Mq+iHZOkVmDsKU0bE6kZNkO42CW3DfPnWxWEtuCzvZzx0Kb6fn5U7
GXYuG8o6w8HWywbFlh+ta9XFn0jEXdAuVp6JxJ+0G+SJuFSeDTpp0bcb08w/gZgv
7SiOXH1UuFsL7om+mpK+UJORJlItmtW5LShldxh8tXX/gTMpuL+4qcPZ76fWPNED
4jbe9vbfk5FQ6OdZuRuOc28frn+PUqOJLxtIw3ERuetXTgbyCHX3wFQ98bJm+NK5
bD6v0dm6bWN4wByhTjvOsCFx+zdYGkT2pXSYjQVslvM0ULhF/dCS6WZWUINsWE+h
o+VGiG9go7JGIA3B2oHj4uMKXrPRwtYLvHwVmtCKnMAv+GdWmpyzzvNeAIZLUER2
eKT/FbkWAja0TsO2FZvvk8zJACwJPOY4Dj7J9VygB4i44Q3QFFbjiK6FUgdDP01K
f8BToSaHoC8DaPnt5+/qbsATKOGhU0/f4bbym10k47fZZkgFzbXi4bGHFMFEv5Lf
I1LrAVeNegOte+sIue6nJg3jWEvu5UH+6Tb3iAJmBp5a8UgMgE1iFceRQ0EDDsU2
bL5f6Wi9Ifhx/HEv4Nc9HUhKRmMTiGydSQlON2dod1IFMedSRFJl8xjWbSFAdu0r
bP/X/2LM7T/gjyuqXcW4AGNxVi793APQ7eLTLHmLVxiDRhrJVfUbNOPX0LWhCqeG
9CJ2RgMxqdsKexxiZ3YKAh2AnPlKM0DFnhuPHpAixXZYYimla1PmUutdkFRucE77
piWW+u9BMBhao1U2WaZ0JBpTt6Qi5wLU86NhvpLPbnm4q3UtoIwSEOj9biXIRpzJ
nMaMdpDQjZQ9OK89MLimIRRT4MmAuSuV7mLNhNX7cHdtQjY/C91SuFOy4ASYFuEN
Ex+HeZoXcmeH4rq9jssiSOE8SC2NzhQDsXrIwpwdHUkdf5w338BTWvYU33M8IwSS
u6KgZMEyGTmLhnpJhVuTZk2H+ufJo5hhS5skZe++uFGciv/q5OjKqPigLlARQV9x
QrSQon7dBIe/3mWT9ut0bkwc4sJyqwvZQl20O4vkht5W0EYdHt+PTuB9AypYMLzA
zxg5pGIxFCe0YRj+UKLedhqCzmePbLfIBIXFIvVjE/1kSGKDBGAV0OzD1D87oFSd
xZu2vrUAPLao5yidpjvYFXM0EaI4KAyVYM9Pmwkn2aLFry61Ko8fgzBfBHHsKhs5
RyFVvnPOY6qoXY2NmhPaXtrdu9WNlmaZrWENZqY9YqLGyAltbLKH+iKnm+k/ydx6
C8xwhX+ZdDM+zhM0ZtOniXjD3XqbEu/PkdWfSwtdGQZBgB8fr+MFpQtNNN85Mf9T
KKfhU4PRHzxm6qS+JdHZOU+NNn86UQSgw+MGyl+8INxlYl2qwkwatneihraF8irb
znTkCkmI0vn+o9VpQB1eDjoL/WKgc0PGqGFdWkEyDCGRivQPNZMIoVLUhjlQVmvf
KqH+bTSwzgsoRch8oxs6K6a/tUlCh/5CR37XagjwMTl0SJx+dWtGkqria3f8ep/y
uYjNLRYHefjZkuCVYJGHGeWHlx7scR0BXPVg4yTjWpLdF8xSD7XXcKNkxCcAYybx
G2irZ2L4z1NC6JKFGNICWikGghR2l+qnBplQFLmMIN9kAvah78CiEsowXmHisJ5V
7vkDWMWOt6gUEJ239iUek9/YnJbVBpsvAuXMWLX4100hSJgKftFW3DvJj9fDG4iU
O6jG1SLOLbJ4fkzu+2nuTFwZQE6EMeFBW03LgWQ1WBDIOtlR9e5QzmOc+ToUsBhQ
dAkIjWT8EYQHj0JlR4xXUqqmNlVjfPLB/Bv3fL8hL4eS2oH9EiC/axinyDAWxnUt
R+mTWla6B4l5Z/llSyPQ70tV1omSTCmxMLBsU2z1ubMMVDKK9tn8ZbK8DZazEgP+
q6c02DQUa4VQaho3qhDcbKak/2KZAVWLIRM1tZ8Fpp9xDccWN92ksQ0mfgbtNQl6
`protect END_PROTECTED