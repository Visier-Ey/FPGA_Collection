-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "N-2017.12-SP2-4 -- Oct 23, 2018"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
A4Qr/K2gXIbbXHzDNye4pyBSFtst4Ye9kxM2LsHbBN/Gv8ZrqqMyr3rDm3T/H3M/
Iih/sCWvAVyWlLi7SdXlC7S40GC7BTtvOzJ5DzakDNjeKiD/f/WUkAQAnvDTKz5m
uyKRi8OYJ7tMjLbHk4hOwhH/APbv/7W56cLKsxqiDiA=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 6080)
`protect data_block
xcjXICTXakDBaYrVKZULAPpHwab4KlmJeTeaghOOWBOiXLKP65+D8j5BO7mP3dm+
U/v3hZSmqAq2rS4fpfFFK4fMJOPfQncI3/TjMnnepxsG153vt5o7I+dZ3e5hRFsj
na5z/huCWFw2+b/WgfxFmFNFDDp15n5kYtF5J+SbJ2upipYmFGQ/AUKDVL86eSrV
u8AVK2LqyniY718zYFgYIfObfeXnvnJsu5q4XVnNhiLA2DQ4JGov5pmtKcbtno0V
zulZlQyk7ZrL7Rn1MZBMEk+X47HORZyMsmqBaDZrHdIomPe8p5+QYSuuNbcHy0X/
86R+FdHoE9whtJDA9FWjdyEfnVzqYqpSbXQ8gZgA4HBgi9XLDLz/BBEmQ8xn1vlp
qRkAx5QEQY0MZiwoBfU049PdFZnyVJxqSZnNCXMmvHsKgQfZuZgMcXhKxbZVZIu9
o3O8QxOLtI7b3SbzK5mr/vVIEWvdYm+xS6+rmnjYoOVPsAXTcISycPG8QhMJrYYc
MCBcvwnstTDYzsD70L8S/A5HGjpLT+9UlHCbt3r6UwL/0dB6EE/4GjZiOJKKV0kQ
lSGTzh4Vov3LZcerp7GtWgOMKd5lJ4z79pM/Oyq8oxwz5KsagnJXV1lYhk3y+JsQ
b2T+/p2O0N4dzheHu0yT01JPj7BER5WHNxRyuh5VSLFywhIrHtRLem48VDkEKlng
XlWaVe4SOOe0ROhXElvY+HsnJvXeZCvZadNnVU+X6UhGIpi3okQTti5wMk3n66jN
J3I6QIw5X7+s2IVmCp4+jC9RrmxAkysf2e0H+PNLACkbh3iyrW9GGNqkJyroRZUU
EKZAinVeHpmifzKXW4f6+FmZp7AO4Btmv+1DtUg/2KNGJiVPZLtVr9zqnVsK3WOA
yTIy9Lvv9pps8ZZCbKq0y6bOXak+yvGoeenYzDUNMrdU5rgLH+gYVbp8qrrYJqZL
jRd0MVp+zWFljBUTMVFV3bG9MDGBhFA1lBNMW+oxvfLKxnOMUB3oAocNDC+Mf15f
tWTppGsb5zxeiOzv041/EzJSLk2cojEXDhx2bWFUcabSJYypmmy7ySRj6cIY3+6b
i1T1ELgrjHlmN3JOoH0m5IjXu1JlEF0VpyLk198SZ7ouLUl/BN7aSYquJAt9PTFT
k8a8C+7JkvIaV9QSzvxEqdlzogYJ2iAILqNANaj6uOESKKfcEOk5IIJJNW3OdXxz
7bQBwTSdlsIXQPdKw+EUtKtEWk/+h12CEhMLV22IBVlq/tS6nPb+hyvhyytLhC7+
/ZgA8gIVWgQCTOAxAH/guy8qP+SvHpO8ZRLSC0O0r6Koh3B2CEjrTIL/H24ta3Gq
qE/1R13e6AGz9oe5yJOUWZihfL509/VVwQMayHTdQE2oehHoAxFGXof7tH0GNe96
oI4pwDG19THedgvHkDcNSjaEX/v3az2ocVusEBIkAP++klnkbF1iSUXF57mn4qtf
72Btk1cTpvceHJx4O4JjzNI5kWwQ4fSEk2vKnuFKTTpdmgvs7i8KKoNmYlnnjPkz
FuXJqjk8tIScLUlgyPz+sEihlbhkBG7+7i9m8GZhBxDszotY/szY79Cgz83DPSny
b+5cwvDyTvhfhZa1tJB9fa9jEoJGYeTllAw4QzUjRhcNbLO0ZmySYgBTp3dHnPYF
p05/gTFqME0aGDIc5qMl4NqdiToa1VS++2g9yOX4KWdGNy3CARlfAOdgtUMU4koV
ROI9TJfcnTqTJM5+FPrm4TS90o/ZF/OLmorlATcJg0KEyRUlDLHKULD5WN380Yf3
xWiNknJ4gyjoWr/8/4axtkFOcYB70av1zIhaWj/hDl0d72QVF7elKYspdHOJtnUt
tPGWelxuIJNxKYjttfZhL0or8Cn0yqW4XNvKVgv5JTfU3SausfN6vj9ObCdz7fmp
r/cbJ3lglQlmNKC1gKPhlV298zbAVxC3dVrEvpcuSF8zcHvgpbZSOz6q7FZgNn0p
+pQ7HUECMSBrK2jMEOHjQMiZBZE2cnpJux86xgcHJ8lOotDrHtstOFqyMD6WS+LB
iet+PH6nr5tAjwgY5Ho1on9LdIP7nG4b57P7AQcvHQVA7VETBTWrcGuI4nTLye3n
Tn68iFeHbfJHYaqTpZ3xeC2nNmd9YA508u6oC+eOM0320WoVtMBrosGCydkJZ8JV
N7I/O+7bKJJ7mfpJqvj44wjvPfCEzUiJNeJyEdreZeqSZPZVnxv1cVKhaztPgDO8
V1AMRWf7CS+SqQBNqZl5+k3x4h2hOXD8GEn/Ah0SAiYzv5FuEdm6YEq43bFhEJ+3
QINKvTIQX6B8OMa5oTky8ctNP33IL5kzMFcuPkalAoS2kgoDaoJdAk+MEwvyiWuS
LKg3GKQdjO95MCudwvjebcS7R7cfkXYrrDwEydIsHwzdQHgDLIxmvroYwimYsWDS
QsjHsFHJ5V/10WFTzhIHT/XXBiJCGuzpQ4w/QW3W4No+BtpwPqKlHYXH9v9TcGpx
F9ikRatFhccYNsGKsYHQGqn8RDSLlDO2Uce50wIdbIDV1eyE/PdRUBn182QcnI3W
Vhs4auhfnTYc/dWIX7xAfrH7m3wvDd0W408eLDpQErDPF3k+9hZXv3JcYlmOd92K
PogDNv6KpLr9rHMZlDWC5PkYidm2rmVxAK1uk5DCMgmKo/DMSynMuR6WwtE1/eD2
zgbp/VnSaQVBrpAjKpLQOxYEHy/D3GAvnqBYlm3+SV7K5BPN+cHtIDW9uDgzmHcF
N3HKnsgKtpPZjfz8rbcIotMkU7Ukwg19m5yoLro0pzjn9lb/z2WnifZcAOgwHPW8
Lv72RAac+PaYTavEHZh/k2QZ+aL7N+C7/2mpJBG4Ym7ANRnvzQQ9JcrEeScRo3zd
NmrLgj+OtXh3yUR7yD2CyED3bEqNlOgVcemUmKIseQXzS2oOCArsxYmoakW693E5
yn4TXQ2XUHh0iYl3OfGJ1XtrtMiqvHnaTJPDhVVRZ3+zcce/N0fbkfCif4X8PUVo
h2zQvjHkxZHvqtLovAK765POkoPz7orpT/1vonXLQG0A1mjIe/3eoSQW75gbijmF
7wrlfhGhAh3InYtP7s0u67292nzSXsGZkRcDLisVOxrADqocGDX74vHe4VNjSQ/+
9xVhO56EuxtnRzW99VBcB4ODeYHQ5z8Jv5ntD7SjyT/o5X+1mLiKBGkY4BPDH24Z
PZEQlSANhUGzJKWR9VHF7R11kabjFxpEFZ0WZxFOZQy0H2rX2SHMiRZUjwJUREfx
qVaUpYhqm1K6iot1UE8T7Qu/l6OeNZ9/+GZTTCOwbJsguIcV1uqIddMOdvw6LACS
jQGPUCQ/BSGOfnojr4cZzeSCYxNgamkO9yse8WHtVDfF7KtlT0Zv0Vd039VTKPei
5sl9JAKAfQoxGJrW9CKTDJ58OKRS0w4THIYGHckOCLVqKEUMg1996SBnRccO7M20
fc52IGii8Iqc9ox7FT1daHaqgxv+fEUsklj5QHuDgJqrIJij+LiSW/MNG+GkGpPZ
Gs0XYc+VGpOyO4dVa8+F51R9pJZ6c+Fuj7Mwg6rj72vaVvLlB34cA7WiBjFdTIfx
et4PCNQ03Vo5k8jY4+QiIiRWLf8hDicNSMegLX3jauOrfE/nbC2fs+vsdnrQ4qhs
cgSZoGYYtx6VdOaBXHQ/o/9Tatu/mrKcsXAUJZ4TLuiabaI6yqqLSU4I0qBmX1ys
TFyNOSIJrOf5/U4upED7YBUzQ6KdB6p4P9+6h90B4BYnQ46N0Utj6Hg8SvWZuavx
Y8B7w3GzoJXn19PXgwMXsdfMwRH3fmW93AlgGgcKWd9HeYEnvHpoGmfogHNBBymh
4zWfEyRV2D26DmqTtQ36WDNZXfF/rRlgAbPTjAcsqMs3mq9i5Q8GhLLn4hqUT8cO
kQrKQK/0UULJAIYPbbBcCyLfrjP2GLf5b1XT1XX/RmlZ/R1hl6Im5B+oqByQheEf
KdYmyWxvujxz8OmKAi2v+h8X68DGtm2cQsw7lJD0UApOwROZK0a38MMzSVf+rJTe
IrRNVUjkid6JinqeZ2j/k3JECLOI99dWUGch3lW2kKue7hIWB3OwPj9KLrI9Y4gY
Xtr9Te7++r2lPR3OS9dhXMnPw1EGErioHcacd+N1fDxm3B7Jxn5nwS2fi7O3PP1q
Ak3/EcmtKulkHWiOVw+yb7ozwsYzgTpNMhratVmBy01RYS6h259lfwMUNFflytXz
y+ndSkw1/1Cuu+f/yA3h/kPjqnUEQ6fB+Z2Dpp/Ud4QTNMXoE9toBvtlVLVl5/Aw
dALLq6BVd97Nj7fzvSX2WvKHKusZzjDoGPuCXNZokAF+VFVgcWbpFE09xmSDLW0+
BFrqw0Q6y5zfUbkWmVL/I131QiUrcdKDMwmm0P9SZrq+wxON6WCt8jjEcG4R1mHF
Sx2Vn5xPIT3hzxvS/LCLvIwoXIsMXuOv/jsDScZhR50LByZrIXqiEVYCVySETXLt
MR8rZkjkHHHODXkP8jyYjA8FGAw3cC/MIFsWRj0RdmYck9j0oJ0PJaYN/E6b7OEx
w+PMMrtpqIIvmmlJI2DUFEUcQ613qPuXT9gbL/RosUUpbELhuZVVdtzHrkeK/15G
GH5RjEA4pIwlYLyIDw/69gPfJ7csKCDQx2zcLDBb+jdcGmIgyMOLKZcRlYj42KZ+
GbexEhnLofvdEtZd9UJM/+e4pQcgx+v4brOA2HoqLm5eI/dSo/9X1l2PajUwdGJ0
k017TIZQEEBjubVjxlFfpQXsCqI9TJi+pTxb5+c06XDiX1bNhzL8hRWfhibwacKe
f39i0MgehNzXQ43GG6k9MLpMMYXs8FyhngxRGMg69th9J/8zFX6dArn9pqnfIgWO
4fOFhFRtZo+2KKh+DRxrOj9/Xwz1sr2WCmstX80JBk7c5AQ7DQkdo49/z1mS590e
vEO2kPBzwLrCDYD7/rJmQBbMWJ5GtyfG+RcDUL2FyYsaesJZ5KWI5Rxp93MCw9W1
hfcDXnYCi4ox/xDbi4F/ZbjNIBXCgh1PySHCTe/EfVXLT7KOp/U8rHGKmShfDNjH
vtPCIwGvDfR9sPOaQhIO6Iek/gCW/Chzvg+r4Oqg3jtsZZdaJzF1WfV/d2RCLfry
qfupsJQm3S86X/u7zFIpXiQg9sEw3YZv+5XxQmmWFfu3sCybNa8mqPhUwjGgTxYu
BfJ2KQKLJ4I5+ogWrp95WoB+OAtY/YknOgy1uCkGhHVJmv0l28M8UJ5WK+JOKnPM
MU/RYyQ7oyVBE/tyRPb0kdU6tsFNSkh+W9hPvqGOhNSLC8Z8eEXRXMskysfUQxUE
xXphEEf2328KQIkMNch40YEp0AZWwab+nCbMIpFKvFuYESqwaj7fRm8UXo1AkkL5
BDZddnojEijFLY+VPINezD/zRNlPD8gHL3Mm5Fd0EyVj8OmOW3DoWEPzow6hvJQd
wW31Nkk1uEz5hIt+lCM51Pg2bRfah7GHS8Ajdh6hG6UaISjLvv3U/WNPmoj2dfEE
PWMuwgTBV+ujMTWl1VEUvATX1KU3LqOZZF8SO4tsDGVlyXXGRpsxa/CXuj69fNzy
KPDlaT0FDgg8ACt7ZtLl46yjGDCfXjxTxvTjqB/Yev/6QSAoT1QW9KT15FJS/TLK
mlxWETJZC6238D7XKkG/wVKzCWUpW2CXdnNix+uBlao+Vbz45e6w4tQiao1QckGm
NWDFMrDDUwIOaBr8ynlBDGHb/sHZBm6G6ukkNac1LZ1qRn4YoosEpW/kTumBHYt5
/6B7R0BlGuW+vLeIrTXNHV1ZhJODTRbNc/WTpe1VjlKShMypcAb/7kep5/+3ZiiG
r1Wq9kgGL45lS6ZDDcZnVlm5co96Sb3sTNn5s2MuDNTAG1JkTXIDQhznVPV5BKYh
ro0jqql8VUFukO6eMSCjDf/OnVTG04qwkQ78lEHGNj8XQ5lSgH3uFCCU9tIRAaGa
6Rj+VxnoupNgFzjmx0r5bxtKcn7saaw6seVlhQS0+uAyjpOtJkCKy5qePI+wl1zB
+95mBsF+IKRy8RHTsMnCe3lqxSwWCHdFUto0n1RVG/B7JNheLHL/yYEJgZ3DEVcs
6b+glVA4P85WoClP2g5+liE/8IkofXs2C8FDXVhfhcC9l/IgtO/eRJsTgYxZhz8a
keQbu9kRkKHuSBb+TAzFCvHWH626x4YqqOk/sxGwKqWg0LFEdoYZZ38fjkxrklCh
f+dFFshK5jdL5y4JywpoyHAxSx9bULx8FFNN250AqaUU2tUn5ukFHJ7vVbsMrvGD
UjvxaRgY7Xvdei3T63H3j7WkF6ahDuXnT706KgsYrXO0cPxeM3m2C6wJsbZUlefB
vrTGjbQ6bdeERG7T8dJvvJqX7ZI3QXs3etkUSJPtb7lfCIUmgVT2AT2947DOb8AW
70G4c2k7Jytxni+WYvKO2hYGMNrv3sL5hJLwQyUTYl6IViO2iXi0Qi128nIP4EEz
YK9GqtSM5ukfQX61SdVXq1S/LoqWv5qJU+mlcNGcgxH/n+MUBDItlaXUV+NkZiFz
kHTAHAhsZRyUi+0+ZpcXZ+G7A214r/tl6GF/1zxjUEx8jGcvJo3d1G00oVC2BfuI
SmgyqxKfL2p3xY1MnztJBkuk4Y/La2v8+d6VdbFRVZsaxa9NO2TYfh7vD1Zc7IBb
6csLG4EOpO+Otb+yCyX1D2tf1gJaWUXDRFs2WLf64t/ghQaS6Xr6Cp6TXzJTK1DY
2j6O2jcjLIYAdfvn8PvVOtU+lb+WS/FC2Pgl+yFQd0f1uobRMW8TMkwkHGD0Blpr
u/FZFhJaWloocjew7bHMISNrvfmmIRFy78mTsIkn6roPm+SVOo9uk5DgA4l2Tzby
XlTbvS6aw6yEbBqF9un/YjIwjG/UuJHjh2zh+/Dz1xzhbZ/kZSlxwIfsDauaVuLa
LYamyb8sCfdtgJHZ2b8H+RIN5KO/C+pIXPi6UQ7E/H6/7z8HMAF0W8vg0GAKq4Sc
c93bIfAshbeO497iW0ZLyt2ql6OoFFl+vPBW8bgW9Fr1+LCsIVqBb3zZLcQGDfC6
oc0A7TuxFiWOhG6x6tIn6FQvPkPFkv0fMy/Oonl7WpuucJZf8r8UOy3K2m9b6fma
yZ4/SC97hOatyM5CvTxxqz7y/jxzKHFKsrGgeEWpIcwwCjufUFVTiutoln4TxetE
jtJrlGcHNVcbgXOYYuZ39z/Jn1yIq1XmrHnnMPVzhXCFUyhrpPze0RhFSzhOmSih
6QvQ1uC9V7u3WNTXouxn+biCDCb+FB1p1r8g9qMOdeJWvCPNqF8D6BP1smEHUzy3
3NeWl6/5p1LbK/Dnjxdk0ENOfyKGIGdb2bSRUOLDofZmEFykyLmAPDguYLTS0xiU
6AWm8Mm/iCez1oDRIGUxNxxMEGgUiLb/vm7o/3rlbNQWLQ2DvCkKMqVF9vRhdqvC
evEhoZA3lfal8On3PzBM2NmLfxvwuZ5CxAZLwPoqop9WChRVgthwESx1o9edoFMa
6YwRMTADsSHQvoyWsIJaR+dCmS4ljKjKsjthYrUQQUg3NwZXTMTWjL4NipMw5yC6
3811XFfm6L+M5K6RPfvxjG2SYtfHjLM1bt2JSvkpbxeL/g84UdkPOXHNLmm0Iuuz
POnnOP/YVEuJW7ASzcTaAR2H0oDx9GlmsRD9DdK0oFrDyH4+Svd9PXf0qJ0xoCB0
rc1CGGa+T3BodDTQoc/fmYw/X3GtzL3fR9ohrwnBcJuKTWVHSziFPbokxqHpAxUD
wNaXHlea4/o+Tl2f8rqcxE0yreewiSLeTPlCyobfzqL611v8ptiefc4FSGVFa0+G
yg+QO/T/x7VIMTydO337NqKB3ZgQdTj8RQsmsUXrxV1fgXgT5rgE2tNU1BH7tAM2
/NFykYxe24NSmZzTx2AOTLUP6mFKkX027Sr3aIpp14Vwj9FYTFS1tDzQCf6JUbgy
MseQMBZGcFJ6U5PHL2mfA1JOF1d7PqB7vt5Pygzb+qyc3VH1wMxMBuGXzrGR3mMV
flq2626N0sA8B2Cb3y33TghnlfwCwa5DlLmeFcbbSafnO4vu8tt0R+mCp+6rR7EV
YtFTPO8gPnphJgKSOA0NWq5N3g40N/U10Q3tPsIOo1k=
`protect end_protected
