-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
--pragma protect begin_protected
--pragma protect encrypt_agent="NCPROTECT"
--pragma protect encrypt_agent_info="Encrypted using API"
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
--pragma protect key_method=RSA
--pragma protect key_block
SVk/dikU5grouctqYf7w16DZsaYegGKWIWXEN454PZZn1CT0qyziRmcDiYu4gguH
Wj8KqPAKfliEpr5qJIh2PGKtQosAR8RsrLPDoXrOInFxm8Sw38DX7yJEWhjeKqmr
48yiVynsa6Xdhs3RKrHyw4dJGIDZYGIENotJo5KorwOePZ/XgVasq9aBF4sExuNQ
onvsWJwZCSfLjqyp6ZcY5awJUXTIdHwtrtQVi2ZLCFAdR2QWHS6G5BJC5EftfBfx
/XdBT6CSpM5+LcbIzEqAzbMRYIRLf59locALqO6iIgzage/OUj5/dMqUVqoglCDd
Auh7Jx5zLWJsn2D1TNss9A==
--pragma protect end_key_block
--pragma protect digest_block
78380AKXLbMFxDlP4XYW5gJxhnQ=
--pragma protect end_digest_block
--pragma protect data_block
nSDzViShdqm9/BRjWFytugLEFehJpzzinwWbh3Cq0HRdXai3P+zYYVYuMKR9rGhM
gBdNluEmcH9gZAhVQGQf6MCUrfyOcVsbo6gvor7tSH0hCuwac3pC9wjdKPn7D7+u
hHpJ9Kw3uslc3nv59PXSEc1rESxNxcCu2FTunzlF7BC2m15H2EeQ838y+xsjAB8V
2PQfVw4U8vfXC32dRLNSYCgxfSl1+I6gNPmwN5HOYYOfyTMcsBFfRBVC5eWoFz8v
sJ7O6Md3aUL4Pr4WfnRa41tJBjoWPdTY4XrRSQ2NnOdGyPVvcB4sZXlnB/Iugy96
60uCScPbrqnRRW522m+l1balufiX7t/lO+KicBSThRSLouoavv3vK1z7o7+5b1iO
eOLFjJPKMuF4IC280XaHdFsrkb8z0KPFZrGrnuAjUXY6rvXTclAS7BcSaCGTexZM
xAIPiyXQBYsdNGNsYsTBJvYAoJ9kpqzvHOQrMFC88tgEnH/njM/9j4p7XEcxbx+h
DmRnMCQ1T1Kumu2aRZSCB3v7DrY0ybqYTmAXgyUnCsOhhIxG4uTZOoqSPpxAl49n
t6ELK0fLtbTp81YZprYJ/iPal4Wti+5ddwMK4MpqV0HZIqobOoN6VzYnWdTumrcJ
gzl2iGnxBAYs+JfWf8a+u/Yq5LI1d7CQ0wFZKFK0ZDL9//WxKklXlQDg65+RSsWY
IhyKdiw+Np7l0x1nVR3veRzhvJ/eyNuNXdSnmOSvN3z2rGM+GF3hKb7v6RWXd+ba
zIdQuet7B4VQ2hPOj96+/4AkoOAPJuu13ajuqoF5vYMtcdRqFnq0TiGf0/2cGZbl
mCPFeJzB5g2VrMvZC/JR6vEtIiyOhtIxsmTpXoxGy424r8M8XzY1wHhqUz/sbrjY
wDnsYbr38GFL3hrTEBl7L/uRuYG6vysViwU3FNNprTAQMwdHOmUZCe7oFU+QZ/ru
+TzJe7xGg/98SgpA3SXeE+NgiQrS3BMheRhOE2E+gtDPDiuFgGDg40DfGj8fbZrc
HKf9Z9VIQDMI4IuQhsb8BDft0jlCUK0sH+NzOBOG2v0gJIeRAR0y4wCB5noVlPIP
nM0GjbDZNfpjDyYetYVN7X7cGo1WCVeb49ByxPYYTmFFqf2NmrQPY0otGxMs/MYB
bXmbszfeYsm0tzLYMAMfTBDW/30udi059oEWIjIMU6aeldUzTOJ7EkLtSyO1ITrf
U3TCS2K2gsxQH4ErrlWvkTjtkE6QIj5n5moT6dTzzZUXKvqQROg7hq732qLVfEUS
l5Xl75+cSLP8d9m7DIsP1N5GBiFLk0B0KypnMF82Mp3fG0nFXG6T5WHYhXCTdbQE
GLcG3D7x11mhrAO4jSvI4ASo+v2NtF4EBTrHq/0Gqq5HUoAUuS+pGHlrs96Iaij9
Hm5mlR+CpnL0Se52U/cxukMlV0H4Vmvn3Kws7vLwxHWYqoMeiqPfK049jjBf3+YV
mhLpcmWz/IZQhJymqeLLOwgi3BvUCwRWKNpqyaFBp+oVebOtRAAQzskoraljWOwh
9Daw6PqOnnK2UsMWJs2YgMs97SlYthKV0pt/jrBLrhnH1nh3BPfAuYj5hGsbt0My
ktVUjkFh3Y6HGyaEk3n0YUGHR5bQ4Mwn9y9uLz6eVZFw1iIXi8bobPhUFwXHTGXe
H2RJbj25R/ubAP7u1V7MXKBIDVCI3qQjKeaFHxT4s8+OxVVjg7D0Q1YSKKn1f83q
+T/zMhmckVqL04wfI4CdTQTNaWxORsszFA5Z6sBatAp5PTIhesamEw91W0s3l0BB
DrEkHPN8+pZA+3wr4rBYbqdb3pYwbUaOQkACBAm90VaI4mR0Y0z9bc3ki0eUbJ9t
AlPrRBmQP7ZihvL9V1Pk8HcZGe/VO5779HK6UjZgYpSS0BAb2Ew26va0TdHkdzEC
aQV60gvDzlGDtgWX/uKblu62FjwQUBgOXdxBEwVucEtQKzBfkzf92CgxloNXXFqG
40T1Utml9c7nEBUQ5KVRQtPLmKtYVNSzDWey7yAqWLUg6tnsn1z5xFJdMWLxgFgS
UYjTRLS/QT5N/n9Uy9DE4ui6KbPr6mHlNyfWbW1mC158eK1+Pgg2IUb+k86JSeYV
w7ZIfZUYYrE3SvvzycsIqaesJyzxfvDSuqcR+T4Q+ID3f5DcKpjF36o/UxMOhQDf
BEmUffnmuXCLinzxaYa6WBUqN4Ii3TitHBakXDEinoWn4UeEjp0dtsPlTj8uuzC7
tZdq4sOYGQVuzv04KYRBN9GnMF+RngF2ikkVJc0z1qm3tCatwTj+K75VqRv0rIkP
T7o6TUZUeLcNRCXbdLp2F37yOa1hQmjV8ehZFOjkTkdIEVnOrtpG5Jf2s9wPH8yw
vIWhQWpe9V7mTzPq0sHqF5cUD09Y1BJnA7nGKvCNeWWM7TbqM3PFLwaf5q5Z7zhL
mc7sdYjbdOC67+XHv9AyM+8e8tKDFNozHwzxkKlZeeCkX/RSQefdI+Qq9qZ1EPE5
rAjFczRZic5hDNqHq68F0g3Uf1yEaSnD/6MOTEt5ujhVS7g4Oq7P8/rRQjA3z15H
Pn8XTD25V4f3f6NoEKMZeZhmhh1d5o89tAiMCI2/AF06QwACwBvfPPLIf8wlD6sD
sHNgF57DkTlYlxKfxejHhaoKJBmazolZvxD60XDYCjN/wmnqak5GdU/sUdlZc3YX
QmFWxzK1vTNliHzeqfeJ4EnFey+4cp0qTqExGSbWZEdjoip97JO0Pdfkovfz0hqU
HPGZUt1U+5SFBxkRcKk/3r7GrDt1Z+VE18YrbIx9/MZteh/gmSSLbd1vXnPSi9OO
YN07wVrkpRMPkTQWLdpt3M9ImyysxldFvQ2lihlgYaF4K7HrOgBhDy3TXts+WgS+
w2kBPbxDNomc8bcTHr6sT46GbPaD45AIQcjN/KTHX0OISu/SXeLwE2eopbx2aN6h
qgO9Uge9IbXyWhFzwNG5HwUenxH38CuZyvHb84LSrbHZpRaw2NzTx544WdfmP2/V
Pg7MGK++kbbGURH8t5ojArYoaRWAvIhIIbAyTcXXy7h/ZmF0s33Jk32FU3JwsQ0+
chL5cgIvnPBagEmpYoFOsUvCaSduT/BD4a7ilMCWLqcPXewEOi2bVi1y4YZlfbqy
3Y5wNS+/2BajFo077rLnkVpyx0YFTy2KCqbF4E3v1lj7TXR0tD3SefFcTg2/OEK+
RJ+8C/d4N/D+HAJFsheyBIxwYKIXkzh9gCFQxf0NfUIsvtadjDPviXdLBkNbeMFP
MVgLbYORb2m3VazS3PMu1WNosDB+4o9vey3RSr5FiGoCqlO7W17GlxH/eSTZLLQZ
5eOZQlcCYHvI0u+cCao2NX/NIJubmzz+GS7q41ypq8YX3lrw1w5fQCCwGZYapgWb
ksmlzdOUSXtj4QbNCM2e42qRLj1QfkueeqWRS86xq2v1joK4kEMcd1DC1MofVizS
HrAoZwlcOL4kFxSg6nim+gjGTXvrr+sQ4NaXoEjNQ8FekZ3LC6kCQGgbYQtZnxlT
djxHdf3POEY/SuHEIYoX0vaWsUr46c5s1HVcOZ2FQuG4KteOaakfeFRHrr7RmsY8
PkUoUien0j2hVHRIQVaktTA4bRdzguGe+gT00o3MM5cKArac3SeWyRoTnhuL2Dmr
W6awbIzh14CodF9PqXlTZ0AScfQmw46IiIG+hKN1/gF1Ku+MV97ZMH+bGzad3tll
S0T1KDPQ4fZLCOg9+D4/95qD46Fi2J7AFYn7eKtB3/ZWmnnV9MdtjvXuguvki6wn
AMl7j5C8gCH1dB/CvqU8nHUyANgXPoRCG0EuHVTHh0aEXLpm9ys2BMfUoHlHjnNT
Ac2yR/bxk+T1pLZzVfNzzUY3zMmMPPx40XtmoF/lknuLmEmK6vcOfGDMkqo2bx3R
d9mz7asi/HyX7YcWcs7xwjX/1TSKAjLnmr/dpYruDm9bIaE+DTR3cLLSe16IL/0e
fFlDPIAbEyyQ3NbFK5fEP0zrYewt529V1Vyx0rDm019JW142TfofPiH9dK816YwF
sFr7I2mScXxtbuCAY3mdJd3clJh44qLw/WUEldr1BGbHy/1thcFK2m+pp4OtqzEo
xymzokxqkblk2iay3hekekONbfwBWt6/0MGHrzAoFmKbO/ydUUgLPtbVibPbWtAv
D+nxjGU+C8vU+YpY/JF5w4Troi8GziE+g2oF9vNF5XXii925GQRK/hsp50bvhvlV
CSSfNX1PdPBVAX04NpKLkrcF13mNEiz+uWCltxOwUIyJ7/lqwujPXOVQgxbLZsOe
A+SqvHxlf9/DMy2XCv63K+DH9JzPV6ALwbmvaFadWljFK1e68AsL5sgWkgQwRjws
MBRY8U6ybptEx7GG9va4QrtUYvMQVF6+fA2GCZCcbYr2bNYKO4AmkmCJjAOmq9Ve
QYAZ1wMw78hL9tt/HsCiygadR0fm6l2vIDMuTMntge5lwIOFW5k2P1oGAkjRcYOL
rf3CCjNQZvn/Ty3UbqIxWwUKqJG0VUxd3FYxjAVT8XKWcPqGt00jLkupRfiz2uHh
wNC4ieo5DXxD4CdHQv6J7OOyrkbExGv8ymaBG1Dvw521GeltQrqR0vOga6oye7oJ
vWYrm9sLG5IF04UGuvFRPtWZ2dbs7SBONyzUqLSGl6+DcpVPJXbYOKuFUpS2yQge
5w+3eEYyOZC/gwZjk/dHm865NFFO7s9dD0MZoRkzYYjuYNfmDa/V3KZJIvbHbfna
v9voj30HKIC4zdJoS9izH14a5CKsGjlhobarYs5Tr1LnlbR3mEdok8FZOt9ANSXH
USWOxj0b5jbMW9id2J3R3EKFz1qJeuOYQ/AA4o15jFGUD68p/u83RQ8UoboToqnZ
tZEEwKEDmQzL7VWnRkY/4c7ZxF8IknsODOW+dueBQqTy8pIqeAU+MiouWaXhg8dK
BjCzqIDA+3FPbm2t+N6ZqIqpHrbLtywfnYpt3XLSljceiS0wojMM6MeXXH/StDSF
QWNpkWn9NZEOVW+8mi/ixP8HXb8m09MXMxAcHq5uqBYw0Pfvo9XwsXPcOE+E+oh1
pnSm7wk9qIcviBHTHPjFmTsTq5S3gaFbOf5s9XOnq2QE1v0L5Popft9muoU7/A1d
3XiSduBdaUT4Kro8mMjyuxLIzz9muevaF57iNxcYx+Zbjv/QM0TzGeWHLTr3yIOY
Bl+rmGsMXrRIoDhmlyBKjuiyXXMDRd4dxulEmPv54q05rb3HeY/s2Znsp+zhINNE
YZydEIEoPDGGTNO8dgwwNALYfnhvmweb91HMyxkf9bLDrDDCL/E/YWoYbJF5NMU2
cpwhPtI+L/NfjNp1+MN6BQ70pJ2WMMiKTTMCC0HaXN9RZFqNVyZj37D4fAwxXvZD
oUz2BJHstt9wS+h1s34Jlokcf0+9SIRhriY9WXfiUHTh32LkpJJDbY20W+6RRMcX
UalamudCrDoLSyr9lmFnR+c43XTmhlbSHoA6jdlqSgNCsLqAep6NlC5ej0zPkGqu
nq/rdYREoBkeMZ7PugNCLv/EHgJiQWJySpovH5HcN1TUK0BedDlQcPgctxo9nHCh
w+1KyLIfjIAu/8I7yg058qRgFvt5SFFat47gxjz3wBiKgplWiO8NVzyjMH31iG2w
dCggpo93ZkrCOZdecyWV6bp+IE8zVZGZA7FMORgVk+drwyuUjjE5d2ef2aUiLmTH
evwJlpryxYbAhExC9+e6AWihiCx2Q+sIzo4z06plJEoccZ2YzGEwephujzXqXmIH
JUUtRYJRhZ5LKopXDucUfgyGJDLJQZjcAawMYgzUfqEj02tbNXXtj30+mkt7csbv
EZTnYuE/Yj9UWohqzcsyYg9hfRdNnzFkvrxvRnADLdv/5amP9Kq+6r0ldGosuZnL
8O9dGdpVZD74BmMFfQci2iSgCCi9G2OfQy0YyMm7Y2Vn2xVXne0SjcM1QVOn3mSG
SfDKuHgweZQYeu3tybKFeTi2i+LmLIVvF7iXciOrmZrE2ghEQWXd8heDqhuDFPzE
/yi4c6VFRVGKl7TGVxNNdhr/vyXMEcC1DEUpPAybJpvyxOpZZ7mk/VA6zc0fCsLD
CHlnypEbw3quh2Dfv4iiSl0Vs6M8qWDbuFMYEoaKBPFwNk7qClF4nBm5h3uvrnOF
Ruo0UUq1155WBF0zzGr0U3z6HSweBytRuDYKxMewDhO0iXTA2QamBUUsA5shZoDv
WmQVuIrrWsDM93WZoS8TId6xg28Fi/HeT+Zg0vSVWLzFhjg9OJ481mbKE4XgHljo
cAMSosRIMpIpMvIRkgnPoAK/4/yKav+nWe2h5VE91LvAz5xQ9zjsRqoU2yRnZ0w3
JPuqOZbb0xyJZNZ5w42OubvZdI5mF8p3J/555ye15kKkaH4oMRp2qYx3j25Dlfby
yrQK2GbYK5nZwMXX4pHj5cnNd153hgN6jLjq7ZPT2AIcJmMol43Bgufh92t6F7Ko
Errjn9j3gZsovRZ96E9b+W28t87wmuQjV+LblR+76mfamchkF+cyySu03OqioA9J
hB5S0fcHJISY+6pA5eYjJv6JKZMBuV8PHlZ72H/K/dnfokYB23KFpVAIzAEP3l2C
ecmLF61DmgE9nUgD0WPh488LnlmxndU6tuLAv6MIp7Lrs5G62u8Qa0n5w0Ym4+mk
9gxDGZkQRW5I6Nbxz856ZGnPniUSpa5Vxk7Bmvnd1nCJ006YIfhZruhnV9U3kL5F
rwiEeRoY2rfl3jeVvljK3yWHIjS4FCPqcqUpSPKWcb6KMlfpT3qUMP53vk84GwR/
1QLPI0ZDQJQRy+FDEPWAVztVqILyJmYvg2nJOnV7mW4wpCAj7snKCrKtGfr+nz4W
Vl9gCyQMID7QxjO27vhpI+E+0rOnIyQdTolj8t2EIWSfOR1QZXZv+uIWjI/llOzz
xul8104m4n4yxvl/6c8I8V6ykJfsyPRezCV3MG4ZEz9QBmchdZ62za/U7nf/I+eM
ekh+UtoaLwUD+VzVlqg3il4i72zgW5KdpZ3ksYvhdynysJW+LQhLF/9S6TSxtU3J
iMWNLNZxfVKbeXhVYd2sCo6BTKPVPxq71rLMImfy9IDx81pcd3SxBLjERH5qMMM9
0sHfLiZsG39X4OaGcoHmlTB6zXKOS6Qgou6u0OK/IIxFY3LwsBpFsfi7506mm9Ac
k1BdSALoxXd/VHysnl7oN1zd+Bh4LGXligQqqg5rxBW4Ag+XOr2GOrbcneFIRUTm
bG9BmZ9h1ytpwHycCI6n2ArVXZWjyWhxhm5Yw9aR79IpXq8YP+gQk4vh/QA/DiNu
szUAPQPU9T6AsNR28v1xj5WUlnMrT7Xg12I8o0RlhNxg78C/Qa7Z2HiZidrpPpYs
kySlElFZEzavPl5iKiNyEpP02L/Z530orQKD1cy46/lBE+JFfaiQoztZtzwvCqd7
5dg0dgbmdWZkVNtB6TBx8W3GamfallIj/UMztQy9qYYfTsjoOUFeBTPbpksx/C+P
TpuG1YHT2FIEx1ttZk+SLgeMVlMIXe9FkJgd/m9iSPSxrwuEb/VTiCt3hOdzZxzm
INOrsDTnAQhHUs9zDq9AHLmA3WQ80rAyo5vjzaQc2WVbzNBMewbO92g5UccBgt4R
XGSt/YjaQOmSuZLfl0xp2gjK+AGyGVj/srGKvkE2zg2RvKr984hVyRzbjq4OVQvE
j+8NC1Xn4DZ6SDPTOX7NPjkJLxBHUMn4crQ+/KjIMDWU1sIkhi002NN3RUKO8RDv
RvQtDCIRMR6uVloTIKDuS9ErdBEKHzOFy7nN0tHFkhnK0TQThx0UeV7wbi5yesIp
yHz5oz/qRvlbbI8ik62Zi7/rYHu38PzVhXt0fV/M0UOKgbOKtvQb/Lna4sefhccv
sX2IWMz0pb7aEvOejqLvg9RWKnSPI4uVfZ2I941ZIiLF7Bke7kWfVAn0NaMxZF0T
j5DDBPaKXZItwcsJByqHizx0A3QbFMeQeadQTuIx2vEIgK7lVSJtsE+CVFM7jkXb
x5P7fSUEZWKXG5jAl1Zmd4mOUPclANF3G+qaySaBLp7l/LPFb2offYJJn85f53vP
6bjxXwdtIjKuxe/Zfc/KRPg9cdAtYgQBWIFdrhLXJUyGA+H0r3MsWmIZN49GxYkm
+2oYcn3ixZgCwkH11bACWFCwcdDGlXY3nC8V1iVgyk5Avy+DUS3aoPpGdjO5TCxo
1fA2XU6iOkcHo3xQVn4SHFyQUzE4fdd8R0E6eaWrDr57Dnm0qfdhNwjFA2kQvAeH
zGyc6S1yTGByVySfejK/GzoPGIdX6xKbu+pAwQCwARgfhxPBSibXIHCRpHQ2Ec4t
uqNXFAKIWYdmeyUAsc3zbDi7IYiXKsWBSPslSoL8Y6ZAasDw1Xg0rjFfDX9bXi1i
s/5WtBz1D43h9YxpLktV/H5g7prAi3v7IVOaoZM+BGOMFRr7fSbTUxsW4+1NSPQc
ufywgGtzT5BFWvTIsHQlrKdvj1e0aQD+oxEU9k+F0IIplkjPN42zy95tKTus/Ck8
C+cr26RVZbQktg6OCxDERYsJQ+0Ir+Di9p4yHKU2S/BD6S5LHOIvEeaM2dtylMb3
hVw1IVIN/xlCfc76y7KeFnniapqRDrLAU7iCU3kRT+2bYELsCEk88O6z7jgW/gIX
p8lGZ7wiy3GjRKbCg035OJ2drA1LepmatMsXWaheSx40sKB6SkWT1VWNgD/o6sOs
wCmKELd/O5J5zzWD4SS/fDNe7fOOcqcYtk9eXJwk6bB6fSfD9pNstgPLNrUeLMMr
yxUxuUtSq1k1FRpp9SvhbrY2ITX097nqwsnkqgESE9dKaM5iOulxzIJL05/2hNhu
676F4cEr9OgVnA+vf0FR+d4oRmtinRawgPJE6PJjtTbc3Es/Wg/iY6RNWkBafbhv
X6fh2tP22J0F6AKs2ah/8hndbL6n7a7L5S0r3o7wbxM24n/cw7Y+4zoQfQLAJ/L6
tw3/xg47xn/BVH71V6iTj0iJw0KWIA5WpFDj5efTkErRYj9UoaTeCCcs2rd74sFI
+e9evsKPKMGoAdZ3eegqrnHfngIFuC/3MrsiGbA+d6V3fqsVhdpcLz2Cl+p8pKO4
AHF7a+dPbOA/WO8niGAg8VZXlUTiePJtbzOORkl1P0pSyoAwhuiyyjxNtz+Su0Xe
i0ffWwiFsPQtHXNPDrqWZl9lSDBi2+VRk8IZ3+PVEsc01CkoECfr4Pw1dc5WhlrH
iNNqHSQMJf2fHvpi/gCiwHe9mKNFtY8aUehLmkSIY6j4xS0aOAnrI8iDmCfj0Klb
r9Vtgu1H5ehlD3jv7znKuaBAQE1v0KlCZFP/2llwTjVeTacG4VHEkdkPJQFSLMfo
oOKz8och9VVCgS0pRTfEfMQuhdOlycxIknNDxXchl1fZYpnzmk1HsbixlihB5KYc
9tQcKZhyjOFtfXVnNoVSzhoHlRlbceLdGmdB+Kji5DDxt/N7G4WLTa0JnqIHr5q2
WW/mSzzaMNKG7ypWM752VesEWYcZIkRHiebCvZY2CFsuxhIyTFdz1+Gh88Smj8k3
NY1tDHmT8M0LJZ5AYXVZESo/dD3ttIlO8R7KxNkZ2jLBXIfZmn5C92d1FCidWfMV
zIQ+mbPlSDKVr26Slbxc4xI/qnYSe98dodsyNntwF+AtXsJ70XkVRIY5Sr/KXL4y
nTaMy+U6HTwuFAQcUmlGNu0RCSjyLj76Du6sudRQOgbv21OGZVmMaCbUIBUjCyO/
Ir9jPebrR9IvTGOuO/L1/6xoEf1OVNnBDmoyYrDv62ivoDZ0RA9skQLJuVTdBQwz
QdXJaHirerc7sfpPD7bNhABCO4s+tnXKG0s90DQBvRFQy0iBiOgwK5KibUbyOx/z
xTKRqkK3WyFvCtrbaPd0NhIQo6zKvGVTT9Q0sy9NJ0sERvT1NS5olFgWsOMNo+dJ
KRoa9TRoozDcw/AOxPa7OVGpCSOQRlUQPMJMuHSoFKgrjzO654voBWk/twn75Bch
YkiTHbgc1kZQSarfLz3jqHnYD64ntbb+7a7QQWekIYwAn2nseS4GXOLslmeH2d/5
xuAS/oZc0ji028UkHO1wDKpj+HvXdya1UG3w7eZuTyoJ37/TVPLH2ihNn7LhaS4V
NVG9FGOng8YppzqjRIn3nL2oAecFPHQruoM29cTpejb7XU0IBgodUeXgXSjxzWG7
+XZiizVnAQervl5qFM4THPxU9xeRRChRYif5W/fkSw8PUtLFp7z46OrBAKSnCvzW
qAiTOcmKIW0poFoSbkz5Yi5ioeyfySLL9zHr+KAnDf3p7fWPUSCQPHAGzBkhxKMM
QjsHQfQRWTnefS/gAR2Iqe7X8sGpa/QbjMj28j47KtEHD0bQT3R1grG6LFmN+1vV
fY2AN7XthBUi97YsagbQCcGLWcITESIR9gZZ/K9iXcraxFu7Z+zR/DX6/RZz8f6s
UO5jK2hOgkrr7kQ6J9Gv5vt5QuY0jPZoZvxMgpgLdl/WsZqLP/MOt7ZiJSpCAyTG
z0IdQtPlou5/4eMTeAqxo2sd9ILxsOy1OvyOhfBmYx5HahWAASJJAPAZ2beHparv
bFG7afs109oPE/1FZz2puYTMMla8FNc9J0L7h1RSBlWMGwjPpzmXHWwsEUJ0FGN8
HOKd2Ly+wjOGwjcuos03gfYT7a7tYH8tjJAa06nWum86I8bzD3D+16SXltsZv43y
k8gAuNuwwwUvDNHd+JmRRvh0YaaUWBCiR1j5mjBk1e7OM4J75muns3vbzrEOI5rp
ibYYvqqn8vxUAUVKLLXTB5qekdzGck9PzvCDs/mbz4by+eoyEAt7H20yjPNW9L0G
gogAIS9bvl6n7Uw/wnVA6ODDW5ixHxjasGsnIUVMX9UuBlgcXKj1v7cs1df+2khf
WEytzqh6m21jJdfWMIT94mwmfwu4Y02yIPN3QCbF60wCgQIV5Yh6yxE5C4dGPX67
+rPQQlYH7CWscSGG6id202zNMabd+CUb1/mX7J/98HAqmwtm5FxOSBcepH9rqGRI
zBfkzWlOc4ya+CVmoAJlRmJ2+Rkfa7X5a3ywUZNEdNof7ufbkANkSKP7OCHtnU5J
seFaXS/pmgCtcqGob5BMWrzOr4kUTtqa1jeX9Nkmm54pbD8LmPAM0ylCx0Wwcttc
Bu0+EfU5vLzIfxdeaSQrqjqF1Uj6FNzwEtQnNuFCL+OMz9KVWCCkbxiu1/XXGHFb
LVaom9jiuF1s6NopJd+c1zOVBjj19Ru8YQqAYkMYlCFD4sIs9VzCsVeNheeO/WST
eZzbloknHn8NHqAGI05c2wuA4zpfKz2+GMZV3jKGr/vdQs4bVUCJOxcpeIHlnFrM
6L1EOmMDO92He+WYLn9PvbIkA4oxSzdWK9Q8h0c5By+ikMASxnCYps5bE2m9qy3r
3JBoO/O0ZYVp9fGg6vhlR1+AKEA3UzMulCP20jcx31wQh4mvXBuuzwzDBR9jfS0K
CDx/bI2DEYt2cz9bc1VeXkzdbo0yAp1xUNtMh16sR0Zz8kSAQ4UfI3jOtZjDS1E1
dev534dJ2TcNWmOeipSWxJmN5zbt47BPB6W0+tiMk/wx0co5te+9mbZs8Qalte2g
Z6yTcD3TeDPAYFVe4mAOPXScH8DwoA1wOpv5uxshrMu9S6yetWRlltX68/I4vdUY
TeQ6qR3zIuw0XR58hgEYJ2gfcRXgl72QSgCPZJgs5xpumtxGJAecvAKiEKt1DjPq
zcIE47hfGD/AOkZ2Fu5l7xbBxfg3/4WOgwxGgvMowu/XomeGHQwCv3RBbKmbqxUd
boxKZQlgLRDLLcmKQ1+VHXhn8QgomWPPkjG/P6ZWac3DH+3TDwumAGIEnM+Sk2Vh
DMdHBpnF9Ujpr/f7FdXugE2LaJFSyuPm2cswYnvf5RAYf1xh43XvVIcgLz3L3h7h
dfko0ssq6z80mCF0WcwOzLkVqu02iY92fOL2Rm9et6dRs55J2q5tAFAodktTd31V
J5qF+2ydDuVaHiL/eiQEv8oCsF9u3Wr79UiUSsx9YsVx0cfU14Go74A7VHlmh5jk
14dZzgJ15LIiouM1owVOabVt/XrY5jySQYw1m2pE9tL2GD2upvFJm5OFX0Eh3NPk
ZQmGieAUxRrUQaitlQ404hLc7QNCCRa7h8DeI2N8hvLAi3tK2G1NpQot91BvmYov
QktDL02Kt0wUSNnYS3e3Qs+PgiIef8rb6uEDS35Ri4F7L/vSagUKcmHunh+PCWOK
+uKYGfymQOo2tlS0i3zpaTmMTjH3cNnbJo+e9eXj0235poiMvBA6H5v2GOPUMBNo
8NGoaT6aX+9lXu9z1JnvA1SjSdPz9JYbCTwiAGQ0AIujBVotp6EGKIfCNc2FW4jc
gDqrUjyAL7ECJmtZTtgpZoPWT+qQ/uoFBsq5UjrM6fPGjXpA/A1aPvU3d4PwXK2y
N5p8Ji4Yd7WHAMUGuwwcFWmZW7ZDt2fwhXYTGgkZPWZoeARmATJgCUxzbz/Q8t4W
IGyMISb35VVxTH2rIn7j7Mr+63gH1P3aAcEAsCcrg5rAc7NOMY1S0bPIkxbGDGD4
mCgkjGWrIz9Z4jcYWQ4iCiVGOdcS7JD3dPGLZdSAuXdsiV4M0muqctQCQ/cEt/v2
QPyqp1+Kabgg4SxxvTLFMJf+ZUH4Blb5MmvY3TgKum7g/XDGSxW6f2QXW2tRW8yJ
+HrPAdWG5CGV+izW9448+So3N2oVgCOdLZ/JjPUyK7v0C76uNprwsH65TUwtOHJ3
CcEkufBGnohqZ+SHea7y1T981UAF7Ze5cIMdDiT7JQW8oCJdKb71o59zFjO9C8ok
SwgNkkHfu7iNIEKwIm2jj2886+dXfNP6dtqn3KLQz6V2QOC8OUhzQ+56PxidxZNb
dDr4TJtPKSjlhjwPHfmDOI+VZxSU9K5pH20p8j6/tB76Ipburt0anzapwRR2ZZOs
8dmj/i0YSeZ7QnHDy1qpuikbTXwh0PUSu/QoCwjmc9i8yI9qwu6qiwmo7F+z49Fx
QmRFSC1XWgGIGDrdpof+eJshm2aQGNdPQd0taYvwkpn3HNamyAmCnS6mPrxkZk9k
CyMSPrsxWvX0UNROmuhjSVGS8se0cB7C1m/9JU9gCM1vcaJj7DWgJAR1kNihOnW6
1Y0gjVEGFphXYopXRIe+mgAZmw2ndeOuuOFAYJiw41RvuDgvVRobIsitlJ/mp+b9
qCkM1LJlPZ8I8qmdNu1sROPeYuf/G/jSUAAGLYphxgZ9i5VvsJl10C2Yfjh/FQAp
sucThABt5Q7chdu78bntzPXlNoI1eRcYbk/L3uKEp8hitBxkc1AygUur/Yae5gZ3
EdEkNKJ1GBw9bcpCLx8U9Qxgq1gq+s6irHsJBKSj5uIoJZhc801ba0orYjk4CRnH
w51wd3jicJe3CwGQ4SPRhgCmzYBYUl/Sr2/SUhgPfhb0t2wMI/gZLpML431DLNC/
ok001m7lRCueqfj0vYYvk0EEElMdiC1i8nH+OHrAEFhpq1ZmFNywFQPTxOaIacXW
pkKBbo03Ij7NdrRoaweU7OUu+vmxTVqtKsw976Ga3crvvcZp8kSVCE6zKrOKLDU+
LjzDvQqp7BibkzEFPGTiutE1yPPKc+x8a1Lo7h15/CfHj1Jm4vemCvbjpJ8z+i4b
7jOYYIf40HgxPM7/bb+Cc+3/OcAjGn2vuOYwdmFIfQ2RTe2Lxl73QpC2Q9q995dH
vxfvADa6Oi75I2RLOB6/gExqTGcxuWCuwoeIxS53PyMihdv8ymXIyyH2muLPm4TH
ANQSgEMYGv+egWpIQNFWL7fj094M6EKTPTycfxGmgvfsFv9njuK2KfJ5mJUzlLi5
SjURPs97Ff1rYdzS2gmMF4+Ej7BSd82lsTWO7cHEixQiG+ZSZZvZxUgZxQ97Qytu
DMtVgLAOWxKbaPlRJvDdNROuTjWlBGeVKthH7qoyLB+CmYFYnpeJ+V+4T6NVWQB8
yt43yPWyxMcGJyOu4pBvs/XXOZS1INoE+gjuzqk8fakxdrGhWPydmzwXmk5L5Swr
Z6EgNSn9U1ZHvDCPC3wVBY48G4RbEn2F1bCqHJnyrnOKYHfLJeTnBgzM4oDJ6Vw+
HcAle6rMD6e6yE/yMqjz4L/4wcsjb6PedXVTbB73N3N9JwbnWqI7Qi3XCQGC7mTB
Kq+2Zhq3xmzOtI2depG2Dkau6wfeTJNWB7xqXjaaZr3mWMWVYs58L+JsSzZgRF/X
dcUx7PBBsSmCRGWBbb29Cy3Ei+6tzE52L5FIOT7pjJKwOOs0s1JGFAginWUh4/g0
s8V4JWfPw9G0qOLY89EDLgrBHaI/NxN/jpB3hb/eo793BJuKRwCSOMQtx/DDzb6h
GHMNzYr/6x9gZ0tNfkPi1h33hp6sMERtLKjpU3SqRxedKasB2JXTwH19p+NT+4nZ
21iwairOaZF6XLHfShLjXxuWtDkaPTzoL9GpB6hmBhW8VAr8IX5aRE3reuYsHOa3
lEyOTlroYWK2v5zwOtQ85dVPLVbf4zIAB1BydRF+xYbgzJbAEIxN3sdE5ezZ7CEe
2R0FWOnlR5mt8i/2ueKY/zx1ofhz09Fz0L8l7z8akdN3+Ge6SP8qwZaYy0/R63KS
9iz2Bs9VTGkUQzF889zP9C4MEJ3Jp2Se4yT1HfmQlroO1MC0WD3ucazDluFNqU4/
ohfZ9YM4dn3gp3u/f+Ux5giDUF66cWYW8Dhm1sjYC+46QHciBCUFrkh08hcAZMt/
IC0dbyuPWO1vRMjhxRAIxwHZVZtv/yFxJpF54tsxZ3fYcWFrPYZqSFFci/rmtzow
bflQWLK2o6gT4IGDipaB5M71xD+husmBiFn5/vgWBH0zK10y8MoXLJOCf8xrmoou
Q79wtJOZ/0eI3JlwTclh502XKuiuYqqduvNoqXquF9VUEApjTr9HIMwBAxpGEqCe
0CsvHekZwzZSpr2hUxnhwIw7AxpkeehDJZPy0yXBDvKJby2wi80JXyzvUTSJ8nnC
SXhriBLbn4QFDWivshLBtn55f7/5ghZIqgXDAsKV0887yUK7CMblOxYdJJRTDCIy
NvUTtc0H1xBIcNLy1w+Qxpaj3aY7LhymDEwVTD4pDgM3TwjUnUs3gr3TYtWwAAwe
W/fYmPeyb/yAt5zZMbLRrHplgxP471XffWkVaxQr8Y0j3NX0fGxWmfH28cxhOnoh
GqT2bcUYVOji3U4bO9yPTUInysva0bPRXOqG91bHjfu0GM1negCahKtT1WMFjDa/
kKYrsWoGnBsmfEbyzN5hY4xZAvlFba5RqCsfpkqaRKZ4YWWHMR+BGhimpKesUhs7
MzGS8+4yMvJ3aYX5+psMPbwVnamW+Ej6ckQteDHXWyqtDRv1UgOujHFuCiVdyQ2W
txyiAwuyIptbPXpVv8ncO7MLYoYAYopuoPJnsicRL4YuUSyVJMKt2CEpThZtiHEd
lYNv/h//PKnNpcgL5dVupr407QRHfdGKeX90sfDBMpQczlIaaKpxZPNllG4zVAFO
TGufc5kRR6eRUOqR5woLBqvCy5I0qJA3mgmi6z02lPj1uka6JXz/LphCjxb4M+Kq
Yb7q4/oBpZroXjgftqINC9LYo86XiAnZccDc7pChKydDlOYCJVqjJXm5WyzbxFYY
ZUbag+KMWP/mgNDAF0bmc8ATDdrfulul+faFkLNT6muhygvsHEu+TXQWcUdDBlV7
i+JFN0VOPAxBmT1s1rrt+RIOrsoVmqYI9vFxhqTZWnRFRUjbltKg29FYGVwT1Jj3
y9DSpYGo6ZuM5YS48RWwjrHyC9rAxHJpts01iECLwAnqoYMu9E5PvtNe9lOY2+ej
v6EZR5SNJdqxKzVZ4vUd+1jOzLqWF7fzQ9x1sCT2QUZ+NS0nT9gwLkXWBTvYbFFO
u0ZAcHMG6zE8Ty5gQ0SuxftZ/m9swI5IalZDUYljV6dBYedinFfkqhDEAML7rbrk
lwKFaYGhUi87OLxA5sil1XUV59AxdEzlz9VqE/yFH9ERpt3xb3GhPFb2FyZ9q449
XJrEr05Zme5J1oNBSlpQnLPmoB0WFs/p3DGe3vEjRYiaP1brBMf1vfjXWkWvvIzI
drb3LTl7p0SwIMlQzfWKOtx1FpR0mMQvXS9aoWOyweumYSNrsIGpF93QcXOYfXH2
YtCXj9KbBliMI2qoKHpD5K2yAIWzua9gPQhYrB8A/TxEB4uJe5N4tkjf030o4POO
DjU5ZtGN6g5+CKgrcHiS7aLXJvzeOpsf+RJw4oHiJHRHUBdRlxSuQlGrYIGi/Uye
WXIHy105h2fTEe6f9xwshJuakead5VCNNZsL7KyUl7oS9JepNxP8P1Bngr20OEMN
iAN1c7payB6fzxsxn8OAR0jo57eKUbw9/yILns3ptLC3/hHqH1AhqhCSWCMmHSa0
lEGII+eEj5EZCBaYY9pI/K3hySHPBkCZjBPmOrQkEYa1AwepKwWleeIJxFGCPq+a
xd0O5etw4HPPShu+YDMusb0isDsZszh4mm3tPmvFo3MhGwkDOW18d4OfxdXWAh4x
I/wAwOPH+Eim/GCmh2oqJTZm5hZb9R9JVDfL9PWQmct+WisBGA4X8RvDdrNnjSTm
H7N+iOQv9nNWIBAbBQEnmLeC14/99bnxT1QNrfHu8Z2TuVKhJxERjVWiJzNRHGh6
q83X1/B+LpI2lLgjFtFM6OgwUjCH4BvGPuRmVQz+eUmwJKAOmshOeUxvHyhFl8WW
d79EtZvyJ7JsSiZx197BazLpPIM+mdI2Ofy845426DG7vRrrtsIXAfhRVQ8XiGen
plyNXE0T/tPW6ZtQXnK/ut8xi4Lgx8Ym/bpy1+L+Vc6By4W3t3W7kxX2sJpSj6wa
2Hbuplv7NtU8uiFL8JWHGkH2FzrOdGxNzH9c1QThiMkRmk52pdwMdzbpeEU9pc08
CYb2Fd+PdenDFfE5q8ohzwLJKwHLOT9ETNaYZw22Mb/t6o0f4mQ2NUKmgysEut0M
3nWk6waldbOm0p8aLOxC30DlHGpNazlrTHouSHFrk7BrhBXYkWFnO4O/6jiLLDtu
BPV2FBAKncetWHjfc8HbKgqHKvT7la1Vy1oNgxq+3j8M/CEFCI5zNjsiAmwQI5ZJ
kQd4lLKuoX1CoMmC51ARJrr1Jx1D3fX8tHR0BjfNYN4re++UJDdNy/HFT5JFPeFM
OeDGXEVr7PG4xISZdp+GirAat+LuCckywAYs8FUJV10bctVZm99zHk69fzHTKUYh
vaorS6IfiNxIRKeKAD9+sCNfS0WH48+UiZCCK0+jIaurP85tYwhSj0YvxjK7t1g9
DYJSRMbNimGJIo9gyIX9KDX2x/OIg8uva2/oaMhOfpFbA5ALovv5tbROmX3fPHQT
SZ1nEJfjoi9AQdOFF2mcknO+yWbMVd9NPLkPrMjA0q1vWtQU82OtaUqREb59TPLi
aCA/lnDuqMQeLrSCh3K9RNbPeC0ft1d8NWWIbQ2SZ9Ui0nmJkBd2Ntapu72s7VGg
vEFyQ7mqBeBrUDZpNq6Fmwpo9/ViCcTFPo8oxZX/KWZ87L2Fx+pWA7vpz8WJ8PKK
lOcTRyzGjY0aOkrZvJXgT/vfABGncyRxC2Uvx9h6XkNVQf+5ZbpCC2J4HlrKbUxO
Cj+DYBlYxyglryVn38hGdmPdMcoOzkcMXKL8ubuFp6q9gulDmU5FSJ3V0FfaGIiC
JLdkYsehOzdkJ3z9V/3EPb2BiB7/KaFzpjKwcppZGYi1d/itR5s1vl0T9+wZrH3I
HJjZEgam/9U67LN+kgziKcPQGWPFiGzjbBBqIKqD+LsAYEqWJbhavqgWzNp8fv+J
TAd66+m9uZb+Yb6tEZgSaEYtZnmzIhFnCoqSaKhnFTBw/HTzc3ny6qaiaaNlNOGR
9xex2cZfyY6pqvjgrgZex4aookdRgXAMdDhMiGflbkdfs0c8aNd95z+FM7iZjAIa
qxdFdBzoxpZ7najxxggvwLRlVF9ySQa17X+25L5cKk+kvEVJ7a44EKuDVcA47FW8
MXElWyhWJTKQpbjGQmeEH7DCxQD6ysypMVwf0jqY7srkAuEj4iAb6untQb4omIrK
sVTqa7s6w9FkU29r+hPYWNoNKUdkz6r9KgqLkLa5IDY6g3ipKzCVGdOb5939w/um
iV56TZ+CDlMbR95Fq8LoJsebjWb0VYr4VH1PS4wvDtop1P/dMa0fSPoHCm/685b2
sqcVXpucPCkc/mDrs72N3AHEivgKb8h9ummrvIt6HrSr6qJARIfv+4PEEjbW6ewt
0rQjVwnyYggmOBgbTP7a8un6CHvIgtw7cE9MZmVUAtMsP+G7dMON+wpPoC/HjKnL
8BuV7YyPUt2+KpuXq1g2yEEyG5sG2tpJ6f2mYY9uOX++yeNWJOBX/hYb5ZGacpc+
BUmVulvxyYcOTm30bwERTEKrQWBQIljUWtkE6Y+iu2xaSaWOAln8byrxlEkMnrdY
vPY5VBLg4JSUl16moNWfkF1m12Y7o2/5WPd3u1Nmr+0Xp8FQyNgwzhDe3uMxnHqs
9cvm7ABt4kb/UNO/2pWitLYgXMLIRzDnTI79MkOKC3rJJ4GxleGIRlZQtE8qCzEF
51uaMky9OChUCw1dB+FDwKhDvFW2yAmw0aDFPemoB3Yd5oTNUCPISLA+zbWvdwyC
rbIAFzOujT9XyPbe1tyTZ1etGhI7nqm8CE0Pq/pfkedIXIoxu7oOvP7TYfbeTV5m
EQo73+l7IHUh3Md5FUGEhOInGNvxA+XyErEiUatwuuse+COT7ZBxmnFddl9GtRoB
G9zODHv1647m8/qFhYMNkZ08tuLtzY5tUjpWAFx45N3CWlUb3MvcQDolcA1uBydN
I2tuBQ7J1SqhEdr0UiY51H8QAich6um089OxdTPRVS0aBokyDWHVVF5pWkiAHQBF
4liBpYXLx3BQ/crEluKCNxgI7wS0np5H55m2rNchTb2M1dQkLHCvwFZSMLG4uG32
VSIidr+AQMNvQGzbljZldJqMmvlQ4IV7EMNG5O79dU83vQz6YhX0REihaJrbqpm/
9KTCMfBRBEqxaF3m8JvvCRsGmVU/bR8c3rAHwM4NQDZyHAKxS9y0ajil+PrPmt45
BgNgu98yuIBYcV/nx9teJJWskwTkZF/VrNOiHKPEYNNP+L/Fk4ArDjZfBcEwNVPL
O00BXE0D4apE3GRUaMJP9XLqubXJ5ihNLyI7AgrLcPMP7SSQWhPxnm6yTWl3qVcI
wp2FcBCHDc+YBB5xLTGmgl8Ew8DbHkWJOlZGHYBoHcIT2B/tejIhegcZB/Zv0tZ+
4EhmSMHnRqACsSKZMYTPVOI1KhFoO1JN+CB/+Ua1oxJ9Cf5UUpQgRVIZvAboYdaZ
6vlfn2322HgQIBykgnJ0cIuj2iyt/KtAc5bNninQLrPWJ5EmpB7TQA16Ayyg/Cfm
TDBpxyz2OVsSGTTQS1RLREGrA6IQMLdlMDAPWFBWglJZTiLiknQ0RNLVRC6OECfe
RPgd4SCtuvIH9XtKdWt8IhSnw7KclM76BeK94iJUxXh2ZSYPQhePEZXz32sXOaLF
RW6XggahIUWuDi0ehtYEBVYmiTQ6OOHXgSHaFycoYlPrQ6Nw9I7eNbExoz9OJI1p
HAf6DrJWbxwQK4n67Bnq1ranDTsPAAZXwRMIgkjcSZZgCEF6UsZ9uTyGGszT5MYz
s2FdhD/cNv1u6lRgLb3LGwMxWEqcU8MuCnxu40FJBCWmNcfk+vFRBR2M+Wrya0gx
jJLK66/JRy+m7Ijdn2S0hhY0phibeRHm89LAyh2ozaV5l3X0qNB/08dQKJPXASky
BJThkp8h1VEKilvaY5Di5Re9WvZLeILeElWwu0W4wQIwWnCk8sMlqL8Ou/9iTuVM
ocs6EX1G+zO2Sa55zoNO/x7wq/lZHP4s/FxlpiNGduCcAvkEtAQmshXKsVuAyqvx
UOR89NaDye8P85lY4I2p8DXKXusXur+3SDC9nlLCkg8jH4rXaQbTGWYgKZYfiL2z
vuUljZX6lh9EzKKXIIhhO7UcdjOTDmDRM+3h1kNPmkaqHFkEci/Y4pvqexetK46x
KYiMi57u74Q+TBdZbEMBq09yUNkhDMmoRtpIYO8tusEMFFRFoKHH5QGRhBvngEae
VJCreq+gamJGnf3CFF7N4TcyCfWA0gZItIh3haozRKu05WOF2brkgubxBRucjLn1
yxbeZ+03TpGP1jJP2Lqk4yd+XDgnsZ5onUAXt1S3puSoLaHpIt3+q3R7vCfSkls8
AYn9Cac1+9+/7vvrawjxsXgwOnXIlFHm+U+E0t4805pKALVsLyieaOOYaiJ+A95w
0SEROVWd/ZHgnMbdSkbECUVo0bMtRlpHDIyp4dcqTdrD4PP9nOoxkspeEIONLoew
l6gTjUPOXt38iBmTnZOTNExS/ItbWn3ZILb8x5y0ybq9ehTU9fhpp3W+JvkazkV+
tt0rdzr5BhyAJ84uT0ATqTMj2DOkHGpRRmJaeeH13XARvOQYXbLDDyINKF1eiHoA
fftL1m8BrwZphWf+ihTBa0PJD/yLVtmTgi/0x+/JZjBkYKuv9isprgN7PThA1WQc
iwhTPYnolMAAhvW4xuv07veF8lOlOuhm5qdcSsl8s9z/ZgqLztKpb1KnT7+A94D5
qtGL+s9afZVNgnRFsQWMcOU3oC2fSbcDgFgbF1Q1b6ZbBEj7mdmc97nBLOW+72C3
4ZN/Io0hyUPQLrdLicjNQ9pTXRwgkleHv3w4FuplMyAwAGyM6qY8SqjQCPc/reyH
XaFWwwTwVCtINGqN09cWKuWsD3bznlA86A+C4T5QJ6iqhL0Ikjpkvwe8HJYsfPf1
9RsU/deDzpFpSPi4hwfsjNidnLMlIyIYrupYpzyHnMDR5tifxC0z4g9qYEn7n9Ag
ESCUW9Q5k303M8gYDmG73WCMnzbtwPFK94nPb+ZGDKils6SbQvtuhWHMbCAglh4I
b3hnjzHMQovfWpzaqCqwIe721zK6bMhStslmBz8Ix2qaCOyxE2cgBPD7Zyy2szTV
BN2BPvJQo3n9jGuRUilQe/iyvzwtHTq97gEBuih86yTDN8xnRkTiTiSy2mJlP1q8
DTnUqx3g1PjplZViXajk++gUBGMgBBjh50DxrgNoLNw8yyMk1PyNKskJ10GFWpcQ
YUwuJAqzYN2CspkIrYn8/QTwt/wOKLN7g3uuUuCdyjunLNQQEs8Dzf50aUo+Nucq
F8h0qEewshrvzBtDgOrRJ06QtetqkinEZgn4FLk8yCeoROxuoIhkSfijLnzJny2r
OAju33us9LU48nZ4rwxLvnCcSiJ8LwAnfeRp6sme84hEcH1VVefuciC44sDpwEZi
24lbjSQvXx9pZNeWKKJghGDKWsiKQ3NwD/2S5OPqRRR7guKLC4HXRtKtsxarz51R
07S1Lpfdnqrf1XQ3xwPjDPs08OmWr2dy0QpXpwV/4r9ESM2rS9H1Y6f96LAVnzqP
Wa1g6MVNylWmmRIXVSbs8WUq0QaLYzNBaF+hdtg9fzbUNoDzratZwx1miGAUeqeP
9HSe6H/nLYRbCM57nhdDvhMBn7QrOn9H2PgElrdPtQ/V2fM1HDxUltU0eqpBQOjV
s+jANVJ+Dq+1lHJE1PZQ+uOLfN4Sy5SrW2k6/DXuuOyRdlCYoZ0Pxs2QuF4jzSOg
WLGO+TdLb35jg8dMhJBw23WRd3rMLuqCQwmBrFYIx2v4wC438b2UvQZSGUswmmdc
lCL7PQA56HqQbdgsB/YLJJDDrhoXY6ZbKTI4jV/WwivFUhx1JhmK1W5cBz81WXLk
3bkPbgQps4nDJy26Z8bszbbHexK7pss6xy1FhJE2vcoeCd+B1e29kUIFjISpotIt
BAdvR/eYBLqMutmGmfn3HcIy60g3bggOnOe5DkISz5ktcJsEsAfrG6QwbqvlA0M5
mMs9CFEujq8MAi19sWOGW+4ZxmNgUZ2Xp75f+oLn5wAGRs609xzv0tXmUWF7bPXk
ioGxGsgVhgUgqcBjFrbEFsRwMYIqfDbljfoytdkKJBsrwO2JZ8Hn6Bl7jRXcYaLP
rf8ezPnW07ZLxr4Xm/yN22TS0x/sAtx7pezqH93wuRPJ9XOhz8MlFJKAX8TnF4nL
iyvosTXJguJnCbK7szrkUiNJJD0y+DZ3h/iN99oxaszxVNwjTuHPdnLXfZlzDA32
mR2i9ybZ35fUzRn0liGvPZe2vU76ofprVtvoDHS/RYLi4iDUJ3N2i4OHRbVrwZlJ
9248pG2/kNvVe4spDxISE5Sy7ZNWxdXloj3niCnWPqVyhC3Jb46oTViP+m2a8iVs
MW0sFU2+bUNCXi8gI277j80CTvgpKvNWlpZSgkOj4sh0o8QbGqq8w0tRBoVPcWnr
Ce7tIjOSuP38nvvb/98TbYb8fLigoErHG7m73KLVTvmXg6J16o37tUrJC7tlqJTI
AKrz8crIHP79e49dwwrCzELuK8LOtRhgAiOvJipfb3N93nYA+4xnlpipjZ8SH6Rx
wRJhbbXp+evWhKx59QfWwRczxM0YzBcnHLbJQAVKHL+sNMqu87nyTRO8QulcOZNO
U4iitXgtOjww4sc+3jRkIVsWPNVJ5iLs/abLRgCbwKSlNfmFxyPkU8cNnguDDyer
ldAOLXRoclFOBEqZqH2xiWs7y0GMbTsPRfloTrddfi9FJ1XuUTW96YJNhA7I7D0n
rQdzjhSR8xarEZ5YKdiAGqAxqMJGNBvZbvhdJXF8RPQK1/AvCc3w0qhkkj3IcRht
E1xYq/azJOX+jXhXxAvCkdSHUGwIcOM/0iFkDly7zjjnKVDpoZabd0IBzXpgwQD6
UKOP/u1tQGAgR3IuiOzQQFMHKjBJUh24m0J9FXHRdsnMDiKeVWqMz/OiRzHyItdc
k2SVkfkUyoC8r2IeVj4VKqv1vbxGnyR0oxOVLV1lMMT4/u0br2XCVtLguXyio7vm
nmP4aFl08WGn3UgLw8IpzlVL1pR3LCxHY/XIjRXd1q8oRKZk49Q9reLgf+BqbFLi
jdGGIsxDgIQ6cECVFtv4M62CVlbJ/YijsShj7mRPHx7Ea7Pnd8Ht4qPKsASKIIQv
Aud4dd+0fiH0oSfBo5+Tqb71IFXPKyCfjniMFHGWskRDYXy2XIQbi8503xeTfzg7
dl3HMr+SQ/8eGLa39h1ej1I02/3rnlmDCOYtDccIaVA91ts95YWtlC7GHNBTqnlS
5R+KDN2rLNlM6+ltavrQMireXuo16X2PO56V07DX019QCKyehRSuG2+fc8F47xzu
j1H1faOvJdl4YvTJf0lykwBlh7ma6d1ViijF4ag/XQfi/V3fhXffRXoH06e9rZse
GqBQy9SGflFWp8VkbzJDS42WEfpE5PSjKOQc0xEWJYFgtUD8vm2ro12YscXEcumZ
QruSAx156/OHdFlhTy2WwpbsO9aUz8UnXOGiZ6XITkLtWUMhrvRaBFNkT141Og9M
P6yDR17xq3N6TjKp9El+GihaKOUE1vkK36cXJLAyHWWRvoAr25+jykncrnqVRoyS
x6vTvKfYwLpt8JgcEN3Yq2MGVx7I9LOZ2FZMVhRNqo9lIP0frMOhIWNUIhJ+/KgH
odarPu2auJCOKQg4D3V3SHzs+4BlBgHSA7Y4CLQwRPsAcQ0aak+s5x1Eo5uHnIuZ
Z0icCK/T94bIRKYzm+tyhfhZQkYzJ2bj65HjGK/UNO07lL9LzqECueO40EmzIrML
uui8visAUp+0JYCS4+b2HN7fYCqRhiBZZiMOEWyfwKSMSBbm3PAacwzluQSenZKz
VwdyPdjS41nJ3xh2UPn91E+SHqPAOVxaWTafXCBkDpbIUVab0GxAoeZKAI0oPvVA
yJUfU/VZKA0EzE3wgivvrD5925TKOo0vLLCOhH2UHiNjZl26vgxLhe8pfHjhQERm
ON6lUsPm03m0hm54Iq6+8gEmioe2kvrz8ScONFt+M0+ymw8e+SRRP/SgrMb0jpOb
DcCtyh8gimH2HVqFaLsJoZ1AHhLalsknqikVu0WrgBiur2nX5tImCBVWHDG3HIIB
YSO929B5NwSqJyNLzdMg5O3QCBeJahpF2ojYjs0a8ctZ5OPpcSKwb3ZQuYRTLcWu
Wo7vJbhczs54N5LGzk8p8xfsviEF2zp7gEyYSzK5/lVYC3+Gu18lwDB9c8b1/L5S
m3bVv8bL9xW9R92eLBlG1wrNEDUldaLrWMCNtUdWjg9BKqmo1xU05s1di4BFx8Ne
qYf5SLSAjpm98U9ju8Ch7lOKIQxBH/yf/LEUhBiYCxTRQmCEuZrtDJclKcVoZqR9
BajxiLYTd4rNm1xDcbGK5CDeyxT9MC43xRFsh6er4v9qT5hMjNfzXDOEDEWz/6fJ
vZZZjnvpS9t3j+UG9aiciTkv9TXG8l6yiHrBGId7+cQYodVZsLgfkUkYyqtKPkyR
JCheAiZ1D9DzQbku5oBPX1Z46ndQ/ZvQwKIQxwoHxVww4ykao347yQpt+EXxvYFq
5eLRMHDFrxbwQhGJkEAFIxLENi6NTLD58raFqYFiJ+mreNARgB7HQpClUXHRGqFX
eaR+w9g+KR1HNImnKbdjEj/GAr0EQ4It2FWvay8JBEqDGd5DOcTAR5WxTo/fyZeJ
epw+EYpD1du6+IQaDk+PYPEOlEBhnmeL9aogeu5BQMJ0K2sIFaYUNa9pxy2dYT94
FLa8cvEJmpZtKarOb9Uzk8g1tT6/qtefeczOBru5xCB+wI6eGLh3xsq5BVScFyo3
ROGUpY2Gp4y5wvPzKui5mFlo0N650ASfDN05A2LAPSqxBzFH915sKLejJNrCfIyZ
6NvC1VUTZQoxVuAe88uf64llX2J0GFbuu47Z1VsbEn5CuOXioXqcD+8lelSs2WkR
Qdz0rMxdj2hAfzyd/6gvLX50BTJxfwsjsKz/eMmRQFRSCe+v7SRQWzfWseY58JAs
OWZE+p9JXvZujAttBRPEtdWr6AzbeBtBL+O6rksRiRZsxK6d3rsjaQkWXnLbq3Mq
rETt2UbHjr5hScRmreHXB9TtUUFmGppqi7+eUHAi6AkzCc6pl/3i9K7hztxpRh1Q
xpeE1po55+rrkQ1uLRiMXOCe+kvgMfpMhybJreygHWYQx4fR0qf9t+fH2Jb8Xa5A
9IaRKUQvrgmGp87+5BKpIAFZLqpFsqKl+x0ohhH17FAnNPe1glffJasU27OAuYnG
rgj5pYKx83q7ggAMiWTh4Qq/bJcMKx5OJsYV6eYnL4+zrW9jpqSYlZH/DMtWQIOo
valWVPqw0HB+viDigboFtsdJ6tG7tzP07czH2nqV0P3LArDP0pUKajTOekBR7itI
Jxl2WqQU4mP7M9C75yo0mLFyEp4VJT8WF6bEwlkJ1KlChr8mbTOyDE1ad6+k94KQ
NNghqaNvZVyjvVJ8BnsmOaKvdCPalCEZVMn7QD9fTqi9eDfo7PepkQlZ4OYCO9jb
dUr58pZnD1VejJWblnaMnE3l29JxC9FHNG8HFJanl7NTS1SGW7hTiUkPBuQE2p4D
Ho3lmN2HtoJMBIf74Zp5vCFRUuH5WVWuXC84xtZU0pmWetc6I32+OqkAGikk/sik
ghTlfFHNOHJJ7nAonBLxiPoXO24ifj31i2eRRKjWfgipZvp98afbF4zMTFFpyRki
nzWAf1e9gkGWX7pZH+urvOPwlL2YaL0mJB4z3drST5albmhXsIiW18M5FuKMsD9v
dU7Cr0TTWs3SqXHqQKiCRXuTRSfgUUhUpWatL9NPKDY3z5Gfuly4eUhxLMnY5Lcx
iL6GgsgjgC/JjQqgKvGOEXzAESYoZvkI1UL+v7RYAENYZ4Yklopl6NWyhzpMZKcH
rSdjXIPgJvEJdgKfEYVwR3XRFyYt84p3Hpw3tJm3fB0kfCgvuptxPHvt/x5XCjq6
11JVP5h8cqBg9zzawzhrZMLmsCEDF4BxaimjndRIC1Tra+DsWH3szRCHWTdnR/RK
vfy76QrFBvoLlrvSlIi8woh9HpX6LWHEt8ZXBfQdzSi7jHtHww0bj8eFFbROkgbf
k3zsF+k+17OhwJG+/XwRvYLHYHrB/XMIXm8HtLT0XvRv+Dr3U95LzIVjSOKkqHjy
L8MGlo3QgCLMAWU63KGb5UuQWeOggeSP4SHwXSyh7P7NopF9NKISFV6Y+3h81/YR
LTgzcS/IK2f9MpTnOqOiow7f8ssxiTLsHxgCfpx4piocvAM0/wFOGUKS9aEj/S90
OAS+CtdEzPeN1kKt9ZupDtpUHtInrMMt2I5VkWGv03hPSYjlADpyCZmPWKtRhw8U
6paugnXzH+3KtYp2I595ydHL+5th/ekf1ojpN3GZisBjiXjwFIDcFwN2uWLwoXdZ
3tKzeA//obVSwDVF1cA8QQ8dghO7cZcxFphbc2Q68BfO90+BL2p5LBpqCthsoWhB
zMEoryA/EqcFLq/SOpPLw9AcQ4lZgAX3to46fScI827JHrlc+Ako2QpWV8n08FBw
hyBTywj0Mms7matOXb5ju5oZrCEG6YMTO3+W4dlETWeyh3rhD0IqXYDx0P7Add3O
kee62dgkiEBZrKTDABKZFxAwXO39m5n2d625M3tla72OqRc1l4xo3iMl7mbb/Rq+
Yj9JUgT/V0qJvp9QjujgaSwjAv8hTn1IDAlQVIjmHF/wota0tNHWlkTSJUtfkLpJ
vdMax9u16vxJi9Or1Xpw4IP/I5u7zmB7BftFp6NN9kGgKXC5kbgJSS9NEqG/ZPJ+
JE0Y4SmqY8vVoyxolOdeYvB/xeJqrOYZ/6qdFixeTrS0E8pHuxWMlr8LtXmUxk3U
f/5RmzvUrCD0Q/beoIAXSECRF8TOXbESy7Lnn6xxZB/cXjjfOuSce2JIG+3SHjvQ
8+ORv6AwDCtNYjSi/Xc8omSEMahKNv+1p+ZTm2i+GgeZAgWTKNZo3cNWKgCX9J9e
YKNK3XG8auN1GDOq6//FykHBZ8gShemZc3W178xLspWO6GcXIdGV8iTbPIpe6yUp
cbwE/eonmqHvlcmwXix3RvFARBw4bDgvsok9xaSsSYcJY2Hz0zm2qlL/2j7VlqxV
O3FDtxB+m+JOVbvFDQef38Yu0yHiiTee320QEtQL3bTefoD5bnoOEK3qAnCu0Hvo
+8k8Ua3PjFbWt+b3A7vuZyMuVTeFULKZorJ5jQZgrGmocBYdKKDxljfXF6rZ64Xu
mCSCN+aIXxMCtEqfZ8MBLiZVQcmpngacyYau1Jy/HrEVKk4ySCev+8YT4PaUXDUS
hSKunsZjQ3+ZuyS3LmufEa+rfSmHyj2MbkpOCiD42u2qDz7XBL5y54O4rKM6myWl
ZmVWx7a53oqafHeg1CvgYIW8Ei0J7DMRGffLc0Jl77aT8Q68almL0FK7wSZdjFx5
d48R/NK+Woj4dQZFdfXvzXMs1TE4Ujdg8iqkfL07F0UeNKPCnq8u5HZt5xP7aU7A
9tLfXkuKoGo8J13fql73vjrtXovEmtBg7VD5+5BU6ygFLcqmyXXjuoy/2MWkw9HR
5Q3/+uNd7kUfR6uxvwX83puoSzuqTWYVCZwMH+PlpnbEfpNJd8Z+WyLrDhi2jak6
Eij7qufP0/vU3kWMAL1a+n03Z0VhTT/BM+Co1HXgrswjjItbDAAPU+TqO0h0LjL5
VcLZBGgegIiXXUXn//32tewnP87cbZ3SUcZlEwZV8AfYnqnZltpdT/3Dm+nQDuZH
5qJ5ReqAuSbIRrb01K+3F2QYijVODYCGZycAT/8g0dPxPDzkTn2x+/LrmNDkOBFE
VoxjO6LVs46W4/TZNLUzTCsEv0vfkL+gWA4sG/WsETk2ZSR132rAovdC2HPb+jE2
RNM8IKGdN2eWtfD177O828ZZIlcANqndGwBr+DO/vf/o78e0Im2YekjfLz7dnyN2
zBqK4hsKkFiGpHT2Hv4SgkGIK8+hKfUw07zPESR2sp99rJagG38uC3IVi5GgXgji
r7oo8baD3HemWw5bJO2ci8uH3NVqMBdMaH4+aLpwLsw0076Gtmrf2jSPvniOPpAJ
OWRdP4Orhiz7yLAr9uvjZo4TPdLmB6N3zTF4TZwkmzRmaTqAKxlp7s7KmPoPg4Cq
ZM3Ux1NmSvoAa6NU7EEl8nRgoqAvAlreZ8XlB4bsoRxomwS9aNwbDM9EDlnnlmcR
CzzUOIJR7/x4PmbL9RfYg1HAsbBLMYsqxN7Zrl6A8GlBlxhGccR16i4RLkpyI0Wo
ndx+W4H61ROVBtxyBL0ckX9CxFBQsqjAavSd/Lo4dqk1Jps7YyzOyX0Lg2lBvWPR
nIaV2Y3Po3oNrzE5GmHhNPJOARffbHf42OLSZFKjh9/zrTGl7pSHRgAIvV2LCGW2
Cb5HAwu47YK9bua4RvPVD/tEPG63efcRQOTZoHIuaEuEir7F5t/hXwGfCqp2sBM8
sLCFg9bc8Shq+pBQlf2bPjf+xgte5UPCE7r9GI38vZRYtbw+j9R6+SITp16hRbd4
7RB0V8J6bQcnXpyYc7DlDxT14Nu03xRWcQLStl0hmwN5eeVFDtPpEHjW6H/TTBfG
wPzVffawQnUexEkrYD44KJ4gBZhBr4gvlY6uU0sHLOOhUnKLqy8uaiZ04lX/++uA
vI7PKItmGBF8ExK+YTNItgjV3A6NV3CUBGtHxj++D2W6rTJ6eCGZH5NO72pEUneI
P0/6Pnn3eAaWUwU9yTZ8GX6M97Dscb63BFC1j1tVuJftJmrw8/W7EiUP+7M++szB
gxXCpinpAx3gZQ+qTSiTKaztU/8kHacaE4mFzP8+J5HdqCFrAl6wOyMO7xCaC3nC
ngoKqtiQdSoDmRqrIcERgTFJXLUg77f3oILIQP1AE9dv+X/YrI8Ceh6cnKCtAr0l
uaKgiaooN0kfuO6f8+cCHdDJc3pNP983qqpwNy+KANhogVYeXj2/WSjbbOWUAJ73
KpGTbtr0VzOllsnIsSXTB5bNBph9awZweKLHwaA6Wpx9XhznPddbMpR29rjc6OSE
HSUkERcN8q7Riyq1SNhLCIwV/0V+qNNJEcitU12G+p6LIGAe5PxGbnxguhjGSzSc
OVwWQDFJLSR+3Y0A8ld6jMMxcxEPfcqIvnPIXUQxMDYaKI6INUtbl3ZeeJd51lRa
vLNAA7rXnsqUAbOxdrLaaBPVQ7hYd2MT9SB4OEn46J/9Iq7URzNA9AiGbZ8n3tqp
gee06YCwMPIziM3lj1QxhM/fn6eMv/0iEmCMtcwjBX9wzG+Amzy3oYZHW9cuKoQg
dZW5tTeGUODtJDQAG89W8Yuz+zzfyLi4iXIGCt2e79QD6Asi/I6yB43LETTdoPgV
dKcRMqgXJUmbZfAQ0cz0nj2rB98Y47fN9VoJfyJxocQZTHH2/xyo61YIIgUda40S
q/Ak1V/yJLqz5T/rnXu7cnZgahDLtgQpsnDQzi+hkliMdYuIyiWDqvsmw6reKNPh
kNYWUfMcbPe2tHXE+pxlWBr5k8VDfT/T0uaNoZCQFfyST5YtwAnZbsNlTORKRxF2
tHeHvnvGOcZ4OJrOrrjtGZBR80mhvP/7nF06vqDqTd/pZjEyEpzvzkKBpMM4t6ve
zTyoi5MdEc9SC3NbrRSQYIh54fwsbwBZ0sMXKbPAEDnnub7jIUT3BXboeQcRhA3u
U3ijoWeqydpTYk/+gUIV7fyP7q+SQNtxCsdBs+Ipu6Nh74Ur2ERb9fFuJqPN6ehP
b6jKL6H953nf8B5vtRMTtqBJrnvhR3UE3NHrJFiBl9j24O6iAcSRHRYc0Eie7hOe
jwtEa3g1dy6134zjXuz3f58vGkgtd5CMPGpLbVd3ZT74n8PoNkRimVh3YHiqp9hN
uh431VCCNc+vZLl8vtCGQxRU8y1Jh/HYMQCtGdpu1jxBcOYf4/oafnw68l2LX5f8
9yrZ+96Fll1Pp7FyCh9yEZr37ZO+sC3pubBp0bQVfOUIdcFkBQtEz2Hr59y7Lbd4
S6UCWyw8aPuwTf0SnwImeB3A+3CQzX4Nt2u1bbcaLNQTHayN7E4ggmXN45yWSH2x
3wlmYU7nl2Qzn7A9+waredk73ZMSOHE3MqNwtWXG+WRpbVkpF7viktLlT+gO631W
akVysAjDkw8OMradv+sLy7CDIgAPo+y96lINZpQTP343FBfDnyazr2Pr5Ccq/E3T
vWbo8T/R6z8Zl5+sIQNitnhKCtj6QhYHGhsllNGXD6Ir/3/dYwB/kJYmpgvAjSR8
T+NHCb7I6PW/pBZOygJBzYmltC0jaZa9wed+f7w5PszE2D7B3pxmMsj45BaoPEsY
cNUCfhlrnDsXGKmcMK9N0kqcna4DESFLLeEXZLMR160xDHlnEAtHyu3ZKu8WWM9U
1XIBQ4x1abDwC+utGH6yT4pxFXhEtGlebEMrFw43ynWI7QKAQL1B30zWwW8lI1Lr
WjX9yCGTqBb2Q0rJ+SZKHXvKI+pg1ZVdqiRR4zSMzt65spyj6Fh7eEkjfukGfBY+
7B1eTzqhRIUaIWmv6/ItwmrVWqg5JEgsNneFgqmw+y/4cGROoiyyJF50uI/wOLGX
3UPUwJybBWevKM9js5JlelE/2RnatTebBKSeQSQPQgIlyEiHfC2AO1qP0OcO77v0
mJo/CQrdJyESLZt/ty5IrsWYlyZaZCLN8D5oRlJnaCjKMdeM8wX/RDJTPaGXACXU
DIVJEF0skhF1HfXh42kZlXYsQfeH+3n/mVp9PkvfR3dgE3IaoedaizD4Oj/8E7Ul
JM19GagcVp+Gej49qznptQo1Wo1or0d0vnBYa8yAzrtUCoZ1rDM7fq3pSCSa5pZ4
02kUFMYWxJgDOVv2wF8r9kXLrSqbblRqvAtITJg7rrMLUHsXK+82xgiXf5s2UoJC
GVdT6hWo5oJ2tPo9BMxNrm0KZ5gZN1WCzrI6oSoG/Gfr0c7m//5oCy1Jb9wAngFo
++rSTPC3fOCGeOMYG8uHz9aY12TW4mIxKJhHXLkKB893Q6859m/wh7Qcp7MHzbwg
4G8mUTZCR62aZi1EHr4xy7thozwTqJQNi++lPg3jezSBiDJ7F3PTyUE1H6QljVTY
QLXHpKFZltIlRNEHQkYdP1yv+o/Rr/Ppg/+FkffZ8CWXDB9q3Q2CMA9dxO8i/eI6
2PL/TO8FabQ7nzNBFPSvI9dfWr6ZbTrXZmkGHzgBwKLFPc44WpHAYwtNECIlGNFw
cjNeqjXj3Is+Ql6hbyzqBk87aLbYh8ONd9EUSYXOEBcauDC+BXZm53JMBX3+ox1M
rN13KiSl/QG+A2/H65gSyI9thMXOxIYRlRap2K0PEmae+WFtqFW2DRV9SIhfwRJX
m3GgK+RJ1JsE4PkKaSsv9LgzKMTPD4anE4DpEfgwO/LaovOL3QRLxtyNSV/IfiFJ
MjW8a7XQpXPOtwlSqzrFVuEQXY1Dl6pfDcmFsbhjxqgSqfsCr0wBsQMzw7aa2c17
9CdM8j6sH/j+I9Sor/mJ51P4e18M9wdjw3wuZT8ooDHApxswq5UzX832LYkjjjo4
zT8XYyeAtHZU0CsepIz71Cx8VpWwCK5Kz8IT2vannFhSDHZwpYXB6MFvOKpZ8Dqv
RClV+u/cCUyoXb9g/b4AQ3bNi9InqCZwzQM7gupcAOgHbupKMsCOM91yhU/xfLTl
XLp1dtP8TcCD794XVdMmggl/Pz1EsHvhRTA3ZYNwQ3+krgqJvDqiyaW/x0GJJc4r
yo85DrrlavasrwMqHR6kHFMNC3Gjk24Zrq2WNvIrjTFNLtQeGw35SmlPdJIwNR9B
DHtiYSRGB1DSbH8caAuOv6eUIYmyT9mxzwpqpWvZfgz3PLwm9jMEQqj/hVRJcIpj
fafZ7knWUDcHcV9x7aB+Z+m74M7tbTR3XDJSK+SwqXCScopLmON2EOQtVyE4L8c1
Cu30DGlawaRju1/8X/VIQRpcH8+kLL4uJCTm1aQ0XIy/rr0sgavg+J0zRDopt1SV
GGHRvgDHzGUMQf8ANCgJxXEmtYvP7d24PGqhXL948LEQF5krxpnZVbhb3MBeSgk0
Q6Tp4v/Hiz6GPfI86XTf39eplNbQxNtfrnUHVlgd9OQ9YiYTqMjdbD3lJ9/vtGmy
EsLgjlPaUT9p+4CiWXpRxeOVu8t3EegjCrmCJvGfISptVWndF/0dS9XwkjgQQia5
PT33MyNUnKDPMtboXOsFhxULINZTbvLNcSjsz9Grb5Nk37hqfnCZl++FpIuMtkVL
5OQhNg1bxQdIINkfQlmAEl4gFRu2UEj2NjcbyHLrt+iXaWsy27EoGufjzwCuxVIc
JUNIW8DlYoJCQ2vM8sGWm1zpkSldVvM9L1i2Pxvbp5GjG1X/IZt90wJ7xuuotEx/
3pRMN/5eUpzxoMaWnRlfH3zt4RJnCprqm6g+4HZmFaqagZY+3oMxlOxfU5XAhKJY
Nn6wGqGZ/S1maDVjRdFX8RZw2+zmIkdbhAQDEky341QBaRcDZrVU/9Nnwa7/ZEVJ
c3Oe38gGWt1A7ozlZKC/iJx9ItOx+XTKnEq6HsNu5eXo6QJtkSboLxZWQqpMvxO8
wfAIsDcIeEJJGIlotQHr5yg4ohM8+V23Sy/sWx6lgmCIqxCHLVF80kavet+veUOf
VnsxOsj6PgdVSQIs/EIppcEUHuLRWlCaxfpoCFziCz8z5KcuZJSeZ3zxLhBD0I/E
qoj0uIyXy7tUSXGsa4Rw4DNilREcsYYPVtXpTShAiHHTU0/9Lg3chLuiQFiu+GjF
rGdFDe4660Efx1nzPvbowc9pHp+kVvOMi6LJVsR9ZuJEqCc+phE9HKcr3/DnjRsD
UQI64Hh9nAkPNeJ97lQ2q4uQj5N3hnlbR7iUZ3l/rJejE17rna1+9FyYyJdNsJ6C
QgTJG0upr2ndKvaOXZnHjfltGVy4/vg/FoZhWQZuTB1HylApmKcV3VIN/yImlzJc
SDg1zdIROijOhZma22+U+kg1/bFB5LpoT87V89xjrpsKvNGhZzsD7hTAui/Kn4vH
pGNGSI/VBnLs9pH+Jc4DX/qHui/c26WgERXxeicFbOIkJSRUhx0mHDK7c4l1vMkR
RdCyd6O7996b4RLGi7sI8iRpHAuRh+rQFDP5wTECnJpVpj+ddI0NVCYzWRSyoviP
A+l/6Yd9CTAw9PTT46dHH0Dd2mCV33RKz31rlhc2ZGVdGMjDzLB8kRCoVuY/6SIh
N/jmukJJmnhXk+RoujUtjhkQjiYHw3CpQ46L5F2UGhNOsENJ6d4wVIL/H/iK1Sia
4CQQ5LWEjc8ajeJ/boGEW3F6a2C6Hv7vy+5PCfH4f+FwB0IFhQlMTyq3I8tPyPwA
AVHJnAzJtSoUA7Y8hySU1ojH2wu8rKBCHk9/TQPSfiTYR4lKdIaiCivxUv3sMhTJ
4eNqrlvhDS9PAp/mHamn5uZICRGkLV+xaQCzuI8rXRckjxpRYUWvOcbDukEpl/If
58xW5qzX+l+sVvKeRKJvC82nVy0WU09FPkYt/GCE/5YNJmnQtOCNWmUi0TJGVarR
UKgZnDBLa9/J/c+Nxfd7A7asAKVacTi+IJFHdixtlgvtH9rMgr3LhNS+bvBLEy5T
jBqlxtXWZrntymVyLyKSZYg6VVcHE1HZ0ThUfnbYQnHMjhouyOVDCAMmgZAekDA3
oIky+oF46w+5egBHP/cMt6Kq1RNnXfcuQ+/m8L234473bwrYgAp8URxqhHAHkASo
4XQjCo4mLd2LnmPZWfF2TMXFXRe2Dx3Q5tc4JTPuWWLY7liXChPZNB5uPFfIhiKn
mHQOziilZAWfXNHcP6JiaIIS62i4R6ERIcc3j3BmyS5ReuSfTVuFnH23FCWo/vVq
c12KkCfbEPYZSFTvc96UT9sWm896WbFqDfwnUjgg5LajPQmuVvzQvgsNibs8453y
UR87Awd172+RjMDjuvaCQO1lba0aXQa2vcd3iWfP3YyJnM61ybtvspsZIsnhebAc
XMEKFldnaWxDS+Xry420a9YzGCPmkMQzT5W2VhZqW/TCi5eE/7yAv8bZu/ZTDMv8
qKJ2cVS5WCNLkyQ3VDIhEYjjGR+LHPDfYkErA91et9LxfsEinaGCYLM2BDrpsSh4
slYYKJlUWhyXedlcQ/UXbNq7FvrnpSSNFndqCpgps3UQKmiK7oToScOPq2QMyI7G
96J+LUjHB9EeJveUCILbPAW8Ovcj/y1odu4CIB4CE0Mp72PvuK0f3ORp5Jb6Oi6f
RrwJwgMYh5Tr9btNPzXpXV2tTdlsqmkHQGfWXcWluunoCUomCxx+dHao5MKmKHzz
JWTJE7D2Rt570ilziN5akCGmYqH6tJJZ5/38q+qcJbbuzwhmSQOML8jhaEz/t9MS
9EP4Tbqq4+gvDWA84mjlrevSb2J02ZXxcpEusN67E2R1Wijp4OJ8HOPVSxvrCv5+
IET7zrkwFMFLpA2DHrGHEhcHASaNBb2pvZERLes5HZb7PbruGRK+DEhSydFUBtnv
dtnG/+7CnqXBknStieNj+eqLTUmINOVk8u/lXLnM6bLSt7hDqFbqE+fTfL3buZma
bkVmiGN6CmehpBpfNMZ0c5ej+LFjDjQkKFoSI7pEsHXporadhu/1Nr5YTdhYSlf0
CaeHw9xtlfGjPxj9B6eox9e+YQxLNPVjUrP0TfmvTs8xsIXJ9kOQSbMzMbWKF49r
PtvjCwjyeCRmFpXBqDYEtBYbKs8T+jX5dyiHLY1YfIttWUraM6q8uRj3fXDaWUPT
94xbPc6Zt+jWXSau4CdjooL2+NxYEuJFfT5muZ9hRTSuNRRyyqSaQ79pn0710zG0
mdf831Ri6cI7dIfzHykYaCUM1ljUuxfQPq6bVh8Kh0TO3Zj4GLqtQIBGflQJMBDt
e10umxnNmaOZUF6XLDkE2zCyMrXQUuU2COclC5dGLdOUFcWMyAqpXgBBESktAS2i
Qf6uhxui2YBMbqIkft8/0LYXtHd0Vq1/qsns0DDFUsgMH4BWCnolRn8dadiCnkdl
859pq98ILgPvFG51hrl61s5vnVtabslW4xuwZoSSpVHsh7aX3u74n9XfJmeytz33
tGWVOgTbPlVFJhGMcSktish+dL5q7JsOLek5JqG6gezKGqaiM739p74sxQtxA/f7
GrLhm9bWHKu94f3ZMuSEIRP+Q+KbAxtS+2fCqGklxQbBcL5LhYig/ccMLna3lWBp
B3lxKwhLP0lMCpPKNlZXcvDwmVUPkIvuhYrnRqr4M4aPA3ZegCI8awqRXpy9jTNy
glslfhyt4lJfTzYtPFHCfsx2limpD+F2tAsdrT6jbZCrJNIVBMOTqST5u9Xfvajt
ob6wwjg1CWhzs2sLuX2W4BBMrhYem9t1gqWUPng+HdmcZ2YubmUFOWLh1qiOZCs/
gskbR4CpT0jSsRECDGoiC6EKdGk/0t2lOlU/OMAE4A1ar5nFML8bsB5K8esHQ5/N
hskWLPpTt+TD16wdJe3A4fXqzlQxLoU/do2ZfLtGKMvAkBumde7AARaMkMYJX69u
QNvgU2DWXenB6HuDrK77FrbzRf0smM5lz7Qte2vM4JQsgQpygJF9HUIYC9uggm+j
Oqb3QdJMaxo5tnnRSnHyAUCIZrtq0XjawHeJPIIBhKrud4iokhGjJKVl0YG8hpT3
Weo+J90hzaYv/SQ9E+YMfgT8SbbjCMD/NKpiK6FeVvOqHxtFn2mtc5aRCU+zEcAP
LRmEFFtrQurT6LL4pwHeUPS757r3PJaq0lnxnyLqsgT/DWO6/Ch2LUrYWnUDJRap
kKuhmthJ0auoxlYd9+PHYWkdYP1AZVhDMYJc+S/qm/FTR2J3tJqoLMH8nZTur4F0
pNKer0W+FC72btuTdJst+7oGS1QzhGUE7fwyUNNLIwNEShJdpPzEHPr7PDCa8qJs
5yXjpNiKjO49tfcGD+49p6ZpXaV9tzRluYhHN75I1uCvs6mckK0cUr7NprFjaOsx
tduRAhIXAP/dmbWmdu6ZFcdFS5H4IE6olVJtEwI26pwqS9RzGe03qig9gHZOhAbd
ZFINC/nfwxizKXZFTdAjw2FkOcHqAHGwZYH8+fmSqvqSEj+YZnlJzmk6/GqXiG4z
GOYpBjhs49Qq1Phat7sA/QTXPH7yFlyLQMKU5VMp2XkJz4kUPAXhc3fe3j2i2CXf
fGVfgjfUzLPa4RK/6TNPmxjl+7CAMhUk4z1d/7XOu3LiBdWEsAMntIEX3AsQdJXY
PprPCwujcTplSHAGefQT/9OVK/Of1kDsig0NzqkakOpts0D7VT0gOS26Lj5D/YeH
j8P7TEYRYCyOtCTS7UlK5Vi6ZaRGM33VlgzORn1ib6nvHg8a7QudnuX4SGAR8luI
yfKPb4oUb/vnXNKNgqt7j77e6PlDUN2RZmpJa8v3EvJFA6zbLR7vY+BLrprFDUOA
fR04iYT6CU561rNh5sGJjc6svjtIHemwNYsHQUfnJuTjo9gjq0nXat5HQ2Mn4j2o
fnvMuxu6RG22yNKow8QRVpEIRgnqX6JaFt5KgYYpp1SzxHYi/3JMV5PM1v6+7Tdc
74hNHHiQdRjO05JGMZ3PVi2LLPmyKSmqluaRXypixn7iDfjIOSHLozUMk5BZOeN+
KT0O9hzYnAGFTSCEvZi1iJAAnQ08BIvsnGd4VJd3uC/qozTbTtfc1f+Y0aqwLZ7D
jpD7XoWS6U1vPeIoKyvZj7dSsVWGhYmsMX1KZTv54lGM7vaLntbI5agTm6gy5mC7
vDfgEiwMmT0JFVMAYr4T6VHhR8RQDF9PDgN+u101GsUGeT/sUv2ApZ8UyIiXa4nv
eY87TGD6E+zeujx6yUJXKOKdo9Tn6MNeGah3E/dMInAAUIAHGWlArJP8BRDaG46L
OSnw6UjFs9HRceL2KutNIkvG2TckD4C+GFMWnetHKn681z5qFttu+v8UKIekr43j
EYUOujd+Yrhubg0hj0aVBgMaCrs5kRTW4NRf6cEH9Z1f5vM6FxV8e5D7OuNG+gfo
5vx7ZKuAWPtrlUpc6zj+kYPp4q5b/D/RH7PydQ8I03vMadKl46r2g4w42S/8RJDg
QZvy4tfVGD2TMdy+G4cM4oMXinKEr+N2nqxZTRJ19kSY82RSSTJgg9WxorLvuio7
VTMfXfgZCknk3KSxz3SyQ9NZ3+7AnbQI2G5NDABm3A0K23vxa45a9b7HA1YlqI13
PEfr3KcxkgKPeA+KWlHy3Ony6VXkaHMTgkMfbCERk/zeb8GYQy+mRjc/R01LByTQ
pIk0Vhr7gviGZ997yWo28wYEgQsxUUsF+8+IK2/Dkj6UPdrbrPfdrqYiqg2QqUZf
TTfW8sg7ehV1RanGM/1yBSZTqRU0aVk62dakIaby5QnXCI8MRyXjfYMQ4Nagpedl
kh0W0hW0SWU2H3UBBgkC8C8ycguFNG2WKT15+xODsT/3HpgOA0siXD7iThmC1wBG
+t8bOknHSo+RD3WWURhvpw==
--pragma protect end_data_block
--pragma protect digest_block
Ny689xmqtRqTyw7p+9Jn6K8fDT4=
--pragma protect end_digest_block
--pragma protect end_protected
