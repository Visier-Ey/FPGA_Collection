-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
nRHvTPtUYnjsaxdHe1qGsqDsX2tHi6fpp/El3NZ6qdu2CZdSxSoRIPgQRatx2fn6
bBFaZt22XqUWVKUkfVvQk8GSWzpFxNImICjGI1/TTya8ouFhrOSENPoGManleQj2
+bJIff2E8TROvOwebVjZOTjqtvr7G9IXNHx7a1eqcI8=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 8004)

`protect DATA_BLOCK
b6euXTNTcAcH/oKTp6bAeciZDNftwB/vp2WzEMJhXXMbq1LEZMPH6uGAlx1I+6ee
bcT0WpQ7zyIq7+KCBwPvWqaOXxbytjfsveMMfaPRl/3iFqFzk3Y69QhxYlNQz67e
G7m5i+UOwSt4Q37XyRsEHzqHUkTX/yQYrcXDodFNwhL3/RlKiEOZS1F/6zUj93Hw
l8pheMuOuiPm7l6DQYG9nnDgPZxb3Xko47aKrBy73kHGDkRbqhdPIkddonMMEYcL
z+fB9P/lGr9VBeERcoEaVvHmoXr9U8HOTn5IQ5PjZSdYK0oNY4G3EKaWD2GJCgVh
zsa77UshQmgciqACtEd3+lKFA4dch11WbvmfWO+oOZX4JyIqigUbG3tu2JymU6H6
/Mwi10H28FoOA3oF0gP0lAgUFWVs0gmO98tMYK8A/BRJNZKxmlzbCWiIjezs9yjO
a/znKmi/0zCL7EgCnhpKwTfQ6/MTdSgXqzJFSCZAQBbq3d9SnP6ituNLD+r8zaB8
wDAvDOTPoaUtd43xMyj2cQMVLuKzCcRNtTo2SUgDkElLXgZV4AgVJPIQ5nC7JOJt
s//ShTV4aBrvSrBjwo21eM8Yxpqji4U6VFK4g2pY9eHdI6H8zzXjjPkbNkcezVfR
gplz8PjH2Njxn9ppFXtW0PqY8jFuX6764zGeFVPeE6d/08lB4D0I3VV39s8v5NYS
+5+g3c1DsjuQFCiKz9gAfptn10hdoSmo7ecGAz+QW7ZfgKfSI6Txb2r11oJRBF4c
HIxBKohxBlJGCNvMjFDdWMot43qAeseV1Bl+R/3od6XPHyV/HOi61FADNQsWTCNn
iDVtK4gaPI17TAFmIGsGcfOBv9zX36jDx+I1dk2bBXQ9q7bJ6LcQZDCSg59QtCRy
/MyXEGVOjL9uMruwGK/PEwRWp8Mi2/x6dOT+d4hqIKQplvWyjtEEAAInKvqsnHOP
CQRjozKM1zd4IHyL6dWVqtj57rOHhxo/UEKNke/Z9GsRQBtIidTwLemhy73WgFvH
Sxh8IMn+I8afiDoh4rNzRAbQ9TGyPTv3xUC4tgnBTOHLUaMTIkRTDWeqJApLExQq
LZuCxHOL8502HhFp3rmibER5mQpRb2R642jj2UT7irrNnKH/mpSzvUtHh6KQRs1W
wJt2yP9Ns4GQ3xPRUGxl1RjhOH1OeTqJkgx+jqkv4x/o0oYT5OSc84fhhakrOpp5
rpbjmBZjm6ogWl1X1oZQiWPT9+vaJBwKSIagqEZBFWUitHAcYRxzlLFnitJab5xq
l34bI6WurkAc3bnohLvM2/RRh/5pHpuo66IfswOqmTxSu6WSUPhW6176yB9qnxDT
9wH58PSHLvUoqBdUuyJuzK3lxyq+xy8Wp6rSdlVosVDp73BiZIR5n73uTxM4iUlD
xJXvA8kIM3pQ7O6FooR3hZRv6y57IZlR1Slcsv0Xg/j9K8Ia1pbpq4IYZyyeUf/F
VDUBi4bS07QggXGtqUc7DDhp8AkY8tmvnHyFdzIQY9WjMyOMgtdXxAuZvt7pbOrb
hlkOq9IaxkvMRMdk4I6RR6ULeeYiJv8t9fEF+h9EacX10vViNCJnMXmkasJ3znkx
ZaTh+dDDox0iuwObudkhuefGGVAb7odSCatQilofx359ThClSMryohS1FHED+1eZ
hWMrJFee8gTEpERfcuRreQQawqRBSMd9QyavOhbDy4bIpgBKCiByrmGl8TMgJM31
nk5aN7siaTpRQWLDhEgw5/NeO4ow1jhkgzKr2+yj02TqUg8QLV1MkuDdAWeiEC8C
7UecgcfCjUhNSvIX3HEG8OcDmPn3oB5zS+4SH76jEy1SaAZePTpo9iYSdnlck6Ww
rvLxxzk0jeqW1e1TcWTHcq9CIPsKTWFSLB7tXZZ9Z8+9t5LJoFMQ/XllvZirD5AP
K01/MG0c0OOP6Nu+I+/z7Or20mQT1+SLJ5ECs/lGJp8HAz53YQKTJJJJ0cfcin4p
gq860jip/nk+Fkh8C7YM+YKVkvmf7du39vwnuMhwbZrTdUBfpVZlEIlWZ5ykyd15
52THy2IWrpwpp8/sg4eMFscq82B/dw7HU0GE0i59HjuWc7aT0Xp88tph0pYJ+Y1+
7mmfF4sb3Ictq3PC2GdNuH+gDLi42Y0+PnHskAbnAfCICxB9iNZ2eNfSFQ8LnbT4
HQm7I5VhQSVAeb4yqVaMWQXCQHutWwv/fWvUqgPLYm2YgrjZDPXxnMMQnAISKOQh
GDXJz1Qz2+pW2Yk+HhQe/Z84o+THuMV+dab1b/XY/6s7h+ToonrsG1xj3GW4rKDl
X9331ndfIJ76UMYYGMV5CoD0vluWKI6KdBho7JuXgAlWniN8rLkRbmeZL4ye3Zso
DgtRgSK1hG6xHWSVDLutvTuSJQnJNDFCqUuKG76LS+ur+fF1n0/NrCaR5PyOwhGr
6RqV4p0Vb5F5vzyEboJESDFbruexVMXtfAJbCQA4Ul1JsrlpCQZs4EG1mksMWP9p
g6QROVbwvF0RJBtSRsxFlnT58+3rnDGJBdhJfkIr9u8Zb3Z6Uaiam5wSy5/VLWZO
sOwnldYc/M/RdrJMpa5EIxonu+3TWCxLy+okGEaMUd5yVbx/Knf9Oo2uTIdrXHP9
AY5wqY2FJ6JV/AdpSk2Idm87T0wFoHZLFrmFzO79CFvfxQwVoYpdLGF8hI2Ffypb
V4WxFKIM/Z5o1aA6CXpVnh8sDevfTY0w0h8/XJHHCvPdpXupaRP+kp2ojYqcaW7X
UZwDkopdCbqPCOKSPy55bPI8ObBNnbhPTDkPQIBM+VRcMCNgFw5PCn4gB8exmWwN
Zjf8bAc62b3B6w5cnWvQpOmyT9nS4Y5iiIuP9ttKLZc0KheijpdNHGAEbm/RfK/4
yksQBlBM6kb5otrxFIh/rCyFkkzEEPkQTO/GxfNCSYSCD3QhC0Dquk0a7KufY5yO
+9+Qm8SjDVWxS5h2E20BdoEqsoP67QAqTQDIc7BjT5zvseoQvbKVMVNF+YJSYhxt
LO1O3uxIGW5BY9uJkpgwfJCMtoAqs0O0zSmIaC5xjnVM3iOP15yOY9b+3IPYnT7O
pDSs4w/n9Zx0LB1vT8IMnP/mkkQhPAAEpIzmSwklmCmIOfAlZnwviXTDCBA+hqcy
2q8EDZa0Xx5nd4+DXv2N71tsJlcnGnRb2N6tmrAmYN9/xkSfhB9OGXn6x51KmMEI
OjgDmCfmPmipmsyxIV9q8/QQ3u1VN9Hg/wTJB5FjZXuGN/M9SQ1I9i2BWv47/u7v
UMutszaxLIOx41Xq4Frylyhli0fXHBTj987FTl2PzWUn99+eUwFo2yJ9XZuIuO4D
PJngNenIVui4Dv3BFK0rnFGfPQPNz4NlsrLBKz2EDuS8lXXfKIukysYN8tCtMifN
lOk8OG5YQahALZkSxkGKz5WEpXIUwKfWctnW7/KdfI3OKWLtnBjozwnij5oXGZjv
HLAcqBi8+gAjDTn+SvCMLwjwAwSCviT/kOYjHYhb++FZxlWdmvoOZijoKSYrO2uF
DXLHdSSVJRllrhO85arx1UjTuWJxZHep30Xl9BDyhXvw20E9kk4VEd7EITJAevLr
8m0HlXFJYXUkq2wNW3S8CG8wwzf9D0RkkZ+mi38SWWbhBTOk4lp6S29xr02a5oHc
o0ewG7vhKCMfHgFR2/++uEVMD57zlnatcgnySION/gLQD3oVTP07NXXycZFwVOtI
DwAfNDz0ydOiDBTiR3LCm2xYlgX4l3ostjJYgHXJ+Du0cLXwb2Iy4hSSzAekd8Ou
WGy+QeQplhY6m7X3DhEgxafNNDYUNf+gP8EFB/j+1A7885ePRCvK7aOne/HK/QOY
BiBSBpDEffR4CuvmLYwkoYU8OBwgXuZbiM60MzX82gjrV/PdZS8Vek4qMMlJ9rad
hUgiCjgUX1zEGYsNnsNZVXrPlADikEfnXIxWlvjrztwYgGR3tJ16hoMawK5dA744
dG/pRalrq4tLQyAf9PtJI5djuMMEoCKVPeu1WVBHJaeLdXFFNe+MkFS56TVWpNVh
vE46uDKNYKhnIEw0+SlqB+OBg4JOcHPf1Y/iIlHUwHFLK1GbJ39kjFPi7UYQGPkf
16QAXPAh02wq6jKbme7x4OpR8jz/yeBigUR597oaLP7Iip/nZq5DPSwuPKUaN0Tm
uxKiopSmPcKOmAKCOcBLEKMxGRwSSV3V6ci/UXX3odBpe2I1GQUmg+joAlSlwgdC
hGur1wFQ9jbOLRC8YkDVM6J7z5Qj4IxrEVUuU00sfcTKXqkk0aFaOU/R1yqN4pgU
pECTtZ6HviHlkdxl0R7LPtzJAz6354p7+s9y4MzdMj8O635sb3JjHQQWRL2tjC4b
h2TIoSo+wA9rwKBRmA8L1SHtO4Kt4JidtxR4j96+OXVZyhhSmvmXJOinTKaOwN5J
xLB9k+qG4Un9pLkpllrDGQCpmSFBj7N7nHqsK3hU9smbOIKG/471o9DHdrkA8P7G
cv/2S1JyiRbdpqZUG2EFjRGJ8P0KQeron1Raygw8Us84LMqSI7CE4Vi1bW43amWn
kNWBAAABSd4EOI+TgBGOGvsyNq7Pcdp6z7jF5yzr/fOaLJQJ4ngDcV2rAFMv92jV
Kb3lIrusQnQPcdtYSHiYS7H8Zmb4CGnnGp1+9rks6i3JxkMtRxKbYaTYHPM5P9Eb
zay3LKZGw9GzFLssV0quVRgz4EuSfZm1EcTfG3wry9or/PdM6wqDZqYwSA3oZ7CB
6HazcVXoJ0BfRNxDf06Oarnsl1Js3sR3szK3z7fh6gCWyge2fZGBL9mT65WWu0mR
UEaKdBNfiMf+fCfsHFRteEmxTyBraQw5ZfJBbiUbJ9sVxJuYzw+co+NZoyfO5GIr
3Edwmt/8oayYevz/xm+eyu4SxU7OOysDr7hiPclyVXYwzPAyqbMv6jpon0H33s10
vtXu42LC/h8gAgjQ+qZClFhkgIXLmTtdVALE8LO8OcQ0Y4xs/sg0yL+2Cx2Onbf6
DCpvrNOqOyH3tiBWP5zZ7NQoS2Q4pWd1MD8YuBvDQA1z762cmOZ4GMHhHizwnab/
8+tnccVlIHkRK/A7jSKUfENmQlwJUDxPvZhxskH21qi16SmANpEWGi+NKqQHUA1I
kWpAlRCtU74idUffQ7o3V2dguZCRWEHprI0zCd9lhWv2dakPUCrXf/AocRJQ9b6P
rhd8npN8sdMhsxxc3k1lMZYH0t0n7vCUiZEEqvjoihkyTpbaXMnR8xO1biUAmTzN
fpmaVPgEtYASrlxpc5iY0Be90Q8FzEZiL3kgev23P6QTOEYrwbnxhSUQVrDf0ziE
amj4+HDoh3ejl7dKC2ZLl3pxB01cOhMr0V12R8C7BymzW6Yf8aEw8k9N4RwJP89S
LoVkaIzY1vMl4g5fujy/bmtnB3BHat3DoO6BdbKiI4OMqZTO1Zpb9IKxh/eHFXCF
BBcVnYBgBaZR+KRRv764o+qMEdmpATO6qUG7ncXjU9jWv7iSFnOvLZNyb+tgMOGH
o+lYhcJRFR7BYULCncJVU2lMeq9JAAuql+WyCZi0AT05wQGHOdncRozNBeiy2W2M
3OkT7k3xyHtyhkU2oaolbXcmcsdbOZ8nJJZ2GWez/OJmHm0/a2fetjpynCQ5ShsY
qL1XPqudI+q23pc7/PlXaR2g9xkYg8CNxn9+D65g1pfNeXDka+O8v6KoLOBT/sgM
PJ6y3wtoTKTYNjJHfqJcUM+iXd1YVI114xmc4Aa7UCm7jmu4R6XXnN0TpK5W0ORY
Mpangwm7kYdCw1qzQ1OrZApuVm+cQScWamBZka/wv4GmR2qEgSnH206EhzQtq7wx
H9Gk9RQ6/T/IpXj58TIzxVf2F1ofmFPOuog5es3q5aDiH4uBw/Ngff1Illpvq1eO
d2v1MzBxrBGIMGBd0h5P6rMp7UK+GdzL3QXLI4bm7yaMa67RRWW0nKWr1UzWvWwa
lp2vsB7mqP+H00LoTOYXcb1/JpLGAcJVSv+g0SEDZGbWYV4cNWhRPSj33wdWszlC
QDGRizXcIqg3Rz2e3H98KY3/xqxius4+3b63OHUwBhG4Q7/hWPv9FnH9QeYwYI1V
6l8iXRUWxIP4TvnfRwEHrT1WhuMPMCJ3oymMWZ8HjgJ/5ZYkHqr+t6GarKKPpkT6
1UMYCvxbKDmYZj8LLx681kgCwKwMI20RaM976riozwIy1lV4ZArmZvz5ZmLCMwSL
nWobJfkLWsr9SbLfjHRCWT/zXuO7MljmTYrn5Tu2j1tOwZH71R5r/q7w1+Qem5jX
k2vvbogNyi+PyP12LCE1au9UMzlBQaAVTAPaa9F57ydskUrvdGCYS2LhEw4BLPzR
cUNhRXSCz+15SZIrc+tjQT30Mj18J6JaUsFxwJLz1CPiBnUeUPipGGzPvIlJHNMs
BDfSlTeLGQJB3NqIQxo3wfLG7jhCIi3O87lLIEQlCsx4VlQR68w56Cf/p1QkdAB0
s0OQ+qmFpN4le5mXj3PgGynePsUjfCKItI1Ba32uRYbKuEcTg3pKsxTC81J8NFKM
M7uF1/jCZ/3feg42qjgptDoINLLqoYvzRi2Snz5/3qb/44Sz2fKumyC2hss60dYd
7pknIqjo05ZBy15CMmJRlCCF/EgPQsM4vjY5kIAfmvR56QTv/H9Pt0yX0HuOVMrh
5KrkO75EWbxygrM9WzA9kx8CtOwlBJf/u5I1WRtcL6JffxA/alDCgFFRYMpGllkb
thGwWL9ISw5DpRYym4dcFMIxxOGpWEunClpF4vDhLeul0qCFLv8KF3m1+6quXxmR
LwDvStY45zQzk6zW2dgg1HrJ7NLY29Eb1jr+OSjlaB5Ds2A1upHUxqP7hkAOC5B5
kBx/kepwWgxINRr1UFXAPj9OVe+YB4VZn5UpX2hpPcEj2Hwu03u5E9Ee/bSNOj5M
V643AW07tvFnVdD93dSZFMumaDXNc1KSUEpVqm24KBfv5etlKUBzmCgMYw524q2Q
rkHbqlPYRpGj0WB0TYnFAbsuldqrhiMXiaZU6nOZWtqe1kTPB3Os1p+i3L0L+Bbh
kqgkvsNSaQoNmrGYaDrCLwyFZieRS2NC4VSvlPTXuPyhNkbg2o7279oCfM3QWMxJ
Q7N9MgSiKjanx8o3HzDY0yeOLP+glffIWZxlMzctqWbxTcTR6H+nCkB03tzHog+e
tv0uv6MuK9ZZbDL5Q5X94Bfsz5J41y95TzO4YPtK7PbB1Wv0VObZ+KYNA606Popp
SzAWXY7PmxxWgaWojDcnln/CvlqNoMvBpRzICjlEmRsQBIPGMSNZVWp64x+EpEv2
16dvREBrJvmycx1igiCFwHvMxxScNAeW1VpzB7OUWjYdxBVJ7HZcs2KaoHVOxULW
dtD8zY8bmtzDeuv3ytcp+mPvMTU7aJ+tz5iCsEPrucd7BwqvW6A6HGpEdnKaBW7z
49reCYm7A2Y+3vJG8Jn9mURMocIiuPSluFxtmUCuqoJk+anf1hQtU62tnw3ETN0v
EHwXtjt4Vse2ZMgOeAbbEGbL7qQMsPJJZmpKxAVEtGI20kmYB0hLdoZqB5Ozc+yT
NS0Eo364alH2S0jfCEXxW45bW+yo7XZfO8EbQV9X0O+it5vBVl5FDRHpC8Qcm7Cm
qrHot/6h+7a9j5nA2A6f5fTKRPH9ZRZ1zrgS57eb4sCdKgFjE3KR1lUx8ob3W5rp
RngPuFgZKcD9FFs80g3joQCc9RgVtmeFl4NN9JhHQseMWeycXQJy9Z3/5EznlC6I
QpQNsT8H8I2MKv5ZaAqJD0BFptEYxN/GCypexziRe9NLEwYGVIYnpfkMnoSdWiR0
ZnMadd+5NSlRsTm+HKmJLRkUuFZsLim4h3mySyRd78iVJahqAYMFAIyulClx9d5b
oNidL8/553WI1dS0LLeN/pfroLTg8g8qHe4yJt4SgpqUfZY/NCn6OMvW/DPcnMXe
FNRV+vkM+D3MKWVIA6+CtwJUqVNgC1Hh4l0g6p3cRRwmg3tcXQfeuAF6U0KhMx6m
at9zJIb1NlEArmBLGE6G9BPeJGzm+zhSdkwy30YxWkaFWKwzSz7zbj3NZuAuatT4
378M0xQg0wHIQx4seysZ/jin7bYWeYLCwdVTEhATTCHkaXB2u1ukMWyJKv7feeym
JB+j2A2ZxygRJy8Jyt9XuA4zFmmc72u0FUG4B6QZ9o1lixks7OrRKBawVi3GZdK4
r5jyseQ1O7fSDDtj3dtvD0602zbk5TEa2Yxv1iq1Z+C4rOc8aIDImD18l+EaElSC
G8D7yiyNIC8NpQtLBoLjuica/m118uwUorSGRbWWDMGBjTVRrBZ9M647TyWVCx/7
5ks3SvYNF60iWQdJFGbTKfDLMCHjI9+kUeUiTcbzWBELf6CB0pndtgJb4XVDuHa1
jJQbskNuuscgBMbUEGF3OHFZgzzvKluCaFL6xEq42/VBXfvgbx6HhSfBevRVb70r
qk6Czqe24dTvorm228E1tuITu0s1RlB8Xh7NrmgqueWOFjsGBd5TBFpVCj2kUZfL
ey+GNalhoff3LTkOm/GJD74OdbxCc0nrnQ2Z25DVGk7vKHx61y7xJsS9TXIKYmFv
NmnIYtO1yEKOqjWPoCb42diYo9j86JxJXXEx1hKzSgr4vE9Gl7niGGkTibo3hdwo
8R4dU4fPczSkdlNGM5+ss60L4tYqZG367DW9x4gpeYRFEXW9pNn0dWegii97KbHt
c0uNdH6TqNIVCWXOqjtXANoEBTunpXJAxomYh24FTfiMUmM14W5QCyOai/FZYY5y
EJF7I/MlPCdg6R/C21K7pDUe4kk8mxrHAL2wCIqEAAIMe9WAepSxO8CeX2PAmPR7
99Du+aDdB5aB8+5kj9Ie5J6ulmnVwzn4D0HcYwFdZuOM8oTXZlJJb6pndnsSi5QS
71gdcgligxzGjw39KWExhSORlxxZmern28d2yK4hJhRRWxTyzRxKbnWqzzNldQQs
4b2MIomTz29gOvRs5hN5cxtNUQ3koxYdC0VIKXg47Wf6aFfVdQ6QO8IQEuBW4xYe
yP0ns8j6mDGYVO4FRZqy1mCMiVQVYfpImd/U+LqzH2bXIhJBsZeS4/4LVtY9mXHJ
+vGmr+yvGYG69Rrgq5zIrGT2p33x05ehZhS0KsfbUtNBiQKt5vfdOypbCv0lGhAo
IEqIJ06oix/BJNkW7H5n/Ve7MvcQZpoSbMTbT+8WioU1+rac2HU/9lDFb+ysyZBZ
Ydl2caC0aJo7+oH0EXjNbMEvrKIi6IBri3VGn2d3iwD0zxeytG9Jz7Dpp5KP9wG5
iaRQCs76Z6wTmLnCaZsGLF4AyFcELZUy/JHgI4eObH5fjQiL/xwDPHlfVL6PA4mY
PY5/l4zP0TOHJnKoAqIIxSvkmQ1rjVgRpaSyb+XRDS68U63C+XiUkcZ/eE9XNxFz
cTSsVjMeqH3N0FbcNJMA6StkdSCCeaknd5549lPJGBEIn6C49SBb/ZXJnzgoufbL
JOruO3tilYTNewpcH5FBP7Oblq7vDdsZ0AxtM/5UeZ3kfoAc7LtFBY6YblyF1+fK
wkuhxDxiC0wZbT7HLBY87H2g2adq6wEKHy+s45brhPdhlxaPeqH2r3/SMMgcoVKp
jFh22vxc7lyCYI1QzxPK9pU4/yLpA62WpmNY9Emh+OUuiKK8zicYGdSXjvAGr9ap
OLw55uV9SJZBCr0+4RNloe8LKFH5/2VyfnIiKEfFK5gmqMzHufif+tdnfS9wKSZD
GkyUbWlEyJNjIvJNQzcjZFBEcw3SlTGIMTOt/OH4VaFcz/D2nAEbYhGQTn63YVqm
onFeYIluQJfHP8AVZwcFi1jA2HSW3ZKY7+gZmKnsyLu7uqV3SI5LqWt4QzGptPto
ohr1FhCxjt54PjDBKj9YXpD8mWZjiOn+ioUROkTSKXr9miESsP1v8vCWF7YP0qRU
FNJDWNcuhSDzNH8r9j/VEU4sk7X1Twe8aiJ9SgsVaq593m8KoZbuAj1tXR3tl0uq
K9xjBFQHW8zy8NMnmBysB8/zJ6R68WC5+i/NxOyk4DrX+iVUqWvuFA+qbOXjZ1cT
3K+WwQ24NQWV14LUoEsSfSjkGJlwG1Uusijzmxh3zG2+Uzd/b3+guu/KZsaz0G29
Jl/m2VFUH9jz/9EyAVN9L3xY9ApRJ3tiRPyldM8C6E2NSeVKs3dbLueDL4sdGSWo
NU3dlTd9N0rXLPkyxYH2atPF2q4vikBXJKJmisnUUgpLa33HE4kKI2kYnzcOwr60
MZ0P4utLEuhP0Y4jrGKWDxw18tHtLxjkKcbDTGr2+p5KywLw68Mslyj5/hdzgqiz
eWStNPhdS/wz/hdEq8De4DI/vAsRE74ixKkE9GYdAsxzdIpveLlq3Fc/mDBaVsJx
vrJqmKhSLKExRsvikhfohmVnAfwuAtf7gQRCY8ZrP3sheXPCR4yBxxq/Ys3Uy5sh
grNZh+GP/02wPpKk6IUCJvkFNI0j0t/9HPJ6nKaSNckTLG6gS01O5wtQyHdkiyjN
6emn7lEqMoDcVKoswKm3zajbAQfHkdmvQGkwr4dDM49mn/e+HLaHUuFlAYZsA7Ne
ZqIcPuo6ZXQ/Fb3NLcH8yzJWiMO4w+92DVXKwErKFqs4JsHsZi2uAZysYVjtrzOM
cxFET1sqSwYbJMQkoeZ5zBypR0NYhAE1/Db8ug/WYNb5RaiO0MrNH+liEPk17+CJ
KmUje/54fURXZFpoP69HEQ==
`protect END_PROTECTED