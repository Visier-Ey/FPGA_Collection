-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
--pragma protect begin_protected
--pragma protect encrypt_agent="NCPROTECT"
--pragma protect encrypt_agent_info="Encrypted using API"
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
--pragma protect key_method=RSA
--pragma protect key_block
SmooZNXlMo7ISCewDqpHe7xLp/4CLaBYkvqhWwsR/W+XuBtwc0ZsYY2FRasPOVsi
cw4bMa+MusLOM6ygZV925QN/rjntN65TMQ17v8OM7izdxjyHNX61xPVj0x9cpKc1
l1yp2H88n2C1y5d4ZzGUlxoZMH5cuU57zZU9ReQzChjP/bW4kf5w7eK8X85iY2oX
L3ZaJRHZD7av66/6tE7otD+E0kR4EpJOHoXXmpPe8d7mK2D/9l/Pib9ECCs3Fjr6
adpEJEFpH5e68i0KP3g0kH6Bn+HsjKovaW+op8YcqOGBVkLVqkLFAWcptgFgIye/
z+nAMaoXuDHJujT8Oo5SMw==
--pragma protect end_key_block
--pragma protect digest_block
N5bI8lHJiaY/Npkvt3j/SGThplo=
--pragma protect end_digest_block
--pragma protect data_block
KslK7HKnRJ/VChNbtuJcWCgM/GMUk6KCBJ0uXVBfzluB0zxfTfKleLWhYg6uInoT
BuJHE/VqKzv6nYHCPRgU7rF+JWWvC3PzA24N57YuKL1LeoblahMODDwDmEfHNBaP
bpq9wCYRPS2KUYEViiKVqQ0kPW1ir+YWPdbEqijsW1E8JFeSgRprFG39EC1eqvmy
GM3+H7XZdmXO3VPKabb+a5TKslfvgghmPWKwWu+EvfY1V0O9VOHp9r+ud4afeMPI
ho6v32itwAwD1s6uv1bO7bP6MArbj8R4rd/J5eMfUJA2P5crZIFnsl+ZxOs3xmVk
X58/+nhyQmizx9JD0aBPR8L1rpapqwGt83gRzEuymi+l3OGJ9723+C341NCAq3kY
OxjhR09jKZQAh7Rt9jPpsW60L8Ww9fTHDhsmrPXWL66WhYhJ5HI2UDjT+4U6Oz1A
nBnVYUcr2WNBWNxE4e2LAJfpOZCbr4HT/8IWrUqzP9PqncgnEXmAIORlfB78qmX2
3GEVCQmz5mATmBWP679n7FFJ4pN+7x+W0fnEXH7UoPWSTB0Nm2I8y+35QfFWJbGF
728Jc+o+I4+rxYp5DouY1pRDQTogCyYNZCGUHc3sk4pqDIJd1r4K7B+8tXTqxXPe
YYEo+xBaesd9Qi3W02KYbCZwywU52lotvITRB620oXqISHr1B0rYHTmFpx4d5pw2
2qmOPpcfftJrQlwjVh5oobL4Bh+LzADC/S93csc5mcrLDMSgHxcbkwrDIqRyJYeb
PmhT474dP8nJQyM0TUAS0hvT9xmaGdL+3NFLE8Hv+W3Rl98M8vmGfGCYR3FAIilD
xPobL8W7p/n71YAh8F5Z3IHaOtjv3wkzArtkk+1e/CDvqeIWkrTAIDiMrYwzgW2N
ruTkbFZgxO/SzHM1yN6eAiaGeTx73Lo6ZYGS9lnwZRwsaZ9ZBSX04qos/N3eS3w1
ZvuZn3SRC3zgqgnHx0lKiLMtWQF0IseerkHKeZFHjxXYRShc1iWnzAG7c0IgRilL
x6TWidjEVUbfOk4JV9UNnHEWooYljWz7OkqMKeXqrAfXTg5lv7LZbVzJXQ6mday1
xYEv/jiYG0EA49ljzFEDxmYxfiuR/MIFDZP+8nswzzxK/iOHHM/KRop74xjM6qg2
wZDrnoFyPLb2PuCw4eBCV4S4UeAbDBj1upoqkosAqDrVNzqPauVqG+yZGmquqUCG
y+faQLaXM0KfDaZnminWmCVf+oQIqlcaVPIAXKBMuCHvyfeTG0iAwTU/mZi9/0S+
CDEPmJINZUVNOJoQyOfcNMciyG0403JV1z/NmJcjQaWRGt/WO8hZJGB2/t3tOvgV
AzKTWzfhEfDe0rZtxVX9XtyE62hv3rAwR+/y/wwXREKhPaZkSCSlaz8m18xl/Nl2
H55+y0VkjGEDCwUga+4qxr428pv9D251YomDqk0z8RYyP53ViE9F+bbloVTkgCva
NfpLL2SV5QZDQNY/kGx02+kkedNMHeVPsXoraDqKKTFM6gzXjkisJF++vuacNsjo
CtqyvgGIw+IKkcX8pa2D32MXPBlwpLaHQ4pu3xAaHkY1UUDWNPXUxNXFXVkyI4H3
cZ5OYVKwr+HJh9bfHL4B9hJpdSyoCNtHf60nnAYSuTYexjv6Nwt7Y7MPHWb5nw+C
anhW1lP5tHD9WJ0DHiUZsCrjiIEn+X/JsLaFFFi51lGgRn4b+dFGUOlWYNdZHycG
nMcTxABuK+aSjp6IL+tPH4E6oSqXUhu4rn5aQhCH8DvlzmVP9d1GrergaEg6DfAn
I+WsmNWVD8642eyqDU1ayrTiqomLnzfyFTmXWE9zotCMUFMsmO724V4fA3T+ZeB/
XMaelWiNeC+v7Kft8GIye1rIwHSpRXsFoYBRGntvmR6nqnZEkzLbxbbvZRYIEO7+
HX0FIDEODj9Pu2dQN9W2ey427LgACbKgvH8RfJ/vz6KculfOMhYtMmRRDD9WgJHb
7a/6tEon8Rmbr1pNM2Lfk9gdLhNgXyIKlmxBwXq4ZI8rZltt/oWzPzv8L+3q/2Kg
GV93MjHkEGIMBcxFWsbkx6dKDszO63qOhGZzoW9Erxmyh7gD/CL9pYBdhDf+EPQI
8eR4ebOFgMNwr7ZBpHI/dmpDMWhnY1iyzOYQOfeTqjJkGkssspn8gjHMuxcv4XoQ
6OVl87WUnievTDb8OZSrL4tPC/8XoxwgMPIq3HUHag7U7ki0w3my7Cab5KQBj5yE
CZcsSih1vMBrlLEzQM46iIo9VoLH/uZ4tS9DE8L3D7dFW7F3M2rhbsZgdsO+7u5H
wSeY8BnThfRMQDSxCMl3leRgqK3NME35W8Z14KiSOTRGjVAhMI89pAqLWUk9y/aW
BVd0zzeKWpsgkBllh8vce/u14uVJnoc9kUDf9mXVFuNHubncjWTQC6pfuH+kiBGS
u7HFEYoGLjm2pwX7bP7KN9imksGZSbJ9szMgCTkxBnSlPttWpG/47phWCCKAW+5N
OBRmgzQNaiBl3m8QeFz6Oo25Nvh6uFuW8k5cnVQOK7mppQBO7+vBA+0gFuiVEvNQ
LDa473QKPskDTamh8+e3IiESxyDNrBq3RZ67RuZV5mxMQxWsS1RV8E0Kr1Am24Jk
TYrU6iDxa0sbzZALP76DdxEulriejORLApF/+w06qvyRjH1lAxtpzJxIjNioYq08
OpwuJ258Wy6I+/EabT5SW3vY10FwaF3aetm4EHyXBQKZJh2/yydDpWnD+dSL9EkO
xvhwBjKYfdwZPqj1Hf7bihO+WeCuypt/HW5o8EAgmjCwKkmb8h+g7iNPwMT2hpfi
VlWbX35A2HIs0pF2Nj/+cN9ZNsU7puXCcIXgOpDC8jbCIH0BPOr373myfLxinM8X
ycKgX1iAm74DLw9uiCI2XtRz8ZV1yB9gGOGSkjc0/pAlRql20B/pZMv/LMytrW+n
0L1jcOA5azmpgQ7EuepDoOiOJKxHcbH4CclugxgEYT6fCbMab1hxDPNDo3GPIBkE
0+mEnw/1LUoqHebQi35fBgcF9/Q463sSbd00dADHcGssqviyf/wwC6LcwHMOt4Ib
0uAqjdjAW4Evz3c/mkC7m3G4yE++zoysCVhCTHBNa2BMKkGEWQreMOjnBsCMgDGi
MXVtoo7jjs90/W3hAeZ9N5o+rCuNipwVCJV5p+RNRZ22pCBH46so6Hg+aB4fKcZs
N2pRwima52nzCj0yT3rYGT18Z8ovyD9XvK2A0mskfUr6oiExNW7q3dqbODLWuiU2
E0c3Dt3lhHEqBSGrBBdp8DU3H16PRvmv1WfYLAVktLFmg4C4Yo+AoPjzVp9xpzDZ
9MfdTCK/kcPXZEXWULU1C9afrytSjSsXPgnxERiqqEh7MBDKMJWOGeqs60R2PMYi
UZuiyMiFz1V5TkUrAN1a2dMsV6jeiisk81pulEVWzFqWdH5oXsB3bA4NTwr7WExe
k8LT2eOzuuO+i36MgPF2rLg7Gf9Jp20NGCnEfeEZ49v1NVRlQTwZYFLaGf2M144B
yZpbMAKIdT3UlI31Rf1vB4Gj7ZCv2MnzZtIIFrSGON/GpeySjTLwyeXKcEmWNAbz
yH5E/UvOv/gjL507wstoi0ILKmPen0n0seaDVYRCUy3I9v6isMDrso2GQUizef8v
1zipms9PxlMQcuUjR7BoW4uUDSMCM4wtM/h9murLpLmX+KghHJqmG6RaSUzsYWuy
JbwpZpUefsvH9+HWXVNVM272sR/3Vh0rI6Zlyd3OExG9zecpx/8ikf6u2tYQrc+u
3LnuJVhAJboY7uwyZIf1jEaHctllaascLMOjMNWiqPKCgs0/nzYYOa+mOIX7e49k
m8+faSju8hkjnhZ4ungO8GPVpRcbfyYxH1lBDwAemv1LxsYc6apIq+PVdB3cfojA
bnBYOCDgCoMHLV97AKst6095fAcXdOtcB5o5qVNcpwDetetejeR9kbRkfpeG0MnU
JhdmeHcSW2uATrIxvsRxFdD57ZBOpwwv81rSHoA1Yq/nfKzcsYh7k1IwRRL8yUsy
9/bzaanKC/sD8zRbxsWypQMacibTzhbvWiwzxQbR9smqLBBoD5Klj7e/m232yIeg
hFw54jBJAeIM5EgWykev6k2ALSiqc8FPYK84oBJDH+EYf3DnKmdsfYjuzB3f9zWM
Vvu/QBcTdkAyqyUO1Nds7Du6IVhkr/eMIMpXNqAjPzlEo50xWe1HN8G+SLkzWPyK
T42ugfysCBiaqMaXTFQ6pu34Vt9ABwT/tmuG/0iw03sLQXdy9GYBl80QtmKvY78h
auQyKSpnWTJyyZU0G70HpjWyKaOzascZ+g2fG0wiMUvgsBpwROK8CYOo7MmzW1Yv
3mtt6I795CfHOUMkcvdK2SLFHb6S2AcUbP3U/uCqbsaCnRNSXpjNawinr64qHaWh
2FYrj1zRX294IH8GZ9rnETWoFhrTWQ3sBMUBwA/kYJA5VUjksqBoR1Uad+VUSa75
iKo9rRLoEJhlAfyobQApTDZFxBoHDhVw4oiHQ/Vzf8wCUeR2/Snx2RN8/unuXhIS
1tMf9sU8+VPbeoG5Jggg1CZAgGkZu3xbnVqAYBLxj4S2OvRABxJzWORZ0/knYpE5
s0Fm9utj0xdw4YAohyn+QRfdC3r7mHjednfGUw+YDyUNE08MOSBO9GzhaNYmf4j3
Gp7hDTO+pnm97kJyReh0GTldEDsQEH2Ikd+efTo6+S0lAdCykEwOxWaBUz1z+5DF
f+XxmROlM+4bcLl26GWeO3ANmUtv14gzovYEYCXIw0DMD6hFq5FRjp31vtsGYdxb
8nwB7zd4X79riMcMrh5/dTwuFThULgM1DjKmvOu43t1atCj6rXDVbClD7JhgzRvZ
ite4PVzDA0hdZ3AMQyLQ2Sl/qpvZ88d7/zQNni51m2SgsuciVUlwQcq6GbQpcU1F
KwoNGEEilRs/dlbIPQKqfGKvMUU22t84Yur+NJR3KDyD6PwKVBzJ2ATh8j/uJ6RK
hS77FWLpsPRy0RVRneOomHwDvkod907mhYP7cSo0toxChr+lwn9dL20YqqQ1/oUB
vw7a+g81uuYfNIWZ3syqT5qz03hM5/PSJSzKzBfHXrUtaBmBCryDlEqUU+gCXxsP
LmUS4nO8r2zXN0/Pf+k0vTCG6RtiR66Uw+jocq+lKtjQX9nUMB5Tf+/23jx5Klyx
yWVwWwgVwqa98BZAQgGlrRMV/aT9ytmLqNiymMBhx/Mqkc7zDdGkDnb79ouOE9FR
ett3vUD73Fr+iINDnwWmEVXzYYNx0QRqU69rrlpJimHh25Cijaf9IL0p+eQHx73e
x81zIJbtHDa0W+h65Tgvxn+kpaBK5sU3Rm7lFNNJEOqjPAV+/YAkJAHIraiGOYRb
BcLnAs70HnjVimbQthwkZoz9zNNsAejz8Vp0kI256lsF434QUZIuYvVcAOpFBKGM
eQq7oTNgMUZy7A2TC0t3uBmLXKeiVgTHrfkvq0bSe96CjB6CoIAOzhkZBjBp0yXp
sSccTdNa5x6yxNcaFFujUUIcto7o2EiBiJOPMqI3wLBddY6Ff0VhbafWw1iNMlhS
oB35FHCNn8XJ33w6ypkAD15iQILyxSSdfGNqTsNe1jnjHt1cOY0jp0zXrF7xpbkC
bFQDLZGSYNEcLMHCuspzr07DjICyZcVqebo81QGe1QWmuORFLz4+ov3Lu46wKSGe
bDWq5JeszpNfcN5GMTYJNYzTBEglszgZupfYb/BYJ8envWfN+5GkR+jSYFSpHG60
lvOC93AFpFtvQzy/KNX/3DYt87IuT6IGT6CFM05A6qYLlFgfFUblzdzUrTKgFIuK
71lJ3XmBrEmiZiUeqNCNBh1okFsFlQiXqK02y+tev0ipVSsehblOBilb6lmwH6fN
Smnpe3LP/YQdoZFjlKqmcFiJ4i7kB9sAAXFiWIJ9litNQhdg2r+Fs76oIJD1w+wL
3mjym86a45o36u+9QDWr9qRXbIP3WU+2pKyZSXXiRrImFN7fEVYvUhJpkh0SsZLj
N8VA4+AJImq1nSAUyMLlSGTsa8FbdFodA9RClqKUeuIe5hi7KHWVmBCGSW66f/cv
deDcOTETgxJArYcF5oO0EXvWamuUA+yvNfKw0y8WAa4/dZFkYhRTbTCPcpxTeWTf
3ghyTw9iizjwx1qS/ZMqoXhcD6drDHmkSWRddTWA1H58Pzw3BK06sdd2tTx8llu9
V+Eh/xPblq0GSEfDdKUmxCapd4uto9y/KdlHxbhCrLw3jo21zVHqD8vIqVHKy3es
0a5eM49UhU4az9OenI0hDK7qoXfnXSMjh1aK0S/knrDdsixXuzzmuS+pOJICiG2y
9db6Otq6PTEnwDZprd1ywsKDi7Oj9YswKT8TDgpdwzqCsnlzL48YNrZcwndgiDC1
waxv+Oo60REvtF6T+t7A2HlMsN9ARVjyMwItWzJxcSCT5PXhjBFIB76b57fBYNPE
QDZ8uDN7YSj1uG+UtkK05JvOz8u+RIcbLhiWGvCj0wGRqqeZSv9eW1Tw3Uyk4YfP
vgTSQo8KrcY62LUjI7amdv60hOYChHaqZh4ut0StWLCuakHsWdBlpBkMSRdxVF0a
mXknSTf0t6AZKnB6TwRbykAZoJA8rBHoZm3340sXpYFTngEvMAGdettOavix4Wtp
DdZ81BXFdffaWx3pRBNVqEVkjhkWn86ELuGLgmRJBUNvefE7CjhEb2oCtJTiMy+u
xi1hMjwkVK3cQnt5+M7VqEeV1jaKpBSyNHYo8ByqH4MkEHt7vbt2r1eFUPtIP+ME
/mvcXbaOQjFK6RoR7coew+6WzZ4JKzEyKR7I52S4qk9o4sxLqsBhCMtTGa6NX4iX
Q8sTBL+ard+l8YAMMmyFb6Q6HrskO+v7c7TMK6zMGeeXKzNzCZ4fjkjNGzajErLa
s8ixhBE5X7C4WDls/QlNx7sScDVrOgozGiY90ln7M8+JSt5SlHlXZKbceNdzCZLB
i8fRu/BadC7s7RgzfVymwY1TvjqqC7e6eL4QiOF4bnLulgR49SjL4Xei6poYpKVo
IXTFZOiFE/tdORZhXeE7vQuY/zSnW8R+foDRSaQs06nW2lK2EBSohIl2oJOGwRQv
JhEpTY7pDuhp4EhMUv35BpWIZRUDbb8k29sDF8yA+ziUBU13r7nrcVU0mkg1IdNO
XujqVA0/5vLAS9tKqBDG3tb/5UcSW6m6wwy35B5QjC/CJOPXvnbu+mzrFyt2foXy
gxEwtofwpoYB+vaQ/5jXln0yclqsBWQmnHqvlTkutrFoIQ94CdFiIPnjQOlO2yp9
Dah2nmOuXecCcb+cKNlm7Sj3rhMcCxuwnhx7AMbMIXDX/GlyBmL9f2Z+AhkxTujQ
2LQFVM6QR350mQi4vb7Z/wJaXXAQZd3+yV6cmqmXCVB6QYCWCMS1awye0OVhLc44
YbxwVN3aA7dQyVSeMDlDg0quEo+uCNtUSwdh8L5rYDi3Ar+fdp10Irq5UO1dnvrs
gZhUYDQZNR/DPEcGTPxTcikk5sZICenrjlhqwse+8E4j4JRFeYy8oMD9ZCuQSyt+
Pb3YuDtQJpcronN/aM+hidEON6C9XmvIL+7LMh3qoBrovyruTym72vFhnonom3di
PA2sjQ9l1CuLN91A8+802S74mVGO6H3zIiTxXAaT/WfFLc/4aQdg3faIaAKT9bTm
1WjabPxnNfey9OyR2FA23Bxgz8z5pPCd0ZL+MOc3mrQAZ8E6/Wk9zePBhQ6zO0JL
au62OI9J9vSTJqkIUEhLwwGPH0KRPrNUuDioqeZcGaCZk2NlVpj5srno3YvXDWEV
mEJaETs7H/ZDYU6VfXyIDE5suP/dD8DrQ5IE7hF95CIzXGidVGOYIFzlXXWEQ7pQ
jmrCfSVrBKIpRh5T0jh/C0isdMEJ/AmRirP4mEZthWGhAKoVGhiYDNUBXL8qqSPt
7QfYrCRQek4Y9CZtYoBlvXWxv8Wo9CcOgokwtUr/TVVmTP2cq9uodGt4gKbLN0Kp
vOA0KWJ8DP+5h2yvBKexvH3hCa4ipNmJFearZlU9nxgFTpN+l4kgu8809pgxmOQR
g2JKaVCCGialHM9R9e8qb0WHYKMTYEPyGpcxlxK8pbHDZonBQQFWp4hvvGV1ZBlq
6Ur0vjoYuCp1/eZ6Rru1mG/nzH15qxNZGBZ4Qj1TC2B8Rn6Uq7H0RlVaTHbeute/
ymt7qr2Szerh2a6HQSzq2jJ31wV0JDZnhVmXPpU7DuXd2fhrtxBiLGhcdQusTrOH
9fGPRx/tVeC7BJgIdbCjv39sI8GAcYHtlzti9dhz7kwqKEYHxNQskSGhbOC0nS3v
bO3mFQW/s6++cpZSZowGVZgcIMU4f3BfpsmBD/MbLUAGh5/zPUBX5i9TlFXunEbf
3GYB6e2+vdmxr4izxwVVPqQMh2nuewMAnblUkSCu+J9YKBBHejPN4XEjMx5M05e8
PUKJYYWzorWk5pMrP5KHCRe5WaGYuU1JMmH+8O5XExDEMDoe/j0wPQrUqaC9IVix
gcmQ+PssRoxdj9CxfVMI1MS+hgHFImAb0paEjytM8PV6jfqTsnaO9qc5+fXg5LWs
NLseAi5CMgvPkADNwBGpmD8ksXGxvNhJlxwOrXebNPkeDxMaMHyB9cCFobDLIeM7
l08JSHb96z7ChI/LaO9AeP/fS0yM5LXtlANzOXnds+BMT4pXVHGGTyjMdnlDfSmj
gWR+rS5KIVvq8PjcTBc8RJCH+939Ye6M21KjMWEvZ/6ensqT/p3JebrAwkD8D3Go
YerbFCUyz09xcFfuRKAzbUy07zBHURoiijcvQAOAd1GP5QSkxlHU8TxgXHWPor0W
stD3rfR22Tg9imBLZvcp9XYq2q3aiaKjwt0FGyQewqnG86Nb+aFmd4Qa0gThmQK7
5xl7fEa0gsliK3vtI+seeiF0hFpghdsdllbFXHHNhwQ7GTeLiQiooHY8fKYnhp00
0nE4aa/aw3te0Wr27QibjyUqGvmHSt3GIA9KkUMxRPx15ZfoUrOPzoMkMv1KHhTv
Z24GE2wOEdyawus8SjiFMfdx25x7DlH3njbWgCSaclT6IXRQEDTpKzxk+qIAU1QA
YQYG0FpD4avLeLNXsohNsN6DM7UwrbKWlCcH+pBrojqOPlhl0DpHQ318yxa6tOxU
FPVCDdZH7D6og9iGNagIV7krU+pRPbe6n4tiUZDK2ZxygKL9KMPm6jfECedXt5J9
VZifhdK+E0iiJ8E9ImMtpfKW7++nsAmQZLEuAcsc5TCkOOt4OLu83WgY047doqgK
qnEM4JiTicyntEas88t1nTfW/AujJg8XWf1RKtWLKD8pCh9BNV7lF/6yUU09liCH
ComTSUnsvup66zGUO8uAxr9hNjzKzWBcbuLsdqqEwTaDlY9NWvP92RFGHI+8xLAs
QENL6tCjmbY9nmT4g/OmhTg1VRFLtEMMvyoHIAT76Yu8S9gpMpM0CS8zJ7lf6peg
b08EQ4lO7moF8JAmf+ZbzONapjTX3Ud3MclDFhPi/yH/kJ1LjzKIB/AUg2PmIpeb
eQmng9NNWh3xesNv16re83aidGwF4ust1GyO2z3ndXhLUuxa5A+RA4p+eZy4em3z
ZJ+ngDFiz7qU7sbBm5kuqcrCFAdHku9/qByN4kIipk9vbUwKfPUW/BVvqLRXuUh3
Q0ssFHu+hkFG1VOjysXFigpRH+2+V7A+g9f+pm9ddnO5fkhZ+MTNtlYDXt7PTEMT
6WkXqyrVmqI3C+0sQeQOHipKFzfLpCcBk2PyIo0FBjs40F0lH6X1j+P8MNan8zOU
FfGcX09u3Uw/CsDONI7j5ZCtsfE3UAeg7iUZZIUCKFclhSpNic0PLA17Gc/smHUO
lg4LpL092nPHXYiVkoCR7vBv6CYWB2WOb+ijqb9n0k6VpzpKsAVfZvWaH2S+shrN
kSHo57W8tBlUA/8Xj7ma52441Ci25N/KAq3UKe0kc5tDFhMJ2vBeT3vt17xXFGD0
b7x8ZXIR2ePjjAz4JhcIvzfXWiGN5y1PwzBdfEh69xOB/NGt/4KTkPqdWt2GKifG
S3s/v/EEZfCAuMvCOTbwpWbHMOLEcvU9au3Zd0GKFFbzsYEi1uMG7i2S3IPVY+uB
AJYvyFcasrPtHq94sm5Zdox3j0nDHo+gtZqOl/SCaJjSGtqKzga+Y41KIG6LrgpG
IoWXEQgR5j00vqcUVa7XrFGKb+kBda1ZOSQKGWdPv+sS5gxwaGqAEpnRC1O7nd+k
kFeWjKjxjTRLQd3RGkAdW56KCThx8td4QZIZQlRX04yvgQCPXPa0pW6OZ7A65AWw
8tw5ZSxh4teft3CtMX+vwP2z3smokNJKor8lZ5MGQ4pJfCWI4ZARuunJBVeYLqMC
xdaTvfeRBgS8Jr0DPVJG8FmBppXFDSMpt5Dog+y6GaAkJcg0HDGX/QNutmr2LCDE
tPgfgfN64Iflxtl6bJkQim3nYrT+5Vmi9eBBud2U19CoBd2vHM1k3d1KISAzCE2j
O/KV1T0uBve9AP35icV4hufYNJ79y1UTd4FRFMoAGYspqWVxfikqCKFUuGbxjvxr
pgEL53Eq/8mHJ6cmEemTzychDSvTQ61pai0KHcYdDkqG9Jk4pDh45o2YXF/Je43m
J6/64eMHNnXesXcMzM2ghYWIFqWEqF6E7Jx4hKSmS+UNpzdmk4M7gzCk7o/kAevZ
IGHN2OIMPF65Ei8PoYUTl0mJytJbhUj1HOl38nA4KqzIgWBHzcw3R2O+RP00Q+Vl
KpPsoxSnNSmG9zz2eZ6icvYhd6Rl4GbVT5FL6/trNOet3VjAEntDdHkAVueEgMGy
vMwrvQ99dJNC/tkSoE//Bi4B2Ldvkp8GNfnibnJy87g1aiG6DosM6tUrtGBQj27C
6r8/WqWxW6vT8Nlv3HhuShCxWSIUNe4NuHVPvkUOzB0ElWWXapuKkTc8TCpzkZHW
3ALBCaWDF6eA3B6pPrLjbZxByyt4QPtGRLDFlTaoWqk7StUdgVXob3KDMq3EM4G7
HwOpiKx3+hDYXKJgJsgymL+0D+/VbrjL+J5ViWRKtkwK8NPA8GlwSpS7DqLVU2B8
98iSHFd1j5ErCN0llAcmGoxZIQe2Pkb0k8agUIEUQdxLGCmBpGohIr3T2XCq3Oy4
AGRLwGJctQ9ySClZeUrHIrjOcH74ZN0QtR0fLpZzdO2Ep4ttxJDiqsXAEAMPQKG+
xRIpr/5aNCq58mr1T2rpCy7U4oGPcg8JzVdL4Ia76d5k9xQWnEppRnYVlqVKxgLf
GE6mlrd9XUEluRd+GHLULGewTXs0122tWalj7FAkrRenPNccCS9cVRaCpmkC1QCs
ekQDE4hm3qFU2dHz7sfNsycx+eKWix8X6AWXHp1y+3nbLzZVLTIOpdw5Np6NE/sl
cW+vwlIuGsoFx1c1vdiW/KcwOgnGda1Ktsz9O1BqN7kiPNLghhdKR3c4CVzyuFWm
1+brnrmxr6XqggPPjnuA8RF9xgeW5NfnNLqEWD4xfEsnn9XJRZZdGeEVM/Hb2W+p
QgEv+oYz0wQHyQFrZVkKnLFP6uJizqmKGDwEVkrkgH/NiKrICG1a0Mn6B5Qe985f
Stcv1ViMiQ0bibCGrHw3qTaoTjcLXzdDEgggZ3/terOrwtO2RKUy5s9KNTXlunNi
h1tIYGefc9r8N99b4iBKu1xs80HD6CBeNn6cp+EwE4vU+XooIOeZFqEAO+asTbFK
2NKl2YVIpxqBmjW7H/3cqWm4/+q77WCpfLWRf/7jNzTkNfj2iGK1kfZPwDlqkzwM
jbg9tLNJAx3v1ONVy+kdPzMHyYzWyMs4gNXRqhKqM00YRVF25QbLRrPjQTyyHYpD
SDWHfXuMRiwQyAgxD9QaMfHUZl4ZM+Xm8t9+u2oGgMeM09K3v+9putFndluviOLN
s1jEr1etIV4itMQOfMjGR4El2QHivYPvf63m90CO4gj5CKYOiCokA/dh56LxzTJP
LafbY2gnQ6b/+TbvVYJ2+LnPiTcGwdlrV1vfZKz/Pu7hrziVBwrSjdXCio4i3bzP
RzQ8hszepLE3oO4isBigaj0utCCE3a7Pn1HqwqBPccQtp4vHkCnyO05ATgOlhDX1
/jKySgyBj74+61o1kqX+OhNpG0Lv8/vHVdbxQWQXjiwepax/yILJhe0gxW2UmgVy
m0FhBGFizP1BQqrDxE6Hm95ssrmXg7Wa4oCZfL6q36WY5l7YgOP2chDMABQpDfC0
Qm96gGtjPSmsPXNkTiDqS7rW5XdiJFBqEmnzdU/qrDrpxdGT66BQKjOSoeBA/NC4
HgvNPcTgaiK4MEBj7JzsLNeodQKmz6gCgd76EOxr19vn36fuF1Va6S54GM5pCws+
dstR6zfC+Y0/1wt2VprEWahXfisQ3/Mn5npCNIj7uwGBMlBc5jIKjMMz0xsLfkJa
4q47lPjwXY8YkFB3eqZ/9UrHSwfJ9UcFtaJ7Qzhdw2jnV4xCLSsB4fkSkCpxA1vJ
ybfqBBs1umQ8cAaHgojtWxY3E291hJeSSvPCPrVpptjJ4uN+7uAHEUS0O7qiwLJR
nXf7kLlFq/4pJu72bPrKMsTsKhjBtotIJ9J1kiwsR6ZVfWkVkOXD+ubXeJUTjeNh
ACZpzJtdYlgo3qTYb/L/lA6i0aZTODhGhjpAh05k72TgMT4OSaJedHJCwn+DxE9p
XwBA3nfGOZUkvcR40bzOMXfk8GFDx6nn/WAJxkQNcAEpm9YPsNcddwiwtWidRs3N
VVPcD7xvH4AqxzyNlHUKgyeS12lYQLrS5J95+zZEMvSj2XkQl788hYyUJeoSP8Na
oZtPv/ToLdMmM66Hj4UdSGFt8W2WUQfffjurlCE1l0Zfb0OneBWudznp3mIt1pno
pUY/iFMmc+eDOaer0thp6VUk9bqMQdb9K3Uylb2Uc2jO9amSMsDj7HO/frxMkU5I
5PTnoKZWn/2gPj13TzznFN2+qMt/Ym49LCGvAeVdjYCvElsh+CjoYjVc8FYCe8eq
IRfYQLyRcrkoj1tQZOWVmFnd61ATBNVC0zhicVfbf5ou9DdE4DcZz5JgMmgXIINs
NvtxilFIGOmFAlRG2/lEA0aMLObQbJM75vWrLRaj90tHATAmTv9OeCQ+XMkEVeaa
pAlRlqpT94QADs82kUr/whsxoOGOVci2HBgy2TOwpHAV9yuKRWKNEC7zM862Cm5y
NbTvvxat3u119HpFMhFTtm1uDTYiFWlkddAbb52wj5Z5viD3kjMfOO2VBGDR3niw
DgChJND5x4WV490n+/cu9V7wgMOxl60q6nFd6vbwao/to2R5rkzMs9Ym4E1aOo4y
1YkbrP9iXEEqwCPSZbj2uqLd0Rb0EetCt1QU1CluAZdA2mDPv6aFuaVgszMMtc9o
XBkG8XprejXtUmmmaGtYnrAoVW28WBc4LQSnsE5o86t9DPkM7yZijwusqD82a4OP
UVs+3+9MGUVZFLH1miakutqsowoc/H7vstp6jCqmhbhrVii01a4yRp8+f1smJXI+
Ot74xWuHDN60rRIDixmdy4saCLnPh+Nf+o3yTivOlV3n/QzFOLU5zwY00u15X8GT
nIsuLuuz0MIJMfgMkS21UuBHRJpq+5RjTkeY36lBftV0Ec6uSewEeSD0gnHUSiCv
c231Cwgm4tDGZkwpnwXzCxQ8GE2nghQ5ysIb5mIU2lFM5Ny1dvShY24/xszBgaia
xK4yAzWr/4cUSH8xtFS5CvGI8O4U3nUZ1FmasiXSzCSnjCPd0wws3QM3mZO9soSQ
blaR1HekkYLNeYbLNVQaZwhOjx++lF1J7sY9loasAmh9BAt2e1sgD7RwKk5b08f+
OyHl34lCtN6rcjUK18wYV3PijuS/AAwtVK2Oq8y9V8P6SFlYmhEDzljwDWFWlnhL
KtX+QYvPR2UBqlYnDhbbX/BUPald17wqGOSaLNiPFLSIiyMBxmwln9xucZiOKI3u
+6O7Rs2jmc2kPgpbjtlV9fr4St0mKm1BSD9QUrAEIuQRMj1h/zZZTy6WlwA096E6
6tWpuG1QMMrenQs4OwzmpFIrdDqDmBLfesnFZkey3UPfUf0aDkb1kfkJti5DWQJ/
d4EOvJ9FhGkDWmFuoxs4OZtQ7QrPDFl/Hy0ZMOaHAKHII3VRnRmWddCJ/WrRG0S7
J6Q9ZklgttxDjRHKU/rO6tq2n6xEGOBvQqwojQrTBskWPsp6CW2yf/AHgPUHe2as
jsPIgJCbFwTj68MrVfeQy/x1DPb6At++sGP+T/C50YUM5Gm+1yTaNczKJsn8jJhh
vcW42U8QrU613OF8awGrfIe6Ar8bthlfJk0znG+IFlkABPHT5gg0c7d67GcZGtYZ
gqC+DUhUSvYzJDRnyFzF1ki4QppJ2aOQSuJh9dMJ/c2zutYWdViH/v1D9qnMf32o
ugCVyoyBwh5n61GW1zZuljc3TSWqFtmUrGJkLQ9+38/KnVrhJhu8A3gkg8Hq4DvN
RRWpmXy+C6DmhLUKT1ebrW9MtXR4vj4ktzJg68+gwqwRqY7Wjm8ixHsD11rRxaz8
UAxy1ChGRU/P29QoPoqc7OcCkSKMdWFdUzYU70m3nnYZWXj6BX7EOEbxC6Akb0vh
+/M/LLhJYK/IhLBDsnkuAYz5ssrgjhcxYhr2QvEgUomYvzyEkRnMl0Hku1szAcRl
2D2huTokcIWVqTJdUuo0Kq73PX+FwX5Q1dqv1HclBLYFUtWq97k7LpeZByIizj3W
jYa777bZTVhx8RXcfhaWLC+KX81XEc/DvgGwuYq/ByUxb49KourL8FpnXkld9ESF
9wwvktCLoV3bTorlXGTYONeOTvO6SzEdLY2mgHUZEBte6jtCJxkvB4K2f510ruQ2
Ht+5uNqe9VDYWSjkHXnqPCe2WODgwnalhx0aK8XYwAv0V5kFzMn+mhimjpIlSY1h
ZPLXOUbolzOUkVxrBp5cXnobI7gVskw1s0VUD8yuHogwKgA+7MygRM3J11AAmOsN
JQ+s/6wY9zd/dRI8JLpgKoZAHtXcdsOTWoMq/xbTE7FWIEFAk71iRnpFBF89s66d
+ATr5WcocD++c+4q9LGO8Xuk07cRKig0Sfe4U5DnSffVF2dURfrMHh8dvcg2atFI
Eh7a73K72Iwh2wF93hL8qIWByiOTZiJL1N6674NrY1EoOTxAfjZ5kxD+Y4GXmWRI
OCIiOBuWKazkrlctkrxaaj7yb4WkXHd9ZHjzQuIDCNOExmETT2cGtR71id38DnWL
0GrI9LjwAUWkW6gObDjJO5ETG+SJLP/F0Gqr+7J0GkkhzauslcXh8OdF73k7FBOW
3wESMamSvUR3QhBjfBDY3O8AtlLGy60vijtRUNBc6lKRvP6JdLKkteMAB9uU92Mq
xIQDUmeMjNcmSCrgrDWYocxypii9DrNo7TIR74tQAj/sbP5f2MWSlc7q9MEBBMqC
fSYlIOfBLow7cyYXt/rSU+NTj00pYHr79s+OL/3hkAnCuVTxoUWXrHECXgMciBcp
yjGXrYaVMAobtt0n5n7EOgLz7XaH57PADJ/i+Zj+GSJeyXGbK4C49XT8kRi4bkbM
v0PJh+u2FMJrS1QuLFq63RCIqnLHBdTToDRpfTR160EqDlnkf5BehnQtOzV7zU9a
lvVZyg5+wIdEMQi7RPIN6EiZzyHLcsQU2FRXyQnlq2Qv3w0I78hVJSGdedoN3DPH
E9nuOSXaYpMf7Ln/ASIeuy+dnPpTRTpshN83ora1Dg03CUMZccHh8k8e5f6jVxWT
/kJNOjQcCf/fKy5jqC/W4319oXOVvMCr3y7gIOUK9KJ5s+cosFGU0hq62WlU2hh7
qvRppco7oXEdlcoheIjGss9BCrO7/oVk4V5+gLEvXktGslvfvSWWitZ6U+l3p5bQ
/I5AvS2/GvAroar4W+n+SJHmvr7qTAW9BRKFWgYAMD/UXz2u9plw0mXRzNYY8JK7
hPpaxxRRPWaZ+0tDxcXmsW6OyKixeIcS2OGVN9nKM/34csH8OeDKy0swXDdxkNgm
hkPWwOp9R41DoccSvp/LmS3PcQj4740CeUk5jtoCnaYhDS4W6tklvoBSxQuhuHob
Ba+C00PkK4SLkVvaooB4PCQxkX31jQrmc5U04kTAzNl4lS9SNpaOe+rqbKRsfYO0
sSoC/wBfNcOwUDY5K/7Bxi0WHeFWNBWAPobSfXh9PpdqkZzHSVdVNxVe39r6AKW2
PjOhmI9KhOHZ5lmb/uBkOQmwkto430SRw3gJUQ1EYeqaivj7vwb04pXkT3Iakf8L
aGajGT6uHYuMV9LBYbtURhNYgXFOJg/QXmmrrYKd32EOa7ZTWrCQU0/25l/mYWpJ
V2FjTmsvuev7dxnl67gFQPEgDnjDFCDOUvf4jfbK9oWV6zLgEW/HXfXpbNaX8xWP
AyNfF6AiE9AIQ4GdLZsu1zfxwgiAHkeHX2GBwNin2jAEh7o4ywy2RAOJOkk3j8B/
ynG8EVxi/N/SMwDKJYd/8HanKM3TfD+obOA1R27nbdpLzarpZDrbNOyB48YwzLfY
OGuO+MccCChOQbAnK1EhOI5t3HeO96w1kw/+SCMP3yEFSI70iIMvDgdL6Vp27Nz6
1b7kpvvwNmnhcaZZ+I06uJPypb8nXjbg8zIrtdpp5QpV/D+FMmvpanDhuXtRhK/E
mzXliBZRq8TlMohdgu4/AMJzgsPXJSCr/5ZhnTE4MmH4JXYYlz68ePNw0MJeAr4o
/bK+8juMAWFtJD1LNlHZ4kdU+YUZXxQqOklskaKcIoXwkoka3PTD0RLP0PTYjtLW
4BzsUTeX/5HWNYB9ZiDa4P2By+dVULhQg+vkKvRE2Ha0jaxQM/PIG436KiUxRh9V
7yAq1fSOp6QwlxQ/MRCnpl8LSZxg68aF7LIzrE4TQhKVAvKR7t04dVFphsWCAvUX
D1hRGMUDOWe0DQoKC3AZt4Vh1nuZ2NNJHZcNO7eVkBKZNnGU3epPyxDFh+wHOYFP
zmhmhnUqIirjrcgsFX6Ug7TVzfN2oSPS+vJSjV5fLdMvJiig5H3Z/q0jDD+5bMDz
Q+sPPvAQIgpNLHXsxB8N7gj0SaDuFELHzSeWZwdMsm6VgI5shCZlAvZDcM0aEDTV
yUcWWlUl4dO4fCQpg+AlQ5sfwLlqIXSUaxlx/ggTj4+cfqts+MZoqm95FNi7m8wu
QXIp+iwNRAMDFrOhozs1kdFG93pZsXeYtYYzOOGBo4wiYHpLH8YT2selAtqNCm9o
S9GzuWT5zm5Yk6yU6xV7+mfarOKs+902gH2/xRCCyR/fDioiUciU4Gq/CUoyd82S
IWzQziAgNyPWEA4OoDCo8YhGs+3FcKhSsbqL2BS8Snu+KOVCvvk6UV2UC2JoaFR0
dX0PZweeqmVvHbuUTu6rxOfkzLFyAY4xKksylo3ph1Ou4Wf5Ed/GUEnnMgnGZ/WF
eY5U+X3MXuhpVzGRxXKsRP9eo4cEyoLOnsiiC3gbL5dHybkKVr764/aFGzeccwIB
+TjuVlM3FhG+bQdZo9rARhhgxdR7cYPrpzzdhSQ6nNaFj30P7BMl8s77RT2Z3uJ0
78xmag8+uveGEM8CPel37NJbIMEpTBay24WsosSqrBzpFFnvxiAnsCyT9QyPa+VN
kD5eIPvEWyvxB+cRC7zCZUzybvNVy2GPrGLj6MncJc5EX+8q8aBHsYBU1vhEDD4Q
pk0mG9zKluL1K//gbcbvEvtYS5yoh+axuZn328bmS0i4V7cuulAESFk5rNLMiD8n
W9jTyQgry2pK2wQsr1AkCw+RjNVNJKkzqOtLQGe1WsMgaYmOA9PFlrvwKSY2HoNJ
UYPWwI44Km3mtEPswmc/mlX9SZDh2rWpT96BaFoL5WUsiAB4rnjtNDa0jOsGQz5U
Qv83+xohoy12PMPC9XWRsW0FPxXmhk7NfnwWs+nXMtsxklAESPg8zKs3j8hsDMQ1
Dc7Wia88ionyEoX3pOZdkV8z72e7XSI3YeS/sy01dyZGesVlTsSWcaC1zJOo9TbA
9Zd9vJFFMFiPELiottwediIj1Y+At0kd2ywLyuy8OtU+63QQVnNZX3Wi6huix811
KstT8tpcZ9yfnZI3pxVFmC7A1k18xm6tV91dQ7gPwCLNF+9ZsfRZqRGDLYHCP6kT
sXV1zJfNQurGgODjkaBRE4pzDs5jhd66idwPcm4eFMDN6wSnWrQgtDKsP4gMZSX6
6y+96LNl6SQ53VlP1CWuISjL0Rka0netkLzguLf5dfCMaK4+o+Mz5REJoPIo5xxq
V01QbSwkwqX5elTOfQ8qISfRpHV39J8TCy8ie2CwbridejnkEViQplFy+79M0qxQ
WEnfl4n9fUnnAI/PEzfYAoRDOO2l14C8k2pDPP0zrQYAOvrsr1DEvgwmVZ2EB0/S
JQFoQou2iNCdFiRBIbvSAz9ZipJnP6LtbeX2JLbDPz/PYGrd6viR3SNSE5HJus2O
VVKMTL7WULQUB7ESJFRGv6oo99DkQyfnxVIaEKsedBsow3259aNDo6N/rOzfs3mZ
GnABcSkuUlOJG+6xAS93R80SnmufWc2q+vgAdjG8s247Q3fZ0FMn7TR0Go8cqrSG
1AGFHxRv+XhFRmCUWcCk8reuNTMek/OdnqefotAUdpWxiMaNTGI8E7/f7Pi1Tw24
lL5InGFBFP5J6LpqutDOBdmRqgh3bbyuNdti3Nq710PhwIJHZkClll4FpEZAB6tI
CLFdY4W4nPCBSfLCSWUBHq+F5sO4kAbu+iKOg4zc8ilYvziV+GOnirqaV0+1bCaI
KqBSEdObonn4cg48Ixp0DxE5SLy0II5xwaFXJhczNBEmJy8beePKBpOGXwG8Q+4W
6eBB3t9wiIrbfqHxS6YUyEYyb9kPqTJXhuuTgRuxWPMvpJd5kSI8pjKR3NG6ebfx
YWBmCs0QrgQ2/9f6ZMPzINljz7xtfz8d/BOJE4DEnJGIVTF+gqHkfBe/RlnU+iIv
Hrh+q4dzDy1ua/hVQ/x9G01fXQt0H56/MIiptRrp2Rz2ySbZbxjzuzjg0HyzfsWi
HptLKiwkYSwvCIWDXyHfUnw8wE/2BQFziMeXUr0T8vqpxoPGztN1htne9Z7r4GMk
MuRcQaIlBIyKG/HBAouw5btvxwPQ2RGElinugTdENwPnXeqqF0CmxTkZ1QuDT3hw
ZB1B5rh3KvJC2wIFORhgRkE3JyZLiU3bvWpNPoHQjZEQ7lSNaiiPA+TyJwwbKPFi
vAFttaMHud6N1f721chv9Gy2vbVhIYS7E7uE/7e+kTKhb8s0OBBvOgvMuvZul9YU
piomyxI1t+YO5IvjF9UwRqBXPikryLMhcad4yp2g+HJh0+kcKB62tauaa9dT//6P
6ZbNfrM19dRyxBsiOUXYPgyFjUlY/1fnlPae6EWXQPMFqAEQXHe6Ktd3A5pqlU7b
46wTu1Fjjs3DBNNWEzVO206RYD6qL+TEz04ZwUVhGyEKWe/ccT8/4uVYRVVMDh8I
y2MCt3BJrcdBhKekGyx0WHfWbS8A0X/fFcKcvSV695KE8OCkgBOl9avwR7YZf1sa
xK5VnZFulTM3jgU48KNqkhtpRA5A52f6tPou9Yswo5YyT9dmWf8qmeHa2YrBngQm
V1/MDH2SG6Xp1vHXQX3x+STmVy7kinA8q64PVhXInKoxrhQqhux1Vv6DxVVrkFbg
IOHVvGKYR+m5qybbehXLQDUBBZBz2GpzrAv5JDyYrMIZd9kB3TP7ySjm58WbpR1h
bFY+h2j40Bk3+E9CI8J6pxzbXpImhs4Zm+IPw79sU5nLKVqTPJChORAV8Gp8fsg3
ITjotGaAtR7oS+WU/Otp+AyEZTgmScwBOPgtda5wepivMKY9Vf1NU+woKvFPeLHd
bJG+B34aPdFBcQ0OiY5I1O4FgKUCu397sDqjPU9NgWqzwL6/oPZIIZexNeW/cvgm
+PmcaHRZ5CXKdBF1QSzfbjxu2LqWTZNFYZi5NR1Z38CxDktKsofzz+Cbe8iPpYE+
rbHORsmI4I5diLJYqvTAlZSN++Pi7rB0IG6MJaehOM9QcDUIY3UQqJk0CkJOowRj
JIvTPrB4htK8C5zDviVhLZYouFM5MPVWv14kwjVnZcJuvXqcTGFRhePoZ4+2wgOc
MIhVu/Pf6KQUADt8lDzGaRrwCN/Iq4fKMEHSRrLGAq7VxvniJaiF/LkJ9aCTiNpn
MXOQIxHg0QFmr1mwK4N5Kp3M0LTgYq1JPyeqAiGhp2GV1oGjfLLy/5mG/TzvkaU/
NG/lrJYnTUFbyuzQstqZWnvS5FLxR66IQQJUdcqS2FE9Mk6odNXjCb3i/GcBOOnd
lcMoZkIwM3p2AH26Ai11DC0qyUQaI2vUjvZ009yvASZj/EOJ/wOtyRUXfp7A4cSH
YIVcysMwYnZtv5IvoOxH8OSJyN5qkMg+ktCrD/9Z/zYI9u33OIYPGVPddxGVxvsT
QPoqV10JqT3u1FEPJx1Qf8XA2n3z89Vr9/ENsRomflGFQCAWhWLleezIJW19DirE
MK/OwmZB0yCmw84CRil5POoJMiR27OEwJDkAY5HcV+Ol11WVRE1lzARKXnp6lWby
k8NunNxAWy/xCyPe/SDK7x9oH4vwN0LlEmEPUAAp2gJzaOgpQpsBUjgZiqF3nTOU
ZW4gPkT7AXU25tPj1+gXCGYyD8W75fCejRcpkY+zF0VFBGtEB3S8QJJnhVgUrSiq
zHDlAUOVsXag3wIR2q0BwT9XLZt3iSTjfTKkX0+A8sZvU8yApIqk/7lF/fhCW+xG
28tgYqjFhA58u8q7arb1n3hj6cOaDfF19xNReIISVYi0uK2DnLlZIWBPKOK9/OR4
vd6ai5imz0f+MK0nPdHzT29vUg0svzxdf3PcXx2tp90MxwTRcju31p/73qgL8XLB
FWlO55SuFeT9sBPz6At41Y7h6DoMn/QB0BpIuK/LYoW0oi6RukD5xf1B6H4Eapai
Lcmqc2r1ETWBx1Wg41v2bMgAyIJ7oYiSl1/9jR0sK1krdPu+Isg15UVdMAIEYJCb
IZZwLAqsdjOFwL0DLdqJnCdhrLFSF9rHScPZxkF/qBzdHUQAsK/YPWLwKU14qgef
l/kFbh2CufBWz22xyGbrmTgmF6JUhvsdPi/R3/tT0cv+xCFIpoV4FG7CbS5/O8x0
GSS9G3vbw28LgBeKbzwYuk7rYlZY05zlaJdNEkbvW4+w3gwcP9pT+v3GXpn/zxUV
axk1NZHEG2BOVcIHK0DDC5BrG0rOLpJNLv6FD/KHjw6Ceke1zUvOCIfJ3jVc6NUj
9Nv8c62qlWz5Yd+/kxBSbkIRzACIas4DNTh/b+r19uEPr2xrR3dHVk5Ubh6bAhHJ
lzKvRTonj9aod+8hSu3KgPRzaFBFcQbjgM96cOO4poJ8HTbvfATuzh3DomyP+hEq
h5lNxDAxxP050gMBC9Ys7zaDHhsxfrtku+7rdtLaZ+w1SnRCrYrCAid6z0UN3LN5
YmCRyUsruwHq4EiyHUMdTrLDSe1DotYLGQU/hjz99UHJVtCfSwvh2yR+X4+2wwIA
Dntyb4LiI5SxbqUal3D4V5AkzVzivKrPKo7LhMPi70SgLYO+iXhkbGM+jeY1YG6+
KF0PQr9g5nRJcHID7A0eR9IjZ0przXtdK10gq0eFym11FhLHyjDzCmRd6/ECAGIM
XfPalBhTl87gjyGNdPN9znm8DREeOOlr9kzSRvVARLW7M8LPlloUAxqksYkZHSXi
3+RdopInLyeVsNclYEb4SkFVrQwT9zXKmsACOvWGLc/Sw2LQ8eV3Pa/6PN2xeUVo
eTeEqbfkjyvzWfp5yu0rMnjq2Q6Lup+S3QErZns3Fgin97IF7N1RnrSJAdGaHmta
QM4qZPX/G05P5yNbSiA975lw5clRGrVAx+CbxLwPCFE+I1sW8csg1sGAu3pM7Ld4
VRtP4il8csyjXOjN2wHMClIxMN4rHaevrqmr+jZyNA8p0PscNC8JzUVm2Q9tbvxP
Mf8cVhxd4xmvfcWBRLGFvc4RsQmoGs2fd5SpRcF+CKhXDU0ZGdFEtm2nsb5iG/24
ez8f5mjYkX49gq2wim6iW6SqWf3Xt1FCg7/HwVtYsky+JQmkUOhDdTUt04GKyOdm
8X0tZ6iq3CQOs4zX77Z+arUY0gytqWdYYkdcTuedCHpVildJJEWrIKGZPfMmOUVF
eZrl9ZZ7186fwtoYIpm2yEW2CeuJYCx+MfjbFXSFv38oilKC3CEqCvJX4oIP28d9
zwZHDheXRnF6XwvXvXnelB93OxOmKdRHxnnZcPChez9ZqDOcF0BnQxqNsCgTMIhx
V3XnGd91sYiRoRMHBbgm0uD1CxXAOLC2iAkYNK1tRe1tpD/I4RfYfBzMTDAseORQ
Yl4l3VqmqiAL0fJnErRJO0CinlHzJ3hy6p+N68Iw06NDYHt7tdAqxAEAis8MvLo0
ct2LC2QrHq60mcajvi3QOtHbdDjEq+ntJTUWKBsA5+RhMbzxIj3KVrHj2GPgeTrF
Q30T9+pES8r+/f+p1BpyfamH6ZWuvq1ozyx49VNup29Cgiqeenoop2IrtM8NTiEt
y16DfPQnZ7NqyG0IKlSoUfiWihxkoR4fwAzLmk/LiV/aGZS2ylGrqFRGORrOcXnk
8IK9OK7g+ElVrg/vvfuF4QXl6nk+CpBB3GSkC1lLub6s2wAdFXSjw5tr5kJ8iLm1
+owqKSkHOZa0gvMqJxhUJP03UUy9K9O8mnpsMJtctff3g9b+IpcR9zJ9m6YLSy2z
hM/rzUp9yspcsQzYj+GYYP/zLLPgmwd9DQPramHDqF1gwIZRuMqdkPajGnWViKh9
8MGVMTn3GmuOqTscAP01luARW+xutBf65LTeNfKooLEDU4ByCI2Zc6VjJSmbtYXf
4ipTWkX3z7GrMgLF7K7iA51OiAQ0ge6xBarP3D3TcjrnJ5ntWnC3Hct3jxBkZPQU
oYc4PG2uH24Jvb+XwrjHdEyVWIFgdB18E8k0udgUNJ9JuPkkzZDX4syiQhgwnjXm
VcUX74Kvs3mkCsOXgGDZdq3qdTg67lKeXxfV2CkAZJA+PglNjVlw9j7bs536WyTA
QJCOqJCOuHQZ0Ep5ptlrkr8jVW6os64AguDsArRcg0jvFDWiQv9OBSQXnuLgwSOW
PD0KznwyKC9QKPzBRPFZquyxl8K20NUSIja8xEoVbr0bpJmBz/2nqJd2EDti9aO2
C15Bn0CsJvFOSjBM1Ojjqs44G2hicNGlv6zoafXlOEhcLz+b1Nk7W/TPjV2+CsMS
lNhZuTPlFmOeeddzAbo1rAjmv4mkBW/Pcqw0qBECWTsYD7li6QoBShwupzooNFq2
20BkSatva0w2u8IuS9D37HkBc9+YfVw/k9XALI+nO5htWjRjuS7zbvWpxF/uCDUE
eam9KCXAfa1Q0bD1Wmk0kqCdWWvNQgtOTkt25bGZm/CL1VVg6MK17GnvH/DjA7tF
t7fHrIoe9GbYjN8t3Wx/yecgOLVh1WrT6tfTUGtoxaGfGjoJjlYoteN6F6j2kblK
DR0EYFOwD/2YaWOxpU72fD8toVEEE7nbgtt/92hRuJIusl4RRs6jpUU3i9v9qdg6
OLwfLg59yeYqpu1MeAe5DfItaxFHW4LhZ6UgeshofWTmSqKRHqxJ9kbtEPFePQed
sILt/SAzChqWkhVTLxw8oksSgmpi3NKFHT6u/rT/kzNqxur6ylJhUzqKVclsAZ6/
HC9dv8Wzx8Ps9JO5uEkWFM4akUeoNSmQaoZwmrenvx17ltkw68Df2ZDATMGVrf0Z
qMBZVTYGpASlZcEDyFR74rry7sqpSS4F2GloUtT4MoZulYnD9zxQAS2VYduBdHFN
KWL6iQj/sf2zX+gRy5oq22MSLta1R7OfmDY80oo7WFnNxyoI3Lgjqw3m6AFkn7d2
00z5RRf489QrLV0IcPU4LY2tCGUJDZfuaQaLhhFnfKNrfXcHlmDJy8X9YVXgAbb6
RzmcPVufIqgsjeBESH6jYz2cQGH6kQQIpN+5jTTA08j9OP7nmA4yWQKyFu21jfg/
rbEr2ZH4vnYXJnMxXbeIpM4Cg91EEMtz11AucFSs/OYnJ8eRPoi6moJyxbX7p7y+
BhZfyhPxhIMz9SjRKcoMlHwp9eBQbBfTEp3MQZ/XNjAy7V4hsnjA+aXzhwDNH/4D
0VudbWTCLPa7vfFfv55ma9KYE1Homnr9h6KNbW+4VTtqMirE7o2PNy7eBl36zDx8
SX54CTK2cfHuEbCRtFFuBuHstN/jwf/OjVaJR82H8rjNgTXpj9hORBayiqg5EmrL
f5VN7Cp0P0L8GOadRhTTu38aqSWX1+pujEQpTUI5O08vym3L/HGjnkCBpejCgOv8
Z5KmjOMRgeJpkzotPpjrQKa3c78CmfmzhXJUSFSpUQ8c7VO290wiDeu07/n+PQNc
n0HiEGhSuOtfYhcL7tA/7rJJedRDHZIf4xbMsGVHmYBDHT0bECxdsVGxguTvGz/v
mah36v+K/d4NuwfoptsQfBuSW3E2Zwgt4ezxSkeFC4beF2K47qIOKHSjLj0S3GKS
2wzzMYatfVGbPrNTJDA2clNITQLCPmyQn+b8FT6336NBrwh/v+E5CW49t9hA6E7L
oS7KImBYMObaYNnui21wMbcyjaePOuZ7Vf2w44Ha8qfHdqnIfJ6Rzm/T2aNCg/7x
jRs9GEFMzvDLqnggpVYASmlaURLeEh0ItNyFlJLIes70Wch4v4ww13yK0GKcJrQd
OiXNFroJgK3go4o/Jy6McQ==
--pragma protect end_data_block
--pragma protect digest_block
+nlgwtOYhDO6+n058ZyAVkB00RY=
--pragma protect end_digest_block
--pragma protect end_protected
