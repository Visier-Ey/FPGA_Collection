��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���d�v����0�i�=\��A��?��� (��1_B�f�	�Ѻ+|n��y��Q4�]�aY�����*2�y%����>��������K������ �
�D��z�z��C�y�B����
_�U��hkF<�~x�ܕ�c����������E��hA<�}/B�2�4|p(��oy�=��[�}+T�:"P�J�A:<N�gIE���@G�qt�?���o��]n�=��.J	y-�]���F`����?"��;�q'�VST����C����V	�����]��mn�1{j�(�w��#t��M���D7[�^��2e�9�
p�{v%�w���r>�Kfn���yL��e�jL�����*�N9�mV�	%�&�j U�qN�lL�ft�b��FmTs�yp.�p���&��Y z|�Dޅ��/Cq=O-��;�w����hE���]�p Q]���R֮Ĳ'?M�U�Vz�6Jc+�oݾ�R�E�â��w�9�����u^�%�A����|�1��5��2ТA��_r7�p��p>��p�T�=Y'G�����4����m�܂�y�':A��_Q�>�T��I��Ȝ����w���Q�|f!~��CJ5^�+���hX-艏q�Ys!^X�gHtHE��υ�)!,�4����c;���v�D�I�>qLo�	����U��v�.�C@Tl��	j��;��aJ����"J#�w�n�,���o���-t�Fj����~���r������<��z}�J�� �|�v�z���J�NU��Uϯ�NGN����p2�f��]c�'�r�cdp����K���$�up �i�Z�G�r���xW7�tܥ�>���4�@'�02X��X�*tUfӑX�WH�D_Ţ�w�=-�-F)Շ�Z.9i��)�� �����̳#�|TN۟�FH�Fn�} -��F��}N��P���0�(���wY�:;E�2��V+�cL̴��_,��I� +-�=�o��#��$4=��*����BJ���jp�e�+�BV��CʍV$p"��2��������T��d��ݰꜛ�/L	�:|������{������3/iE	�z�5���xJ�&M���^R,??O���R.%��5�ONm�vF��ԧ{����$6��f�5	e�EH+otV����?�J��Y��i4���v@��ZS�� ���޸��i�L91�s*���R���շ�f��A'
��SP��-�J<��g�n=a�ވR´u���OD��\��� V΀�Q��?Q��}����/<��V�W:��_�n�3Z�uY��GF��w& f1@v�9���lK`�wl3�
�m3԰,y`f����@�����m,`~���OF��mܫ���ᶃ���4��� iK-��l����sh��/p�^�M�f����%�3+92P9�'�#�x�� p�w���J�4}�����P�\������|Uc���zq���'_9��q���4n�O}�;�~�=��8�F��fxnv=o�vgXc
��׮hdX�w��I�K�$���K��������q؊n�P��� 3_]�¥�
ֲfk�_a�z��ʇ*<4���Ivp�d��oE���HO*V�t0C"�YF�a���,X�2"��A�1Q�@\�%��J�J�p�Eb�X�G'7r6�����>�m���WcԴ4�����WQ/�>�����V&�[R�h��C�Y�T?��k��rc�~sg�F����;�^��N�X�E+7Y�\-�
�vv���I��0��+�� hc�nc֟7[Y�|���׽�
�ԠU�yޠ O�n݉ǅԂ\���F���԰^*���ڎ&(��7��g�V�ۗ�,��W]S<e�E���l��?�[F�C0��x�'5�޸������uN��{*���gay*��j�q1KU�[���2�sS��t�}��zᗒ��8�	tK�Z��Md�<2ͥ�����h�/�[��EAø8ة4����m�C�Ws$_��v��� �Q�0��M�Ew���J
@`��u�>�avZ�5L�q����(:=��B��}9�og6aS�*�V������]�����.�N{����8˺%f��Y@Ղ�m���U-eI�!�G�������B�4K��G~ˬ����e������x<�m��]���?�n�0v��m8�I�E�����O9���$'��(M��8��s�� "��Y���[i  �>2���.�i`��#$��"G��@���S�ې	�Z{{���/Ǽ)x��c8���nِq����9�Lsr5�W�Z&���a�4X��Ai�G`U})4����q�>o��W������ �q��@Z'�EN	3��}o��@����j����1���nK�7����{�2�[~g���~�f�������wa Á��TuK=8<�DE3:�|�t9��WDyߵ�d_U�h����%k����x&t#��0�9�{�C���=J�-!�u���?�����������qP)�?K��.�ݯ���p�,�\Lc��L�
��\�X+����D�
s�z�2l�*�4���o��rVb;C�X����sw��/��vG�"e��������%��4;�t�av��N�m@zV�ߐc�����kqw1gK���w�������/�­�!R��cL�mw�A����c<�'Vu%,�!�$?�T�L��G�6��|�i������Z��ʦ��e��u�蝛�׭�@J��fn��F	�c6	�Y*֒���a�-�?����a:撣N�._]�*�O�kK],Zm;���*��\%�H~Dn˔9�$���
�q׌��QX��VH�LE�d�@�4�h$حiaR�� b9��d�_-��MB9�N�H����P��H�.�E�O���ؘ*6�Y�� ��VQ�o�֏���qo�ߒ�B�)N��[�vv�5Y'���_M�.^W��ܹ,z�ga����Hb�J��A�"�}Ll�$����bJ�r`� R�b���Wgd;�B AYWv
&l��|8�+a��%-��}��eDhG�kDd`x3â��t���d ��+������e�3C<2;�l]���%}�����!l�
f�N�%�ȿ/b�bT�ye|��n.^ߨY�-@|�s{Ko*ۊ���I��mHXd��Zp �)7y��L���O�Cg;Gް�(V�Jn�8�+���Z�y����N���&�A3��G�TUY�)S^��<���Ũ���q~f	؎/��<��ғpg�7pv����$vqo�M���B����xW�y����u���8� �P?A�Z=p{�+�m�q���K=�����?���>D]b1�t��R$��=���]�U�b�C�<����j���rwf��[��jz��e�m��37��2��4�������Y�nhK-����o޲�麸���fTU#�6*w%.�&��� Ɋ��"m��
�y���ʟ.O��6��˯:ې -�\y`p�R�������a������3HW��j�B^a~�I�N���Q�`�*1Ti[4n�V�J�'~�Лa�������?	��Z�B�c!��x�Ѥ"$}��{WY��cv�M�9ž׾�M�&H���z����(����V1�#�[�NL�e<��Q}�}zU@�(_&ʘ�?�� G�Sf^�3"�+F�V�
�a�{r�So�&h���M�E����r�2��8�YgN�ؑ߫�����T����*.���v�{I#�0f+l`BT���W��&���kF�Û��fiH�;�k�֪�H��ɼ���$��������	)^�{<�_��C�Q/ ��ys3�n��m�5	?�3͖5�f�����TX�9j*�ɋY��;9���u^���hl�:/��ӌIX�:�D�ʰ{���_�NR+��_��֬Yް�v��B'���*H](�Pف~�d����^��8��	�0b�S�*w=�۶�q
�Q����ݕ�/�/a�V�����y��3\\��	���~]���L`�p��g!4V�^Y�/A�a��z�%�ޗ����Sr��9��b��g�	��|�g5�_�I[��N̞EwFq7��!��h����,NK�K<c��
)G
�FܐZl+S�1v��I����Z��\-�]�Ͷ��������Ogt$U�;�,�Y�� �'6F�kRM>�5^���\o\��â�$Ω«��rO�BDCJ�轨�<"��Jo�7Y����n�`M���y}_��>�#?�V�4*�]�("���beyq�f?�Іoɩ}K�ܒX��tO��Cm�$8�Y�^9l���J�Ա��F��B�]o�����M�m�{�p�Ɨ��?.�6j\}�
^���}qF����Xz�+��K��v�ySh��߈�'=�Į�O�pA1��/8��@K��.����?�:�bX�	����x[�c_q�1y
L҆K�7myʴ�����#��0��Z�9����1�BΘD4��a
!��g/�]���V9w_�1f�2��ޑ��pN (ay7�� jp(@ְS��/��j�z��8߫l1���IS���g��N��yp�:�"6vt��b�ϲ��� "\'!E�8j�`g��{⻮���P%�ͨW*�����e�>R�z?{�6�� nOR"�[��F�QuYy,'Ba�>y���W�P{�	m�a�1��)Y7��S�&�)�(R�4���6v7,�_^�sbe��g-���YڢJIi�- �Di�4����0{{�1/��m��4��Y8�0b�]Ѳ����c�8J�p��9�O�8�����TGUQT��������]'�
Ǵ���td0��F�q�ɾ�gy��)���N�ٚ/uۻD���S,�*��^t2�\���wM�=��v	�������~V�y�����H�V���1�.x�TӷO��C�y�7��-�(*=���a]c	�\3�ut��Q�gv�.�\����u@��ɩtN��.��6TM�8�	>H�t~M�(d�5��D��0<c�z���O���7h+L���0o�"o�R��?P���ؙ�HUX�uU�S�y��]��׾���v��d���U���J*<�bo��g����ُofx���O{LZ�34���@�`P'ۇ��x�7�Bj�t�0}mk�a�#��Kc?�O�Đ��-���^;�W;���4�U�6H� �c��,W�%��
�G�Ng}��+�E��ʢ�$����6H�2ޕ%p�h�^p�	�(��m��'�%���͓B{KP�u���p�pV^�����A��R�S�멹���u>*>�� �ni�;�S�W��Ϗꭅ�Ӝpd�y����|PA�5!O4 h!�(�u�t��|I�<� �z�����\�`�x�8��Ń����k^ /X�����Ւ��8�~�8���nF�w ��E�:��+G$�B�?ԋշξP�]�"����.�� \ OQ�z�혂6���ݏ�����\(�PBOR_�0��}1}8��,���gI�v+��)����)ejQ�������U��'i
P��m�7;�j���[Ć���+�9#/�7
-��%��u�/�\鶞2�
�e�n���e@+4yQ��2?��==���O|�*�����	2=�$���7Ix�����.�u�Sa���ȁ���m��82 �K/�5���?𜡣��QD�ͯ������;�s��N�ƤӘU���(%a0�ޯ�o�x����F;:x3hw��鴩�S΀_���#�ڂv0�"4�U�(�	�ү������	[� ��p�ؘ�>�pt�"��V��33g���W��O������t
�}�4y y�ysj���X�8.:a�A�ؗ�՘^�I��*���]0L�c+������b���0Ф�EK1��ی�#�E��]�N������"6�Ů�D=�m��=?����zS��i�Q��=�t���2�:�fH�n�@|	����x���f��9�u�mvO��h�dV��i��&��u�N�?}��?�6�
�x��*&7{V���*`#����lobR.j�H�)�ݠB���dҏKG",�[��"���71� �8#��8${��o���s�%^��4L��E�af9��O��i�!oi�:կ�/��5��c�T�О�h�~����#\ [���k������[�aDY�����y�٥�U񧁔Tߤ�>��	����a*�
�M���mp�G�3ҽn������:Y���HVv�K[>-m����� `�$�2�/t���on�ic�q��%HL'�k7.u�({V��xL%�6��X�o��H�2N���_�0��Y���ߒ�5���W���q�p1q>Իo����$n3��s�A�7�C��2�bJس�K��uJ��l/S,ԉ=C�ߛЊ{��'��MAb9Z�ߥl����n:�0"ʘ�p���Q���r�/u[I�cIצͤ#x��U�.�N�"��=B����:��_��������I����w��������]�?_pJȘ>��GC��T��Ȼ@ L~�*L����Kd[��G���&_1P\��Iel,�lz���hב��^-��{�7�"��|T&��o�s�>�g�+��+v0�N=��t�������K�[2%���K=�z�@GڃO��v['���0$����d3D_�/�q���O��ݓ��X����/�*�c���@�2J�Yh�c�7اȠv�hyv+���J��:��9u[� �Jdn��8{c�6Htx���ogv��>z�{)�lZM)�Y�!
 <��qw
�$���%D�#�6=�Y�N��c��j8�����~
d�pr	Y3._����%;C0��/�弎�����C��6��������q-]?,g�TK"�4��Z�e�Cש����t���-�B.��_B�s4g����!��1e�,���a�!�v�3/ h_�,.n��EcZD;14�JXT�����qtN��e!��i��z+S�Ç�����u�7W~��E˖+�ȋ����ʳ��Ѩ�v��vţ�wK�j��4���I�O��(�o�>�FJ�"��P�.�e��߁��j�̶���+7�P�����&�؃�!�(��=a|�C�/�,����W�n�V\�yj<Dg窤1U���wN�9i��B�����f"'�?��`�,�����{��A�����)��W6�k�r}rzW��W)(2���l��h���&��wG %�j�y��v�~�EL�I����Y�2�����Sޠ�q�4�e��g2��:�r�Ou���?�W�1rHK'R��t��D�����d�;���m8�	���$�Hy�Miӎ쐐���?�V�V�:[���X{�J�R������jo�"�M�=!ە��!��|Ʒb���#��^�;�
��9^`�r�v�}*�'�0�Zͦ7�K�!��N2y&W�V7���歊?E�������DcΓ@m��r��S&Yz}���=�YH��<_�1U��}��DZ�HL��0�%μ[*����L
�<N\�L=�����D-�)�Ԡ�+kO��F�u�-���n�"�Ǒ�k�[��0R��&�M������'�T��t>`J�%?�����$�/#��դ)��HG�Ŵ��n�p��P_�q��+j�ӆM���?6���СE������8槻�V;v�< �+�$��YN;g���@�����J$�<����܁��X{�IO@�^z������m�!��e��^j��W�mԛOH��[��2�d�P�&�v �N�r�v �[�л�$"(�q8ͯފ��|$���b�	��i}��w����Q���)��+�<ھ�������'r\v��T#��(��#5�ê_	 p��X<H3M�UaI��^����@���A�4)�"h��3�gi���? �y�^+�Y31���E���9�>��4�����w�!�����϶������!7Nh@g�Y���q&�<�P-�4���,}E�S��8b���H��@������]/>��H�Ƴ>���b����I�0[X���U�� 5L��3�4I�� z���+V�4�^��VXS�T0@�k���m�B��%�d���\�e��l�Nvfo��R��E8a���©�ʇ��z䁕�����ɵ �f��i��E���p����)[f��I�lG��� z-�I&�f]���
�J�ʡ������PdޮHU*����L p�qI�q�E���n�ҿ{ݼ�.��Aq�
ܲ{������(#	��Oqj�@�@�n�e1���G~��+�&�٢�G���穹u��TA���"�#߾`�H&;}�����-D���-��ho�d��Jb+ޚDmzbm+�A	WD�/37����9w��#D>e:������({�+�^�P�~�Gs5���(;E��}p��@