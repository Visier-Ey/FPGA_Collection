-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
--pragma protect begin_protected
--pragma protect encrypt_agent="NCPROTECT"
--pragma protect encrypt_agent_info="Encrypted using API"
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
--pragma protect key_method=RSA
--pragma protect key_block
bcDS0lOCXlDuYSBwN3Y+zsHkjgRAz87zvs6soJHGicsZ88KybG3OKOAaqWsBhKsI
V6b+SwKfgu6OJdMqpUw2eDDgcVI2qUmDBtoz1lTLi80FcBl7YKOUxyvuZrbMRV4E
Okdyu4C25T3hBej9znrrqK+ZFt1/uFu+gHbzEv3qL3LM6sXcJ6jR019IfyZo7rYl
8halskqUavAlYtoCoM7jElR6KMMQAvoi5riaASoxFE4VLMhaoLviL4s+af5Expub
bAJzKsg1RaSngPv9ClxL+eVvAq4RISev5Gv6dTxMtVup1AyVbvlxiqx49r/JTc+G
U8wFtkB/qCDEXqopXOmRQg==
--pragma protect end_key_block
--pragma protect digest_block
NLTPQ3VZDgGt0HZA78vdIFy2Y6c=
--pragma protect end_digest_block
--pragma protect data_block
KC9Q0SvGz7CDFrwaYx+/R8pHnsbkVi0BjOac3u62t5O0nwcU34bxKqVDFkMC9GGG
uoRsKI4ODHmSOfU4wICn6AxY6jYsvfWUwoA61mckoL+arUuw9MiNNKltKQVGALvm
Rrb8K1iNpx12HVsfBuaXL2u99/iE8zW3n00FNMSg4fd/txyW692DhuhKgNWiQwj5
XYPPOmyX6L70YbpjvtOJySEQJPrzYbrlHlQlXEwCMKaXW7sLkNc1mgE4xREe/GCR
lwt3/kLFD3GNP7Tyy5MXPUuzhuY5b5gC91V8+frMOj0zqrxjS0HxZf3gpwYwQFCZ
1YXfLEZniyFA8NkdnJeMW8LOz9B1e8JWfueyR5uTuYHmsIPvxG9yvcFOC9W8juMW
R9+PxnEfw9oiH49ezihUZHMUGjTcyq62WQKfoVcnc46ZSoV1wnlgzrRo8nJDs1io
HGdYuzlcIwwQyMQblc5AMDJmU+d6KQaiBkRXPSaYnxiheXlgAMxe9SQ4u33y6uER
uBv5sksShTJv0YtN26lODpCxu81buF6YtslnmQqT7f7Rq39pUQzqih44EJwkVFp1
kXcwmOU37qSgtV54JHArhnaFTJJsg5lgky8lmHR4HKyX0NvlSja2uIYQ0ZdmZb++
04e5p/9czoiNK69xTTvHjkiQAEXDuL7SuhVK5v+S+spbQP5wgKdxsaJK5j0h8Gue
euq5UOAZCrrkuoWCZHZLZQ3s2NYwHHie11VoVOVZNlMqubPK8462Nw8CgCSWxszf
XZTXcpWCPx2grxNrufgfD16u+NTargxtywR3ObraX1ZkM3eFds8E+6qJkHrON7FE
zj+PPNmUXnBxhCeqbkQ7whXV6uS2q1MHjNUl698lDSVT9wRBgO6xMS6npXArfaDJ
7pIPWKtnwrPwnmJRmA1HxRHqMquW9C4l/LQl1YwrMVU1pqIQT5+oSBdhNCklfZR8
jNWCMcSkkMuPhC9Bn87snz+jDglHGeJjTX9RuwA5uz64+VekykwvPf7JhNlgsX/s
6oPseN67SbyffQNFKlg9rcNoXIGCGBGlmAR24L45Cd/HSTysf9Uz+bA5IHCQOUPw
nEuPGLCLrp1VJSSqlU/31BfSPeG9mkl4wmeifC0RrecLJdRxM6KIXn/Xr04DrzCg
9WmVjSfNM6Vp0IHE10DAY9A6AWsblG3jubA6jAMjcWStPajdma2F+ih7aT56+l2b
W8Aua6pJEOH9NHrADnigqSX10i6omp6oDAqfxDy22/0Pstp0IsfF8P3CWtI0S6bU
KLSFNxUkb4fF8pFJYV/GSFyMtyxOAUr1viV05IMwmxMJWGKuXGik1IezobeXyeXw
ttazkCSmaG3aFw+0eJ1dsLaquYpLhpWMPzEhIwFfQ2pcMDtZMG6Mf2IDNCez0R/V
LoFwK/bir8Xmh/SlOVDuIaL1tCyFOt7IsZRUwjtSbRRfvHDmLccevdaFL+JXP0Js
15rN5mFaVoWTvtqicRS8vBj1ACVmF+bUVxJxxxfm6UtNOUM3VsQujzXD25beTNWN
Ahu6pqEGAm1kiqfCnfZSFJh8TIc6QFF68G/b6rWF9zrhC/V4M00fhe2z5PtpMzJ7
/DUk4vo/8nfyBz1escVWMHC5j2rtsk5GHVpNuz1guIcFwot1tEVjgeU3FhrHy/p/
g309Bqu7iWVf3lT2TYbpRpe8fB8vlz6v4QQBoGTXFQHm2nCSkNjlP0/eWZ6R6XFB
+sbruFX5QnHSXC0M5coNdOpUrxm6bIEAkp9watMjGnLrzXWIncVnBj+7Re6As4Rt
cMU3qnRKJgNvWby+YegxBwVc7pWz61XDvHgroBN/42hhRx9JhKMd2N9ElDjFNjX5
0Xl4zAwH13b/r6N/VPew/lwy/2KVtbVX/EvSzNZj8l9kbHJEyntGBBWRU+QYVzRC
Q8ewtTlVfenRflT57mF+Oiqi45eAw0I7Rtrhhzbs8xkwoF07eJM6ZMlvcI9dPtfM
tyvQtckXSTu8Cfj4vIqDl/OBQdCrOY2FsPqMVhoFdKpMet7naw8ltZ3Te62VCoiO
0mJ25LMNbZ+4QkvnhU1ctJnOIaxLLpFEAeZ+3bswiNj9e4RXfY578h0lHbDVkueU
fSCIvp+XwyabnLNkhlxiu8Fi5/NmcZqwcjQ6k6tfzHyhC9/7oyPQHfaSWHPmMnzg
Ibrrl70CM57owUwEdc/B0zHr51Ibck7YwO7TbR+n0AYJCCrY0z7ftweEhRMyeVtR
/f/1CY/e79vbV1MWVmmDhLsWw13V/W2H9K6ZHbicIFz05RGh5kPFreRKy9AD7QNk
tpJ+xAYMjQ/qcdTb0RTdKbAe/jSa/T4TpydGVVKZ7ZCeBpscLuM02zEPisCMgZjw
qrlsrhyZSXmB2srJJP+tjeaIZuQfxV8pMGGeZ5teQ2XSVVjyiZ5xJZfJZ0ASdfRj
5DX/cdLHiDaG/egPz3qHlFpteeXQoYlkZ0xv+bx53PUZrigVPX9/0+V0BN0Z1LRu
L0+A7U/10hGU0U1rDCVMbntbPwy5VZ830tuk3xfdQ4/7YWzRGyVFjr0lN+kIWeFh
h1GSLSIiBm7ABABksd874Xqvc545M7BWZn1WPVgNNTwI6v68b5fWOpx21hvmn3VU
xO9OqKYh8tYv3spLn8lzMUMWRS/e8P5l0KdOlf1mcu89dyMFtAFPopNiFKoAyAdF
NnClF4M2IDS5gdLiUx9i6thQ5m84LmETnxwBs8bpvsN7tOf0jaaP283tvryjEL3+
c0bL0sUmc/2QVHbw5SF0tLxVo2UDghSTjPxS+pQt/Zt9VNXvM8c3mdu9i9usFNE6
LtEij2y+Lq7pti33XDiNMJtAfLUKoI2MsKQHS929dQo4Jhkk1kiJs+Rf6cnZZ90h
NrBEUl1zVXnMEJsVoNoMLMGHELxV2p8bkAs5JanxiZmG4S7Su0Z/aqRRxjU5Xxar
DvgmH9cXNO4ht88SVB4W25LmiRjnuwUam1nRzN75NOkhOWOJMHdNoO/iNrKUXbIl
3ghFWkNr6MqwJYq68yG/hGftRoxyjsWLIRVNtIQoweoiMZU7sMjDEN9beAgetOmc
Ro7i0z4NW94v9bidrR+MlZI3U84DOWCmPjiVHmr3MauB7AB8aAhlxIIEFsFG5f62
jocEveCCFesvtWpS4e9cTzQ7M6obZHgPqOjag2TwhCETD+x/mY/IrdX+kEbU/eFs
mdVBvOg0rAxZ4N+Tq1ec9qJqkT/xx9J6JTSbp4vSibz3hmZWG9MA/v/CdjEC2q8u
Ry+3q+0m4foxxEZ7qh1T0on/cnsrdlDh+ryenHdZBeuZhica0Zr1e2KEhnkkFAvc
WusJWOue/ksN1+ZVrfQ0+Qggsm2vfAdYhzSI8oNgAt7B1v3H8tCOBGXTUq/pnhIk
P2mfjVFcUvmw0h6sBJ8RaWgmA8Pa5F/fR9PJ0hSUaP5zxcukXD0lPEZpD9HMmVRe
jQFMipzm/O0yoeCqPSHPzpJm772OivgbeAvesiVuE+XwBAcIbdgzQHiFBRIj9R7u
FrtRxfPlD4J5c1ly7APsoZ6Uo1/YzCyPRz0q5UHnbr8+q2dIr44+xa/iAcv86gfU
/B4NOAkzV5RE+mXUVHnmQYPkUpKQ/GMEP5IkiCdCMlwXoj9SoByGEmBz2f3tQwjK
i4/rTtQQnApchVZ9OVOY+OKORWRYi+umC6TBE9VW2pSM6DHKueKeoTFh/dh7JauE
2+oC0i1yGFUEtHR40skPM7sUeWHvwrlXvzbDXtzpe90SP1Ubi2MWm/2vs8PiR8rr
NVtjT+x7P6uAutQC88KMAEsofWWHK8+r1sy1n6/5R6NXTpfjaCuIRGNC47xh2nDA
S7np80oKbpOd/p6BYup0DKPyn3ubPKKSLLDgEJIDReHBSgv2ti5GLxm/Cx7VmPPO
GZs+5UzIacvMCg1Id6wY+XYnM2oYJSDG6ISTr2yWoNdzxElEZgF13u/q0o4PFN1a
2yyjMFAzO0/mzSrU5j5WmAUCL8mCU8XHyT6yzBrIEk3YPDOXMbuk6jPeAkA9tOOY
qkh6rH6z0eMNcBDi0mK71haUFt0dnjv+4/YzIOwCPFGG/71wQuX1STZXhDZp2opA
a5i4fNqoCvk4LdGERqRDx1XFmo855Ua6ytSD9KEbqCJ/AliPgkzAAiYztQBweZNL
CLGbZCfheQo/z/budlI7XZcexaEX8j/fcRIA32rxknKkoomr+Dnz577JvQj59aa9
4/mM1JCth+QqosMNGiM/ghQ0cxOZvtjOw1XBnsyQkmeCUPeOo5XkMYlbwdg7OnXe
c2lNmoN8hYA5zH7/uuVnDMxaSTNNI5wMy98qL1O0Jjhu75uIC7KBw0nzBp+gYs/3
+79b4SxnVj5xzI/T1lMvvcOlnL4wpqg+Igb+KhEqk3wrLX0FKZ2yIzXRNO3c6YA+
KeLq3HTkPDWwZskUXTvLkkG3ncgPtU0hYPLWVRRo24h9auWJqxG4vAoDumMkc6p/
5hxxRmHrP9plnxSv/kRzGz29YPHIkltTa4xu30/mZph8BoBy4AKOcwCSQe4ttjc4
3l0T4SH13xtyj5W17ZabzvKJrEZMj0LFhdWTWxQMx1lyw7H/FqvMenb9ra37PhW9
G4csp5u80RHSHjOqPVFUrm9geYqLGcMN/f76k4wsHxJMVZnPwT87cdbhwf+jkwm8
YCLn5AInnMEKdgXA6b9yjniXPkG1ZeH23HeV/9leDQnHm5e61Bqf5aSki946+GWd
bjyMN88Zpg75JzffHwsoGZJ6K+kCBQI6i8K1LufILfyQcCfzBhgKibVNbYd+LXsY
U/4YXFv9uVaiLzzaMH1cppkC48BuFvEKLJeuxR8BrgvQZxaUcJo4UpgCExLka3+1
MyzpQZh0l8rXEbOD5PHk6+MzvsST7+roDcargmr7rfYJIjGG7jVoQ3aYCeOPB5hS
Eq/xTXcmewdTnEIDCjoPJCUhF4Vgr9mKSLD6SHzKuOQDGD4bQ31vrZ4n8HXzWtMO
yiIqJRqnZ5kw+zDgM+y3zLNMyQ1MAcAHMa12lI40ZsJV3yzwApso6uMjff24439e
4FpH4E09ELMnmwU26oYqT3o/xFUH7eDzd204RUd8wAhc2lFA0xeV8HsJXJ6nJ+y9
Na+lzmL3QTjlSRbdrdMrd6vPwWebGWeSAB1P4cAEJa2zQvW+0WH36faLAz7PuX3B
33eJEFnI30Dv6Q5+e21CD9Zx0LT9nCxv8+v8MKtJAXbrgGtuRUXdVneR9uJuh6Ca
2uBEKSuZbSoMGHskLFYslQMAs8TG9UvpJ4SMxd1oEB2G4/Yc9YKGvHfHJ6AXz0bc
n8TyhCmGpkxDNJ2gQXHM44hw+3RbLhiADoAWn5PoSczJuJmArrnKNPXrjEBIUO9J
SeAOecCMUIr3cSsCT+vA1h/z52QWWAufwdV/we/BCluS4AUHknLA3gI0a6EzqpA9
mjKQhXW80bgTarZtlLq9o9iwb4GCtbsWv289tQpCBaH2ZdAerdyUlhMbHaGod5U+
YnAedVqPeuak8/RkFdqVhr06cKzAtJoUMUAGQTv0kZeoxbK70ktAtfGei5K2i1T2
UJFNcvMyPYNZa9W2WI4fByfU4T9uxJ1JO8xlw17RKpVRI8tde/9gNz0yAAqNeXRt
hA8ukA1h8lgYl7XUAKgWrshQBzZw/4ztIJBLZ0TYSwQeAqRJmCuHKcZruZzjGuBm
HRO7dQ9w9AgaGTSV+mG9wyMlgpBf5MlgjBqnEMzoTtH4k1rd/oxPL3l7HRd+H3b4
wbTT0c6WzRjwk8BYETG0vZMqaa1BToTg6Qaks1ZOJ1/I8yA2wSqu4WphD7ulPoen
Gma/pOn+rwPrwdFJzhDq2MWJh29vW8fCIHALDowAMJzz1qTtk/EjVbpc/EPf9rCi
VZf69Xvz6pM6JpqcDk7LbiEq7AY+DNBFtkNTiIMOFWy5TUmNWCswKSF5guafZ/HB
ykNhvPvmOvq3iS1HtGDK9PJP4K9F5rbYRhkZsyRDstZJj8/6Q1zl4/vg4oY+7VUC
ioLM8HbU9N3NobRS0ep4gM3yVCgdMlQOSjGJMWWX5RHUWRXyBkRqQoP4uWNtIJHR
La+mEwIyFzxqg0EspOvIEx7rydnhxSr+FqsPO2Dc7U33i6s8fXLa+knYo/1+T0nV
nvhlZ9dZBdpKkF7+TagQFFN1LrwY9IOC3U5ckeu0hGii4GxqBJuf974E9oB5mx7C
7u5nAvfjZD9MvDFIE0LAE71CpTdJBQBX3Xo+mNfurLVnfCrKKSVs/KiP9tZgglJQ
BBq3xHRDDcMn79Sk7XN5BmG+LWSYCiZTvKC5QjiS1/1c2nsxyb+81UIztF5zTLQL
5u5Xy192JupwPr02TMbtALcAw16499GAZmLjplV6geObyIEiz19qBUakgvs08L0b
kCQw4matw1GEfEeNzZw6Nrwcp/6MX1G8dWc6Edmajc2XckFX8NT+HCQ8V2Zpv4cJ
HZ9IWTGGaJROXraebPou6hhfKOpi0q1KRxASUMnj51d3whEp8+zKle3d8ULoxjHK
9qTb0QmffBqjazIPQqHEtz63TeYDlndrWOtiwY5G1lqAT/4czm6fYBQ0lJ11z+Fs
jZLZSOB8EIdxnLKh40UMu1BckTgYamKuBzolEARJq7tTgX7tRgRQK6tjh0Af+R+N
nFoxO0R2bxFIZjUxOVGgZJZOM9hMy/3w+jHvSaCJJM/GQpBGDcv2/+/dQwjoGqOu
dlJVUIrjsgeewzttJq1JAzGdwgabjJjWOzvPVhspn5HvXRxAL3ONU6mtRowyo8El
KgNikux0coT92vCLyGXohTZIkx5c0jseF+bGcWS0R0U+lLy+qrRRw3nZytRRIm+H
uBZEiJStL7J3TipoDbkTMX7ieBErkA3kOb6c7IPoF2/iHgSyCjG3lSi5A7R1hhd0
+KxtQU8A+VAcJalFx9Iu5K2p5crxgBB+Lot/CXt4ujZS8Sg0XsbA40LKoPWmX1hX
q2AjtOAym06mJUnM46FcAXF1qEYvEUYDxoQC/MWMWRXDGxfEAStzZmWIZj/UdWqx
DHdEHsvxjbgdt/JPEbizrOyCw5NQnB5zZnwVqVn1nW1IAGO0vo1zzVyRMTnyyxEZ
8t52oIjX/ja8yikFkME7a0OwRLsaHYGXHtOzSfNk15YFWX9BwakOZFuwQ7tHvGl8
R0zCHNuDXwjwdNmKqGEsuNoUZNbGQDABoWvTg5HncEsoO8vBMNI5HiTw4dJF1lqT
2b053HJGI9OzOe/VSzjCfIcpZwwSvOFU8cuSIYrUaB65mcSJALqP1pru9c7mQlPJ
ml3Vd3N5b3PYDWyT3lEyyR767s/2kZHXE/w0T7FO1s3t92GE2gAjhMWQqtLxT8Vz
RWdzNnHOmQKAkawqiJ+SJSSZ6hu7F0ATWr6sDBIM7CPxzlDDyA009ePgoJy6oXag
XjNCJXdxVxS0KM2/zQTvRSQNn74Su5aOvrPFgzkdedoQ/u1iPGhgyMroSJ9zMGjz
jWnPbdmf8BXgy5//DHQUCMZLETb2VJ6tX4dh4NGZF1Q+dvuo1ItYimcD5Yz/HA+B
b6+HosCCA8TpMAz8NgZB/hRk5vopUGaJGRqELzQ0rxrz2jpEXMeEn7gGwGBjqJPr
6f9Z2itnfxTO4eKBWQIpZYHxkWIld7/t/wBhtsk+2D09nu6tysgVXvj82EvJzwZW
Gbp8dDvwQ5XyNnX6OZSfdVsubUoH666Jf4Tw4kBOuf4uNGZhVawOolBitdMKQvRp
LYLrGfNmr8Q6Y1hUbtGf/2OjQbDkK2RrZh0YcgFc1oTBlD1Gji/+RfRfc1TVaf4N
ZS6a6C0XdGX0Kh8zboOyc8eVrh/zaXXs6pqZnmn5lbfUPEd4BCIHyU+bo7PLvB8c
VTt4FRMP6PMZbGBbnr37feJLz5VA9Q838ey+wiNVp1IRFATCN9xBfsnCXKEAwpGz
/dKKzL4uhXgJdk7MvP8mYEIUa1m8YHAC0ywF48NcrhBev7GnAc8zdA2Vv2RB/l/Q
ny/n7af6w/pggvFvUfHwQ7nz0GVyVphKojrSY87ktCbOaqJ2HbWbIvB6Qw+ZfEhk
TJ1D3cuvLVj4Lvx0J2/gnyCmnrgO9wrRxBarJNG1dfSel6lbgLMdo3wdugoxgGxE
vqBNoJzj+aaInklnwrBeBxUuG07nrY4+CWn80Aw7TQ1SuOlc+icmTSREjjQC2lwH
QOvJ/oZv8JXYcTez1ShOOGXRlJrRlgGDbfpRf6EO/YFvTk3U/hnL50SgZdDMCViu
s2k6J8EPdQXcEtC3Nk+VvXOgH2HruBZAECOJ1eKT0WHVxblnS/wZLyOjYuQOwkGi
wBClgG02bjlL+3Fnci2Z3ghR2G76BMXws2bPdxHrPPxx//wqs/LmBQXoKYtd5s8L
crm0Jh/UDw7Ehif+zXBSFkbulbE6PPXRAeiSUx7IKxACBsHbc609XqEHo6xVbHuQ
KC6WhYAisZ2EYXveFdVFudwMo0KugLDqhqBIdib9i7W9FbbZGtS2M+VB739hlxcw
3tIKKuD3YLviSZCdxwG5wmgqVdc5sHI4dfZ7qoF7nkwBprLNW5TeW3XgUDGxO42P
sLRt82CkPLpK6esSC4LVeK9bDwqtD3PN2u0/e6J3n0hbUBQ/k0bB8Kgwl5olIMIC
25b2ziC0ColOwZFw26tScbsRYfCi7NBhekdZMGbeqRnSiQVWVxRJHCLkIocLAtcb
bPK/SjLCYWvbKnUItj8vpeAUI/kj0beGRigXeDwS/QjQH2j07nL1hPkalwYAh1np
OXm3agsqtzKCFMEeUa2DoL8bCf7gUpq1OCxKKCX94HUjkBweNVEbWONqL4nXQmws
TagfpbfPY79OC0ccVMQl798FgoxdGXCki4DwdLpM2oQWc5YcnOewCO16VsVqGDKi
fWZD657wyltMAPWXQME/Gndt5PqCibi5DH1zOcJ4f68Yu8m26+YDWb3CsVK3iz7j
XqtZUikJHXMSQGp9VbCUvpMR6gGbJadCGd0mmlHUWC7kaS0OmN/mT5eYk5DCBEh1
xTKUQ8f0QSOkc0kj1fcoWSuKm+da+saKF2jN9Z7WOHbnXpbCKSffFxSxDvm0nKV+
/yTLEvTCc9ElVE06F2zmcmeP12Sz3ozr0dz3d7IlCwyziKD7QxvYfJOL3MWZsoQE
jEgEvrNtnADYfSghPmeZZYriHE8xakGB7LMlVQZi+oJuK6+cSCOzelhZOegXwN7r
ORZe33k6nxK9cDNyT8p1IXiNb2ZKS/PY2wP91CcuGtAWNg43T/u2BDYGbNgyQ0qz
VnX4XcsND9fNCV9GKUKJ71ekz2RaiN5kdj+X+0x3gEV8sk1P4sIRoT6jYleGDUNp
+tQYsEdvRKzfzuE3Hu9+6NGbMbyo/QbCnKMihg8MucTB73/Se4hsglNzoHo1dwdv
Jflw/rotihdB9pqt7zon47W6BQtER9SyxCewB+LMQmKGyg3XqyXGqS7mXkKLKHQ7
WsBSANWsI/vt8e+MRjBu6yuPwcNPlY1tlpwK37GkcaZqAmVBDrJ4j0RCux03oyn4
hu5VXeX2CD630LSKcViYJIyIx8EXQ7AC/5BMAUSoYiTmLUS6/XmoC28be/70zkBT
NIw524koRmKCGT9giNQVn5F8ZOneI4OT8S0OYByWNAw1cm92jqUNUCLvwvhTLO74
1zJtdicyxsDv8sjXq+RficYgbjqOAiZFZG8my/nDLeOjYD3YoF93gvV0hveivy/T
MgThomMClDgsrf4a0hxuUDGYVkmLmtGNaYRrzG0WsEugpZ1onDngR27TuYQlYf8i
utZ3zayR3Nt11NYTqYzeX3Swn+JvIWB16gb6/v0M1b9q9GYylmQgH7cH9gL5g3vt
t4FjbKJtnI8SAK/shnePonVC3FIyherBnqKdbohdpuDfxPwZGDOLLL04lS5oGMQR
qi4yVedTp1nqzxnVBe51DYPEc/bFVxVm6mG/CS+M5/PVxzVUYr/N3FPQoMNfz7wU
SziozyrAZDlcgP1XrDQBnzGbWAiZJURGbmEzH+TQWs3wDog7JwJlxsTyrhu0glJL
wrm9ESHq5SibvJaSby854f5iSSbZTJaYoymmRTDKviu6BVktrPVW/UXE+sAEBZGL
YALH6vmuaTmcLYtwAu5w2d9sv0A/ebY4gRKgyTpKlIFnppF9RINqvubch/+VvkT6
fUsVJiWwKP4bw8ivb73Yzt7jV9PavUzH/dItI721V69THuIOCIlaKYp5H/DII4Jv
fo50pyNj6Iob3NZ4DLPovzaRl/yrlECReZFJ4WG1kMYjLMnaR6C5jy3kV+0KJejK
OKMR7+arfPHsprN+RB/KdTiEttPUV7EmOixgBsZlMv/uGjNBWsZlEK4ORZk/ZKZj
s7vqkivR3RK8mqf2RcUpAjmFcChHa8iB5uYZlf2oUfepXdctKzIwufSTzTL1gfLJ
Wt+U/UfdwET52+xnbeiPhst2BkY4kiRsS5w1U11g2hqF3ROpVLK4ztaH9ZzEPxJT
Tqb/v+7AVyNJOXscN3Gg3fmx5KUM/mtS1ETi1leJrNYpGXP4pbvv9/2QON963SMG
PmMMzalBlaks7UTBMS+D+SUYOufu6A0yWifxQswQ0gwpDE5Q/D+lG5nqI0Ozzyl5
aIQpa754TZseicvWUfAcC3R+cVJ0CCMTh1mKhc0UXE6Mf+ElvaDngZWTRNefXS/E
ue+dgTtg/zsfuKNUEjHVlHfaAyYTpT03DUMLgmm2RUtEVhefgEcibQbih181qheL
nJQDEj9K22IQU2UxDSUlbJQdqb6qQ6t4jzJ7tfWj00iK6fqrP/OUFNPNd1Z8hOuD
CdW4amdeOcHUM9b8pb6F09kwctPORXkT1O5tYXGX+Lp+/rFix5I0IC6XZJR51y4N
9L4DZ7iN62X4pMFkoM5uIeuK92evXHAGKyVihaOuZy5FX3fvelDEq7uim8ma/UCO
a9TmhDpioRyzpWQ4csjraNMyObWu1ZDvx+WKE0AbZS9fORNObrPOftV6aOeaYj+F
g17z+nRLH5EdsGsk8rgRZVe4EB2wch2ZCZqDCzEO7Yg4qui6Tc0L//Zp2ZdWtaVs
T74JXNVbOJRY84riFNzziPEwVGgyZWKHwiJGcjtUCwijaqF6h469glWfylo7IvON
vZFe+YAYVX2uKSnQUmJdCcGWEi49RJblUl9oCXTiAzEIxtlNf8VJdEKdv+oHwnT/
hvtBw1pF9q+0AV7KxvZN25URoXfneVnTU3NN0wO1zNJDV9JWFgTlbjWPWYUwLg9I
aY2MXxNRNsQcHn89WvXHcQUGmQgs1p0MurvhtPyw0TjPkLsH9xzXa1EcRoSuwCtX
7zKHdcoUHdR8kpkVPLe3zjNvVw4t0vTcQDR9WhTuw5hKOoEhxOdiZcyUzLYMgISo
bdUucOqJ1egvjCT8l97zKPoT39swMhLmMzgo2SqtXU+EvPgU/jqpJEf+cC98gPhR
m5BxMP+SVTGMVfqT2zZ1MqHSlFTYZHU5IfdwoIUh3f/KNQwWW3Z8yzkKORFk0jTi
Yx/Ltd7G1JMsnMj/qhrvAcI3Ul8Nt5K+LJUvUoMdoz2ZrLflQwWAD5DpTwq7vSa0
gvnhkSAhr3oR/lt3+FiLlhKyULq6SnJrAtq09yBLbT0qDbsNj8oPMWmIfqb9/Rsc
tkvfmIpd+3WFV2j87kDpZW5p+nmKYMDtfnj02BTDZAF6cRZw6JXX4YeCeDvNm+66
7WKH3nHa7vewvuE5u0YKh37dGfAqjfx2lAakKn3T1XrG/lceBmXMswnEYCPBIBYJ
+sDoQhTlGSU2YyMyAJAwzqEf3aqpBgas5uSRGrJ+stXicCRjm2fm/Qu1JmbL52lY
S/pyXFWLWz+oNWsryUd9Mrnj7T1faiNN993vSrh4k5c64/BLoT7VnL1rLbUtEpNn
PRFuDwt8Map/h3IvyUqvGnTLBgF9ZhKE6UE9kg3MIPnXYddj9N+dgpT0oVY+bp48
Im5CWYpEJNe/NButbBhjO23kJfz9+vHXdo8azGCLgcbPwKhRmOx8j2PRnsMWsLqW
eCVkfjJGA61rb0sxq7w7uvkkNQEJtbL0v6KBfZ6h9Q5+8JL2lZxGN35g7+K4OtFU
Q9Q0nkf2MBMhCYKSmeDBqp8xl8uXkqWXp5CGpSlCKB/SgTXkNi6kSuZDDSP0CJVF
aAcC+ZlQ4PQ6tUzH+Ik4pj1TzICaYgW6w9URUNK4lnPaJoAjM5M1OX/Fb2FE+UCT
MtmDcauobkCnBykcJu2G1yrw6BEXoB1yXhL8axOKajjLIqwPePVoJrG5uUy3OLxD
RXaseQbiNiJJRHgy69g5ItytCPYQjKaAfhTQzl+lo3x0vtDXFrZt/gxh9cNErqlZ
4LUrpJVAflJE+5oLYHnuOOratT4f9IOFx+EAH7lZJ9L+XP00Hs2AzpMNbqI8b+rg
naBfp6er5ykid6WdlinfADWRSdKUGUe1lVAOtBa7VZ0ufFYDJDza30dCMKMteD+T
LfFEYdflWFYQHMKj7hUqtRNOby4Tt9dyzRVqrrlt83Kgp8eewJJkix3zozofGdrD
X10YyWMZ4zJw/gbEaXs7JRiaYKWsQSrFaNLMvPsYpkRBBPNoivtACCHTDD1WbCG6
gJY4saI9fE0/pj3kxV5ob7SV7r8loSC4RLN+/JMS8XnCca6RF3nhtj3b+kL2+Ma6
FaWQvw2ulqRCuVgAa7m8E8uiz5hHD4LiqZiK7sp0yYV74tZNqF3lKuR0xll1dYgz
yBGpR4vXtSScZYFcoNhbq4oU2TCEDkNYJQ3hnj1VoekNQtBhZbXxcJB9z8za4KFV
If2p1pZIHSLRkf07i6uxF3Xu/KwxhtNEmKH1yH38VQNT9MK3nczREZhREwxXEBoc
0Bdu0hDTQVyvCJ5RHVRzUxPKrm3FSMvryKMMespMYXbkc5WkjvwHU5HB6wac3M51
lW3uCzHcpQ6Lp6BO+o8ro+JFFwNxcQ4Jv75JH42VtBjWNZ8Q8aj0F96VjyWJegcX
zalh98dExGzep35Ru9FGjofdELG4emgAV6zk+0COpozErAG626Eih7eKZbsYn2vU
e5v1t8eGiEgF8WGWtasPiAOHdUoaG+/5X9y4gcyMA/s870sxS9zasgG86saYdgit
UwBaZJk2Tz/5beZZxniC/3QM32Z+2lhrxepy+/IcWti2E1bI7RIIdfj+XgU1oUWC
6nikv7LlNXIlzgN/alrnDJjjN5vAKgU3X/CTOu0aAyggh8tDwHT9sp99Me3ll+Hy
1rZRoZ60f9tzrxZfZCYTrvi7IO3SzpwcV5MYkaaZ5CMtKyCjx2kzOu5Taa8uI8vl
RefqQ73vDWupejsLu2EZ6mDCIBPq0mCmLgXGnRsI0we/DT6JVGTk+PqZ7J3CXpZh
eWkNOxkYh8Sq0KVNMvq0JwRpvFbPJeUtBnzcJQlVRHCvJah4UBeNI8VaIjb8ZXPc
MBSX5vVBW+xHeKhpGYVpXspQCQN4wFflF4SQMqAadSgP+s/eOx3/VwlI0QFYzMIb
i6b7+x5rUye16Omt6k2yIntgVUAx4OdmzwkgariBYx0VxrECvXa92S+mG2qOSJOy
V88C6j//Xtf+cDjwOaXVefMLuWg1FDEfKc+gArNFUysSWBwaHS7uAA5Zr2S6lfJf
qlbQr0GANAGbOsVqR3K3C/b3suRDxfJRUpMwM6CjQzQdW1LmQvhjieKGzRdNr8Ly
galO1gA0E0BndyCch/tk7QsmZsdBLMAwQ1yk32NhoysD0/qkSZ4v7CokxK8VieD4
3CtcDKq76/qJpOW65/puDm2CP8nE9EDMLscrwPadX4UWcSFy6deGd+X79aMRDUEI
Plgii/6cK2tw9Ya6zPsGudK+CxNT0f1HbUJa2eQxr1AMa+5UNLmvOfTpvYawvdsp
VJ3wjwvmVHfbhZBprSM/ChE2IfHSeoKRRHWOT9KtZ01hIvX+Fb+z4kK8r5DNE7W+
0P/eP9my422tvZQeoWA+0nHBSnFTU5XSbN7Mi9RU4y914/in4ipsIuZN2tdAnZg3
kqX96kIrXEIFBCHH+IAA7kYzlK9S6l26I/LJbN3pj9VGzQTbWQy94PmFmBaJ6DYS
fM0PiaqU8CpqeKwy/lJEE4PRbfinmJbW+r5SFKBcFbThYMxOhdy5SxVINYkH66XN
U7kSUBSo0mbYRtwNdkrb4HX4sZ9nIaBgTfPsb4mSwB3m2Xga+HUgjnt5S0lI68b3
I9Hc4iqf+w2n7ekmjNde99Q/JtZQx8II8dxua8LIX/1+qH5SazzyBD3haRkivqq/
0c6I0iWgRPBv1y8vAGM3MinFTzvSM0t2DqLs91tVnMI/uajZ6B6AsF6Rfhc0JQ8z
iiFOJeGf/trIN5mgNvTfKYUfnoAE+IsFSHkIy9VPRp5GMsu/gb4H0v32euw1XiiX
FkS4vLkSRVI0E795MMDXBywIbvXCToyWN+xGtZc3Jr5zdT5PHk/D7oUshhuNonkf
jhS/wGkueBHKCvVBoUB20aE8eT3VP82RIsWVgQdKBwKLAXjjunAG6N/eeoQRaqar
OofzgWkFp3FtHJR8DsF2JQh7VNWGmDK9GXkdVYk8cbSguQBEly1BCA6bNIy5RvzV
GhfLKBD6UgaPrq1os7OQF5sPS2RX/h2CjL6rfeSF/zXw/R1mqOUa7b7kCKlOS/9Z
nHnRkIfgJltEo5uI1ZOgxbRzv8WzlzJl3Rkf3IJudirQwKI3PMwAOmuSpQD79MNt
+VyxHhrvard/aJmJMc3nRJJDpxYycFXq6pkOSsM4itEV92Qhtd9fcQc6cHRkh0Q9
JoprJIiw2qcQxYe2W1EkKHOUl2uA7HFcX+W846RV1x68EoZ1mdKzvL2dwHGBIVOi
zORJFHG0hpjXFnJoWdhAH0PtOi7gRnMWBSk+0sf/M015+S5Z5bjd7PJoC9SC/gq1
XRpmHCHzphze7f2uBK02d9kGd0NMhpWJRwT5GUuNcK9kUSbJSZRFK+ofFV+XnMYI
g3BNRrfby2fUG18fL72bzAw/TFwmIT7wmzg9iiJniFXXq1i6Y/P2Sdme3CqJIYRS
/hrda0K/ukNJkxaHz/QpvE6KEnYrqz8wQd8MBh0Mg/0WfE+h8IUI/qfBbGNwqpOV
NIPLXlNqozb6yAeSbN0jTIOUv7RCoRoGZJWdJZ2v9QdRByNW8/PYJ94Cr/RXunbZ
d3vRg1AlFH0Tgi3O29B7n32bqeHT3M7XxQwvaby47pG1wfML01yPimDFps2MaBNo
s7anvLmQazeuffxr7tBh6P7SFsEFSMmWvm/QM9vHud6/UfQ6s/HD2rpfwR0qaNuo
AcEeLhPLFUCWjSq8dLYXuVcYjZLF+VqUvoHiCeYRs8SH5IzW0PNt+x4sngUD03nL
Zqf9Aj7ZRJ9bJBPFql+EqahourzFBzaGVZf2uFdKDOsAfIG8rEFBnqUF1+VPwQzp
4342up6f2ZWdbwanG9rd4uzB9c0m1JgWSNLeWJzIMSC2bDO+mHz9EA0OdIt+xnnS
YTlT9iEx/cuaFW950dJdDmf3e03U+Qp+f5WWkP6NM6D8/7zuLVevPnbMeXgi6siS
AvKfg/jHT2+69tSk7IeiMhJ4cFQJwFUZLn90hObJz6X62xrSyJytYIkbLSKsLqaO
7t+C1xYnjxqfE2mI148159us9F3Si133XT43iEJDNBdN8tfWvoo3DVZ4A4RHZF39
iaSnQhYVrAwNF/xI/PgR8w2VultIA0MMwd9Vsvu+PM4VBQ5ttbSmdFgdueC3fmr0
tj8tC+lfiOGB4Bv+HPG+ueIRkyIGnuC1ldSw9ev6BPnOCz+GNLwHniFqzitxT+NM
GFMhHntyhxCvET4oJGZNql1yFUL78YH6PvnGiul1UrOAY3GrlPYldUwFc5uAVfWH
xMwbZ7VA+vCovyUU31sGJ4RA9rJ83HRXwBsX0yyDKbxOyf8McRnItxyIKnjnAnbJ
NbQTFMzIocnMDQUVWX2kBjiJopwZeP7NeSc7dwJ1WDMOP0bTlVRShIrRrw+2vh2O
isKX5GV6b1ZcfC/M9pRXMjnVeMU7uiPjE9gUmldUAqGFAyihkElK6VlR8SHR2D8C
hVR4P34bw2ciiLzoaCulQyDY0y83/jiqioVywDYNsVeZvOv18OCno7jhcKSwTFdT
8N50LxEQxzim69duaWnm5PwAYJ0zAhvVU5A0XxVj71qYGlcyNl/mB3IF62DCaHpR
xK3vuITdvS2EnzjSEAFB9uQvCVfM2TkLyHNacZGqSAz1lEYz8ipRomlJD4HkLDjD
kJ/PJS35XrCvTBue39vKJebgwqptIP92fA7R+k66AJdDKW7xZTpfxcN0T5uRps09
z3GscMXw9Ta8+B8ZdQa1Ao2Vtrr+SHRGeJgVM9hPtNbk/ZAlQzrywSMVhp45WJIT
cJ+bNQRMCm+k54rgSNFjyqVJS03/5+PJUTsnI4Rf4vNQRJ5V4/+Vbg0dxwM5e79D
--pragma protect end_data_block
--pragma protect digest_block
bpWw5p/IYMy8/CI5GFSSuwZY44E=
--pragma protect end_digest_block
--pragma protect end_protected
