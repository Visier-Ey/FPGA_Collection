-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
--pragma protect begin_protected
--pragma protect encrypt_agent="NCPROTECT"
--pragma protect encrypt_agent_info="Encrypted using API"
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
--pragma protect key_method=RSA
--pragma protect key_block
ZMUJtvL6EixKiAn9GoYv7X8ThMHt+lKWtyMLH4O7uvUd8IM80uxHV6rv9WXck79H
FKOTkZHLdfQjD5c105rXfacnDQ6z2n8vLDr+NLHclncoh7+XaKrQN+LBl6TiGawS
tFNy6AOtoKCOH9Glj0AuY/SQ+hO1MvvIotzssoB4aZpLH6S2jOftT5M8ltHK2G7t
/ac+hrTgct+rnqpuG8c7FBIyQkPH8qnsz8O9yEIM9eIPqA6inpi73mQt3HlHrrUQ
GaoxlPqWHrbDlPODaw+SZFEnzmQe32e/JVAIuOg43r1Siz7LjnIJ5G+rt4bVX8/z
S5wU1Lls9wcR/u6C4vg1oA==
--pragma protect end_key_block
--pragma protect digest_block
CBin2t3gBIPdBgoUbpYxIriN2qw=
--pragma protect end_digest_block
--pragma protect data_block
YYpA8qD5dnxuaMolSGflctTaC6xPIxjO7xI7Y4YOgT4iohcZO2o9Fvre3FPAbK6s
UlPKNJ2a2ohjU0z/BW8Nak3Bu9KaK1YjCGQUDUluqrFSWNYrSuWN1JJwbcFWjJBI
/2R/+9hm7vwzOzb0vnDOZRf9yYnDtF8IaQ2t/ZjeJwSAXnUsfNajjw9jRjGTL8R7
Tw8VT5ih17ebY883iJ8iV1v48mvMs9DDhFd4UyvXGyKntfpoPntBN9zhAs6fN7Qh
/PvC2Dj2RQgwpl7pJXRZTSiHHe9sMLoheNGXPqKkpha9leS/3tNe/e3Z9d8xEQ76
3XOQUxlNiZyiOpeiQ0b4PTDDVER1A6T/p+LEhUtA/MtgwWDdXgdqO8op/HNh/epM
ee9nScX9hCCv39qmKb3XLi+Yc0m2pU6mAKQ2WC0sHIrvEIrD0HKvHXlIRr1Lv0ev
zQ/6tlUOfOBXG0WDT/rfbsZmYrihFzwPLpuq+L+xwHFSDgFfYyqLaOA2r/sY7cF5
9wf2ORupitaNEisHjvpkd2MJmMlXhuOPUgKss6mSCiUTk6U0nIBnIrjzQLXFpdwT
yBDYWWlqgZLlLysVF2O41h3QLBGfWfTgfpKx3jycOCME1HYDJ73IAFu2AD2GvNKQ
iJofBzZihtYnjgrY5MQUoYafEblkqKPDxnlJMRFBhGDrzhbz7qn50vxXLn1Sb9LN
CQFBMXUYN/mt5x60mQbJYaRY+zcszqJuqW8S9JIpKMl0QagjvPo+tL1mW1AoN6pC
KbvlImXV24GKgaK6Ebml2UNIMlgRwFmHeY+3xiabHJtY6uVa2eoDDHYPL8ivtyfv
pkTGlGRv0n5Z2rRc9i3Sxf0RVsHfG2+4n7EweOwU/kgoZeXTMpxTP1UP811/4UOl
Zxxt9i7j/cWf8RxYF3h4iRLdFrxRR+f14bTu+srn1Tk2JAYaC8xHU8i/N/DvQrkK
eyTASLl1Y7q9pI++mh60siAVnP2Ub40tkDaKpFi0mKO4GBaZvvPISeDHwDKUIE4A
yuC2w9/BVJzLFC9Jv4CbvgvM4Od/95hqVYQ5NV/KEaXzFif9r73gczYOcvW1D8ZT
KGCo9x1nwu5Cc3guQCg2UlnpL0TjeFPFa0QCQ1kKFY5L+kYNOfH1j5KiETZOc5Yu
Vb9nZ1iYIKD1dxigMdRZXgn1S7Ki5N2lIIYscRlSkHrIRSOLvezj5a0xolXrU3aX
dZyWDyI7Hr7uQBD7dYYD+fjnEQdfmJO0UlB/0U5d2KXXrrcxMo+GhAMvSvhoNEos
OEVa0AjtwChyFQqWouCgCUCwDahl1Qvf/ce3Lkon74J8LbSPgWLWhjP49s/8qO4z
TKCBt8awajjeyLPbO3M6E+nPjQ1+scDXL/YmJdX45Wp106jA58B6tmLpqY9D3+bT
ie9+HeDqYLW/UOtydiyEl2uC01v6+v4GFoac86dbsrMfJ2jSYs+VwazZGt4Fh2tn
3VMPC1q4J04UhPCdd7MjaZMJTicArOcpt3i6SeSr/mRchDXIQMImf+AalSD+LQRA
oeZ2CRgKsDoGYnk+hqPk4kWBe71xxT7xCAyAJB5TRkPFhiA9sMAVbcgrW9xXXmCf
YeaZH+RsjkeCskMDydyAfixp/RbekgG2zs641fmOfI+HLlloEEr81OhQkb52TUe1
lbjyY8YUI1AJSFpGH/2n9N7ekAFefn0Cf7k33FiCj7QD4Ss7/52b+8HynM3cHYNj
rmJm+ttQAwJmoLitk3J0PBfvWMYlkm/7avq8VCAF0bJv3kYSJDmuoepUBAuXG9iN
HdVPSlhHUxa3i9uyysKdnDslRn3URr53ycaBLW1NfUJxOiaZdw/9ykCsPf90SHW5
SdgIpgusGv15kKvho1bOfQXixzthxcigdHFRL9BYaaKihLccqtX7WDhWLy/2F7Lx
AyWQ4EfkRYLWIYo8QI8a/t9SUjAVXj9T3ssMWLR3Owjutqkr+Xn968USPaSzHoVB
vG+1GknASUksWIMwbpoPCsX0YhF51omHya4iBtfxTe9Oeq+pwHSgu8usacXJ8rG0
8j5X+ovUjDosiufF5q7mkZ+V4bp7ofYIG/xHDRSzj6z59/M951e2Rau8T+0pyNda
x4fb3kc40jUlrSjgSUFPjs9W658rt4nkewTZyANL1t5i15UpFuF7eofDZvFSdbCv
92OwaNwWoBFAOJA6/ETPD0ODFm/MeJxqoNgnf5yrQvI3GLScossZt+zUD0znskce
UPEOVijEg++7UBDUTnQQ5SGZhL8l6uBjHGalgI6fE3arUR+0pcy+U8CtPIEbi2T3
dXhmmlNmabW13WG3nSeAnuwA+GYa6cmhdX/jwDNSGcJJlMQteUbikONqs8kertdJ
Mhc+vEZabmzH0vUja5flyx9Lf59XxdF7UhOKwkeZg+Ja5Un6zJn1TQXfPr+oCPOh
gMg6qR/kdsMy43qmqrQFyUEfp8z9AoeM2e6iHc7bzst3cwTjtD5soA0jgzSBbwBi
uPvzPVp2+DOLpiQu5WkPi1vIUT8ZHgnI5KKdI0O0UBZFW5Senl4RnT4VJcKXWmpQ
Pil/T5txo3jj6b8sIctUeDblqXJA6SgvRSk61K5so0OECwn0tH11vmlptHh2eG/P
CMcakGw5DAmQsVHakz6cNVhwZ4JaWPqMGUVWEyPdsW3xuL2EPPd/20q1YDu9OzmH
wek6p4DMCUycJCWmeH8vtDaxPqTMo/2HxGRw1aPHSMGGGaSWKZlHqGnBaAPMD12K
oktZ5vg+FV5D15c0nyrYsWINIxwUGSciWzJ/5CT9wZvZReWu0+EWkMLyLQsA60q4
E/1ENBlPifSPAdH9qTu2bTHeIHo+5xZTE+gOnx/nmsMkAkCiyQ1eHExG9NhRHj/0
16nZVUfqfsmpbcGQJf/uc2R+O40iJUSia21DxoRHJ1poXNeRcbKm3NUDs5NsRwij
wb+sa9dzY0yXCH0Vq+qiMSupZeTAqd0tJyqXDn7NfaxG9a8IYq7ZXPyuWiuv1Uul
pvLEQyWTgO7bhcUaD2nXcnbAaln80VeTmU9q43ChffDAWHXJUoriXUpF+vTNwcU3
vPHf9Y2tjDexBOYEHa2p0s1NIVrdWzVh2tZQmEvO9KLJweG7zbMMXyiLRNM0KLAw
BxxsnCWKz3Dj2rp4nroasb0JJI/hLjIo0xBOnhT/gTefQP5FlmORRqz1PVRnnjFI
9Bx4UjMGOJf9IM/xtDzdEmIZR3quZGZWkZ2qnqVtiEJbD+sRVQs44UBLuUbxbwYI
FfeE65PRrkd37/bfArclHdawMum1C3+pDIqPuIJe/taTNrYivEk6gQuednta9gLU
Id56NH84eBD8Nekg71gfIrOrIVUvdZ9PVMxpEBbKkPKKbzmcoxaJcPXgCGx2KYPh
3fTrxkWhL3udC6KJljpI9WSYc+2RD6n43s4s5NTvuw+Vx214rkXTGzG8fW/3pLre
1AM1RG2AvNfMlWkauGl+BD6tcWSWZRkGJUOD4gaQtRAWESmESSPONDP3LX1eKH8T
f4dLVT4H8sobpTndB+GbEHu0IndA0qgI7KVYwEbTr2s8LdlUs1SBfpn9iAEotoKV
b+Ic/JgntJIuYCma2Cy19W641wpGyRp/DOFoSWtleyVJl+8V7t1VWfLptUYyR7r5
Qaw0DK58hYPtopsNY6e/sUNDj20yLZHx6GDilEOMv7099CSQb2+V58vAjvzH18Jd
bMztrjGcss+olqiKcWG7Q4eKF1m/mGkB9V6aWfDUF0lzI/0N7WiK5ZMajQIbT1B7
ufdk7O2jBQHA4xwn9YDanOsJVeu67rTR3SKEYmx7fH+UWcbpj37RWlSsr+lydPjX
JNUC6Zfm8N4bW6Z3bskFEYl6fONJDp+QKVQ0TpHXTqWRsc8FRNbTbSp0rc7b+2t8
JMRzIQunYoORQEDu1SvurZj+JNtMRRnQj8Tj7Q2S5FAsCj0mGxLvygFjLe98Q5ax
PMK9eDcuBUmTmKWQe+4+npOUZVX0HBr5YA+SkrtJ9zjrmheqnrvml5HLQl50woUG
npwVUxHsFNcTaSphmDOhe0re7QtG1yk87d192KymRY2h9QUQe1YiWgG8ySmqj1Vc
h+C3pvV+4srh3teXJa6/bSVTdEBI4Pr5gX3Kp0YQG0hfycN50iGx6N5Rd0jGhyU6
1RSyorcnHMH9gsOqd30U4k7oFjGpq8IN7XWoQtisICs9dLBhpqFJZS9DVVw4fijj
CByJwPFHe1WmV6zw6cpOAZLiMnUensSPMgWoeUaVNKkRa7caQvX4SLMmwakH6Frg
yBJQBl6+GE52/5mzZOyd68u+i6D951VRJAZbJ2klGUt894vg3+ujIr1XBnNZDkhE
k/H9GCv4F2FG1jIszDoI398KuE9JD6W/hC7x2eCL9VyeGoKaefuaFPSUgH8W6KH7
10kJ8zFF595RG9NKwBJZOH2PFwyMr5ENOI+a2tsjRBUoUj5KIMe1HvWfoz396C5z
pqBzY8ArFpTPiizUre2n15CAjyZdJqqrbCqpoDVbYIwxNAeiNidv7rKi3N/YJCKy
y5K6pIRmoGVKYMHRRHACW+9+Yo/SFFJeu3zJvVVyqUwPW8h+MqJGN122JHjrz6nv
0hUKXgTCjdHI93eYAqTSHeJVITOGDatoItN4BveTB5b+BAXqpboVfvADjrUqm6/4
bQPi8+3Jqt4zxgn2dCr/JubZ7Rvpsm0ETXO20m7vHpQng9Ckx8kEuAzBxA7bS5Z1
GH8iAvK6i10zqZOWYaGmYDZRiKuiJU0rcHL5pQdW51hKWrgfGaHtpmqdq2R5YH4D
vl9p7TDlL63enzvH82EdhV0/ueqS7zYarUgGNOwm7VKbyIYBgZXGr85HDKpjWjOl
rsEuI62ELrVuRMVqQbFnnT1K1AG/8vb44TFtvwOwCxCnmAXpDfb8F4RR/sKN3f/0
mFSu7XBnniSxYIFKGL6Ivu+AyRC5/onMHCdDyeSiOm2JU1V1o+qdDFUA7mh/dCnM
Knr9ZDF+lokyGcV/6CIk5AcDSJUDZOuu9gcICom3UVWd/GYa1HEM5fEnetM6rOrf
XPp+Lf6OX/hQXMp7YAyxo96ch4JBTWBYfe/f4Gbiqb33v5Gyy++0RLyf/+mNEr6p
Ij7exj1plL2Pmnh3WxuzEw0M3PWyoQMLFTjmZq7q6BedN+Dt9GiZTJQ78+SJwB9I
85IcG9h22M++RxHv+O1YBK7O0gJjbP+Fgfhr4KeCBeqAwr8BAD/q/Q4OpQCoLzj7
/Y72qgrvg8k705NWyQJrim7u0L7YdTGf4hKdiUefviS0M8jgZ0kRBewMHDY/q/J4
Nd3uR0jfdHT0CV596ej3lKXzdZqN6VX1/skmgw2LlnlxDCIsPa+94P1Amncsh8Qk
E4piREV+8WgpOaXzl97iTmvV1bUSzBboY2gEKYqZP+ozKHleYD6hAPVQnX62v2++
ZciU6spfLAq0cwU6OmGw7VJhhN2XMtAAeAch6p2ZfJ3ZMshxFOv4mgoOjqv+KJON
s5BWpUEhrdj7z6+j+1LKG2BfjKMgpIL/kIl1mcWHTlV5/l36LvD2hvwrhDalPG7F
98FPfRg9wAga934dOCfFMEg3SEloaMXNnjo0hiOAj/VPSA4ER/gi9kvakUBYnZbK
KdNBAznKX0AB1aK3ka+6nG1QsS/6Atmd7pYk5ziCbKRc07wPk6BUeX2gvDF9OldZ
xY981cS5vAWFFrznQlBy+pIyTlZrqhC7BDadMYbpUob4arMcJbYiEfRpx6JFTaZ7
WKAj4x3n44V04YuC4TvL6WeHLNRH0LyfWGMwBNEYE6c5esKyuRAo1aVZH6SwT61R
f6rpBp+zrLvgiFTIfMQjR7b3CkDnam1KQO4HtaUed7JWmhPJgxtdaBFx4tC0oxI4
k/jElJZfbAZy5PcbotVNI0sdDI1IGRQkBRMHCaBM6x8WPWffLohRqVJ21lHlttXB
vRLeHrHfJgbC6UImIAQrg1WQsdyMxU0W+FCO+hPulOOPcHNrprrSJHsM5jg9XK2u
3WIKj9eUn+U9c2ANwlfuoiXmEFMz46Dt6DbhvpsJgEc9/yYNWMM1wbHYp3BKt3xE
nviTDd9MWW3+Qy6wwHa05eiduAhRRY0xrA40+INN/1ONfGoMUzBp76sZbuFZczzK
QLEfLkR8GU5bC03mKYFO1ANMqi7xYXFnr2zFgCZGRBM0DPI79GldDjgVxyzqyuVe
FvFBITH3kOrXD/bNsKyEJL+fz5rrt4e/jdC5F3a2NO6WuVQdLfXxliaU2gJzgj0o
Y91usX34zHW+tiucDfyhwqoTCnJSj143L5lxms79iPoJQ9zVRBs2mySTMO00jh1U
jRz35PwMgrjfSqE78b5xT2/VadydlyBkAFx/KqgxunQmlx0FWBolg2D3LRz1zENm
CYg/C20zVrZaXrUg3LPCTGno97+RIYnB0JlDLBt+NQYDFEKaSzq4gEfpFa9IQ2Zc
64goJSsOoieNy1UOsEl3YyyfCbsm7O5DNxq5lmISpg0ZoqKUSvLa5+R/f4Ns4im8
iI6tuONzRWy4AH7nPH/EtJBzWbjc7DcIlpBuDTZJbaXou1sbh09p8IObTv93ZxoX
gBzsU7qDELEgHkorwvlgM6y2UaJD+TdaC4HEEyilyNUtIddaFeFGvepfjtPQunoJ
eWjX1amh8/P9qTJeF8+RcuJsg8WGqStk/bmnCdoWVP72XS401fNSZ9g1b1ZS9Uov
afWpax2EXw8neljoXnag2X/ZsilDkXr/43XdSSNWWtbbStz8Qa0ZnHpa/4qqPbdy
vbazT/yPUyR/43sTsyvGrSUt194BQuJWIl/gRjTSWbZ2BWlxJacxJaKT6AFppEAJ
VguK2zJz7U8Z7Ttb47glREYT1zS799Llhi8zJXJrHKJK9xJK1PjhEANLUMjDt7aV
9CRXyJ33Ez890eQZtOrXkv5xd/+E/Cr+rAUuMhWOlfjBKsoL1XozJln/hq99g3Na
W335WCB1ZGKJ64y0W6uuWcX7tH/FjY3xI2xSZPcLgbaJhVH3rCxcI4q5BWwAdhv1
VV42jQ3XziYEaPYwawi/Nd8XDcMKGW57m0kHws8kNP+qBS0yF5XbiadBRnZ4WGMG
RnTaWE8a29X7Y/fkBq/wz/BzHeD7SXV+DWZurzrq89IE4B0BNRYnITXPQO148ony
uATh9reG0r+PEaAg0d5yvNRs4DIClnBArk5pIVJ2tM5yUma/u73QIE4lPcpOgpy0
6cJhghjbtPcoLx0hGQ3Z/JDjuRfQttAQwveVWSB4BegGdyn7fqBAmMRdRjWv0dsH
jmstR1Xr9LJphSWgLFDDM9G4AYh0uCKGOEmvgQCQKYSTsb1bAzM7CnWqwoxyWiub
/05bCSMwJ7MdKZzFUSsO8jzzumh3X27ScShC/HJRMtu1AkoXL2EukNECWngcfHmj
ekAEzIHrzc7xcU0mDHTD+QweqPIwlqLsCdDlIo7RYq+8Ba0E0f4jWSJKXI+g0MNV
1U3GfVyjY+S/CPipFmnF3Bd+cwJ6cwWOSAnGVhdUGCwjKky8dvbMH7/A8DpbriI3
y3eCZh2LEimB1tgyWBZJ+KMNRFbDdAWxIyr0MNEa/VwMRg9FMmEizSRBu0B1iRom
Uqk3Srk1AWIzYCm5K11GABsxdkb5QNbPs3kzgqR8CecChr+DJsciP/x0RoWyrKPL
aQ9iD4MBMI4pFS/LHZ47tx6HJbQqAzYww2OAGxIpU77U+FfLFYUUjeyGDXsFKnMf
eWGklM8F1zZz00S+/KIm42WvSVS7TFCoTUuSqui4Ouaj6z3y46BgBS0qfUXCErCd
GSG5AHigpdoHCsXMJUUlFLwxr3gSCsyWpZaYiKQeKiCuq04JyAEJ3z1WrCpWvtAz
EHJbSfCtWFmQjYZAKtYwh7fjg+cGyb2u9dwEbUMh+7dKLjWCygIPp/Xc0W9knPX0
vWZfvHlGzFR59OpIp7kd7i+yDEAllaSaDcbiP5slVBWGMG4eQfeLL43SUSjRrBtc
e2z5IaRKongarIJt1pr6dHStOiWJMNbn4w2PWCBBVrnwW37D3fb39hw6EWGf8s9S
f45OEmW/ib1euI/kr7w+qiNXw0n5gSHenHyXHY6wp7JLMqu7PlMqu7MchY175n8v
AVk0fCEG8+qI3f1O/2lTs9DzQ7eubZ+Uo+e7pJgsEAHd2o4oSqtNffubNuYivNyl
xG0fN48y9yp+7HplBYk8UaNguUYdgRxYTFHWSJutyxJxP5wxEIqJ1Y/BNoemmAu9
FvMQaiL21lGJ9Y/f1oyFUAE3DjWt7AMLQWdl6Eqo7s/VuMLt2NqJT/KJatAX5+5b
DT4l5w4YvIi1/C1aHdjLp9bVBSwM5ZRhsyMzrQoMzpwqdcgJQzlwC+OfKJLei0A9
N5iqUxUyUxmD5b6EycgZlnsa9N8OJfo+0kik6Qzh3xep7MgHFYzQ/ibAeMIyf/d/
yh60VsKS8xslnGT+ksJPFEvUtrsKzttPMgQP46mSfJIkqy/oySsXzdlI8V0qY5FY
Bvet9AuzhQmZXfrEXsaW5es1YNx0/1hT/kp7gOLMPUOHMYMY6Z1jmEXoKQwnsivT
9VD+xs7txHFmKl/ekSRCdymax+s0r/9D5sFbxZP6H1BPvx/btg2yzCbFisPxqCPu
D0n+I0LU8RY0yffOVpJzdTXrr+e764Ay2i0GrYfaOP/AbfEfGdFpF4mXQRdQSxub
w/gfOP8KP5VNk8cc8iQMsHUfHxrIWvabVp5rT+rGANPUHetnyiEUCOG+mEmP3xFY
epym9/a2dF+68eiiSJycu5QiEdqzlnzaIYNoFsVRku2K2qt6sAacqZGu0ZKDZpl9
y/tiJvH8V67Uv0kr1R1EBIrorqOxXXM8b3A4aTL+pqIi2TPTn6TzC0hdeGHoyCWG
ietff6fsmzj2JO5sfbYFcAlMBJv4BtaDx4JIW4d0DSVNXFiEs6+to+sPbWn9mIva
TCNttWQXxCcWXYlLmzj9CzMjC5ssQMDhiQfVy3ALUdcqKd+klOCSaNtqsotPA7hP
1CGnvsri2DyfxaLtJCMicVwi/1/sf3HbEjlJ8J70Mcjoq3RQdn0lkC28ViAbIaCY
2mvLIHf9VDbu4E0ab7AvPFgFUzJFUNfI4TCdH57v/ixuxLbEFvcA2suh5MUoWbez
GRgM0mYIK8mXhdZRAUM6WPJX7QzYDz8qS67xnRmZ9901uToxHeHSlTe2RXyIIdXd
faeXB6Scw3JmL1mHqvrIbXH4sg0r7Sie4+FuIP+zxNrLVglMIT/3+LdqNXhZq5xG
gTz4ErjtJy4Ylg+pRpk5ixMVU6MacEx03leOEXZFvYSNOWZ3pbmY076PN4af4i1O
H0In0toP08nwItRONrzCxx7ntQFO/f9hWrNtZrk5qHLp6FiP4A7z0OpcPgBA1MXk
v7rOoF5ViJ0SAcwZLz3x5gzXwCm3naDqCowASt8yFpwY8w7OgpruAfuzdHMg6wfq
HQx4pX8d139xZaXDZ6WkyI0rAbzuqSdVx8CzHmZC1+RUzYQmMLgLq+ojUPV6/ZpU
xLEz0CS2yNgaU5Wu/AvBpRQNqDlXE4Pek/kWpnq+jRlYw6NYcFH97etjG0QgmEIi
jQ+YUzxIHLmUe8AeQHpKDJeKzhir/c/h68hnZAR1jtDdtMb6VMKxjU6FNCOyEuWK
hdkmCbvkDWaMcyXPWqZI9tNq4w7ezTJSFm3V9WQcRhWyjlnQWJvky3k7bc0aw7I7
BYi1++/ukiITYNw/pu/8dBNDIXNOtM3swMc2C+H0g3lJTFpOr6jYbpPuMnjgfmEC
Li8psmqBVNryM4QjqsS5rXkf7w9p3EWLk83MVhcBc3B2BJn0sBQnWmOiS7/HmUpe
gzBKKxtH/3p9okaqvUfAV/xjnRzBWSGFHpefh7tx2GoQ70gfSTSDL+dzTvytBoWO
J4MXMJ0dcjKgS6BJ5Y2WJqnifcQjaZCJjZFjx2429Jo/ohprd8qMsQmOd2ZMmHHp
ii+PcJhcBO3M1feY7r1cEK94rJjS+zh0Sbyxl30q0lIM4sWGyNcHc0HFEJcO+DbB
oJwlrM8DCtY5WBq72pA5lcIQgK513wanOz48ZJZn5GEmzTt15efxBvk41IQs5g/n
6JbHwcHGMf0+GlBDqsF6eY8UQWBFPb5Apg3Z4ZKOCO/8S4z2a0vR4l9HtYTUQ8HQ
1KTnEc2mEBUJmcZ7Z9FJy6YSJjDN5nuLH60rrXPs9MzgfjYOUX1W1dQvQ98Iaxbt
SG3B5+exf42QXxbSrTA+pHQk/rTtx8BTGmeQtuBKrNBFruYWVaIvBxKVXoUAAUXp
MRQsheb2QsdBIKWnYk6egGvWyN/XH/PYKCOBgitlmjCujkUIxyc/H7Aa8SOprXPT
Skhv+IhmX+b+EXXVqHnqmXqxaAK80I+Cc6QBlqCvE9ETywGRHgXzk5A3lWx+PeCX
0ppg5zFws2Dzl65CHwaKc9zsZMg5OMFXNeRRasi77SYGlQUDCJvErqfKMrdr7Umn
rQLi9Epkjh/zj5qj5ub8vrAil5M8nysUAS7arbMP5Ku5t2jcVvA0V2+wzTjyNJrj
nZg4uh1U7DHGiiIbBb2rt7udmzLNwaGTnfob10wXfnuMTjL/SeqCuB9oVb/rP2Zj
RBghhw8MfICRxW96SlQLBuXcb0bxet2b9I54oBvtINTrz0ncVk8/gsJRTBQU2Smf
g+b4lbZSO+J5DeAFdapZj9LU0Zija4jwAiMFkCmtHZMMLVtHkezhie7Yp4bW1+KG
OPHEI6BXgS5sbg28Seh2rM5upEnT/gay1W/dAZpL+B/HnIULS8dZQH8Hq0P6CjGv
ZnrpU7l9DrHpwtINYg8h/NJzoUhu1P3RaT+A0pJfQZtGOKjyWjs35gSEIi+x0Zns
CsfcAIOvzxCMSmUB/yrt1lYoq3IXUkJHPuagWnncTMC8s6VsQOvUa1PSQxAP2MqJ
RTfKOiz1D40hZ8p9NLRMwpEJNuj9iZEltB2m0dFtiO2DVbe22G2z65MpfMYxBDD2
Kf/Js5x3g0M4HkDsWKjPZr7o6L5TRTiw7LmlFtbMzYD6vgLt7n8LmZnVOiGkZzUP
fyRhi8kyZw7TEdAAc6GstlQzZz1lZwMQUf65nSt1jA3xPpCECN3MAXRB0cYxS9lA
PMTCjZNONuz+h7pyHB6jZn7Yh8oTv6obgE3vtOPNP7mLCzRW6/B62WZElXPsXiqr
GOBTiUjSWGhMEo4wryW/6vLiEC00jW56TkLw6Nda/R1f2uvpLifOXWHiwJwRKEfd
T+bJT+mLpBcYhwuLnbfQpoogQ7egN9LSf3y4bPGu4yKMIaLHeJAtDWus53WdViid
L/4iJaAeqpWT9hdklf7djuBqyZRb93QiRivKCxL1aOM1b79RmbA04E1GiBncCfHj
+wi5dee3F/xwUi0/lRwOh2Hht97G/S3BgyblTNjf29tvFrNE4FxNnISpXsLiljav
C/Y/fC1SHJq0mbtBDwAkTzGZT6gTjX7qOCpTxveqqeJWIROFYEN8DQLOyXeDYo2C
XwLnFC6i9f83MaJJtkSJTGrzzP8/V0k9Qv1IpJFwgWZNeI8VtFAw3fXHgTUGGpH3
k9geuf17pUNhRxTn8y1FoOLShS127UENDKzetXIkweskoI4gogBdFLAe0vgiAy1e
4FIHUd6sy2em1Du/XZ86+fViZK1BSoxdvwbttTqe+Y7XjJIRsdfqdDJf4wZzb1Vx
8iNX23QA886qkKupOVaPzp24MIEz0q0+uHko57Vz8o2UjdPygCVxmG/FCHmMEish
qHCDUr3Ag8c+qKxgSNdLYsSKT9seLX35zEpm2BdmiPgoLf+dieVgU6lO4JFszh1c
tUCnGrOrwdgq7BB1enrKxl6jh4TNyNKIQ/8RodY5VfBjh/rTqxExKOR/N0MrAhI2
6EKeb1cvy2VEPf+9Wnug+Kdibmzl6WYSkznXXr1RaX+QqRfor3KLelqoB5vkPBil
0LP+oPMENz5dffD/04Nj2GE+ICUvnkgGUU9DlHp9WgabHGa3r20RQZhbmEr7uu6V
OxXQGKFIKpYXZbB4yUjiUeJckpzqYls/ZhRnh2YL+UHprIzriiHHNXISumQB+UZ6
2XOSrJmgB02zX1Nq0bAG01flf1pqbZmlPQ7T+b+AxBTHS2WnDx0nH7Fy290E5i2s
2O+MAFINKtB/amEspEYKAz9XYUfjcwSd7Q2vrlIfur2MHmgiI0Ll+bg9KYz+rHQv
lsuOvdEAFM2M0uVrueGbyL8Bc/KdpjChRESA+wPponrY39zg8sMRJzmaywyLtsR7
/tI79DRsI7Qi/oqVz8+elct6TIpsiHSuRUcItT0UgK3I5SiE4ioSo5HpncKEgC1t
cS4/y9C9bu4P0aha8Hs+HsRzjkp+02dalwFl0Tzne3uKsjRxKhwlpp356FLxgq/v
izHjVm0GX2n05W516nZUuuefgx/JscyAQHkWNW3HPOIqoGrwiyn8VeF/R5hJ7Yc1
2cZIJXfR3qpR2J+3c8PTaRBJo7lO28z29blbNkV+mqx1Wiw5OryK5Rc7Q8hpGMYp
xKPNoQTQx08stIhTouQyQhCRW2PRsJvyptMI+KhWXcX9yiaM6t1tXuBA9VNZ9+sE
acZxojt9zvRgJnOmgE/366HnmhNI9FFdTJu9cCCLuqUnk3oTVW70F4sqeo1eBT3d
fndMcNAax7VRvcejZEB19MrlCA4Ai2c8zrl2dc8bR+K04MaGecYrUPquehnbMf/I
cg59jcTzZReygsPSSntDGYOIxgICEt41eZqDI/S0Iq8933fX1vKif75g80Af08C7
mpAq1Jo3mUgetlEoRq218qWK30IFmklSxZFD+w80U4gQQh7xXiNvGlRTsgfSbiOc
y9ImQlOtqoUEpyXL1i6qfn/GsWF2M1ijTrc3TefmY44=
--pragma protect end_data_block
--pragma protect digest_block
/jTBWsdUIVpsqpfGpdjzDAgzgww=
--pragma protect end_digest_block
--pragma protect end_protected
