��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���d�v����0�i�=\��A��?��� (��1_B�f�	�Ѻ+|n��y��Q4�]�aY�����*2�y%����>��������K������ �
�D��z�z��C�y�B����
_�U��hkF<�~x�ܕ�cޞ���c��v�y�?k	?��m'�67@9%����-RF��g�ϒ���ީ��W��?+ �r��]h/4 �SU����d*�
�����1�d˂�b�V�f�P�(��-{�q��R�8��I�˴E��+RH3�A�`80Vm_�����a�+tӟ��X}�]�70Wj�����|�ު��#Ϫa�����m�A�)�[Qav]6K��}k.9��|{p�'
ʫ.�~�� �ج!�*���P�bC��E�c�Voyiҧ���R��h�m����d�ƹhu�g\@����}A�ٞ�����qw�t���4,�f��^w�\��}��#����bpi���V��{��a �����!l:,Ɩ_"�4�V�\��^�a@�����-�6;85y��S�Ę���Ҏ1#���m�;@�gǧ����]H��̍ �$�6�uq�6K�O9��{,z����#�n�k�A@Oү��R/�vV1��eYK�E�B����4�:���ҚMZ�Z؀�o�:>�|�6d�4��0�q7�/���g����@����Z��]��8k�V����.��SU/��Ǒo���t�������:�V1MB�S���Q��)�g��~�Y�q�K�rc=��?'B��wڜ{TP�b��^9Ya`�wr��m�>xAǖ1���9]�X𷩙o���"VZ+�;/�Gs���ӟ4�Q�Ⱦ��F���>ΟJ=9S&8oH������|(����ȗ�L�ډ��Ce��.�H��.��x�"d;��"��*����܎��*��Ȓy�~z�罭��C�"�N���?	���6P�{���|u��&D�ȃ�D����2x�����'�);1(�U6��z���J�]��ۨ͜G�ds
�V��SQ�B P? ��;h;5���%������JU5TԢͮ������բ@�����=��ɒ���S	-�u�i3�ss����:��ty����3Ulx���r��v���u�Z;d��M��W���Qv�l�����%�J��:��3"�o�Vbu~^�߇`����6U��\t$CAD�-�TN'Ѝ�6��_t
Gb���B ���F�p��Q5�`�H������k;�'�=o�\<��L��:-�x8����$�W(@����l�F��a4�tv�ѽgG�`
' ����%A����33\ƅF7���K �>U ��#��߭`�������䑢��N�h�����[ ��R�O<EМr�>�O�
�G��1�vl�2Z$j��53����Q���Q�A�vt|p¥s�9l4A��L���ݗ�O���.ZKt��`��SEA&��L���b��5u�KOΕ$������ƾ3�lR���D����]�ɤA]}��&����h���]	��7:��,.��ⱴ1��)�J0�Ŀ����S��
�������؍�:�ON�~��k�0��Ͻu{V&�_�"K��U���H9�	��}W+���'�g�VJ��YCy-�Khr 6�C�ZF&��뻻��`4��Ƣ��9h������L�s�!����́�)ٝo/P�ji�n��=.׀BY⣙'c_��=ce�l��f�]N�^Pr��X�kç���ذ��ɓe���=ਿ7��$r���/��#�a#���3,a��p�	e��ASS��Q���C�X	��g)�׻���5V?��"R��ˍ��S�rl�T������.2�.�'�zUu ˢ6`ȊnόH��u+��i;���.u.�Ga�vzN�s�ʑ�ꬑ��z~�K�����om� �g�ܚzǥ�H>��T/��d۝�dh~we7Y]93�Cu�z�N���bI��M�{�Y�hm��J$��f8�6[W!��
�EgO��[1�͟�
]>I�l��ԇ^�`�*h����!��ֱu�����(\��<��If��q���P���(��^~�q�J�;	�-�m�ː��p.l� �p�`aW�$���d�|�&5�AYK|�!#�v�ĢE����d���
5����9m�R��\9�!P2���Z�˾�+nLh�+)?�� �p��N��]��^?�+�[+�s��J(��n�$�+4��X�´��.�#�?+�MG��W��ϊS)d�F��ùMGi�m�u��#/���gm��G:�M\E�/�5MJ�Hh��n�#�F���$�������&ȧ����ܴL�����̖=]Zȟ��q��9� �����ݥ����X52-㐰����VOOH�r�c��@�4b+|0!�� H8�HZ`%Zw/9q	�}И2�D��m~o<-oO2C+��ڎ_���\�(�@D }a��&��I���C����-|2�)G\�ѫ8նr��0Jփ�|'��dR�)ߋ���u�������8q�p���m3[.����a'V��I�%l��[���a~2Vԙ{R�!���[�����'����Z��G@�;�?��k�|�����t{8L�ӜR,AS�^��m�w�*} ��zɎ�4H��UqCxc��Xd���l��Ä�̟kI�zJ�r�����6�%1R.;���rP�ĹV/��!�L�=������08�]�Y3r�йm��:���v�&-�sz�`j�lgv=KqV����t4=G5{��QJ��Y���oIu��du�U����_�m��D��[�"��42屔�s�sB�B���R�O�¬A/O�,�)5��g��,)�?G�*�ǅj�RL�0�Q���.?}e��$�|��Bl��,Ԫx��B
��h-�P�~A�4��3 �bC�R������`ƓS��`���٪.<�p:��~zB̏>;2��<�IUO�2k@�:�L(��� �W��ġvu:���Xo�52�-�;g0}BOFи��ћ1"b��|��K�5I�):X#�y8�CbU�>�����X$�L�Y��=	f�x��C�,
��a�\z;Df��7]T3L�R�ˋ�a
��`�r�������
�Ni!�E�4��l@��\g��T`�黲5w�	 p�#Wj���z9���j^�=�`�W]�<L�͍�Tsx�蓫�&�������0�<(�w�oY ���=�4wY�C�/hu_^^[A����n��M�����-���9�Et�n�1 -r�\Ce��U�jѶ��*���|���^�[iȃ2z0��(q�?��O�ﳡ�3^N�Yh����6���m���[���W\����Ⱥ��@\Oߔ�7p����-ؽ��V$���Kzފ��KN6�����S�;�����a)�㾴�J�,�?��
�ָ'���0�A~ց�15�Glf@�8�Nڍs�P�k��i�"��r���F��؈��˗�t|")o�\��/<۔�b�� ���a3�x���ё+�jk��}�<l�K�;AV���"�c6Cc`���{N�}HFS\g��	�G��g�jRi�J�^����7��g���l��@L,�UA(��UR�q?j��O:��w�s�ed��$��$�e�:L*�l��I�fϦO��I�,���P\8�\ {j�����s� �˾M�ݮ����;����w��r���un��F���
S��o�%��������W�G���A�����ܤ�`���vд�F�9(ogZ��[�˚�=Ń��#eٛ<��T@�B~8������)����A�l�<.�lts86��X������^E�����_���6�!^�6�O����x�@}T ��-6����P�_�cՒ��D����o.�JU8�݂�9'F����
]�6Ac|�uӤ��M��H��8�߷�c9�-���M���W>��H/j���Ԓl�4$���v��Ol�&g�t��*�7i:Zn���Nl�V�f�̺���͍���W�Rj@�Lܠ��� q0v�e���	��17R�Ҥ{_���fF:�DS�1�C��k�� ��[�n:ߔj�:Κ�!�;���u:���ܶלSu��##ˀ��n�����.=���t+v�<��r!-j>~�06�L�]��/&�Q`_V�.�x^��/}5�A� �04�x��9?f��ϒA��*3��D���ҹ�x���yO�xQ�pփm�/�1�]�_��|������3ƀgoY���PhN�p<2W��#��˼E?-I�7��6'�I����8�L��`\�ֶ`�G��`�h���A�Z�?[1�MZ�2��`%ҙ������a�X���sJ�VA=u�0��w�"��Pg��RP���ݙ��ޖ�7��d5Žg״jh�f�9pd�E𘲹���.U�D�WSer�ZhLd4)�W��3�Q.��Cg@dzH�g�~�E?F�����mܛ���w�WX쒐G^���Q�c-�iS)�g/d`�A}��
�����*@:c��©	_���`�U�g�r��9<�>""_v�0���\�1
�r��"+��j����mp@a�WS%:=�*�GApr`k����	��Kc���v���r+Ȣm�F7Y&�?�����f����Z*��tYE(k�1�.�ǹA���঻w #� V�¹6�"l?��5�������j	�?���!Ƨ�T8�HR�ɻ�iL�5�� 
%9��Q;�wt��>��1oR�	���˔o�x�t���C|+<]�'���1m�Z�����K�)�kK??��aQ�����͒�_qeֆz.੩����]�Q��=�,b��ZlEO3��n�=�dd%K�����:�hӞ]Ϫ� ��Ҥq$���x�����#@�L.����5�	�#�3�w���?s��I�	zN@٧�ؕ�ɚ�)���Le(z�	*�v���;�J���~t>z�^�Zl���r�Y�20q�A�[�B<����̒��nJ���Y���z��î;T��+�~�@���[��`	*F@�CTR�1���,��&Kc���y�}��E���C]�)�N�R3���4y�f;M��M��Po|�M-�2�Z/f�6�;�^a/ɂ�=�l�
���t{��f����c��o��ai �hGjl��SE婦��>�>X����y}x���j��p��\ji`�&�����,�"b�ʙ�&��t�5/Q�ld��酞"hͬ��.��X�:�Y�x������d��<m�����),\��1�?N*v5ap�6�΁,J����N��@dMHu|�xʐ���U�^d��b�$�����BW�;
�:6�q4��v�ghR�J��� ג_�:�bH�%�k�CaQ�/�CW�P�$�Q�M�,ىoΦ�����Dώ?N�����^w�rSbk�T��X�:�w�-a�l$��X�����{%�7�@Â>��Q��V,^�mӨ��$�U�p�hL��Dw���y9��#W�vy50<�S��ݑQJHW:��J��D#N�؍)X�Zo�
�m�Q��V���mD�l�k�I,�R�w&��{����~mw���vE�3,��	�)oL���Vb��ܬ�i�/CǬLl�}��3j7�U�Y�.��#O1Ǽ����4�к�u��j�Ţ�昄ܑB (��ܘ$P��&@N
�"ɉ*���I�{����^]��Bw��cv�BaO��s��+E��oX�U�' �%���5�ŅO%���.1wG-J��`��wh��tR�z��Z˷eT��IR��6�K�d��C����)���벡c[TT.��:'6���"^^�歓�@�I��yAu�����*����Up`��C��b�{ʺ}�o �1��|tsy�c��[���p�=}�t�Ǩ��*N]����*9-z�V�\��VoB�%f���M�c���-{�j���!���-�RV2���?URY�;=�dl)��s[�BY���.�S�u�_�U�d�3��(
��|���T����<�YQT�L`�^��&*���Y~Ѭ�:<��n��#��f$�F�}\h@,n>I�D!A5"���(;���S>�����9���S��FЪH}3L��u.��=Ьt���<�ZX��Sw6�}���g��}��^-�_5�4ouW�*\G�ߺ���i����:3 �*���	�=F����k�L�$q^e�B����-���T�H��7��ĩ��&���*#d��#'�o)�=��ћ��bKy1�|@�h���ߚa.u%O{u%�/P�����/ި���Ŗ\1/�c�]Q�0h;���{+UGH�R�����#{�X����^g:�o%>�*^��[ѭ�[��ɘ�<��?~S�)p-��%�b,)���ť����;<pE��I�(�!�/�5�Is�?�y�9f�Ԗ���������;���|{�y����9���7��b0��V�Sr+�bW�>p�qȕ�e��N=���zy��C���C�K�_�q$��ۮ�;�:��.��Lı�m�-9�W��'�r�����e7*�pj�:���@i�!;������ $�� @��3�v��������pk�ț$���j�XT�\{Ą��S����*��A�ws4؋&�Fn��׭��qW������2�ܐ���j���S�9��,N:I|��t�����OU���r�ӷ���Q��3kk�P����Y�YQ�QX,��
��&7�Rh]͗�#ISY�%��I#������+v�\k�"���XN��guτ�d�}�q�pb�!g���K���<�-��np�D'{1��beu���y|{�}�p����2�h���E܍��M��2am��	t��&*��i���: np�1�����n�}" JԔ����}r�~�rp�tѱ�=�-JA�PH�!���xK��G����:E�\�zO����~ٜr�f��^�=��:'�v�^ük8���ȷ����y<FГ�����:(KObj�@ɥ���ܧ9�`��?�RuiG�>��%r`�$���)J�]��E���t`�
�Ž��KZ�t c���u1��Pދ�ܮd���aio=���Tq̀�Up�V2d��hK��n��u��Nʻw�:��z>�����O�u^eIÀ���fD|�:�
��R���\��I�yg�|ckZ.��VF��n{�#>*{T����/���n�n5���L�S���U���z*g����{��þ(a�9�U6�>_���?ya�,I�ܼ�7PB�ϵs;=+��%V��'��P���|�����O�ɒ�����5v�HR~!�k����*�tĐP:dA���/m�%و�X۶�h��f�|dY;�꺦�����B����uxf\B�"d(]\v�Хi�O*�+�̩�kA���zSY�訏�ZN�в�������ژLքTp[*NE��Ī������!$�;�����8��,t�>�Oy��l߀h���׮v[�s�X6@�la3-^�EX��� ����"2�`&3Y&?�T����\���!�U��f�yM< ��b�T�rO��7�}Rˑ�1"���h�k:�$������8�Hwr�|Y���(��$����m<?��QmBȣKܓ\��R���#�?��Q�n �6�t?PV0�>�s q��}��>d����C��6�H�I��e�	�"Тs*�G5Ǭ� W�$]���K�>D�pS
bɠ�|Ɖ�7A�*_�wY�T8A�C�+,��@r��%,�Z.A�'x��O�Y��tDX��|�D6��&j{Y�oW�Omm�JrD�}|v�H#�����A�(dx�̀5�����֏@�̭+@�G�^�2��Np�6%P�@�X;�x;W������]���z��7u��/�z�4pY��:�δg��Q�D[�������T�~������l�CnO�,6�S�!�pb�j��7,ָ��BR�Tw�?�.bs�U���u\�b�׳�~r]>���EF�K޽QeeLc��b	���_�J��$_��.̻��ޔ�O,��6�����)��*ė�إ1r����~�.�<m�-JJ�$�_���U`*��`&]����s��z�Wdۜ��5�L�p@xH�����H|,�y�-�JjKŻr¶��9��Y*��b���di�X7���ћ�]
���3#��⭷�7�̱db��2j9����Iz�ETtS7&���.Du��p���� ��u��>^ZOt�^��E���Z2�� +J�0'�<?6���r:��;��j��P䍼Ŝ������v���F,N�Jr��	/ �U��)�ȥ����]���i�F���۫p���1��0*�} ���\�V N>���fTsm��R���7��1��[JtH|z�oZ�WI���7!��BJS�Bv����ϓ�D�Nnmԉ�s��5G��UX�#]���A�[�b'����Zĉ\ډ$aJ�ʐ���.�9d��tq%M�A���hR����1�hF��<���G�\�d��<A�z	�ԣ��6�l��yu�pF�C:A��+R_P�eF9m�"�>$$gp�wJ:a$��5����r�r�z��9W��.[�FiG¾�hV)J]'ӎ���ǌ?���6a�u�[߸uk���_X���"ˠ�X��9f��;����Fn���Z�ܣ[�͒3�J/�QM�r��E�;P�7M��;�-��I���3�g��"��QXd��B����H ����m������o(�-����e�idAIi�>���{��%������gd$�O�Wcf�!Ò|�)B���E�@*3J�m!�[�&�
��>�1}Iʂk���/�&��&۠l9�w�����J�p7�`�Zb�4�+����zcH��]0xj���hK)��Zh�wܛ�ɨ�o.�[11��L����^�ר֓Jt�&}�a}�?|7�5��
zzv
���l��a�.D���p�{�<mD�͔ʩ+�)}֡3�#�'F��t�G�k�s��$菃�ҐO�0��M�r@P�<���ѿ��N��D��#'O�u ���W@���Gg�w��܉��:zr����xԝK��u�8o�H�G�1g�>m!��0����d���w���%V��DnH�sŹ�c��o����c�1����r6����Jn ��_���P�~.qW���W{4So�+l���7U ��AJw ���� �鲪Q�nÔ��:��4}˭E~��8�ޖ�ۥ3�SN�mC�Y;��p��H�`a#���DⳞȚ$�B��X�5uA�*�`VTT��_�`�	�Qo{�R�OaB6���Β�Vm�v�0�"�� �Vz'�?�	7�%��|���}}��a3�M��!�^BwDfӺ彙N&�!�6��B�;^x���>�]@�.׎)[�@c���˙��םp�@�<K��`@O�n��&�JW'��0e�UoB�[2�$:eO&e�w��ْx�6�@X춊�9�a�R��/d��A�����p���C�N'�U���x��,y81E�b�q�ꛃ2�2+�ҍ,��A�,*'�Dc>�B���f6��q��^$[�P
i�Ď=���Cpl*�!�����8\���Q�q��M������gV�a8tp�������]&��7k?Ӂ�Wk��Q�I�>��(�L���:aoe��JE�z�\m`&_`LIm��#���>�� $h�L	�O�dʣK~��<�Y��h"!U�|�Ŵʮ�m�Շ�'ER��@��=�nH<N.-�Ŏ<��Wf�VM]��IE-�~�b;��󆬊I���.M�pE�1\����p9�i˱����b�Lo34ckE�eI��U2��́�Z�>̒w.YH���U/�󊋂�y�(�)��C�0U��8}~��L���Ds���:*���-�n��μ;�%�$F�Q��e��*M[���]��n�(��ȏ&��x,��0*"�Q�| �C����<�޼rcŊ��]���e}7m�"�A���x2\�}�_lO�ˤ�ҙ|&�Y��hґ	�χ�8���KS#ɳ���I��kؾ�⁧[�k���خֱ�{�!l;#-�|YƁ���m|3xd_7�6���y���N��n�.���_���,h�Md�n��ǝ�y�J��Q��{��^ِR,��!��	�i�X.!�����}O��e:��+\j<���Z��P��Q�t��(](d�-_VY3��=[�D2��ᆨ�7���n�*,)��=�Cz��^�g��>%�� {�Qe]�T�bj3�{ڳv��z�����V�e7�ǆD(hˠ�W�8ܜJ�V�~�/��Ra�(��]����hVf�C_�)��/�w�C��ޑZ��׻�������e[�J���qkW�n4�C�9�<�������2�!��+*rPc�Ϡp�� �����������Q&���I�P�9�䜤%+D������}��z|X���*���^D�N`�?)HP�96u��*"�B\J|���� R��H�Ȧ�p�Ɇ:��W�灻����lA1����|D5��.�<o����W���"生���̾=�V(A�yA{��XBJ�=��s� `\��z��p��(H>����k!�G>jTPtg�eH�^��N�u�|�.<@K�\�a��I����ѓC� ���+˖�����'��Z=�F^�������7L��+}���[��rKi�hg�)����bi���%�k�;"(�)R>h�H�s	�gMR�7 ��6?�9g���$e���Y&Y\DP)�.�=J�� �Hj	�☐��C�𲰿�2-��� �ٺ�-�tz�I������˧Q���`B;�	w�#&�`�0�z���������D�{��>4���7�a���K����
e��Ep��5>ڄ�T�#�3�AG[��;©
=y/���5��I�<��&���-��v�o0��'`��+�
չ5�#�P[�j�j�x{g�d>�|��Iỹg���ؿ6�d���il��?+��@�F�C!�F��T�L�KsS% ޡ4#�\�L���}v�մጵ�%�~<쏝ZP��U��,��ʛ�l��?=���!g�Hq���d'�=�(q��훟Lm4H�����x����ߖ�Qx$����IOPD M�l�9|�5�9*�nMLu�{��j�7۴uiM��X�B��;'�$�C����~]�Z�q7���,*po�A��4���Ԇ��t�-C���rko�F4���ڴuU�C�Ӯt�J���%�~d�}�������4}&��k��������TR�t���J�iٮ�{�ki��T����kq���:�����bjpP��pLh ��m�<�vdV���}����;V���j,�d|���C���P�w��a�ƥY��! +n5�@�[��1h�X�>���b�?7�`��{9{�`��`?�Lo���O����}yRY�\!�Q�{��� B��g�<ۧ|Cc
� �����0�t���=K6�~�l��*�&���i��z�!�(o;@��3��7�m�Uq�����C�-��_4s��PL5�w}-�N��-w����p��)��A��]�9�qP��֪m��2�G��� ��xjh�a1[�����~JqZ?�6��$����xFl���a�P��*�]u#9�/��U��Omh^&����a�_��L�7ɬs���������9Q��"f�,��Eƶm�������+h����P��l��ĔF�x��؈$���b6(�c��ʑ&�G��a4�C�����h�6^Ɯ$�^"J��9�W&��	�OL�g�q"��E%4�k$��U��a�-���]w��En�QB2�X���_n���NL9Mf;=So7(g�G��u��]�N�`����<`OW-^iȅ�8�p��yc4���j���%&�<�na�8[cA���������,UBm��7�`��"��5���zX�ä)��"�7�Q�/��������&���ɵ�C��O3�Q�-��/�~7C���}���7�=�z�E��%�M��:؁`�y%@�7r���ͪ�Y�d(gk�)�h���=m#Q��綩E�#��a"߬e�G��,��Q�rJ�"�̑*q���������>�+����/�?s�${��0k���ԉݑ��Z��h$�sS���
�=q.��v�T����J�a1Ϳ�RbP����;Je�v��ib���ޡ�!<,� ��}��k�i��~+6J1����S��ĽB�������W.d�\
�zC'�EroEM���n��wHd�l�q�%���t�@��I�u�n\�7�����2�����+{"�*��-�D��Ȝ����wl�xЕ=*�J�Μ���ޥ[ ��]����H�f2e*3?����i�V~!��d�y�������Ӯթ
- �It��@����� s��U���7�ȑ�_Pm _�^����	S϶B=ҶL�����Q���g�eE���s,������0�h����k����:��\g��_I>�#���y�t�>��-	�ȶ>����09�KG��$��YVQYk�>�f����n�}ț��YaZ����>=& ���8��*���_79��ܞ�1Q�qبPB~��Ӗw�sX�1wֶ:`�:��*
��K/	
�(0��������� �<}�ш���-�R��[7�����v�&-��A������!hOޅ0/�=�+2����>�����J(� 6cU����%¦��{�l/-;\������Zߘ��	���ɪ��=��Og��+t����>/�ާ��I ��#�E�Y�L�~x�S��ҳ-
�k#ZOC�f{�yQ�JR�^��ف�j+Rdή�̑}��.�sg�N`�z�b3������0�)�=m�&~"N��M`�<I!�Ԭ=sM[y|+�C+DFkg��5�2���O�o���K��W^�x,���|�2�0�&TG�h��>ݺ�q��G��z�9��.�Sd��m�F_"w3.�6l��jo�Ӷ�*?@�*S=�ħMObH?z�<8J� �S�3NT���S����Z&���UD7]�C�[5����0��V�U�0�#~�mј��2��,���۹=��t�KB��	��M��������d�pe�Y��_��J;��c<)��c#�p����)ꏕ��
i��~3AvD� V�}���w� �#]$�����E����1�� e]��`�ri�D���Ww�p�xj���Ӡd]�MϪ�ř����|�%���;<	#֪�=� eB��Z�]U>C���Noh��_!�ϻ���L�I�,\��@�ӂ�o����Dc%D��@��|��W������R�~������u
�s�b�v�����CTL)|$��~��541c�!�A���� �����q.l��p� �6$�2���"V�I����V���C�\�uR O�0;�����zm��]�Qx���8�2C�P��j�쓛��ӻ��ݤ��P���M�V�J"����p]񍦙f�	������4z«��Nׯ�B�X�`唙�F�>?�k���݉'"�R������g�����;ИqS�'{���CKՐR��1����|����4��w���l\�;�t�||�J�%��,��O2�RJ��d ���)?���-n@_3�]�T�}O���3,'�YYQ��14?Lx�{��?�Q�v1�����/)��K��ʔ��ВB+;v��/伾���?�b}�-y�_�o���s��Fl�He��w��� �ȴG�LZu�l_�Y܄U��ySWG�a# �7��6�q��p�D��ooY���̩?>{��/���h�*��-J��]�m��(��}F��[�"}�:7G�d�uI@�r��$1]��Cs�Eq�u�[.�cK˄�NK�d0@(!w�ά�V��,���-SEHA��41U�5m�i�eW
eo���\�}ֳxq�������a/��v���kT� � 4�N��/w��L�X7jOfR����e�nX�&Ts_�Ͻ������n������LmxZ(�N�u+,��t >��"^��i�%��bxI�!-��!�5��ӟ�d>!�$\a��D�X�%�&ɮ���rE1�[��^sۙ��T's���D'��vӄ�ͭb���E$����A}E�0�%�V-c1�,|h��o����_ow�A��1�$���	}��&��"5�:��%l���T:.�.��"C`�Tꫲ6�i�8�Ë��1;y�lm��н��R8	��6u?MB�b7ڶ�Z��7Dbn�KN�{ԗ�tI�3/�XA�j��Y?	��.+̍�uq/���6e������e����� L
{��Z	��8}�Yh�i�*�6�w�dMǉ�.`O�
u�e&)Bɨ%����K �FLj�*�ԃ�"7;�����%����s�(w�w��j��B� �.�Ab*U��nh8ZZ���	�W�O���XJm��;i.��[���7T]�G=�6H�O�N���Ə����<��cy�JX=�*�BdwT��	f�81Y�/�𦭵�jTF��y3I�.��t�ʇ�VL�;,@y��V���p�C��
���Dگ�&���&]���3�a�xr��Q���>�<Gs�4�{�PE<e��B >�_��|���DKT� �����0������6�ak��t���zmR�z]� 竎@�=�S�R�@��R� �q��P2��7E�.�����֏Ӎpx�e���@��I��"cp���?I��f����'��y�N%Ѽ}2'w��a�G*�ERP��47��KZ��b��o�nK���J�������Z򕺾�,#��	  ��J�1{*����`/Ie�O��Tj W�������RcC/L�_``ZK^޴܍Ӻ��Y�4��Qi�6�x����_� �Ԅv ��E���B�/�qfr4۟�?����wU�[�jv�����gc���>%���i���%���	!&cg�ϫ�@g��s�V��O[�2��A���� ���-n_V�&d���}gq;Q��kv��T������Ѝ$��[@-ّ�9��e�%wK�b\�
U����<�Ҋ��If��O��Z�3����u��}��`�o��ty�����Z@_�ɸ}��1�1��`�Y�������5��U`�e�J�|�1���;�E� DK�u������G��iG�݌��yC8�G�~��(pp�d�Ť�mk#�T��ߺE�d��A~��B�����V�d��?g�.S�t'��O'��W�k`U\�ǖ|�Ha<����e���_���py�HwS1P>�`�5���k�àK�)�5f��E������FUQSݦK�� �n�ق��}l�b}��&v`�����[��-�m��cT?85����T���4��lUm���)��L��j:�ym�`ضy��(�!_s��7�Mo"n1X���d�I�d����bMp~q���c��5J�S��-� �Vx@?>1�I��(�Y��I�GU���+Uu�C�ݰ�P����C�LB��[��M6�f
������*�!��_Լ��v0��+y��/?��nKN��7m���n4��ĸιI��*j�\��V�c�[&�:0 ��G5J7tƊ���讲��f�)�Ć��&.� ��B���Tĸ�<���hZE#�!c�juA��ˑ�
*x���@���o��
1���|����㍢�\�"��xԘ��)FS���>��U
���U �;��8Lu�z����ބ��8�����,���"$�hD��m΃^�r�ٙ�������KK%�$��a�/�d���4���3��Ƌ[�� ٚ<�0r��S	'�Y�>$�M�������xML�s�o��Ѽā��E��c	�V-5-�+A<U��1A2EjV�N����z�7M{�Q��5ʤt����#��."I �m���)5�U��eo����qD�,�Gݻ��o��d���S�������
�Y�>�	kJ ���!�'l~-�!u%R���p��A?y���s�a�hx�X���h���cz�}�� ��9t[��i�P�V`�M�
"��ay0r��bZ��͖�� �:�;dt(4�=+���1|�C!N�<��G�t���*BZ��,02��leW��o�J'|�%�X�ՙ�5�"J�`&�!��; ���Q��]PY6������G�����q���h2�Cq�`y�E�!��S��f�"���s�SsTij^Tg'�<u!7��9)breh��ʥ�s�h���5�J��k����0�����n�������Vl��u�{˶�n�=��:dqf��Q�M5+�s�:u�P|I��oգ�y�+�=%��2ɡ&�u�j��[�ւk8���a�%���f�]y���M_Tl
C}�괞��P�$���]3+7��z��l�y�h\��M���Ba��i5�C��Te��W��r�@h����~��S>���Y��i"��ۻ�'���y�W�ݰ.�;^2�zT\���Kޤi�����h��}��h���C�_�O���ln@��L�G��L���M�3 l�_�!�l��T]���;��6�3<�ɖ�LQ�����ũ�X9v���Y
*��&��鱫D�39|k��? t�˨w�v(B�}�-�?�K����@��k:S�75����I��16��P��;0��e�D"�uW:�.����5�j֋�C�^��2~���'U�I��c����8x����G�>�\X#n`��s�y��:���e�ܗs��/E� �L��;ڙ(b& �O	#6��J@���6t����x���~݁i �5"�?���;dJҶ��r���ށ���FR#���tjd���@��]��>:�\��'� ը����zrG2+Kʺ��SH<���R���)��č����E�j��2��s��e�lw5��Q��+0�G���jD^�� Ӣ|�O�zD��ֿ5ǬG�cB���[���)�k�N,h��� n���;�#'d�v�	]n}�[����$yK���Lx1�j��d2Z��0��+�{n}(Ǣ֦�c�6)Ɖ��:�"�wu�ѓ՚���:�[�X��I�q�n5��t�� �i�
(GP�9�z:"՝���v���VJ�ِD�K�ɷ%{<֨���Ņ�M�1�<�ֱ�Ao)T`�Up���	���2pJ' ��~�'�u�'C�.KGr̔��9Ì���p�Q2�,�߽���a� �og&�S�jK_��L!�	�$jk�p2���x��o&+ M���p��g_��#G��L+��/ݺN�:rk�)闝�q#��sYa�[� �&N���SR�ax��dzv�z�`�P�5����ZL���� 2w�<��X���^�J'�ZNjyX��ĢdA2�i��y��P�܅��t�����x��=hK�SA�dn� o��E���g"U�U��Ԛ��tbY;���pXլ�-}�Δ�)��L��+I���}��M�u�Mn�̊�J����4PK���@.��ڕeٽ3�f��R��'�)7�p]�����b��q����[_;�M�����,�����8���-�^9p�ɪD�%TT�AV�:��E�KĞ�
�yU�(`�����k��n1J�a�׻����ܽ�0�jr)9�UGZY[8u1� ��~��^�Q�,��v��߿�s�n#��7�%J��4_B���j�q?����"H��V�&U����Y�E�*a[v�(�{�46ME�fi�����el�+%C�6�{���w풧�������
�W�vZ.��#&������I�Gfd���۩eA���q����(�Ԍ�Pu��i��`�V+$|�yWN��WSڿ�֪=�B��k5�˺K('��b��D�J���K�٦�3ꯗ��D����b�D�>�����k��|���_S�2;f�'�t��Q%��peC��e�k�(�݌�{#��g���Lz$�˻vP��i�u�a:�i���iG��]�DD��ў��GD��_�JC�ut�Ikp%��8'{xД}��H�R�O��7C(^y�i�:�ӂ�i�P��b�q�h���~X[�bl�Od��cAPl��ZlIe�^ԄG�9O|D��*����z��E<e��-�l�ڔ�*=C��8�6V풐ˠT;`b*���p]��ҏ�=[��Z�3S�,U��*D�ñH��PBv�]U9%<~���}�P�҂r��7��3����C[e�=�x�b�_�p��Q��%��32�aT+�/��b4���j���8�U����Yع�z��W6j���W��z��d���E�����[�`�Pi#��TӇ@�Pϐ<��{����7�n��S���\V��NO��
�Z��#­�b�Գ:#�-��/_Y۷��G���gh�m�T/$I�ú�2�u�a��S���Yt 4>�����J��}-ӟ�S��屿��8�lZӄւ�K���dEb���R�����/��+���P���C]�l�g�`����E��.*J�(������iHt�h�>�E5���%�EN@����ô�U �����?��^گ3������|�6����b@a�p�0�iH��>�f� �I��9@ĝ���Xw���v�V���e0[?�֣��2��MI�Z��'�
���&G�lp�l���0$zߏ�g�^�8�ѩ�Q]�>�ҕeu��%J���ʚ��s��wi�D}x�̩�=z���:y1�gs� ��y��"�ߘ������0)�1��Cl�_��w�����
�ԳB�)-�� &�~�I����;kw�]B���G
��3���D���-���Y� "�f{@13p?��2"Ow����W�NB��\����y�A�>�jȵ��ֶJ����u����u=����\8'�z0�#��y;B"������r"�W<����w�Wo���yC _��ыsfZ��Uz^�+5�}�Zx��"~����@���jG�� �JvIU�_ɼǪE�FL�%��S�7��K��aU��@a�cB"��6�6�~Ӂy��qS����)�!�	}FF����l�J*��J��)���h~��[�Q�&k����	�Z� Y��e�H����⤲#�'0���zW�k��J�1O��?�u��jC*�x�m"[�	җ��r���댖)X��������vم
7%|��d[G"�P��=��Bq �4���u[��h�\��֓^P�_�ye���3���3nDx�� �A5����B�b���ҥe�J��զQ���g���/!����ݲ�\9D�y�'P��щ	�����&�0=�P�,j{�r���_/o:���R���<�J-t�:���*k��:~��� �n���»Qu(t��tjyc�4;���t`Tg���"����q�K�:׌g��6� ni���j�h1Ro��v��<�q-R$-MOA��*ޱ����3x�?y��ʈ��j4���=t��j�b��F2h�&�_J��j����W]���C�j��<9>G	�i8��.%�RT���Ȑ&��%!ED�"�4�~����%p�{�ʘ���sY��Z��H��G���S���ŧ^U��� 
�~�^���4z�����sZ�����l?���^Nb�c-���FB�6/���2	/���y����z���p��p�\���9���I(� �"$TB%j�^	�a����ݝRZں �\��,��~W��{�gm��W3Tmĉ
'��{!��f2�X#G_魘��Ư�#D^��{��7�'2i/�˙k~�h�Ҭ�:�`)���3��{�Mu�̪S�&@x�(�M�\��菭ذŲ���C�e(.l�C*�y�H�ʻ��V��[�+�q��|喇���BQ���Z�PÔ{��e��m���W�F����n�cl.��K�c��X\I:,i�NC4r=*y���������+�%W�W�I�wi���L-ʷ�GC�ՍY?|�"�ل��`!�N��'D�榶��|����(�:��ӗk�WgpC����m�����!��ʠ7*�$��;7eT\��-1�+PO�֋�݅�b�_���������=�a�(��j��D�f	��+�k�3�L,���Vf�.q:�y��W�D��}|��[|��/��H����f�PS��>zo��i����r���Uh�fM��J)8���EOy��%�}��kD�V�[j�t�JM�s�$�+@շ�ܻqmѺ�v�B����q�|��
Vl3N	�8_�9�/���P$Z�����Or���	 1�a�������>�~�uv��)������1�
�k�������.[���}<� XxD0�}a\iAs�2��OK�������o[S�R@���a����j ��}��Mo�����6�~n�[$M�c]e~������q�]A��'�ȯ>Iڍ��<jW�l!5[�]O��)���#�8~��n�v�dcb�^�����r"B�/�k�^��,W�s��%��A�K�TÃ������a�M[����xc�x���WDb��hS��t	�^��F��3T����5dh�����g��Yhj���#k|�C���/^.�Fd�������=u�ѷ/M^�/�����?�<q�m,�,+m��`MIi�����es#�Ro9�G�����!�z+�E'Ee���h���P(������UhW8���x�>u�V{�Ճ(�WkS�L��6)Fd2�ʻ��u�.��j;�����m(��P_����Nv�����JD�o�u�)�o���d���YFS�%G��(~Xڑ�Қ����\R����I4FYb1�L �	�b}�b���u�}<'��<_Cy0���ר�#6c?[����g�Zk(f-Co�º�,�nڵ�z�w�!"w���2m�J�ˇ}��83���h��s�+<�CV&���3����J�/�r��
E�T�-�@��������z	}8�&��N�]E�f�I#���Xu㞃�� �m����xN����\�HC��4I����þ4�u��-��U�A�����W����䁿���%�ba�)S)�ť��=�����y.*�J��D�t��4n��ą��!�Q��?T�C�r=�b�H���[{���4���e"��8�y���:E{Q��Z����܍���U����!�-Kv�=��&���-+��$e�3'%�f�K*\���6�lV��)����!���(��jN޿W������%�IG1�7	ʦ��
�n��7gȬ���05�?rb�gKnw�G�۰2:�����l����0�����p��̴��U���<%�j��נu���`cx�$��w�y����EU5�- Ii���?�63�-=�а�t�(��؛��ٛ��xK�o���1�9�I��Z��ge{���%�.q�����@�@ h\,�
H�6�K��5É����P���g��)���
��R�hX({�~��d`C:9N�y" ��ÏU��@�CؓĦ_͈���l�_���o�s�>0Α�X����<��(!2��4�d]��]��B�z���^��G��Ҩ4|p�5�7�#����š:"I�g+�$W).>r��@��URo'<�֤Vl���!�0��iNl@r!t2t~I�v�V�ښ�$�?z'���+ᆵ�g���TL$X�>�NӔ�Ƃ�p�kA~&e��T�l�Y���mSg�Q�5K�շ����'iZjS�}� *M����r�����+>�o��q�+htZ@2�Y�S�VW�Rٱ����teDV�mH ��
:kGg��5Z�S���B�s���f>o��w8^�����7�����}���]�߇�:&�y��0զ��{Ք�A�HQύG�O�Ý��a�M3�(�������K�Mq徚!�4 �MLog�Ɍ��z�d��~U�&`I7�1G(��^�������U57��o�X=)Y>��y��l�K�۲�۳Oۣ�)Y5]~d��*��K�J�]je)�o�(��bC��FIT�%�ќ�8:��<���e"��s�*�>Z%��KK �﭅���}�.Z����2�>?
�$*er18"��-_&�_H����=�ǚ�}���L�P�ޟP��C�x(�z	U`I��g�s3#w�_N�GŘB�A	N!��,�ɠ7SS���VLچ��u�#g��%���h=�ׯ:_3O���z���{\{
����J/���ѷ-.7o�R���$��ͽ3;����*����P����9B-��:t�#i�PmJ&�E�+�UY7��UÚ��P���PL|bB�C�Ý��^�T�N�1����P'Tܥ��:���U��t��@6���/��ƥ��=e���H����^8��]z>���Xg:��p�Z�������(}����
���WDJ��J��.����_3�+#��M�ģA��F�Yb	_+��L[���Ճ�
���iٍbT������܊`5ħ!��A��h;sX�*&��׻�O��t�=�m�{S{Q��?����*�M����O��
�Vo<m�c�t�[y9k��s��爵m��`n���"Ț�$��X?�m��i�g䞐���nZ��N�tQ��n+w��L�NY�w3�d��Vb�pg"�<��Y[��[�,4�/�0��nE��ZaT~Y}5/�o�f����1Yh^�"��G�-������.��C�'+md� �뚄�.�>t����w��.J:����3_Ml�q_�w�����z�Y��&֔�@� 🅶����7&��b�f��'��3t��ka�)�B/��bu��>�[e�=����D�Mi�u5�IEl;k�,OCk�a�	��/"��7��&�*�ho�O.�����ĩ0<.�!�²Z[��ҊS�ړ6�1H�e	C6�]��k��Y$��;P��Y�hٶ<��)I��&S��I#�E��s	��d�����?ߨ�5��u����h�gu�Dn�
�u�ۨ1:�h��@��Q���e!k���CVk�G���L��I�M��C>�i3:��'ҡx�L&b�`Y���َ5����Y��c0�ĸ}j�	��0Lb��������K׳���Ƴ��<ݗO�=�����,��8���u�����]	��1��DJ�xswtM��>�E/�e1�CF���0�~���]2�r�b�B�4����f2%j�(�RD�^E��^�2NoU6"�9��|:L�����߹T��^0�/�N�]z�>H�D�����������K��@X��b� �ګ�^:	��:iJ�?Xڒ��#g	�����y)�w�=ӭc�K����u����$!�d��H�%��U~U��%��l"�Jֲ�,����pY0�,%ig6�Ij�6�U*lt'֩_��Ajʃ��U
�>�i�L	���X��sCn�A�5��:�6��-ϖc�f�u|�\��I��⼬5pK��(j�3'�	^��A�T	&�Rc�	NC>��5ɣ�N����w������+�T-j�&�n�������W�A����I�