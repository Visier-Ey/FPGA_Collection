-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
E+EisLz1XROLl+EzDXir75YlKGIRDUCkqVKUo/JI6sjI80M5Z0+CmliAWfCKwBiP6Y/v29cvt9YF
luPz2Wl4MYU8a/v+vBSmju6/pc4YkfVt8zXXJLZP4ry1C0amR/JSwdMs4qOHR4jLX6L6j5IKrOf7
HMS0xSYW3zi38p/2wPQff9ps9ufv9ux4VBlxHp6WatCicUfxEXJcuesPUnOFYj+bthzaSW8mUszp
VmxTgFjDYWVQlsXEIYBGbIC+0mLXXzNpQ5oodhOtyqXdBnBrQUeOKgzKn1NlbfSRQv4uksOrFiyR
jsJx9QE7LdHh0RV6sKj8I+jiOh8Nv3/4LFpfew==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4192)
`protect data_block
U+J/u+7cnm7gS8xrm7EZ6xH9DFwi5n/3wchifI4TpZ4zTxZ1C67oyy4nh3c9sYzISMB7UC6Pvmvs
QbkvyZ017C8q9vJKwA8E4xxezIsxsWtpOFn6o/D53zfEZGyMeyBsDFue68JHNKN3lXknelUS/VKj
TKLf/21jkTN3vmEQ7LWey7WQPiUpv33iRjGSYYK53A+82Lurqw/2FjXfvpcuJcgvZVeT6GGi3qYz
dlEpSQJ83/OLMMZ3Bj65bV8B1YSw3Klg0eVUbp3a9EnmylgItmXOg0Geld5pDh/3oI6bn0EtnNLH
NbgUvavu893KMxBc/ox9fVuvzxXOwLmOHuGgRcmWG9hNUDd1lxCWMESp2tz258vvL6JDHotU+EgX
ZmUlXoYz+H1/+jQTRo0IU04dbefuxyTVUqHSMPs9tsWhm72f3dE+cS/67G41OsOYGBZth5i9uD5b
Zem0P0AsWcaNLXaAnX0kKVLJfd8ektkfbRnI00qdwMyvZTgKDUO59nPpn4+J0atDZvj3JbeIbOCy
/RUgUM2OxBuNiokup0EjUnTUaRnJVL3tfRHJP0mMcb0TYejB68yzy+Ko0WOgO6P7g95/+qGUeqqP
ogdL0Q04o6YVARIfcmH6XyH6Tv2p4b6Y03jGGLlvcAMBUeH5QuJWdXHChshHQvNo/Uc2doyHDOEK
mxl995nQYSy6RCX0wEJJeZJ0GgWrV5wtpTyNOJptrjDPHb4w1BasR3FH5nAtMT8rnQRX+ctKDVTM
7d6WFD0aO9sCvNNUQOB32tJMvJnzfv+8xx/SAqCsOfNkumDwRdsFQgcLr9Za4wKwodVe9McVZfLv
XQ5VKgq4dgGDgO8VA+38+KnRYDBJxj0/mKGMxlm5zw+B9UfqYd6Pl51qwfxddAFLXjxVkUN6F65/
+BGvMLiSa2Ruz/AX4qSkb9s9UJPc/KYhntfyd0dJYSjhtQmDsLtBEA7+apMOm5oo0vZzjqoFyjwP
GoFC9Xo4rD+Omuouw1k5n/hwiTu1nK7WhKS2NqoHOKoQQElCySvXSAD89YwAB20WAowPc4HL6vf9
PuDEoi1RO/Y4obQ3LFqJrLr3NzGBqRFwsiQVVwj5OjQPn/NHamNqG6LfME57NhwZ21R4RIVbHGx+
/k9JipS/IcJJzRZUry+oMkpYB8suTbqCR0L2dhAGme53BjTwAIA0YPBn+osnLngAy81wv5n7SiM+
sEVnTgOTKGwS7tvA1WZZrL+iGK4SF/HrITPBr7bI+VrgPNtsS+K+76UaoanuDe+RoWdjk4P2Bp/c
yEjL2GZ+me7VFYoJoEbUsAb722GeVHSDiJMU/zYW9OJ7p14b9T0edz4OZIfDOazSOejGfGn/rSOy
vYIPQjjy/zB1PnyXdcBaAFyWMKaoV43o/uHifCQCeLALfJBNHPwpUrYk2jaa1/2MCLS8R3PB2Os1
GQhtTEriVtYbG0Bab/kUvraM0C1dvMW54R82Vc/Qm13Zxk//Eo4qmkBzvBT+j9j2CtwQmEmgeUD8
z4mUboIILUjYsXU35AXXXHe5tuA3SIrHGDubWqM0nK2mvRvCQGxuPsdbadXiWUjnt1whJ5ddb2v7
m5eIL5KsBfUnj808DoIWtLUhqxlwDhTVLU1Fd2CJvC4f20kdqv02WpjzUbqSWaluOWa2XXuk8HXe
9ozvUx0GR3MhZl9LdEMHP7oZoIY/9QHnye2JFgWIl8DmzU5bA+azKWZFLRfKBElhpOltoAiG1xwA
6UieToi3rL7JtPqOjhm6F97lsMMIwXrfB5OTi8GoSPBY3CLZ5XmMX4VYNemGiP/uRsUKFeTFB7AO
Nl59ECsdZx0LQdrcxWbbayNTZU0QjZFB8Q/LWcGxAoVFPCidywpOTf5swhXmUcI8piW9kKWOmuU7
IOW2ZPrLinbeMiiLTT4+X3JTThwFwuqUDouGYGc/SKLSJdT0Jymau0uK3kpUa9Qiu8xirVg8ZIPN
uv3Oiw6tej8coeGWc4y8O8yzu8f7z/ysy8OIVpVA4h2OpuugwxXnRysmbh7YFZxca+xOxa/N0FKF
qI+JJIDsxO62/1PVZ6fU6saHcIO5a/ucrUgodU1abjZpIxZ6igVoKKifKwS6z0R6pFuzmcnmJqn7
Rg7u0CIsbjZnkWCt/TmumLHuZgwoU/26Vial8z2w2rGPXq5IBQNnlQw2TErs2hvaUnnfxVvU0WcU
OI14+IBbv5Au/8pQWlwgiNa+37OFNg5PA+Tjd5avEiXhQ5Nz9gSfcXhZWUx1/qXSkrcpRlqVLo7T
LVET716IH0TmemiZ8ANbWGudp/ru0bn6QqWRgTwVWLtB7xgKfIQOJAe1PufP91KbIAp3Nmbn5ub5
ak0FT6KMLsmGfoMjYNE5+EejD96Cmo3Mbr/6FE9VeT1W29P85fzgi6AzUoAt5Qe41paE8H2G6RGW
KdVSBED1YvZqnGte0TSOHIuLzhPEKwiLgmDlGJh1TYZfMilbNOygNujZb0qB81QvrKkKAELvd7Ye
7C36pmzckOsUboHA9x0647AbkE4ecvw8CtEUAbvBPvD1Bm7ER7mHUxe0fUwuQrxfyoI+vP9vrMED
dJCGNyi2EN8GRjbUI4pSo6hBD0/DmJFvaPPvtUYq+dOo2NllRoDMG4c+7fr0gXhWHYsXUzd+6K5R
SmklFc5fILJdtbEvdN0Zj4F4EAmu+hLj4OvzgR0Y+QcFtkH5mPDlS0TAtpJPtr9xt1yCxDwv1Nhs
GGCC2LNcLFvu+yq8BeMlZsi1Y+x0bl0K8vM5UGY4OKDUalDAMMLGe+0LXAQ8LyyMGYXtmakXj3ub
/h1n/37Jk0uSv3Wxrtg4uvi4d54VMT5yiOxwwf4UAH7gm3WTjLlTEP8F3Nne5Vn7RSKXTN0HUI0o
TWeqoPVaUZTeCneYakOq/8i0be+l3F5WE+35ScKhHKTbSO0SbBvf4YA8hxEc/oLJ47N0hG5Pajy2
x5WfAJVetE1ZzGUKTLCW6MO095fqVNAQSzJL1ZNQBG5UMxqqudwHyYMXCRE77fmzJFLaXV6XfQHB
B2O7fRv7OUy2pXAczZ0hRfhQTxbuCJh987jo41qv8SgpuWUGGLz6cWEw2aW40+FI1V36oS4ii4It
na2lG1j/iI7B0w8EhSZDM5BFZMI3JRMrboc8enClywqoCyhZIlJfBUTtut/5S2jDULX40UgxLobf
cVhaRZj7G08+JyUjyJGPA0sGdvB8nbTF+v/2F1lvskmLKiNwn5j+yB82CQwEUw/z8Ow+0aveb/xk
p5fQuGFAS0jmhzei/TFL1ZIeDx44szTbUUMWqXFEanE7rnSredp0SYb/o4B3gHvucKXI939inrYD
vpD6y5YN/W+vOqBeFDso63KQSeapEoK3MT6lOWt4DyVHh1v7LPpvr9jUanZEO74FIaGF56xHP2aX
htDQwKFVHuOW3VzXdzHsznncFhMHsK7ALKO5zz3YVV9jHG+U/nvkVI97OcE1qk+tgk9WtsVRtU8b
EPIb7xJHhJard6ty0w/8+N7Y5BpRF6CWCijIREPVQbv1hNgzTdbNjqwtN1CDabyY3PLgE84YaviW
qaLaotpaOmmuKRY7tj/bRL/QXhcDNFgHbsrE3li2MaeKh6gVXWMmwlwtjwryTD9vAxkwxiN+D3Xf
Gvhz59mqruVDkvWmGutnBDtEb0hI86V3KYTkg86fm+7BTFr9Ll9MBRiSCklX+fF1wUQCkgLF3VQq
cnKtCJ/z3wcCUZbNlrnRZSqDESxZy40HHwYwsOI4s54p3XedtbJaNxsuonMd3kx8SDobH9ch2ZxO
h5GLJrapq3E0ug686SFcjrjQoUEMnyfGVa+vamyhZyp18mWpQI5xcl2nyy8pqAd/dokCw3fJsaqx
GRWQr7BUlGjhDsvp/6acii/DaKLbbmBB0qKQfld94Tm3AJMb2Wse2r5W3iQ2SpxynJDL1+khuLdn
4B2qKij9OMRsqD1uzrvf9oguti/N1RZJMJd88/9gYOoridDTgEZyZyVsDvbpwG09tjVoOoz7GAQQ
dbNpraA/+xg1r0H25gE9yxkMB0AIlg2VXMB+gb9ayCXRxfi1J48Ju+rN2vSBkhnYcyI0m0vR8Iul
v3Jp6MbEK80QXWN6wn5wC9YHyoNqQPpHrFLx6C/nl8R10SYV35HuBSp5qlKK+eGRq4IMzmPpO6qi
AfAPu/mJ/0L4tRalxKT5+5bqVbQ0hRUEhDu1CLUVbKroDoRYU198EzU8k4hpVdKL+L1URnGydL4a
E1PWl4smRJm70Y0vdx0/ilCNInIpC+W7HiJC0mQUhUvBTcU+ov3/gCK/v0MNfpRkAC5TDCRLnKdY
KM6xJDeIoXibf21zP6OJJBVrAGBaH5w7BI/q0isGxB+cB2RcfmvkAqxZCCiXfc3WBqBGH7LusX3B
Y4A6Nv3m1fSrgUiC11FXN0dRJIkrEwa5lwLNWZDMF9vvZ2gNd/Zpesh9tLYDOB5UaDgtUXUu7v50
+9G5vyhWlUzBGTX4IDCTORRHNb4i65ar0YsXL5Yk50+M4aQo2X0bVZdpH1OBIkowg+LzdIU58djW
XiS1vnGAU12N7xdFRJSEad9luUIW2rgppNvZvp2fqwjTbBAWo57OSWfXcagNKcqIFyjN7u38wSBF
QcmcK7knAt3t5g1k6xOBME+1jF1WTCcMuzN9BxMfSGdqHkoa2Qr9aRftFT8EGyMxuLDDZWCcAmO9
1dxuRQxPeE3OBqNhaHuOoHGjCKf6qFAVhxAyTQlsgZ6eVihH4vME7/YB03a/RAO1lUSKTcdVt0qb
y4UZFhAQ+7LijTlGwy5+MGNF0vIBnMiejeAiP4jWcRNGgCch3vWyUpkOtJQtvhjXh7Y4a26koU6N
81bOyLcjfpY8uEb/cO/B7ZJIV/pwn0kXcKmCDZfLYwPWi7wU0c7WTvdRiV8AtlT3G+mF83c92w3o
03su2jIWmVLgdePAghkd646HGl4hM6XAXVFge6oPMUKmP4PmT2WuESSmPeo9T+DrU+XzG6NAa7N+
+RTycD7P9vsj2JzoFGT9vCG/ACPnLWVByP2GprF8nAJ6CklJLkPHAjmhytntDB57Wc3eY6WQd1Ut
T7VUgJozCq4uO9RK2mT8pDySHhlKKyHgCJvgnlhL1QRr7zLT1/ARw5totyOTufCpNzNm25CJ8GLi
H0WCry02iLHqPyPMcB2jdwUzrcJmIxlY3h4HnYhoZXHD0T6Xb6U3mPnMOyVt07c4IDppLl/vy03T
lBwsmz7QCgqrsNAcQj3Gk05Yky8XZXj5BUoBNKQ8vPwIeYrFN+KHmaRCgdEDMll7l1j8uWWHsYPH
tlztiL7DUm6X0prx1nyc/kJfQhnwnWmnDNV3WnidC4Cjj6/ju7XR+tDpCkpXx1Ay2m28rdxnaZgJ
SjEWyU2VmpaxSKlH9V1LNk+sHuuA9ZiMy4/e4fYiNrcZtZEURHDoOCteN4moxxgcjpcZzNg2F+1Y
REEVxE7aiQRhAg+UOUWaw6zcJxdM3lAIbSHFO3Xnta3z7JHmNTLFFmYxdusBNoqDOUVR9mLndJ85
xjT4W9MNw+mThCVdfL0ZY+XhlNVqDWATBwhgI7JmIQ==
`protect end_protected
