��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���d�v����0�i�=\��A��?��� (��1_B�f�	�Ѻ+|n��y��Q4�]�aY�����*2�y%����>��������K������ �
�D��z�z��C�y�B����
_�U��hkF<�~x�ܕ�c�
/�Ast+�t����h��'��2�C�P����d��K(t��F��2����(3󜑽�-L�_�6S���c�;i�L���P�0 m��2��x濚L��EM(����im+��_t�p�A��ѵ�ȍ~���s���<�y�-a�U�|x�X9�������˜�a3�7�0�-Bڻ!!.پwV��n�l6��j�k���h �})'9p0���/a�]<y+*9\{����٫.2enpm�F�z�	����t���Q;ȑ��1���z���/$�
����>5������������H%��q�*�ESl�C�D��������<t �U��
ȝ� ��؞h�og�S^��?(�����HS����P=$�>�<v���,�߃��b��NO��û���8 �ON�5Z�HY�J�|�]즕[�}�S2�K���!S��IK{?a�Nq����	�����[�T�$�VݷPE=���k���r}KelY|na ����m��9B��ƯӾU�shưa��E����w��à�{N�7�;��H;�u @��=:�ꖅC�_b
��z[=�1��8�ky/�����kW����S	#;��7�·��Y���c�$���&�Ş�@�Z1C�;lk�oȖ'*����]�c����l�qɯE^]�C,�T���k%��/I!+%�'J@t��D��p^H�qG{_���5@$��UݭL0jN!ѓf7r���fIL}
��E���h-<����ȱ,f������iM
UG+����;1|�%I�P���k�^9�йQ;E.�F�m��n^KR&�Qs��&� |����J1��$١��z�W\��-������V���X�V��e��ǒ��v�m8�?Vw뤃w�~��--r�8{*�@���i��,=�����G2T2XC��麰�)(IP�H�B2�:����̚�x�8�t��n����=E���b�m��^]�$��cа��6��6e~��R��X�]��< @��q�T�|�,x.:��?���ك㙖7�0�UIE/ҫ�<�j���9O'rz{vP�w|q��7���%^y��}K���J=	�e�L�T���Z���X���B���:����	�4��UEǷ&_�sMaH&U�g r�8��Sh�����:���dY\=�
\��,�JG�P�j���a~Gz�c��N��\�HwT����˛�`������^�a���L���	�_X��0��vp����z�``�{��Ԃ��%�7�S���vY�9�'z?"�b.��q�V3뗃`#��1�������������6�O7�<ML4�q�P���|��h+M�0d*� �
�ZgE>�)�|�ߪ7��˒��z��
�F��7њ��Sq����ݸ�����:p�Sӵ(��/МB�B��29K����z�Ve��R>x�E�Zi�')6��(���C$b#&S��x�#s��s�5/��ǹӷJ���a� *n��N�:�/��n���:�*��X<��B�O�N�RB(���|F�����*M��䭞Ɛ�^�N����Ns/�VV�ʊ���fW=�������#_�J��p���� s���I�w���ds�3�&�Gz�T̿=�Ku׿�6B�2���y����N
0�ToD�#)Vy�Մ"�|q/����9��O�o,��o�t�V�zZ����֣���R��S�`�R6������u�Ŵ[DLd|#�1?�����n^s�P8�-U���������Z���Ͽ��^q��#��t����l��a��	�=��{�Y.[�N29I��$����*�P��R�u4OJ�B�6���+�<��:=����g&3��	�ɐ�&-����W:����F��͋�3HC�ј�q���L���V9��;��P
q���sl~7g���&.z�Q|�Y�c�����4�;`%�1EN7V|��6t���x��E�SQn$�u��T�c��)�G�z�=��(��C�4��x��|n����I��{��J������,r�J��
_��V#C�'t�Xҟ��§�vM��:�J��vKh�1�#�Q��5���93mQ;������q�������������AI�V�NR���j����$Q
�<���Z0��@C�����8u��AH��\�V���];����1�<��9��2��9u}�(�y8�ϩX�Ic��I�pz��aD&�B֋�D����T��&d�	pZ*�9��܏-ޭk�A��%sh���n2�Zʒ`�����ʾ��q����8�����6�v�
�Ap��>�
���zd�� ���.��t�U'����E�����R�j�0��� �=��q숻�u�z����gK	�fx�ӒBڴ��S�^)�F���I�/���)�u�W��c�Su�.؋�W�o�Ngf���>��K�?���lKt��JeV�MLg����r05pMճu_>����p�߻��!��$��@�7�p9�~��\���S�����~�
��pӶ�����#�G�<�.7
��mĲ�5Ѷ�:+9Bje�8�����
ےN�I4}�^!N;��SٌJ��-��w�����xnrC��$j~O�z�L�0����ۏ�G��q�����b�:(�X�S{� Y�׎�	��

�>XL�Q�d�i�+��F�
�u��$� ��b��+�?�؍a���x]eЇ�vzm�E��5Q	�%^�tAZY�)�6k��3�"��e-������"+uxI0Ҕ6/Abt��!��y����� �<U�A�������/�v ��� ��O�3�Vp�$�z&��x�ʦAh/� 4�� ���M^:�C�]�>s'4��W-
,������P�Xo��~�?V2�&=�U芦�H���=�oݘ�L�'a�Ӎ��+�
]�]d 9�h�a������?U����ZĚ>z�i@B��`�����k��!�����׽M�/�}U�i�x6=�TFx�*Ԯ�O�� ���t���#Y��u�h���
1��Rŭ�y�rS-�{Pi�ՙ���k"!�˷v���^�إo�߅B���5�`��? �}.tB&�HZr����+�]�O�+�#��?�/�����aͲ�ۡ��%.^�0MJ��!Be����9;:͢��j���V8Z��uh��L1 �zAl�i�|Hjn��� 3����jxj��Ǻ��|�(�7J�j����x�\�jɡ� [�sv��:�i�Ѳ���3�5̃���0x�vb�K��0(�ZB���[����:������ i�|�e�eXM��9��yQ�9c /��N���g��9��R�v�
Ap(�NY�D�}b_d쓶uR������o�����ƍ40H5��:�jT�Wv��֨o���d��4C����e��W�'�n�#b���j馞u�v��ecIؓ߻��ʛ�����[ܨ91ȪV��اz6>:�� �CL���'�uf�Hu�b��{��j�Õs���2Y��(W���{yI�/�P�ַ��5:��+=��fO�5�2����D$(v��2�"��R �hS!)��i���`�?`��[�	/�I���UHb��M��ҕ�VDP�Kp��Xu��8��&3y�� -�q�ϚSQ�`�����ӿ����������8D%	��+��	qqC<V@#��C��z(6�x�!X��a�iJ.�_~㷰�&e���~_���@�i��>�o�ϸ��
e_�k
�wG�d���C�q�n
ќH9��E.x�9.t�I��]�)��x>���.o�ֺ�aݎ���s���(6yǦ@��2���1�,K 	*�g���J������	�Cr|I���ՕN���yu4L�誈�:��������x���D���x�Fo<K �?����S��-��]W�h���Y���w��w��i�#~����/pMg=�ӌ�Toل!�F?-����gG���Z<��>E�8�wy���	�N�A��ƃ����!p�l_ҽ'<��9��0��\xs�8qh"-,�e�Q,�(sh1�j� >)�	��S�����<����(aT�T�ꌉ)�m���I�7q���!�K|�'t�=01!�����s���(Ix��U��-\�;���3K��W��:-$���*щ�>���&l�A�A����zrR�c�������ą�m�� 0���� ��qE)@`O�L�	��v�-�ðm-*��P���cv�L�'���d�/D/�	c۰�5�}F�v`��z��th�9��vj@��"��}���1��PtxjN�j],������R�������|Z��3�W����N�$�Nn��;��9)l6s���!^j��
)����q�P�;�n���Z{�8�G
�]��-��x'
Ik���-��j�Fa��B10x��UbL1Q�w-T�r�r�K��嘗Dx	g�#wjeS�^�jJ���0�(�1粒tF�I�у߀�c�����=��ɱ�*�ًNw������'�`n*#uV �>oO���MB�����S�q���ʜ���	.�s�?�6�Ǚyx:�lXn����bD��v�Z�	��+Vy&I?��� �>����t#�nǵ����Z(NV���������n�B夼tf��)����>�u�w䂫M��C�M	A�L�6ye4F��$��Օ �Ly"�1,�P+'�`�V�)��;��{N�7)h�'J��9�V��	��)U�Rz��r�}���F	m� �X�(��V!?�����8Q�qgm�T����˱�Y�'(��@��˜P�r���N����(�toe�v\���6���[Z�����\�V3 �ǥ%����A�i����;�E�����M�\���߃�Y�NQZvz���^Ga��:�8�R��6Α��ˑ���BU������x���*��W�O�����L1�oKJS�+����B��Sp�����Ux���<:3G]`:���
�k��B��і��d�@ m�Q�O߳}6�Cem�=� \C�L�J����é���q�Ղ�su���c�KY8�e?���P�p|V�����X�eu���W�"g�i���X[�0�<������E��
�n8�_s���3���լ�H.�P��mv�@����u2�"|���{����^ֵr��j=�0���?c�F��+�Io�������Xt��U<��f�ݖЗm�1��/+s���PW�`!������ H0|���io�h���C�