-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
--pragma protect begin_protected
--pragma protect encrypt_agent="NCPROTECT"
--pragma protect encrypt_agent_info="Encrypted using API"
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
--pragma protect key_method=RSA
--pragma protect key_block
VsKMv9wsaBbshnT0hfhR8G1dOiPYjypsfFYkKuePZFOXXArkrzAiEKmG6hsmBBhI
qnH0ueokwy+aG6Gl17HQ2XAttVe7h5PGoQl1/O6+Bn4cWoNC+95pr0aVcboUUwD0
laMVDR94X6h2eUvFOZxkOFznI+6mDiyogXcVTzCa5IqOHaCXZbQi1FQJZmdC5cS6
Yd3VAfupsTMEd08umo17BjI0GntdWLnNCaPMQczAzLDwi49pKQZskhpHDmQPCSKn
UlANfgQf9gk4F3Wqqkqhd822gFjgMSvgxSq+gTvz9947gI/FkAHUUrO5XEXiFA4i
lirAaN/qufEAt27mwSnn5Q==
--pragma protect end_key_block
--pragma protect digest_block
iv7SNvwIWhKoH1rbyNaWt/XwZeM=
--pragma protect end_digest_block
--pragma protect data_block
4/AmLNixp45pV7GsbV9l9KluEFn7rEGn+Ae4u7JBLH0ChRMJtGx6AT+JHwVZgGve
+YSvwD2kmnuVNfb2fSf5WpNXQBfLjbZIbfsHdK00ozn0UnDpHycjgpyF1rQAuuzj
J6/earb18T5U532ulsOsNobD8MWAFIe5rsHv57N3x4lyGW1N+dYknxaljq0RhIRi
QhztnSBMsjnfg7rmOKKlH96YZqKpm3s2sct88nf1RcBB0ViOXvSNtOoTBOb+GlDD
AvPDXjEECTiPkAtzV05WJzq/d7Ly44SaOHsmZJdMEAgYNwARUdfzNe/0WfqeT+bf
IMiZ8EhKzaQ0XXQlzTFWM1tv6oNWb8+P7z/18Y+Lb+ONyOPAVBFADvDydJ9nStpi
SJ8ZSm0+sgjGB5abwY1SWdcgInKVULYQ7TIfqVFrQtVu9NXa/kfx5EpaKEtViwHW
BxlJa9Pr2cqOk/c1pRgtwMtAkgwEtlZ58NHbUhf7FZqZRw0j/NwON3GfB8oIJUo0
8AWGJrSsJNlAd9XWo1kPQpaXfMeWWk/dn7ND8gyBAZoIil3faAVcfeiWNm1f543+
Wz9mPkke9l4kvRySA/rDwjM7Ph+9QVKEebmstwXeCcA8+XwLmq+Am4qlVWJYVCQP
3LoqUT1+UbdwjMn4E9s2bzNj7m2gxH0pjsRcSiwTvDTtcCQ8ptanxAksTXfTRaMP
WZa8DvoxmzvPB0FAQWSS6slxiPgmeKZknyBUPCRZVomDHxbT82s/SN0iOoL4cklN
WMQZlLeQXD3s/qeHVmBrZolm0iJzybtEZcowFlA/PExG4ljvl2POz2a1Z7WJd2mN
hBPkJSOsBp52rld3OuQrHYj6BnfJm2euhXNpbznbHyfydl+Hpm9znnmWiKStrWWF
OLzAY6RHu/UVJ1EK3izUAv1ISdFBKkZQFIfr1FMu996HPEzbzbeorODIOpDEHVvA
pxdEUFMdt9Oo8QkbhKVCkTMhzi0NvMtfNptvSdFPrnSim+WlXN/Fn8QVv1IVk+GT
HrZqI6De0aIVLqHfTYQoVjXMoXpDT5FbFWN9CjRL1GlxLKRNxinoMfFNDg64HMu4
2TVs+NzJlDj+CUptEC9xRuAlWIAzv1uqeL6cUyGSRXX9Amo8XUhQ1lH4P+N10ANS
32ZjgCpehBIF4GYa9mjgiXD01v57bIKTT0nyezrbYjMU1y7XaDWUdMDoIyfmDgnn
+cMBLZzJQoilCD5jyURGmsddeXTU6lRObiyWrzbKPjVg6wJmofOmiIdTFfuTrbOj
SleWh9rbiFPqnB9MoCNOdZK5DVS/qkqeC4LaMw/pmMERSwRWLG8b0ElbbRu0HXzV
M1eifatAUgtqVMlaFJSVY95tKbIKGpNNGLvuiC9dIwWLZBOsOTr+Auxk/8bRKDy6
wDXSfz2TJpbHl0hrNgfbG6GYZuoFN+dDHfvl0Wr/uykXY+4HO4GATkEomKSi9fMX
nf8xjC5/WyoRtluEKQLuy6PomtKw5Xvr5UeGb61sAH2Ic1ny2xzUU88DaV5UL/x7
WcjPninX+hw4mxdVpXeZVaSVJzxeIDoLWrjS2WCKYsIvfaASXSGK7D5pnZN/3W2k
mKQVKnv0R0qABmBEzv86SA0oOVWBRgl3kG1BOLWL4BWoz0IgETEKX/5kSXo7kP0X
NJG9w0WvJV6umCPgwtre5Tm4XI4azAfOl5e3VrdUav2GYkR8HTTeGfoPd9IK2AkW
Ne+yQ1dC4E4UMyUKF9iX+f+Z01vvvNdY1jix1sB+jH1u6T9cCT73nLVlM9t/KYks
w5ZvSv5CFKMFYa1RN7m4LVdp2vtMbP6xToenti6wCpE4sIGCHXtv6djLwgs+Fc8f
PMrxZtf8TV0Bh0w5LQp8ZwSbkJlpq/Kc8EGTOaXLOsTC/fGobqu3x0Hb010sgFsU
gjf7bvcS2qxfunaooSzVevQfEAyJ5lQmlb7Xon9C4e/wsE+kKelvMj/GDRRwHcGA
059YdApqbJz8CHE0GuJN9T9k13W9yY1UEN/CEEfGVYbKzScKvVhmCeWMqCpAas69
gH6nJFyABUVt2RI19xyghTF6G4y4SHHrlDR1px2SLKHVmMGKVRHrSqXxB8XKGyHr
fK8YfaH7RN/CpRFe801Q3HMgJdc5vHDmYhaEUMUfh3Xlboa78seL7yfm/zUCoeQg
wVKO7XW1DUtBh2FQGMuJBpmlfw1PVKMb6R+CH2KInGlM9301LjvwbwY7aATe8qkP
x1y61IVZeCVPgY/loFnAmZAMM75jmmd9sDVmSam4cdJdURbQX1iR/X8HsLYwC4z1
P3fBodmmAZa+330zY3TiEJTf92tB35HBZvLrGUFUjfKc6rDYe49FI5daPfGEmUnr
rgZU+7WoxfmNr04dJLHKES4p9E/Vf3j25tmlhdZnd7XkeZtPJBJDc1IhFMqa0alI
nNJOwiACb4kRFqSC1nw101ySQhS880i2JnyxnFFU0hhKOusdwZMx3ypXbbIsrF4Y
xHe9ExIzxxEd4ybiSMk3BVL1Uird3EkOLx7BefdjjP6laBq2obvIIsoWiYAmyyWx
qKl7EJppBlS+JKrZDiK46izn1nCozfWSosARzttJgHoMp3ZKRhqoe/zyoZjQxkcb
KljEw1WCDKnhaUI5Kh4wOje136meTwrBL1qpU28A3u2wXA1JH15DY6uyQBHSXg1H
Q4h9ap0WyY9AILkuDVask8jqX2EPKLFPpLJc7x7y/vVKcWsD6FwrnjnD969mdZL3
CiEmPqx0bCtFP+jLgMn+9yACFiuxhR4pGHI4//YW2eqn7iOBdiHK41qAZAkZNyo0
9A+kqBUcdqnMA+qoDj9kZfFpj5Avowg5wYyYsT+AA6Pyn4Le4Ihfwx1dEI21R+0p
HJrnhbB4DvGBVZPjLE+hYnjn1am2INRmbC+7x7vlWNQ5MacQMgcupXVCLh5cVyCP
UAQxrgpAoJlV19SxaEPZGq/9VX71aKlvvTIckaRpXWgo9H/zbjEHGylh7KRiWWbu
IO2nUHeXr+5zHK+aC44tdhyQ4qaXfWvw+GoZasYsSiTfch/Nc3COY9wfxmxSFqAW
uGgzPmzqQARrlk2X7fCbYveCPilJ2sN/ihfQ0bTymqQ8skVun/iqRwxoGEiSb0A/
uvywoZw+KlgD2DmoIbwC3YSs1m0bxTfsmjlKfAzNru0gF8osdxRKoG2i0q0MZE/v
ebpLKTUUlLPZpE1nkx8Hhi+E2IfhycOAyBEQooDVugRaG+U1gvKEK/KVHhSD6JNi
koOZ0gszlW+LExD7SquvLFVqMgrKLqyIye2yz2QTYGW56ZCCjr7bglb1bjyErtr3
WBuOv0OXsvjf+jZSbv/f8vJVemYKwujubFEAIU5VU80YFN/vYYgqvMqt8fZVLEia
2IH/tzHYGYtQwJ+n8TzoZB5PHH9Fz1MuQjgNRq7dooXJwoo4amtT1LBXYU8UwN+C
cfIIueXqcgySz4QK1UduN9LCudGVirAqkvt3VBNobojjn1CZxESgRuxCClGWieR1
GMSdJoi7bMJKuRJ7N2nlfxMDuRPxMx9ndhSZ4WuTcICWXECQbR7T2ceIQCFmhWMO
ENstCm5yPzd4Nwz6gHI8y2reWTNGxNkiTUbLT2OpzONlQR+Ol4beL4F4ayRHyZV2
pCKN+T/3Si/7nMqRkAfm7I7U1EzT5h4d1RWpm/AhRwh3XtNDjcZh+9KsD+aFpApY
c5VLJTGxc0zGGEPjOGxTRWipbqfhZ9O+APDS/9n/rTapt9enAsYkO8Tzburqrx/F
Xq0R1vLbVlW5U5OHk863nCZBXQ5yh9eJIz9bzsgYnQkoouF3O4mD9XYj0BYjqNHi
1zv+PmodN8vxHVcIfPO0FJq9+bAPp3pIGoQHjCVgeW3bQG+l80zEOTueExIj84lf
EdO5V11UWzeATo5FGI6FrGe1C/3RIGCFgrZUw6yVxQB4cpz7ZYCMl3I8E/H03cji
4U+vphfx9imL5eD4yi3rO6/eVTPvGXtGb+CKALLjGPM3kZFyM+cOqXkN23g7hwLX
Z4qYHz1wpoVbk4tCwt6B2su7ugjj/7b5NwekdeNp3giP0k5p7yBsoamj9o34uf6t
KBMz9tCmbTdyhHQIiaawIC5Ip1htWVMhbJkw5qrkEcv84q5Y4daMa/ORHnXYUaeG
A+1ZiRk+xfmPNNHkS+MZ/lar15U47K9aq0StfuhebQdzs/84Hfb7+hOJo8S8WmFL
RgO0MLsf4wHzBSjdgU/n47rzYl3DFWD9u6bxHHj6ySadMZ0TdGPdhC7tAfSckdmX
y0DCFVN2vgbL43ng5ditCCwUbw0TjBjv9sHu3ekrer/+8JwXrJW3F/aWshfO/gpm
PSSdPNweHJyYlORpOM98nltvJL+f5rbPSaP8Bnx/dzY9CmlQt8FD2Nq2XSGiKtSK
FyCTQfHBkfV/JiM7TyCSTDkV6fwuAsP6wxYBL8lQc2z5QXDkfiEq6O9qIHg/XndD
t5NB5Mh1lc1hRCXNNAVumBl10sUk690tNNIBD1wArjWY7W3QIqjsNKPvj/uBO7h9
ykzzWjI5kMcRwqgTx+zaBmoTd72vxOyitt6qR88fkVYB6rB8PnZdRbJJyTKyGFB/
JcyP0vzU1Sj6yy2wQ8UmfQB5acW9o1EtwyfJqGJs0Pr2+xQ7tNxow0rT1jsLhGff
L5FTlrTyyTZEMy9euQomXI6GPVMLVgjESi1HyiEHClAnrxYmU5wYJ1q9xkFowNNl
7TOwaqIaHBFzQ+L1s4JVXgsoEY5+N/PdvWCneF+LLUsp9yurUcGHsAoD/rLzTpYx
SpExYrGontWippvf/QfZpXK2lwVovuFlJV7W3i2w4kuNGH6fB4cqSdCEArOkBag5
DUQJ8SakxQxHQwQinvtm85az3jYBS0TcMnEED/luYN4FxQebK+3zRpamIJY4j8jj
ttXI0DkXavM10USzF6m89Dr4mAQunlnjBB5qrFHQMI7FxBGrddbArt4WRDpGq0Lp
H2NWQx7cfTsyldD1WeqEADPc7NsrG2itd6MHHcMk45EOftvjfXGlVWxaiAW88LC2
HZvp40rU3S61ViChRHK6lnlg4+ImIjF9SwScli5WwMbP6bcv2soJ8KXRtv7d6wTO
BHSJPAYFt6T1hFTgtuieHntZ8u34J/uTvUqJGprRKBzC5kPkTqpP26ZB0xnKxbQO
urnuay+mapRalznITuMYvcyD2ExXU2WufPESZJNhea/GZ3Awxy0KvBDjpNPqkZlY
NpZH0JUmocmSleRdjx6L8taZf1yNkiquXHIncclhTjn5xWiDEnvsJFAyEj4KrXe1
ymgs5fLxsNAvgY2/HyBjKgytHWrbOLVp3Z4JVhZoRBFXvJn/NTLkcrn+jPEAF8ss
dtuN6YF6EGlX+tpeYWNbu+N5gNVQ9vt1r72pe+8vNHZ25041rkRq8bBDqglef11i
bDWfL/+aWm0tUevaGJfZ148IoPKJvqYPVMp1wAKFPJlpRP+vINWyVTfsBxHtgKrX
ILjAxhBr8VI/XBS/W4tH3QIcAfDlL0UobdzfYo1IQG9ax7gv48tnRQBC7jzCbdk5
NR5PKnoe9LY8gG8hA39pMx9T4cA7viy4zZXhfM+AnE82rP1y0uRPJ3HqnFonAUgG
gvAsgyAjbqDK/PpX4N/DWINGZjaasfBd6DObm+fhF1WDFKxKOyHbLf7giufaqxng
6Zq45vj6HXvsWWR5ccYMuLxVxtvCB1UaKiJgbn+3S7uu5TcpgJexh+XCyGot8zYT
bSjlawMLJOMlceMmR0fQDv48D3yWGZP+OxuKw8/f8xkbBqKfT0B7qC5IAwqZLgzO
+GJtJb3FznJ8a1AjjOuI4RqWhi/zRXEAwpOr9gypiHg8ouvLwiTsOIi2uWTiNd5y
RxKWAMVjVMhW+a+iA62VEHQut/ksucre2MFDALNnasabz6TrbOoWnEWcVODRJ5fg
G4oEHynOwkmvwSuRYwl4KgdfIqhi1amxRNGODc9Z/Q+QsK49Ihta1X9pzvEoSh4X
UCZSIpCdiDQymXlbegF/K1EVXI0v/f49CKY9m7kkheJ6BG7RzpXlMUaUQTq7x65D
80T4/VJrCJHShMV96JdMvMOYHyK2XeZo7/wHa1EpwsIi2KVe6pWTKZI+XLH91Rre
bg6MIEOmcyn846vUqb/ibbepEqfpgSxBCEiP38qbCQ+Y1SxMcrX8epMF6DUnY5w7
2pFcJ6W4e33veB5/b7JZ10EZCjGNYwKkJnb5Y0vTfg7uCfXxnMF6sc8cF9zYywm6
r0iMJEnLOYYH2NKTUehr9U5wV/CEJVhawHUzQh7jXmNTARyuRBcweEleccpBbHEo
pLs4vbMDmLR4VjuxnSOSM1W2OXjUQeZSjf52nLO7B+2U6FDdazfCQJG8bvoPN7XD
FW3wEcj5pd3IMq/Y2uzJniwjfWA2PxkVmpqo3fb4bW0hw50hk0MoX2TDG6INFrgH
4rJlMFQS7RGF+EURSFvqOg+6LicpqmzayTM0cF5IzokopqugjwM9HuyVNOYRefML
SxhdhdeYnebbSXwLlIVyYwIhIbfpQSzf0Qu6nKhUS2vmBjJF9vXHc/Lf0FZrX02b
I1oTjHMhsR0y4GUa8dFNJQMYOl1cDscDI5vrtG1hZlsnqkOWcY7r++BWBaqkdxo4
dEfURL3I1EDoGRSKfloZkUha9croRO6qIYV3XiT+N52CdVa41neJFCOzNBBVTVRS
EnMDqv7R0Xv6pHf1OSQP4aXVFkuIn4NnChPJWmkCNQTqcPHUWlv2tkquMHG4hkFI
kucLDho48cl41FFxkek2LuJGl7DWq2Y+b+aw8H5rRJNAbdjz4K8OvJyoRZhkrXD2
kc8dbkQ65PL/BkAGOTNSs0inDmFgJfcsN5K2gyGYSQCnOtQMECAUL+V7UGrYThwm
zxC+ToiBFuDqjfqkI1QwqFV+MRi3Fsu9FG+FCn8zMRxD1nj5yl674t1pgnjtl0j5
bsikGDoEbPbZ+FiYBSXrE1ITWaNs9zy1g+NMVzmhgnk74rHUUMe8cY0wqE4JsByN
h+826w1zAaxtv6nJOvrhfupB4pWO57qwlYPvmAoFmjmCJfhh9+3Kzxmg2/cJhrHv
gG1zMakry8sawQhh9ZZ5COrs4BPIDmJfHlDMa2qXb8WBKjyNlzmMEJKNiAOVKck6
lUHld9k6fhAnyPZLjmCIP5rPaBEg59rSo6VFxvgaJvYOQZMRzOoxS0Fh0HpzTs/T
v7Z/Yx8PZNRS+dirqyXKnhK+b65PXOcb4UvXliCtVFH477Hc/dTPRem6Lt5VKAvu
DdxYRGeuUBPsolOSN6rrMKEJ9cmG3FzsBrPHB6E415gidPwD2v/i6QFaXY/eZ51a
VR+JB8r0zxEP1yy9e0V10VK88yT0jVvyCSdZ3YttnO+Tmop0d1qRqYESC0WxyfPJ
yPpvLXEKMxEdk/kr5dF9MO9OUsnjtRhrf/25IT3dKdmoeEK+6xORqpsms528BC3u
lDxc/dgw7lVa/cSx6Jr6ouyXVYZ4Pf0tAS/Af8gnTDXV/F8BHc5AwNzjdHZB7gu6
wXWGKqdXCRZfI3ONPLcWIRYJhnfwfx4MvTeSY3xJCgJ8CzeocYIOzvLb6JYmpeSN
rRt0w103MBWf8iqn9WNIORuDBiIg7DKB+QdDTeRWADDsFGfJBl+fdcjkD7UgGL3y
lYdUjloB0T5R0+TrKb6SCfMxWB01zBpvl0KmlNXb4Aizykwzbre/WlMAAHBB8KmC
pylhZpIRH0jn5W5IAfwP7KkAxZfOJFhrldtUSLFOLiuCgafal4W5AYvExjjhvTD6
ElTUfjl6/mxt2fxhAAH4+acHeDDyJ05v9Sfz8J5LNuCw5w5DCI/K4fJDfTX9qmE+
gafnG9dl4X0nn/Mtn3V+3NSg2/vhJrcn5JcSLobC+USIQPYZszX7k1X3EE1xQJYx
fS68hyHFNrXua/xcp4Rtw9m2V49uHdWJbWGcFujlzI4vWh9zB0SVRjAvcX+hwIiL
IvRpBix8Hg18wzHL7KP2zV2NWlZoH4npNMBreDICIVkqPJTOFXOF+p0TbE5dj5oI
1CDjq4E8bmRg9K9E6XjPTTn83B1AkQMm7M5HstVMzphj93KiQIy+KwTXFCUsygtS
rKVwInQWj8DQ57oN+W+aOFxURzYrSD2/AgcXflEpzbl1pBhuO2wEMSII57aVLQhx
6t3H+ZSsF+4ZcaDgDCXg0ebMgrzQQEDy7JoBKv09mOR55Bg99WmRGybOJbABCf9P
6aD9dBXxp5iuGy9K6INd51gBlIRB/+SiePGCWJ40zPZKhKbSTzqaz7ETr2uZfQKJ
mbJ5jmWelSAwDGGxu7kZKoCEsNzbf9TMkVIiRMc+aQMtHMKtJeRgc1aIeDFjBmVo
fIt68zZLsV8uEAi/+ikd+GAmlt0/e8WMV6e0POcOulT9XNR8nrStAR4oMBNNe9Pb
V1lowVR1XFdFn3C2R8SN9uJ5h/SCAwuCXka684zoJhord/4uJJAnNoeD7Tc3+/j3
PVBOD4MBMYOaix9U54bBd94Qrpvf3u/oXhLwxoOssNt8HDbNix+Fgk225iNkJkNO
zPgbrc0GsN2kiVVywQlp8GXjD8E0rUUVmXwsu4Z/Uih6a3X/LgQqkfLwkJtsgA57
dkAoxNxf0lLnUheS+Z40TdRi13jsh0NskbxdDoYIzhPebhNcCkcvgbG2x5kuIaLx
GGfy7SWtYBdY8VdnGNfcoDtikUwN9K734DRrFGuQm5JwiCL6pxJclBYRpBYNXhCJ
fLHzC8DE3djxPrHAvZXvpOaVsH6J35obiV15WKmI++iJPOapKhZUEBxijdEd9kho
EcPM6hE7HC1vjdzFAJouQy7TCeOtjSffFy90ujVcd486vvutYbtTRgFIIn8skPy3
AvKx5q2tNmsZM9a7SjH/6S9fU6TdUVEE00JIAkdNyVF0aFGNpS2aSs0SEp0ADPym
lU0VI6HQxf6r9MNnb7DAloPgp3VQC10W/ZJpigtOK93DD0FXvwS3MYvSpbGn9mrZ
ZDk45WE+kgEKEmmcl6TlecfYAn/aI14hdoma3BhL4TbuYRxAvjcXWGdAYvdiTS5R
cNCdXUwUPdTZu8lvZl+ed45tNkMOIEVALIx7JAbDWfBNVtLWuxTOojgKxUpzVyRN
+icBsTJsVENcOjJ9qG+5IFrNhF13d7N2aopJhsrxDzt6990Pxm7NwXzMaK9EjB1y
0T0/x2XnCDx2U7+ZDbkr2CniqYlNE9vtK0OvN/H9W0ADSczk2CZE5CokYFAEPjoD
JHiKB2mfxMyulwfXsG1XMYT60QJU85krow+LigCaNXm48BPJ2mCFDzrYlI6bVN85
D+OnGsvIoRnF9NuBpPeOvjIQpZruGguyne3DJlUezoJ0hhYRPC1Dv0MNTCCyOYIc
Q+FlCSqV9Cpo/TCN+F2Oz59SBQAO/88VyXHTi6vd/OIUp8Ol5v4gXFZcnIjjVMCw
Y8gE601jLeIjIlyAxjGtcBCFZ55S2+YnD8Wk3joileP7MkgCOpRuwcIv22p/Mev6
SsOET7JOrY20n+lUZtVwBzwQ8wqmzOduLGlf4g8W/yuBmR13A1rLil01ewSmiKaM
nHpfoSzUA0VV1tYEW1xzBgLLOXkAfe7QPH71KEa04lT6nE0XmP0IpEtEj/erPr6N
kPMEhaA2QJI6rkD+jZajIx/29gsqS8bzOiiFJabKbwR3mz9E9U0PadK00S0TRuIL
M1xsdCRNg8Ih6L5aMPF4hF0uVRLxKae+KSB72pZtsqcOMheiC8yuHYNIWoR4w0BO
Ttr3bxEi1z24SMhEJ4N0YVVgXrx0x0pFOl8CVnZRPrWRYXLZ3Gcjpq7S+GxCLn6Q
Q8l1be+gSHjQ9BtSVp9ehHEfORCM8X9es2sOpXUPo1tLAfXMupVWQD6i6lPWaKbF
5z/9RHs2meavhzQulZIBfCuOpux5895tmZr4TLSXqxsMJ6pquYtmvrUHgjBn86yv
kB2ENkukdPl++2425pSYbrho98y2WRA+JlOmO3Rcvw0lIAltdo2cc+W8uMu/0Kyr
fOUzOdndgWl/3aL/rJ+H6wR4niv+dngb3i+rgJ4yoGQoghN93NKVGgmcU06F+20r
M4WX3oou0JRgZlc5lMP/xl3qw1T2mqoH/4qjBb0k7+nw40XdLx42TvQcHHnPOuJ/
WMA1n06/ki9icqJz8C9DMF1hBZ19W8eOtcQm9NAb3Mr3cvowyMm8ZZzeKO44V6jk
P4RJvZLyfLBV+imfkzHJ5kkC9u1VXvdkFcoPhiqERUVKX5NpJ8bjmi6ANjJ1igpM
9S3K/AaUiSjZZlCGIqxqS2ldpzZ075xdt2Rr2rO2+OdQo8ssUA9eY/DqcL/OW91w
j78wTdkeq4fEX15N11ILXWbyBCopduHucsbYa3j2mZ47uhnwxMXHUfk+qlGeD/Ca
dcyiQuiCpkFFk6v/mKlVgEc/9TjHErRhP+xfqd5PvKlTmR8NvmiMyd99lixiCphP
9M4or1i/PNzGEOYZlaaivXzg9DKHEGNjsNUqqM19zxoY4uLQ2yqZdTGFu8LDkGaz
rJdpJ+QI15yBDI6YOa7jlvgQn+GK1K1HBsPFFFCybxE/4ixLKnCtsGtgFAtuYRbW
BbXiwq0sEx/QXeWN79MQaVU5KyXjIgtGpar5d4DaevXDXsw9wVucc8P8YHMD2MwH
6dXx8ttA6q1QoV/10Nej854FpJDRQuxnDseFYEoH+FZGty1Z6mR/AyDaMwi6hGDx
6HKHJ/JWxml8n2cZKlRn1pexqM6+MKnSaV13Rf+cyxkvqjqOLXoDAkOZoxg2fJt4
R0PPDVKoQYs5HEZt614QULR0Gb63ra7tpsycfc6uejazAiX7+0pYCQxNQrRj2TfD
UbbbIr9m/o7Sb6tpQOKi4Nm7SJDllLm8ovTm9x7q/GtR1BYFrdgk0I00MwdUyEGy
gUcNlq5UQIEqpjcCxzzVCCirwTHEs7swdsqPBobAtcsVMZQyahst1xbvWajGJU14
qqyo6oO+CxFCTs2xtB3lwsZb6PrDTLh344/+5KHmrl7z24jmwiNsOTQ4ObAX4GNw
XS+a4O8gkeS7EtOOkms7klDx2ws4iOymgcjWZvw7j/jbQ3xjrAhVZIELmKUj87sJ
ouhJoTy7tR5RADSEwEzymKDC7FAm8qDkvCHnyfZJZiO70iT0BTHuH4eP9tDZqVMn
pS5n/D/rB1GpfdHu6ThPl6Avm5YIuXyNs93lEVjzNILAUaxWkrRLqYvdGcJiXu84
CT4NdU45ra2gXUSTYw6PnF9AkSAAUgmzF6iPlXaycGx40/OCZMC+/lb6wxSC+qVP
trua1Nco+45VUQMG9rsGOfvs0kE+8sxBNrLoidvEE2NHVXPYq/cgjSpCQgoUpV6R
v028LDZObMjmq58afNGO/ui4Ur9/3VxtpM8X6FemNLwzI7R2+LoHAeB4A4H0YA9z
5WWZbFI1qJ1iEWvPd4TCmmGuZj1zL9JZMtWUyo02s5q5TjUSgWkLaIXdArzCTlAs
1ld/a1Jvb8zrFQwqLtCyX7fJex9KZiptYu/P48eV84BnGQKP2ucIfq4FgJnBPJVE
OubEnOe1bJdY16cVRtBl5VsYKDgAvWAzDAy7hRJmEBjDG8rSTVP2Ej5Mlt+WqNPT
VjXNQKhMc2gFQU0TLXGPaIEinuqR+tp2GKLpa+0jBxuassP7BbNVXZ2Cg7tXqPgl
a+Rc12R76oFIhcJ8OQ+f5j5K8Difaj/r6zZKhVzKlyX9o7ghNACTtv6luLywsRtv
37f3JmLd1nVCX1/Ha6OkhuONHmkMeEI8+kfieuKgK8rW+8GgRe+se2BEbTGae0C0
EDsqhWeTkTnF7Apmc7J2xRFsetYySXAmo5Ghq+fL3CxPqp0hhn66swFM8xKLOZbx
DTFTBCQjRU9ddYTb1jhk7x29xVptQ/oHfGyNLmIyRIJnWN4LUtGaZYA16Jk2Kbnj
9ePaxMvi8CEtiVQZtaN6M1May3j0nihOI8SG3lUcF+tc7jfJ77C2eaEW41RVMe1Z
HjqYOZv5dBkdX+9L6/pciVZg/cllLoM8aBRz3SP6Bc+dYuLmBv9SQnYSyUR/JQuM
NDwm5gAvpZT4VoFEMrNPv3TcJJ2OVWNl+Z/h4vTOXGrXQD7eg1pSuryzP3ziExT6
pT9tGui1/sM97AkbsSzVLD9DibUv0STo8DIvPD5zPDHfLCYPHNo7c3ZNmDjmBPkA
7ohLlvHvV8JwANBAiEMYyFsbrsWSWS0DSOBBsq0/F8/oyFNwAfvjGZy+96GvdKXx
Ap9HE0z9QRPTcxvb52w6qgwuKpRJQ2cuMvJcbsjs8rVPZZJ3PbNXij2CJxHukLlt
0O9xvG/8SM17XQzksMosPTwH9NIqPUQgovP6ThEDFt5/ptERQ+V1pd3zt756Cp5u
Pr6ZpsysONAoOAiSCzMz13T9xX64sZzJ6xkbOhrdw/UoA17FYOkAbpgtoduTnB0x
tyrdf7Z6Se0RRaLGdDnoBwIFTRiJKsnK52MgnF6PVIg/Lo4T4/0gVjp+BGbvhG39
vQwFX05Dg7nPjlTCW21iQynOH0ZdQvSuGo+uG0AMlla2xtWxH8e9uH1kHrqPn5Z3
csW6OZ2erP05CE0vmjQQjkeOePrzkozJuOrCknPHQfn22J3XpoenUvlXKTo8kKng
kOGFfuAxnKHe5JzEqechMiB3ZECCSnlInhncJkQ/zZkT+G7S644KDF822/ZC2hxt
G6iI/c/NqS96TMwk7ZwdBiB095ZPbnvqMGXcjhk4z14lbDnp7IXeppEbxq86du4t
B+feXxPJk7kK8s5iz3dbTMQhSAs1YKwIxVnzuJHioi2igxNZaI7uaZZmOXdojPyQ
NhjddhlKn6zmk1JwaMDxV+pXl9W9p/c55SPM7jZb6HjWnmR8zzSwhLgHLEuuNuKC
loqPhTb44FdeEpcejO89RzYwAp4kIf1gE4rEAv47wGyiyWhtNQvGPNOsMFuih/iA
YGc1WpPpD59/7bwSeYsQUg/nPmIqWh0BgtYMLJ59uFPM2TJZNX/a6EA9BdfsSB8v
VY0FqHai5+4l21BsRarE+hxXxN6S3FKtxmamWuyuWJ52yUS+uZOtGB6phAMY6E+g
PC7GLXP1QfhzKu5FbdvGAHen6rPq/hnXe+5CCa0/biZNtUQByGKvtGq6Z6mUnwG+
UEZA/KxMQzThazN+tRcdULtzfGxPopVaI5jaURjZTOMFwMpLAb2wtaJekcRzijI/
8fKDZ1idOyRZoFiJ/Uwgs76xC1TSV0Dn+qd34TttnVH1kCEWMujH4XGGvcOmRb/r
BVNpqi+ETtQTVXZY5l/t2QKMDwY5b/pN9viffBjwR+j/JbrkwDC5mho8KeqNHgXK
xY8grwx217fWVhdaj4u7Ky6rNm/1tkWHiVWeu/ZtblJBySxE/oa3x6gjvfhT93Je
LBt4fL4uusp/6v+bc0uRpBKc3HD79bgPEsFCNb8J1Bm5RTjJzdl8eXydxxeHRZTV
9YGOSbyM3sntippLqVJe1In1w9EUh1wCtq1ZrACeYEPACU+Q6xMuGqJmwOOuhXQc
Wt+7JMvydOQHq/hcmKXbOE1W83KeUxuHVaATjyynWHDSSGK1C3oHw3Znjc7gqYP1
Orb6CWCr7RxoHKXOHwWT103bjrtqImqPF/9uSZL8f8euvQsowTGjx6HIvKNSvDo0
WoysPtZORgY7IeFmLOJKgTdhAAqsEWIym/cqPR+7KxeGZqi5tCxMw0jw6hG/TLjH
3xS6el7LAG3s/B3zRuBcZPUkxS0gxYIoVMnJ+k3jFHZbREdCJymUYhTsZ7nHbHgC
QofhT26dENF5PmSYDUEBF/yUxbBKHECtLYAN73Qn215CEz6XapujKC5bvyGKRaGp
ho6vsSxZM4H8mnQo/Ry1ql11eBGszom0ief4uTMSOnoJ264HElivS2hVHy4fulVH
TiSrYwTidEg6rrHgCkWvXrXFyXN9SuSZnF6y7ZiTEd+D4WSHOxSApf7zrkf++ZnD
lqPHyThdoursJGj7QpLae8Qmq1VNYZmAM+F19vVOEgGyKJPlSMCNcUKxhoMURqx+
2JrPYdnYuJmNtDPfirAq6daN4EsBFD5D8DitlgdoKcIeAB9bjkdGGawOPTglrIo6
1WML6Bye1U0Yaez90l5H7hNcbA48fy58KlDhEoUGfxwQtilG74+ZTYVXO/tcTe9p
fXYlND5FHF4ciy8wk9uLtHl27yrcWthjCD364foK1WcEqGKtjNRqXIKORkByH6w+
vATJmOA/R7lLzWg2rhwfQzNTnfLODrH9wd0wDJP24JotKwzNu6pr0B4V6Ithbfbh
rD+12QNHEmbuGQMehaovl/ZOZSjUPYWtKeOdGL8BQT41Jdfwl2/51YnetefohdBn
vn1AltMT9Q1gi4cdsS2qoXWxdBiTZv2w5aKqzfkU/T17q46pUWhlNJBNslvV/Ur2
uD9WbIRUiLrKtg4qsHVdHSH8hnUfRGFatw7JDnY55/IQDbkwzHMA3882ZzUDAbOt
WWSjpflgx23YoNWVWXW0lOttm+v87EYQUJhNjafb+r9g/a0NzPAjFJaEcU7GtXK8
/XpcyveEfOF2yngQvdSId9sAlvYmbut4TAx77b8osfqfYE7YwHjKx2PjJ9H1QbMM
AYAMQQbqTp77SkQtRawJUWEE4aNEpA82wrJj1JiCutsHRMpKxanFHI1BprTxRGqm
lVHCYnOhLytr6xllPS9OcjBNIFqaiIS0kJLLfPOwPoGrgphYGr6WJx7VxaVQ4o3h
KWZnxvGt6Rq6aB6cg7D00RX3mkOtXDXAJTjuowYBUWHUAmZEFZhR6TuuQ++cwteR
VmNaui7m8K5RE7A/VUTE9hcuvhX5WL5yTYbhX0tfZcmnL4UZ+4Rd+ONlxR43zQHO
j42KGQ4LHmI3zaZje5K2Nfrm6g7BT5xSWefCNuZ2WDmw9tJ4iDWnu0NmdKUkKsW7
Ain2SiYIzSSe0jTpJFqBQ8R46bLRmE9p5GbQ5oqJAVQbfbUy181EQ1ox5Ecz4wBB
rJUUjnZv75oyFL0gmDnW7TUawJKvul3dVoHtkyGJ+BCl12+94IzXu8yjagXG4KbF
GKQOJvtASfui/eZNMGSGmgUnFre47fWNyNIO7p9x70qRqWzcsipEFp1pBZArdTpt
heoe6ya4WsgLX3DkunEYJ920ubKY+yzDJePHVz4RW7isq3Ju1VnC6M11j/bP8TqE
Pr3pViMlx8qJI+qHufVGnU9iqJkaGB8Wav2tFQfptPfGLHnb9RyEAcGAfbLjLCkx
PLvi2P98FJquHURLzj9WntwgKMk3D2Oek1iKlb7ZbzIgMHx49kqJI2UnRERxDf+F
glvifM0p2Dr3BRsobLDWLRpQhHiPHBgAlTpEwQc4HkRD2fwXYjiyJDmWjm5kzhxW
BQS+QG9Jhi4ea/FnoolMjtmvs1ZxoUDqyLgr8fb5bGlmlg8m6iN98aZNv9fOqShU
P2Sz8Ya7FLZmd7LbjfCyqkbD/3Qxz5uidtGSqoykP900G7uoDXvKJIY/HMp367jc
EzzNXp55fY/hOEvNEI+HTMA+kU21SNnBJ2fMteXimzftg8dv+hv1Xe2dA5jcNacz
36Zfkwla64OBrDDDw9G/zj/AtYsSo+g5HSSsdiK8bbTroLy1PbU+R0TnodyY/f6t
XsS1AwzHs3raXdj9qt7A/18fImtkz+HZ6ICCUBgAZR7CEcUK3H4/Nsc8dUhcjsmr
lJAj9pcqDFG6kXHdvCI25k8kUhsfYWdmqpHk2dwnLE3tfxubQgytyFZtAVCHqtKC
OwVUQAUws1vrd8M5Sb79hRBGwDwPUolICndslFO1+Bwy/+f7uYiG67U5IV0VCyNs
RMS+k1B1TOnIxU3i5Et88C6Yigyt0chhK3HPJ7F1m1/Q0NohVleruiSJl+X6Xp9l
7CEedbq8iYrBZrAfRdpB3gvw9xyA5j30GnjvwxPTO6NkFcG9yWWt/RUQ3FzEtuj8
oYHnRRr59xU8LQnSa9N8qvAUk1cAWkVDWNc1GPifyRlnI7YS9N9nYuWfm+UDOVJK
b0Ltjr1TNEPkWVEI75Snp8tqZL/oTsQt9S/EpLkk3SDxLzrtDyaFUZ90VcnMNkVA
xUa8yr6zrq8Ls9nPlfm6KmSpAB58TKIawiEekcdMZaspcOl5vwUI0J4T0CfxYgmO
hY14Wwkh9TBQoZkTtlgXHp5UWVXM7BBoA7vyc58ZBdXEmey+Vbz/dfe77JdsbLm0
kEuyvWl+f16PuP3VLEgbR0TLohdDVVxQOgnSVP0sxPl6pJM68bKA3rvMo4mqQblb
ZJZq0O613g2CQwefTr1nU5j/y24PzuiTJZfMlstop2Horapp/+FEy9MrOQiTzRxr
YHC166ESQDA62ZpzTBi9TB1n/MtZZwaXJ2JRRWdJXzuoIirCqmnIcRC5dQWCbyuW
pzxWn1BFNV73FNWmXe6j8umUTPvhyKaFTPWad+brtkaWqhjXkz4m3I0HEUFvLDD1
5YFNwDsc4+J1yfPSHWLwU8jWfQDl/OpWXswlc7f1CQXj6MI+llGnE1yIIX4RUMmI
bTRZx/kt+keVt2plcKTmP1F4+IBugmoLkZQp27YLFsEbuQTJhzPsQRBpLNLuCsqk
o6GeyTI/mlsJ+xRj8mGlnzPDfK7VM1mLexaAkxAr4Syx1Gkk3IKexzu6uxis2KYm
jrU0JCoXDJ1/AR2rHxkpfFtdIepfgxr9/tXxaHqOelYG4lOv5qMgtyNQngt0x+6G
TySZbjOrfLhD0izJhqUREsBChX2+ganT/MU4rh+g/abelr8rZcwpMo5EF620U328
7C+j2Guz9H5wG2Sa0AUja6TCauizUjHnp+1bsG4wZrP9j0K3vIrUSiW29Z2bCevg
ag6T4ugFyHjGbMzPRNMQoOs9/tGab4TRiT7AXQ7ouBiJpmFqHoq0AcHYASj2vSUu
Juy99J2S2G4Y5J2zwEM4HK0sUNQFo1zoagDMUoqI4/yDG9jnD+Kk0GfbehE+fPGh
GgN19GxWfv9b7vKslLvRBjnUKllgb6DG/V3gNRS0JBRtms5rR5HBMudpExZ1FsXo
+Pg9tVNw2wpFArv5e2R+HVSxKB9mfsjI/+IEJO867Kzb5CD2qo+RJcJJ294F0Ent
3v3BVK0j4byggGmHPaZfvARDBvBoiXFFYzlkZyuy93+0bJKgqrGGau5OPN1qc8yA
7cI2VCPiKb40hm2Lk0bO4qgKHj3BNnPbMHns11sDrATmqte+/5Nof8HY1py6s6Zh
dagVZxq5oGs1xAAJ0n3ubffxZ4B9HuoZLUV6sflIrINxWw7Bcmc4B4DNr2nDwvne
pbO8pdR0z3Wa/f3pkwgzldfC1zE19BoQCfmKtY361yv3qf04KV2BuzHxIA3X5UhV
JSInsEd2vhl/CojWq3IPXj+TPs7R9MciECqhkOAaSAeiG/rAxa8GWPUGkJ4I9AvJ
4fFstQZ7D+fwlhBAmvH57XB2lQdPyMBduikyIhhPzjssf1Z9F3LGXa47IXWvOKEM
DPlHrBX3gbuJCJY0433RqlO0ZavxCVlFg817orHSwivz8AH7inGij0bX1U81nkzI
e2fYqD5jUl1eodf5ImXKNLUizN1/CL6Ovj55eu3d0GiURBTJWHB5tuj4V1GJZdSp
Um3fc7ym587xe/+F5hn1YP7jqcOxsTwUKtkE3t5R2kToNhfG2HAS0bUInwuagWOq
elEwad5GfCbdHj5GBD5OFNioe+OX5v3O6juNe4/74tAVOo17T0nMVNEkhMBhniaF
vf289yoa5RV33PlEeZkZQkB5P0GOhWaOobZz7GtBxhBVRrNS4zark2Z+XHrKXcv9
uuDqKvS3rFLuIz9lrYZuHKP90LyzushI/ZKsRwpf5l26DiCULFpYb2hvklpJ/tIh
ps8LvSHa0HLO/kLB5qM5H5FWYoy8ZWEVzssEDPd5/3vT7e1VMaamJHQhVMTuzTOb
sBMQZ7OYSg7i/np+ojNmgsR8/Lmtv9emDEs4gDQ/RI8dd4jM0gWF7RNltiSjaYhh
kEkNrDQjD09Hdcsp76OfikSZovIOt31pKalazwWEmpWG1AjZ/x6D+GRRty7Ils8Z
ChXEC/NJDvNYURYF7KuIDA766b3I77HCEBbe2G3WBrsw+n+4YTjporKcy9eH3j//
0J4Acb4/AUKAe9RYkZLydcmt7+SYZ3AEQhHdwmqo+AFMCjFM865yrGHEkynvi3Jt
D9FLbBc9OM1LCRxVyXJpl3mkstX3jWYyQFn1K3OcB220PAcEMSTTxl//GfT9TQ/c
ZWk3YXOTlhu98oSkyxl3q8NtoKsvJXtL86Q4fIZI2OxN3qGwnHAqkp7qj22XYetN
SeKX8Q/hTA0xrwtUIZTKN8z2GKh6djcrS28hHXLtp+ve4exckypX0VjD1ZFAvrWf
eaq+Yt0McsOcBiq29jbr2uUx62MATBjzjPcCr764qW0iZQweg3OGzwLuvpYTl0dt
lKsvpBXyndjjRRYTZs8xsMCQvCUUccQIw+LJFfs8Md5a6HJuUlbqRLx3fHEJA7Cl
dTSfjsUAUK5eishCchZjBom2J2Wr6sgRtzJwOao/xXyBKXK0C3i7yGfcsB6ToeLR
UCFZo25N5AbSYr/NtMkSLvLyk6uAOI/8xnRwMBi9Qt6/c8QOy+G7ur7zoNP3/l6P
y1+vQdK2qOJGzCgqQ3GsPL9HfnB7ErH70P/F3cl7ZZs9hb0Tzo2SZo56+rXPcRMa
EN2rFB1QEAh4KTHHO+1xiDGbAcUh7e8sjBtV88TRYJs7JmuIrpZCCbh/xLXaKLv6
UOS8RAJpYtPNLdkpQlJzCDt4r9BT8N2NLnZXlgL2J84KiuFhVTC6GkbyIHnhb5Ot
GzKGWZhRH4YntMiegxuDNR2nKVkFFMOymx9Qtbw1+Tsfhn3QJGFyisyW+5GK8YQ6
NlwVyU67LoPZOz4IJvc19jJXIZVLiCZeDbNCt57cBh0IcOBj2fQ2pCyItGYi/9Gc
D+k6YERVPCzSApRHRAHxwIfEXeCF5pKD52v8MKmpjh9+nQ3HrA5lv3wvX5ZkkZOD
rBEf1YpLPfu0ug1kelSv6Lo4AjH/joPG48W0QSqEn3gcZ6WLbT+al8xp9dF13elg
/TE/B9W29NhLReRRmmichfs8nhPfXJUNXP8NDF8AjqhHfL7ci/75ygMFWQdNNX64
hRXIRCMxu+sBYSENYReoc6ifzDWYu99cRWDzYWtFlPB4NCa7T9zqkA79xvFHVieu
b+dJlU8APg/2pRFpCnXkIF8/6NWM+BI50vkK2jKIWMrAgyke4akBmhshJQx1Pd5y
1YmXAC1MimiCVxRWzJF6O9q0+NyryHfSqzO50DFREDXIhRL1jvbRrPX/k0V9Vnvm
st5E/HowhW2hQaVTSdvkFmQaTu9u2NVCYPRjNvYYodmTfEuj/IX/q+SXhNIoZ3mh
pBiCbO42AMa7AHw/6W73Ja54NEu/o6tk7X4+4trFZRrelVzdE1DHEAXmiY4n27qc
scEIcvJM+F2rHt0wB+OfF1p4FHEJWJNA88RwJ6OdMjNLN+wG9c+FC+EDcUroR7T0
5K21zYJtJLMar0EIM9aUBrS1DKp7mJQ6IlzFEhovq7QB0jo93Yl2uMORphjitv02
khS5x66AdKGyOif09DVPogUSsL4qfVIdVTToJODhA8MBNuxh2nwpGXm9+6CgPdCq
KL+PX3zQ7JajHMiHXLYXb6BOBCN6zDG+To8k1KSN9tZIDbe+mBIsoQCWaOz1B9MC
c0qGHV1lPJScygmSlTJQS4AclqpXwj0+JSXEO/wab0WGjJOaIhu2LbIo+/1Z/HBE
TZjWRofhkLi/2mAJXjdkT6IbOFjt0lN1u2za701CuI8QYEpL/EXYy6BHIpqmJyId
9f+KbwHMltbyCgd+0PV16U+BDs0Xv8/hADyfYPsrF41E4nrA+C8gj2ST2GwlGq14
w+5UNDYK7OmnkutHX0vlE7CqNB0tcKyxjbdkdvGawZd1nJc0Hsgect6tTx4SX7mM
pXeMCJAEt0syL+YwT8hHFRcjyOxB7k3eA6bZPifcVuzBRkdoEnnNG1l2Xw5LFsBF
+4NxY76tBszTNqfivDvuiCCNjkkvsXLTPbL9HooK1nkKszYtDsD/8+35nSZKRVJL
IIDoGgpuIEEJkrhxS3l5xdXmBU0x1tosAp1UQ1/7V/nBT3KdmH4nQ6Y26VyceYaI
Bs5CNfpGqg76HrFr+bTuUP5I8+vJKoaZ+spn+73QosB4uJ/zvS7svtucT2YVBdo7
4PoHvnOVM4X10m2V9SFyd1zc6f/lqr7/TvjQkqLoSziXFJFmYJV3PzUrB6KADjvZ
ccfKfQ6AdZl5GASM+EfRwSJdqcqYkRpRl6njRwPJUNQ513SvXhidN0Mx2p0PDSXE
iRwqEFoz1c699Xt+QYZ11+g0dYFw2kIeWodlbMNO9Xq7JZMou1u9TsdIEQ01awCS
t7ldQrsM8wzGCBm3Sk2JpcxgmvQghI8A7t9VcVXiM6Z6sMtL92gW00+Qs/I6P0LZ
85dCmwxmoYnvVRXO3xmB8P7P202h6dT9jCMozfZb9ZWkh8L+jdnTaNj0Go6z7Rw0
dHKnzBpZHp/nCn/rDpoGVT1WVEYd4qSqV8SJgr/Dk30sIn/G9SJEx4oWT5q9He3Q
0GIsgKfxXJAPykfpWws7zbumXw/7vcuTWgl121rnUFtQbV1V9jeAM4m/m1zcXU0U
h5KbQ0LHpqRLAeUO3jEr/eWQJPDN4ZpPd9t7IzmEBCZtaKnXc2yeuMpAMoTHYlug
+xqKnfqkxu+azGOxuf3GijlrfIEbw8lqn8UXCZIuxhZbpCKnI6rK5AMMLkgrN/bJ
f5F45QOjc2duE1C+dH/0z4ynY0JALPxKax+5Ad5EYNrd87Ti0r+s3QAOz94HNVGY
1Zf/YCBig2tma9+t7TsM9n5gvAq7+wTga1LVr902Dv1MU2LjpEaWdMGHffwxhiq8
/o5zFFJ8wHC4Qbpy0iWupq0Qkdp1VgaWK7MH6zmgDYRxEfM4RlT/Qj7S045OekYC
ZpKFe1Ku/L276EzNQ2/nDqbtOmE3XkdB1uLoaTZVeQ70f5lEoaMz4plTDQEDctKd
w4RWzo3HGI/Ck5e8SeA0Em7vhltTHRwxzkDjIQlvddZYkUOxv8C7A6hDPfzKAcF+
0vcL/oco/bXJO8H433QS4tWlJnv5l605D5nf6vuaS35QAAu455BW/ft5bq21uuzH
dKlGPg7zNvBDKnI+7Fm2G+D4u23d6c/k/Uah6j2uXZq/VQwLRR2c+DJS8DsrEJn7
awBr1rTt7Qoex5E7dazH1k7OINGzloCfZ7ebzkf3XPXTCpsTXNQNeE0NlbcflFKj
Ky/TzlcnpeM6pEaBfmsaECuUmu5l2IOOh4T0nG9WNKnvKApgnRZrNIfIARhGl6i5
z/V9c5M+mWGwZU9jG+XO+MWOOrEbchAtLIHsXUA3OzzuI1YQ6xJ9H2Tiv7wVyY7t
3EKsgmRjBVGR7VGh0JSoKA5EjB/pwxxwY1ro+QzUWftnjuESsHeZStcdUTosCoVo
E2LNoTOXrZVXgf5tGc0hsm7w5oES9iMrzCTLBV93HVLTRz4VoAmb7aehkyLvf2a5
E3/vD3LuvAKGnXRCDNdVmlGaci5CLgaBqcwLALEyKPQcosXiq8Qv8S9vJmirXlnZ
KwHIeAGMd4ZXHRmOPNcfXfiOAx0nfmgMSu+T0IyGoCmJv4m1ktGg8Jpm6zQPP+/z
o2stIBZ1JHNW70S+aCMj/7HWnKDUp90yJQmeg1UsXuIp8OchRFZg7fX3IfwsezVi
JCYNGoNgAboPxoCTCQPM2YMuAD5pWDFyXF1vY0EmPRt1/MVN6sSLfrrzllBehKoB
yh33A5huPuw765NdmlF8NQUIkUqfFXaQlBWf314gUxZwO2TUq+8gL6+aXMTKAT1P
N29t1Le5CRwA5K28nF2W++ExTwdONRtMOR7YbB0UKXTG6g+Qqb9rHI7JEalDBkJL
w1pZHvKwHZPa0A8ex6AmoJfIvuN6Q0/UqVl267DszNZ0D+5f71V6yCZlMGpoo6pP
2+34/18aTGDYx4ws1tyM/bqSR0XtrIPiudyv7InxZQ8FvNv0UBcN3Abt8CT/2BJK
sDUt++68uJnOtOxcnpnKsH9edv70B5irODoRKFCaIdzhKS7zTMgchBs5ICCo3Uc2
DAbqAbN4075OYhmyvMc189Z+QJnwEleAGGytDSLJJkvo2ia0uLV8EJuIyuKM6TvS
D9Pa8LiH9TmlJyj0uWaKsR59PA9RP/qPTBqMk6cxL3rtZMMsa1K7SrIqf3pVhdZh
fPGOB/OOGNeTpftOjDSPMzT4MIdWrYaIg9GEVVjloeTtyrj9cFaWlgx13R8owQ2X
FQoLk1gWd9G3Zx4uNeD3vCHfl/syZpDm5aqlL66YQXa4mJe6ride6qNNTD6Ha3Yt
V/9OsFKQ/U5veEZ/GO7KYbZ6CxLEoU1XJOHi4/NsZSO+pJ/V3xgmlcmjuiWw1WwX
ba1LJU8fO0M/O23jmcZHU74x2Y0tS3+1KnPxDDjkXGFnyF9GDQ67dd4bNyWRPAEN
iHyJMu9gQRvPiFU4KnIY5c72BInB13nCOYhZElgR909eb1YfqaKzKmP1eURHxDko
QMo+oR8uMv5Kc8I8u2G17ZHZ4NWwuOxuHh+x+7VckHNezFsjj61Ul/sn1GBJqdNd
2JbEYqfhIQcLzpz7OniZRt8LQ1FtYxb8XMwmsS/Kh6NfN12FQyTVx71pPbdX0S28
V3DVSFaQYhV5o3UBfMU4RPHYF9D8F1eChFy3VsBxw293ozJvF++kxdU/9/eV8t2g
ctejJX+8RdspdQC5fY/ho2KJOkIEPthdG+sCNtsbkqDR9cJjo05FVJQYXw3WDKJz
yQZ0plvl9czIbkPkUMko/OyUslEPS8BDSjNhOoc3LEYqvaXRBbqqN3tS86VlEsbE
ilXrtu8Wy7yW7zBRAb9lftJaeED9dZ1mATQEpJScIaM1n+w2OCG0cJuCLCtp3sYI
ZHTmK5yZgMrAqjnoxD/tnW1eKhAR7ycxhMAYh7efXPPw2T3A43CJxPx8daAMQwbD
Gdl76bFGJqfNVSfqKAD8kuLL3Qstc10OgMG03zSEhU2OVzUFVQYUlgjrs2gJ1c5g
xQmPymTZJO2fBsqffjvMWharQHzETyh4kMu5Xkfk0YG7oznXJjLf2f14eDNP2N6U
rXcCFNqJQCUIAP+jqImlpXAdCKNWTLibVAhoujNTwtUCSbpa4jIhpFT/hmyrfOxZ
ZNLnWFyBqS0btCjvvdxIl4tobIGnwa4xLPa0TycBD9UEADhtaywu7QU5FSYhRWQ2
c+YI2v0wcAv6+mmqHeJ4fzOoUs7CN1qrXwHwK3i5QNza378LWl9mluEW+8uWisiy
IdMeTdcTQWJo1uixuW94GUpHUF6Yi6/ji44ljskFKaK8NVOXK2FgLizyQxsWhLKD
BI7+Uid089+rpavrgaMxkosjjzfi41sRsTBjed3YLg/+7a5FueYTOBK7a4CjADtc
Sx8v6oJpHUu21x+QJNP5KzlSZwv3VRW//jix1TdaV6tgXPHfd0cI5Qfa0uxofsF8
zfi+CJJaXNZdBXfy+HXYUxqATci1AWLZGP1MDXBNIjpiYAzueO1wnurN8J3ozFL+
WhCcGL8LzzlkSSkHKpCWsH6q6wUbgtexrKZgvUFg+RriYn4ga//IEfayaFi+mjGv
fR2wL9sfmlrMwJQLBk3f5AzudYlevtpGQMBJidCgaH+isu1vs+hm/7yxtsHVnnrT
joMDo5S2WIqTdWXrD+9wsUmDvGC2xU2MV1fkS8Kg7+tI2dsDQPpnBlYNlnR6l4Zy
ikCFlvM0vhYLpB+4ufqd2ozb8ZC04bzkWh1XHAGOWSnaE/mbLeSGmdNnMAlCu0Pn
CY2zL39HXR9iuF1T9uvGDJ/x3jjgk9cYrkEdjUnryL31smEO3jhuEVT18SpJA/Fc
RDd/BH3+xqKOY7+g0pTWjEibuzcAxFPYixs9qcbqVDqriTUSDNG47VlOkSH6A6c2
Bqk3KHNKN/IduDaczpUjlXAr+ItwupXWHKFmoLB+p9jZz7e9LaWS+1cpLUTmfddG
IAoASTw4UF5qXdSwudd/bvnnGby390K4eONBCJsnCeSWtaln/9NdVtZBDtb0GAs1
Ua1oKh42XrQc2+Ih50Jp+vF8yBkJbwMkYoruazpeGPxbikQL27xHJWDcK045HLWm
Lgyp7cUIzKyC0JpLd0qcQ1QHj2zhjkYW7PQbVYC2ekOcNaHQup7RmAVWvN1Eb586
8ujTUpY+ohKhrQQSEJB53AkJsgiqRrnTsmYOpl8ozipcr/QkeN8ybtAb/Szj+ZL5
HmKcXkC7QMkPMvUFcmnW01CRlEw/bnLD+4hVKg+fygaIjXA1II2Yp4noU8eK4Lbu
16BzHACdmeo9lUQUOBT6pD0vLuQksSyBiACOqcq14Jr6WQgNkjxKhgQ0SjKiQdu6
HSMyPcijXV7SnwPva6d1eV34TZl0c+jbVn40auPFgbBdPfeEmADCbmXfhn0tZvtc
Jo8GlDzMIe4VVE4V6REu2Um4bRXo9fzsUO7TGtocWF02vpXZumFES9p7DEbFTDGx
Q2ajK8rq+lrl8wTFh7GRauJuvHMv6SsM/bQ0hXHo/ChspFii+GbwRmGWAkXg9avd
rjqMlFfRp5fy56+bcFgHKUGM4XBbNJyp7zRIy6Cq9Mlz4fWkdlaSc0xD+gQ8KlDj
ldbnVMfaZkhO9BCCVJ32iFHQQCf/OZnTVnu7U8a9gZsq8+ZX6fMB6+aWZUpXwVWw
qTMvjWIwKedySZwUAyDyAMgZJEXHTNsS4Njxw3Kg69eOtaKYqAR42qnWIrdqZ+au
toIdLuwz5/mLv+23gtymnCV4W0b5TyjxkD5i8Brznt6Ki90ojXLx5xl/xBsLImJI
PGpoBxSmvVEjD3VlMRaolwNOtIO0dKs/Ct0m3FT56hq0/J+j0MwbaUMGyUAhSN9i
dWsF/6kFl0Ygi6aTXuqfdDYpxQDxktQNtiHQfgRUn5rsrsJIsJtPJnAVnhVNKs3q
vp9v9rO2ViYFJ8FxgvI2oGgqbkU+wHHY5RJ/7ju1gyfYRfWUJmsWzm3cgLRVgHPd
oDCVIUWmiT8n6d1a5RGdZ/4Pr0LwIDs+U2BF8UCBP70Vs/PS72+oPnFwySDMQLur
3P4A83TK+aH7uSBrHsCC8J8nW2ADzJc0bHP2NxbAIbmoLj6JmFCj/PoqRen1kOp8
6cVm3sGBH0Klnl2k37M1SEitFLC746AHTJEPYR5I8nplpJsA60kP1Y8K7hejSXpK
amyWBx8/L4hw2fmddu/3W9aGe3kKOaRgySexT7pOoGcyqzRqyUXWCgDL1HkRKrMY
AuRuElc7dOxJlUKJePKH9XEiI8zPNl6eTqbcKWERbTv7vDDS8EKYrSe/U5XfFeAL
wofSkZxFhxwPTMGIhATK5bB+UqeA7vXoXWfoYyAqQ+FyUKVijCOgZ25HbVGRn1V9
9ddXiptJh2nGGrOi8zCoLoyKQTm8AaFKhg+cE0PYaAxOIm2a0g3BbFq0MVOHb8tK
dybTyTmib83AdWzwGtJ08k/VqZ7Erj/aaiUb5pCI6teh6vabISi7Vbx6bIC5Ob2+
0+aqc96HMLq8KCkSskDowFZzSU0t0Vs7bt+6Hipg1zdyKfKqNDYz/AH4c/wCo7Bm
t7hDApA5RXzPog0bIOvPzlIrFi4l1l31EVIsLCaGBMGzrWypuTCVgVti/U/sPW6c
bQ4TGnBb09YEEk5T8UloKgP62swrbAI+2tFolFf8LwR1pEMdUJXUte6trNTYe5d9
+1KUbkhokuWzvtkMr5xDjyTTX7+tnTt6FbzlW722iavJH1HZCSRp0VO2DbLVmMOx
JU+nNXSeC01uXo31r09BcvgfLV4fpjWn1ZSdumVkarEqYTSkE3kB7qTTjehu2kpJ
vD8eFuRCC/stsyidDud72TZ9+78HKVUNE4Pm59E/27Ow+TQQgAwvoxaVSwbgrGu6
EhK/hRaHYZwV4y6d/s28zDq8ttUey7vjAIug+nS9Nw7R9Oeogpf/Q3NMoEpqbLzm
4j/9cn8IqKYjp0SM/F89l7iLeeFRgt8+mvaPTjQPJ8oBz2UMl3GkrzNS58GuiW+w
t+N/F1epBOR/sj29xnTrCcsllNww33GiH9BXa2NiEwlSgyPezJ0ADuzcxL9E5LLd
8zQ5T0kqv0yZqwHgLIYBoGDHu6X4dOqQQr3EQGGEZn5Npx/cXNo3X5/uUkWq4F4a
8BmNVAXeNwwP58pYqsrFUdLQsolaD5TVPUAf0RjaUxM/fjm2hmkJGea+Ifnd1+9W
/FO1OIU6/u/uDWO0qh4acwZmPyf3ZksNBRg4ME/4F/19QpwJlvW7uuRi8rNc2HZT
AvSwJsg32gIYElabPWVht1FPfI0ktVNBO4ubEYT9KkwCF4b7F6X0aIjp7l/XKnht
khb4b96xvKrOcwSDulMm0xee9Y6zW+9VWbAkfQ9emhRKIC4Ymman32AbxzLMhO4N
JRGhjUaS+YShQLtfvND8+4dbfF2iWeXWqUpLgnKPKxgbir866N8DlKAbmVZ4iPNI
599cCPRmOS6x5UUK4xeXZjxdG9JgGnCUZK1enk2nHoKPzv4dkYy4963LOvkxamP6
l47FRbb5WDM6OhGXaK7GjcqqWJHpolUOO6qq/GGSqi13UAxyl0QlmutoFhxdq5QL
vInXwzTpl4KwAGoFNo9fUz2nA6B1ncEEsoUih2FuxH/d11d0vy39J57W4vIxjaKf
rObidK8JRFYNRCp6blPWsL5etr2pcm5ZChH1WmZCq6LC59UkEIxaDy336cUc5tYy
k7PwdBpXYLMNvUJTW+FJa/XmDgXrlYJxh+Z86v8FW0qJhVHgLDbmV+bGPN+AT/xp
E0QmwgJDgERyOS5NmK3agpkcuyuSPPJ0ByCA/aVlh54L2VOBDfFknChlUpsXmzYD
mkPHDpWlGR6HoiXndEl7Vx/Jjl7bQsyeDYM/5EzFyldqsRnxayVSTBEMiCzJha6+
WUM2JVripJaRFlWFy59vV5r+3CtuyWy2EGyCvgaIjhv4sR/9KY+8tksKlCBuukSp
KVwh0X1W0/D7Zj5bzIpCRup18k6YFf57lI4uFfXLGGY2XwHS2MHGiVHtT1iF5rOj
lhvKndKwfTyYNfYaq3s93DnVuydyqehcmhGMRdrDQAj/YHM8SbJLA6FFxgYyCUqO
hiiqjfIUcEQGvGqWaF8UiMYllX6WFU1vJLKHyQdTzDpzCzObrKIkqL27invUGYCx
9S3503QjLM9hBxDO/F/aSfrPcoNUT1rSBOggBdBoyamOrpBuO9FoDEdvTMDgRhN6
uA3qai9zGTrnZiI2YXd46NGCAp5RZ4kXtHreMjd5voakTOGjYrja3yE+Loo/z+pY
amJgIecxuCiL8zHW6yJtK2HJ0S7xbsdM7iG6la1u7YSGeMqFZA68g0kJ2ji/wZbM
LLHIUmUtcSyUVIIHL6eydKIi1m8deDC2gJrDNih4HUgXXu/uFgbBZ2PDJTehj4Qc
mh9FmWdsA/3lWGgQnvgxYa/LAQJtTPqJqazfpOfiBwg87RIreOZUZEl3kEsqgK1V
GLhyc85wV+EepHHQHg5Tcex2S1emHsMfFuhExQzGYq3ljYtIsi6RnSEvPM14920T
7rGaCuCPKZrkPPjGWM2wsD+WS5FRSICHdV82nBEVp4R/jbD/N/hUPfoLlf/aNOMP
1iq8J7htkuKfTI6a1vaGKIaR0CtlpxDqFX51V2UtWEgYtpuLocC7lMAYCWcVdYJs
RSbMcyT3bbzSJ5MR3lX/a7TNC9Honk61aaW6VtrCb0G/N6y9jD+K1WF3uCBShAGJ
psk4FsQUgfWdV8iCVcaNP1i8qG7o54SEAnLDJz/Qz0ZXlWs3P0qVjOCYDdgwYd8V
uF85kNwCtfuVVrwz3rw1Eev4tEM0BpadCkI6yFvVoBYo60ys8ZwLzq2X9lWaIJel
2JssjMT6bF1cNGoEMBienY0Vhi0MRUe9oshID1QTs0DKJs4BfkW2Ate6GDUoTAeA
ru4efdky3umiiA94HycTpYoKEvAxVzVlQSVRusuulCVNdc5h1y3fBuN8/ijRi+CD
cHl5WrXLcthGGTHipS0SGsQTgiy2vLEb36svj8KJRVB/ysaULzfnES+0EASs69y/
WC+n1nUtkAywqzdo6Shb3YZX2bUKP9+jqoqdjOFnGUogGGASPcqfrdMxAQNVh1zS
l2SsDYTpMedEbD4V4g5Lqm03rP+jXerELrqeRmci3aYlf9+HAL1JrTAondgrUxGC
a8ATbu5krrjIEHd+VRg++0fzgJ7Au9DtjBlt7wWHEnqaG1AUk8Rom4AMrdiqZvzw
oO59/8hYEmYyv0gJxd4xZgy7uYylADnRXq7gf9PVh9A5zH4j4jhJEZ0wyY5JfJLS
axrt6UZKP3gsSCTza3UZ8tqoM/n70rdoo1efjQNus1X6mkiZdtnFZ0MfNqBVjD//
9Jod4qowy582PEKqKE8ANjaLQh9y6U86pHhzpD7w5FrDOM3pa7pU6+LX6nRAnRLk
0yuzilaXAzqvmdH5wHlL5Fzd4KWVcP/woSpNraiSW0z/iwsS1fbin1ccxoFEGYCb
RtKADl3dJ0nTEwg7y7DL5muB8VjGBSllaEIMg12bueUxszy+l96CksaSnMgxRWgJ
wTk6/yfyFvjom/bLTd8jnDWVi4NZTrY5NIo6ImLdDJAEZlp1/4Q0B2a9RrD/wVVw
sAORVQK0gJHxngr08IFnV6MrqX3Vrdm5UGnoq/5HjCcavHKivsE94ZFX9WfUbTcD
MnLSQTmgrEtZB2m5HFkKk/i7p8FwEI2Fv6UWQ72N7L5hlKwqGssJy64pRlVIiZ8y
8tW0cBDgtIYcPSd3FOhqvzmDPiGIogG0kA/JXnfns6K+nIxA6Z0WG6KogWT5oWRg
3C/Yp6bQbbUZ3A3yssFZN+oMslf9PFc4iTRpIeIwvDLf2J6uV9qh/qYZhK9aCctL
xdyLgZkwFVPzzc53Tx1EQDs5zaN54TRGjjXEW+CINMB88Agqmt0tBbjOIMzQDDTV
VHXOTxd6iUvsD1tlIzpnNtljTUqPCNQkis6dxrqzp4Ksl8JXN9D7RMOfp7hw7+vC
uoeyZP4L/IXKEsyPLk42MN0wUXKgMV6RFfPUil8qfShbYSNMgu4u7mWmHVYCU4Qp
PgtynXHzvTJTz9SnR8z3Gypl4o+O2dGT8yE4jhqNj8vYqfQiSlhEPVvTEEQJ3WpR
40BSkb96/9NlqBOY5FS1unb3/t1sOHH2SQtWRppH+4gx/KDQHi3dL+irFUAXvM5O
0n9QGupUbMsMAXJVSOlwyL9AbCQXz7xhKVaCse4wQRDXA1ZELLbgr3VBr016Ln+J
TrMiVCWbhpqqX5tVjufFlIFO0gMhQdN4qnxgZHhMxSjjzWZf6NhWWd6kwf5SblrA
dVoW5DDbq8XeQM/xFuK8cvNDmluRAYuOClD7j+26JCCNnOOwcZqHew+nBcs4MhPj
QlykSJUh6pNV91bGr92ykyK/QQI6X/cG7AcRbrdtCEBCLYRz8HYmFBgS0C4zYAb6
2AOPLtwdjsVFRH5g10wHTxxvEXsY5wJ/pWX7FQY5XC2NCae1Hye9A4Imt/HqZycW
wadS+QWbAUAHHjmJ3/uBnbJl9wYy4ySKFd6DnEy7X0yhZuii7cOPF/blku6h9qhO
kS4o/StI+mg3RGqJMy8NtdcT3nWnoAf9Zb3LNNsgILYIh5pU69ZWsJGYMBilyPwi
TXrrkhd50MRxgunzqXs5c9GxVPm136gvcYzOR7b9RV3CWXK1TBN0SbwWKWHgiM78
eS9QcTwyvB9lxx0d5l7vQ5HLYnvNjPoEJ6XqCa+t24oH0WdWQ3q3+yB7n/WdbEiy
NRLrqQirFmgQV67lxGhTaFowa+M7AB2Ng3uZToSDfUgbL/bU60eso1IDouHw7N5x
gfKRMtk3w6AiOOVA99l1v04FP/whuGwhrfTb2NcAxi95TZ96bfzZbZLQYj0M8dZZ
evYMklA8z0I+VgnGpGebcNm+cFcz6ZrNGUVyXaTKXHG6VoqqOKv7RzdyUbCHTnNC
I6c+dSUsErqNRRs2xMAfXhZjjsJyWG2MnUBEVrOLyHrVl5mnfNlmUt8L5w+ncc9L
bt0UjFOMmr1Ob5WQgWfE2oAvPUy3CPQrpxMgzjGm9bUGZjPNVMMzjIBjTBa56tBh
xhU874reC0AixPvd+6yXaGZWahhRETvJweLryXo7DSQI0GME3rLqY45E+zC6ZBx9
+IWuGnwC5TWWbkafiG4iC7MG6Hv34IDYWpkQrb+Ab9BMzmSS+DBpHCCdUJhqQYPw
LxKlp+EDolqOjBxkWY8dYMBiHt7+y3m8jZ53iyUK9CclnUYGsZDg5jFArdgewShk
U/w0llnnLd+qUicX9KhhJZV6T+1VI5hwi8XUL2HrCs8jiCY5heUYTyUYXyh5prHX
xhcyY20iPTAeg1pLCp0FTVyT8WZHBE+Kw4Go1+SWoZ/eglMYjUdAZMWW5uXA9sIr
ueU5zT/j8vkbfV/c7w7qJdO2FOPGutSM/z7XCbb01pvwOdxw7aPXJooQaJH9MFvO
3sDCpSwcQfLBXLkkNfmKxYNUb/8/6I0BKksBmLX1ivsmdzfZOXkUTkpLnXSkVfbb
rzQ6/EMa7hamp6Dtvj/X3jR8XdPj4cDfkyv+XYgu1UlYnfh30ru/7xC65Tti4oZY
iTEq5b1DTDQEjAqbxlVfk2pUo2ts8RBXkTNPnfpCt+aZ05A6NBWLVPMbhT1sQeXY
tzuNLor8j03I9zWCebuvXzcZbChv0ck41RIH4iaPIsc+fRbj7+C35cWAgs86mH84
mQceZc6r5n/oPXL00yDElMX5JdWg4+WCWy6nii+e+aZXcvdObG1IO8XxTOpB/amF
RCvEqPL5cZZmZ9sm8kEZMnj5/F7WSfYNFicTenI6YxLXOMmM7i2D+p4WaMURBW1r
49r1LU5FsEpLGMi/HVe17gxwkqE8iUH7VBT/ee4W4dgpUzmsx65IDfuM74i262ZC
nOiljRf594uG+wgssVgxJ6NLNFTDhhk61UFEdV59CTJeNhDyWRR9h2ZmJu4e6mfk
vT8tZ9p3rSRY9vTi6dzoLILtxmLb0wrdycKOSVHXotF9aouiCuDQH66INyRvwFOj
GJXCH+GvwXfH+cTYcXplj7txcJTd2bMrJt2QcZeYkpRf5QNGGuiegGOQ8n+ZCVoW
6t+IlYD97OIf5urFdha1FJPbPcLsW6Xh/sxwYQo+khzlY3gdG2P8MOA+lDfVBlde
dMhx+tDC7GdaiBp796L/4eXRtZZtfUuSnWvA+TNMXMhtRxrF2pVmOQr3Ul+ULSFb
3Hp/oeYWJcsEwG5xryRI9dYlCpaMDe4a2mRrOoF94k++CiohikwUQgg4jDFxxLUl
A9t9PGtvFc3gBwJk74MfskzurbeCypmucPcnx1Xx1zqhdNrb5X7ZIIF/KFI6PiZZ
kQwqsHegpv4OMiI4EvYs5tGXpf50IGJg9n1AtFmqstAq9uIabBMhH4jpiKOELneE
e9LZzhHzFkVFH3S1e6+uhuIHMF7j0WEGQq2jnRZLWuL/jjl5/zPrmR+KDYjSCfzQ
JTPHAqa9ilXyc7V3NG9T8N82kZkqWRxQFx0ugMZ5J/auJ4J4Ti+TM2ybSV4lL1yR
ihSvfnYP9uoQBCzk3h1Mll4bAt6/lLfTeSy83zCrNFjIb5bZL8WaGOzleycu0BCO
AHDHZ4xDbRWjASKS+tv7OqaUKsfWG0KBVxXvcDyX9aZKEZUzn1kgT9fPJ52HukFA
Eu5SpDVAIU5AGTRfPNa4GBbA/tkUAzHCU0irN0SjyW3+OaCglH6vF2oMlphnsyDg
+pz3SY9ZsHLhLrF1lQb7xsjWhqNSsbziKxCxFHtRIEhGRy9aY2O1BKMB+B0Yp99q
6LE6hQzV9DFeCdcZApxcUkAEIVPoT5v3aAsAjZwtuwGXa0dmyGQqZocvj54CyzbJ
DqacK4DI+JEWcVt7Hr9w2XK8OIPLFR7YuBpXeE6LvTjoUbEwmXTuI2VQ3WN5RBb3
QXPL6AMQ0uP2AhjQdyprk2mYJTLkifKyvj72Ejd2MxeZvfZSOmZfTND+t2pFHjS7
pVGlrzp4Dzx6GW6moz6mco0Ee/FU7/UhNKqr8rBBM13HGYfxhHDL4BykC+lLZgJv
WKDNjP7yOePJOWvp0Y4w2FAHevrw12jpV2mvnaQD3zgnSsOQ/JGmNS1qfdxSHIud
4TWpVJ02NHlOaMy+sU3vvZzzSZ7sXWVjs0gyph62wJKYu2MwHxWfOaXdsy28BHb7
qlwkN5PEa2UrVzFcDAThXJ0YTkiRyz4BYp/lfVhIuyIvh1P5DmuAid8IF5zptW1i
VrFRIgD0z4IAnYEG64VEqKrxC9xmZsfW77I77w9+w/4v4KTFNKzARHEG2XsmTqig
jYTp7YTrdM/OPtCO/e8rfe1urwZzYmTGdJa9ijdXG39i9eZ/pI1CozlFcQZUrv+5
Q1aNXzDKZZYJZFT28JtOlJ2d5IpSWvCSY4cQn6F0XovB2qPLViUrZyiiG/Grh2tU
9vMFoZZHB8lbZd/fvVOUbKhpVWzJk4EOvIAZLgjfBDORKCW28qJY1wcqvg4tojP0
lESj3smPqRAw1spGrPEAd00XrsOshyE1BSdhLpds4dNXa/xjQEQpOVdeDUJpYPK5
eusKD4SLktwntDAUlrMeXHR23BnlEqb/S9xwFtVQzWrfpTTLn5dDVRBrVQkPSJuk
j7HxhAkXkfVNq+a3BQ7hGebo9JdsmfDckQoXIeoI2H+WHxanDwd0r5piQiSRvh31
/89SSYpRzipbB1DNzu25kGCCuiJStHgEJdb4GrFObol48Vlfd4aDqOf581SRc9CY
vOztIR6Hpapa1RMasn0a1ZLKsubi6k6+0H7qsz/4jJ1E8MrqTItL70PlwMmHLqUU
qP4e1b0kpdcPPb75kmxl5JUcXNjd0wcl/z61BQG9eLGnZksPozfyTS8AJclMMsiA
AOR0oC1Uid5cmme2nsfqE1Bc26lVDYJ+FTc3oQzmgZiQHego3XROjWsApum6alaH
aLJ83pMG7fXc9zSB+OAv8T6Wy0RuGiS7zsldcTUAtHoVwDPGA9vG67vVlEZ0yTIG
mG65V3eTSFLEUsY2HVJ6yDq2UE86+JWbt+BkfahyJ4T1xmiL4voUtoMzc5/0hOA2
QxB62A9UY8oeyEZeHDA1v4O2Ig3DRi6e5DImj2r8bdli7WmOorqXHGMrqy4540D/
/OQF4RCUl9iR4IJ6JhYpDyXbveybBGNGU5NEsqoPzge7tTDiFKtdUSw0Ua/0m2u6
wHOKy3Efiu/UYfYjlcSDP/e44jy5PslGS77wEYsWjp1WFeA4xOHvo6VvhKmn+VU7
tVYCVe0Go7dlD6cUvoeQ+lS4nHEqryk26Zeo1eD8NkwWlMTF2FVrSZu994a1jBWZ
i9X111EIPIkqSwmKMQjjeuSsJQ88jczgS5siE/IAwgIoMvnmRVq0Ap+a5JyM6T/G
z41ssdl0NiBHDynz457x3ixKuv39bB4kqrgPrAWtWFbngXd7JGEsr9UfiS6PKPCK
1JMI6HJZ/vzN3gcMOHFQN/dK6Jhi/cW5TNZXjCizW5iNM0eDv/LOVCQW6u44pkri
Ymg/152x4sQZsYsL+vFo7BNwGP4mD2lOsgQMeH/Wkn3HYnSroNUpBtDu4ga7yAGu
bSmb7Gu9ikxGndxAn80IiXwRq9gw6UHG+Sr+UAzOsB1H9/7ORsFVVUqFOFwRlZ99
Y5wfZxSM/2b2aqTVurpNBOW+xHL6BNyrrjYB6Mdv9e3656NAZfdZhpJf7+XCZX0T
WB76/5wI4Ah3Ddmb7jzYsNJF380Wrc9LdnDejtARtOG4bUka/fzP8gVvmvfB/hHJ
bbG3IsFnMV/+eTy6SGK1qWnCMk14w3W+rekQeOYF5ASiIak13v/AXIBPnDTBvo0I
UeEFa2JZkzhe/xSyl3eqE3IkJKXGKAaitPbybW2MH02YZiXu3MFYnFkrvrWzpHCV
Dm7xcV/63h5q/L3pO4ag9kRhKNFFZRdwB3TBZAXA3Jaw7IT11O1dlvUge4JV2WpF
7uXJoJXrEk2fpAMlzn0yqRrbrzQ4TnTfNT4ZgcoTp+VZegzRayLlH+qI1cs0GOny
ja6jSEqOqLIvrG1htNwMoxTRDI49+NMKdI4tQY5H9V5N6X+3MLwBphVq8gDZWxRh
2wGfMQa/0jUo94HP2EnxFL6plakf28IHbpx7A2SzjZETdC/WsvjpBuOpzW0svW4Y
sKOHSytAx6GU9NclDfNs1FEPeJ24aeftI1CtUEXcqNsZIirlxXzckIJ1h9oHLyjG
bxDuGMqE7pVlTlMx573WjNp73AQmR+zxC7DrvtXWPjioZ102wHc9EIfJu82B3okZ
jCiSfyK90TX2eKh2t5jTJurbrUiHeeTDlHQgOFR1hcUJHkOEvXhuY6yWsFEKBzQP
VyVeYss2WLeFzQXU8VuzLjOsiVTO8L4dBWacVC5AE02rncp7qsDzAo55iRgPxWqz
KKzwgTPt29rT+vZYZH3qzsrep9XwqMwkhvno3o6zACHzVibRHRyg2sTyB08tYp1x
Z4HqUhGbfI/PA8L0ANinFuCTk44x+Kttmt3SBnjK+Au+rJWEKtFnU8siftxL7V6+
V8GzVCn9FbV1y/uyMJ/+E3L0nKgL2nny9eNGfpiP9ES7InYX6x1MSSCtI2xEZ1RC
OvYuM0Vnn7c9/aim2+Vm8lKuk1rN1/fHEl+3YgF6zh/K3fTRaKn7LzcDdg1hXhxJ
hosSlQkjcMEYIJU/mX3YqwokE4SoH5/sZz/OPupoAfPUd9asg4NaDbZlkPG4hugv
3vd6aQ1JSecSuVDekDU71oMoXuaVrVtI4DZmU928yHTW4rnpPzNN+8cdvCbOVBVh
IsCrjWptYSpn/nPNNxpBnMRsWVUZVyxKaakHZ4n62m5/+PQQxg5VesZljoQfXw6T
DGkkK+z7d4ShGWFJK4uvMR2bqc9AZiQ5MNTZYoiRNIbPjub0D9CU819lMCkNOWW2
3lwvzMT9sIIEVMFZK7L4pxOKEgpvcLTS9XWM3vYYchRKQEQ9HkmlrTCeXDABue4C
RKibgUIOB61ScISAGrZMP6ZDz2h2PHn8zTsIrJHaw6JGrTokp1iw8dpQhDzK5R7M
49FiWaT83x68scSYKZ7sNE17zrKpVB9bJRDqbWV0IGVJ1YnzJvi4SNiBetsUop8r
ymSj2J6L4IeA2lcfES6m2rLnEtKLGeDaMyWAmugR5UTzWIYdUUuYHPiXQ5qTfZwG
Yy57BMEv2oRCFrMp7coCZTCOEZZWyCKccG6m3AdD3eYnHgAzq1pDolLHJi8M+qnj
U8MhXGnMk3t9Dzl92ZxYehC07+CGTOvGiQypT6myIWGFSjntjsB0dUJEJ0BGf6Xo
pUPf0TqTJyUJjsLjaM3R80GAS6tI+JCzuZdbxZyb1M/8gP9gB7NoqL4tUmyw1mtR
ruOmpfCEQibKtqp6NiHfqqryoszdDkPbGfJyAYAabandTq/mILsUTGt0uSzwkLfW
9CDcy1XY+uRBIwL2W2L2uUqfGH7FOY57LQufn1hLM7eqk2MK6ySCcwrWAdgsszii
rs83uWLsV3lfKb5QXq/luj14qqkFdh9FwXlKg7t4EKgaYNCVzAmfQdDCtbWomEwz
YRmx+yta+c3DGq7PxBVX0VHkW5sR86rmkh8oCkATzvbPm7ARqaGlVdYyWPAMC8Jh
QUWb7O7G4nM8gIotB+RPftqEpuN9MuRn/ZBc6ZL+NDsfPkBqQ8xFnV/GSL31TIW3
womnJVOQEKelNELOTZpFSwqT0WHFvjn9jXX3zz85zrkVgH/TkwIWdi5BOOkJRUTT
LoW0fdtnL1gd4Ko0puOCMdUZ2x8zW7w07zbEyxdZAk5fC3TrNxKNsoJhZpoxESki
g2TVCuDAtMQyEueVoC76XcrDn5HyVmth7YYNyh5P1gWNIPgq0S6+fNlGrj+em1Ge
kfqMw0hbM3zVu1xNoaILJSQKuCr1oCQFXnxAGuQIYDrD4l+zIw7c1UV+Gs59oAA2
/eqLSkH4aQ+wIIb8V6VoX0vkTab2LjgUPXMW3Uu37IJo6uSrrWwHqlgUJJ2g2Pks
SAn0Gz55GScj1Gzs0PI681xLAK1c2NORS7gRIX9gbmA1UeHhY21pAzsnOy05dEa8
oSNz79qsIk5uuX6r/7VWv14GJAT7ta1petJlq1hGci+8gtA2bJtlBROyO88k3MqR
kazjbBWGEpShXIXSL/XKy/7b9Tb+hZy6Tz1UC/eNhhmmjvn17aGxZMHHu8ZfvFRu
0ThsAFcRymKDqFFZmjmKALbvloxFvv37oIN685seYSeChP8G05KOP7d6oJo/afcy
j0dk1Me5uX5qssx0j4opJrewymcvOO93ag3sDcBB5NSxFc57bMQloM64R1FT+NtX
0VXBVorldDkh3WlZSZ3fyJ0nfD3FmqZQN7WpTlWCKrr2RufJHFNChYlcTxaC60g0
5P5e0HqoWWSn9gJoSg+M6CwiAva/mcd2jD5Xn/eZHK0HPaLfZRwg4IF0JmjLdYUU
GQ0huWAoHS0dt9654VgQ0v22LhtXkSAZHaK4B3LGZKspSIXxjyasXWjLu+NgvVRu
7uqCDBCBarQLzZiBFKLN49U6k60EeR++Fg4SbW30qFYbglNokUeV5gPKX+viYjLt
RrMeGhUAKUuSsvBdKZVqxvJT3obg0k21eMsRvA4o1hoc9mG41HOIXEQtXsXh3XKX
HEqQS4XvPt8ubSYySzkOnagkizv6SwqDu6XIKA5cVmPftIlQFdu7JnGFdBYRX9bx
MhH7Tvbsv5LxYMQy02ndtHQV/+DMhu1F4jgE6dSfHLxuwowKL4d5pPvCqdBM62TB
skrUOzoqRm70VP0VUD1ZaWlx8Z0/73QZojwqoBaoAH37JpBh+Ro6lNHa2ATggkRo
xaV35edty1DEWkVSwEgSI7ZmVuDg+g/zwWtwEqlUT3o7o+dX6wrnYb+v7zVcWUc5
2k5NPYNraBKfbK/a1DhIRQmfmAuv5MGjsDHwJP6w1MlHsNJqivG0A6oPX58/SstS
8ZG/XTwMANcIOkicFi0EN7/clEitp9pXRRsQGbNT+TzYR9jZesRKPo0sbg5hShMF
4lnViBflBeJmcEUR5WSrAWrD2wH8Q+yzXeTnz5gqWUnF514nAfbTes2LgsHRu2uv
KmfkqYAoEQnzpKNFAnCyBWM5/i0EvwwFFzJuSULleSyj2rGAedhbHjCKQJLB+yJL
8KjLSbRM/c3O72clWSt850MglGaWTDjZTNz3kwQYuvmdEh67KRcUgvF+PsI9Zeev
mEGowVijckxgAyfhtm12qdCMT3QVIOpOAGSkLsl45AjO0D/n/AQY14Rwbaq83yQq
PK9QAYzGQ8pzrbFWOODAWYmJBQlxUwfjV1qx+LZJlJVHg1cKdiJKT1f05VMcKKFL
CLxR7RVTfFZ+OEjZp82vrUi2e6flp2i807auSofWrjcNWDbhXAB9QBEIG5WQCSeo
LI3s6P+B6LJiGPedCEieuYv09RMWHs+HMxSy3JojYZM=
--pragma protect end_data_block
--pragma protect digest_block
LnoOCQ4YLbCVHaVTd6SREd8r4V0=
--pragma protect end_digest_block
--pragma protect end_protected
