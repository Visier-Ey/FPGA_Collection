��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F����_�)��� �����7�l�35�mr�_.J���|i����h�%r�~t��Jz�jݸ�~p7�3wJ<�e��Ql;�w�I���=�kX$��QD9�*�C�bB�wl�U�3��(�Ueưh���ǩ�C4Jy��R���yqeq(4���'Ԁ���_�d�ȝ��m��D�`��h��"9���+�G����	`�U��G���^�
a�i�W��8nN��Qev��gdcX��btA`�bG�װ����E= �����ǿ㮍��!z�Ϥ���|��!�̾�� ��)<�΄r�6�d�mS&��8�[N��WqF���ߚ�h��� ���/��$P�:��x(=JV���a�~����Xk��������7U4����q�����E;/{c��V�bD�E�st'(1v��//�̢�W-)��#��)�8�:9J��3�ŵ?>5��m1�������5+sԴ'z��($�>0*���Oh�xsͦeM��?b�U��*$���H���A5ʋR�ݱ	|	U�Х��SF�1\�'�gxW�[���6�Ǣ1~�g뤿���Ց���u��ư��y�{4�U�Yh�w���?�r=�KT��l��/rgr�o�*�ǯB��YHo6s�eI�/���HEҠ��Oh�"q�z�x"?`]�ڳ�C\��N��!�8�*���K^"����?�+p�f�c��M�+���>�j��<EX£{l�W�
��jrD}oP���K@]�Y?�O��-S�օ+�����׃�J�����As����\+�$1v��	��r~���6��hu e���	6߃\ڻ"���6�ܮY�x�?Aj��=�۳,DV�l�Q�'n��lE�+�N���<p���$�>�h�q