-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
--pragma protect begin_protected
--pragma protect encrypt_agent="NCPROTECT"
--pragma protect encrypt_agent_info="Encrypted using API"
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
--pragma protect key_method=RSA
--pragma protect key_block
KoM57QuunQtwYbR4tYWaTFc71rx75xKWQ4Qk5aaGOR53znE8gMlPTIVUaPdYEu1v
ZGtZNBqr47OUiREa1v+7gSHEuW/e/xq02v7WgI+CxeaK+01IZgjEU+TRxMiCvF0w
uQCGIGdIytXZoZC8xZZqQ0ahaompqSLafaIgYhmJR6yoqunMFnLpjfJk8gRmr+Sw
lhPwWF+YF77R5PCqOj+3QtGSkw7PA3B8HwJNvEJ+edqR6VhdmzNouC/MXzGH/26F
q1maUgxKxDJ7leXyfYsxfMhsQc+XBIS0nZ4ktsL1loFmejW+WqVidx6hJ/UYiFBY
iYspipwoGrmRddcUd4Lscw==
--pragma protect end_key_block
--pragma protect digest_block
ikR5ggghFraz66kZviHWJ1ZeC9Q=
--pragma protect end_digest_block
--pragma protect data_block
xlx+tJvCywYaqrG6YmLOsmTrpswu6uJJGpQtqO7a8MZz6YcEleaVNsW5wwW8Qcap
kkOWDi2b4rtPXFXAheiyU4hemYbcB6iUdViUJ0c77hX+nyg+adow+jFy2Soneakp
FbeCuy7m56YrJumzp8Ti7D3w7F9r/+Nqye75k9YK78J1lIkUPBWmBQ5WMJkSppIi
R/rPX9xqlzNYKGeQTSO+VbdorcYhTe2nwFLuEOt1EtXp9Uc3HI5HE3E9iL9LESAo
F8F4wLYou4RjzsA/zvlXANG8qUvlOkdk7GS6I/7nK3T/K/719DlHNqmDAKWI8Lqt
nfpJwWNiC5AqXyhUGyQ7iE/0QBw4L0gJDudXQGrr1Lu3XxrvXCqwOVxtASOGHZME
j1L/tOQ5bW+uslUvsZNcGySsd502XVtuADdxAZAiH2X7JcDWUGeY6C0Y6ueu8nw2
s99FiU0pvrIw5mPj6zVDn19PmScHjKMGSMjXSUNzRVqBVLhRj99NNvXLEQYSvzax
rt8GJiThNb4j9G6js3oiVKC9phZysg/cHwL6TgEVUViORfhRZP9EgUsxrT45nuuP
FjymLMCmDddggAt3BT3QBxQWDKGP0/T4plux7BT2XpVAOmznPvARgeeBIagnbMZH
HHGdhPJXqsP2rCrI2GaFvxpLMRP5v7Rgmg+FNK9FO+JTdhHJoGlBqmrLOWILUlN8
zTrvv5wOLdOdfsI61XvR1oqulsTTb9kdBjNeF+GMnfftNbBevpCapMsqZpuUSEgP
4X+u5V5HqY8Ke8WgWW5iMv5dBbWlhI6S6WAoMbqH6yRj5JoVUyu7N59LADjMLbd7
qCzG38YXy+Cz1jNGWbkFYY2749PR3ClNFlrP23tQz7/2MVAjtuxwR7powRRda6Y3
xDfl/MI56NfgFyMeAvCRIgi5t0h+IAMnHcwXeEYvS7BwczVOx8ZRpDU5F64FZQDV
Rep+2MGe0MqkIBxxTDcjHuz/PCkALqFO5fy39PbtSpNWPcszS6tDlmRr4L62Nws0
WyZsisrXyxmBvjmMY8SibSYVfvXI3ipy4dpuFVDaVcCvogSTXg9kG01YMskMsuhL
ZqfZrkSOrnyWChSSix3z/1BRZL0tPxbVFcNK1ImzV0H3ssAiKcKgM9FZ/fpnpQNN
i2kvVL6JmGfYumYoOqG1ZTseFYhqyaLyOHeCGo1wTE+ismy5sczXhuUkik5SK6Hs
eBENhrpE7NvXf9toRvYKVqsX6eqGMs/Umn6a3r/8FRgI5+fuEmg8aqLDlhl3z+Sh
EcGkJA60eNOuRR9YbOII+UYTZlM5byB+a9fUgV+snWWWMJGk9dhZLZo08No1/XTW
kSph4xs3l58mkc7f/TxnaruQWO0wTpHMjo+hYMhp/btHZhSOjFRJLBPa4+3ZNHdS
HbpRQxScwH8i8IprcgYr1Mnu2xqjNJqlGdlDXUl52HbZpwXmObqDsffc7KiMoRfj
d8vC1LXGI76bR0W+Hk4cIyElLLz0nNEOsJzTFS8Vfc5aqqxPmVagOCn511bFDOhI
+lVf/YFRF6jK6O8RAXI39QRBt9R6gc8zbRe/9wl2fwCXK5WqN0VgXwOahrEXNr92
+4babiJHN07alj4SfanoTse9MZIqaGKtcvlEv+CdDuInberuiRkASkgMHR4Uicj/
SPZqhfjbjzk4zHjjfR54fwFXCe5h5cfRg/N9Bc1DVt7vzfgEjYnFYYVliFdzG+WC
k7rLj5bTEtGQGd7P8dPVlaLKBj/AzcDLpi3caAdVSbQajjaK5EGsNvWF56qU76hn
KMYYb0Qzp9IiVG+zdShzyGwqj/5h2qWb3Ey7fL135VZ3bjKr+k1+ADxjJOROS8py
j/+CipgxWwB9hsnlxP5+8J7t3fwn/WBb6wdfMGoBocyZg/A27+KDvMQJDBz/ZdaB
sZfhjaE8Au9o6imAq8vu+oxNo+CH3lFLQzLCXTW7ERP3KKo/sc/BGEO+eGDdmSV4
yGOJUaICz20+PX6NJe72oARf6DtPbsnI3H8mfjmSi/StCDGLvLtzELZGrFI58WkL
8Ss34LB8aBoLQz0mlUOnVvTwC7cG3jVxxsHFlGo+ZJpT4d7DRIsC9QOaVfl17L3m
d+NSMZNNtm/GDwVPeYKlw6CiJceERxGObByZntTRCFghHI33DRX6MrIPByI8alpO
HD9Kzp3C5HgN4ZcJpUilDW8ZFUhae5/arFP2tiJrjU6w+aZ+nIE+VSbqLeDEXDvr
XjFVYNEQQkHsqhMkZfnF4KxYD2NM391/yN7OBGZXODixxsZLVQw+H2XrJK7ORtcW
EHeUdXk3CVprJ+jcax7xw8Q9aJYYWUE1Jo+uw9m1sGKn71OzAteSPpUuSL3v0Pot
4tproKxeEMV6QMbKxoEuo+QS3cl3wtvCJJuwtQhah9kD29smETAZmRCfFV6uuAiI
PHNotNLlDDv7tN7caaPomYglxeMOYFvm1BVfgV9j2xxftYGcbqYlhF/Z3CQ1pBLG
sVKwKHGt7XAz9dY0U+qY1gCCoPPiZJhVU0NTtqWxqv2wMnYShxlu/XU+hBGGGDaa
jkdvZFtXFTw7MIcS8Twq03KvKgi5Fc4thrXbuGU9jFUF92IdvU0wQVhWye6z5CtI
ChKY+TXo9AYg44USAaJzkUZe1NWrWBCnI0zK5nGpSKE10SUt5WITdQQqgqJ+gPus
kK38K9oSnH9p67j5rprQ+Q5kAwRzjBGlr+L/ydWz5uU5nNC5slH4thQhEA4R2Wkk
N10XNm8+pR0oT/IRlZdc9R63HDmWQH23/Zj7Bj/c0L6jjK/9oFftcXz93ICDughc
IGYpCeX+/YekK6VPqiSkD66EzaSAaygJ9W5mnkffgkdI6QHr4JjFMIuh4OZNy40W
3F9szY3g8TIVkF10wbBJGfpd3UkuaKu5MVWhNVWERBPn6jjzaeaL4PKRfFbDpC9f
UIqo5cPBPMal86tfJsi5SD4Oh0UOSSWoo1p/nwiKJyFFYTrPhQhrQuOGCFqtNCjk
qyTjA+VSHgtVS/jBVIoIGDQ+NY3LQbInW/AP9gXETDskldU2jlrx7Y3wCSgrjH5I
0oWxpzQtGjL8SwangB2Ae/TAnLx8VSV2kVSA6C0Lb8PfyZcxWexUldfaLnlWhlLp
qWAyGrVzV1V5Aw9nax8k49vnm0XLpYrojiM8KC8upQ7uLgLZoT3uZ/X1wM6MWLsC
ne5OuMgV+h/IAKcZC6yhqGpze0NvXvmplLEveAbHJY8dZZ/0lx+ZN130Q0Exm04O
qBjDRLcFnRNaQy4YpKbAGZQEVx2+ZDkqrDMrVrT3ghtGlFpF16f22ahBEBpOI/X0
y2vRkDqV1oofrc+A1IwwIJJbV4O7jNKG5FAeICaZKBDOyYVBczaV95BhROsMddoY
IQQD19W1dAbYyJNh36SMazJJbipAJTpbvtQ/gvMy7oFNmheIUS/O3WFHl6TT/ExH
Mei2xeLLGpuvr95HTAwp1MhVS0t2UF5eRvq3Wx9nPHlpZ+04nddPTrOXojUGt05E
bgWRZ9woCkjKhiJ+xI7Db2aE9lUgoT+Ofpt9oGYbGZgrLNABsHvx/S35thyz6OcL
w4bc+r7aVV/9RYrhpi7BpbI5QCKoHF6wLAYuXaCu/W7u4ozRqLPf4Uj40oxaI9J8
paWQxWS0fBARktw5v5D23arV4VAcSazb37rXOopG2Jrfr/9oJvAGdQ3a/8j7Tw0r
pLKb3eO/l3+yJHANROHgO81aHMx5V9sjBOC0ddWJpUlO26oTZISKE+vf0mnSlDq4
OFxaSYL+qy6oJQzLNjhSox5+arn1jn2x3GqPxrIjMjN/0H+050+AUgznnJXaJWI7
GnEkqlaIjCtDV8+y3w73cJb8IL+t5BhFBWeGaN7ZK/jYqBOYQjovIbR3y2blSEr+
xQLShOkIUC00PB6W9dVv/ccdOCoAktjcgRop1Ttr+k0mrUr146VN2j6QVGpqJPqb
uBWOxfficyPz9J1IuRFnBhCR7thG5ZEi/f4XcDL0i90KBkbuIW4PG3KJRkqU4Uxq
Rh9/UWM2Y+DDStLuU6x4rHcb2Co3oy7OciPeCYx2T6N/fpRoCeMvWFeL+mH+QATC
C26OnsznXBP3272KxjFI4ReWOXMR+Xcn5ik+03kxHgPUJJdxdZKJkN7VbGL94QWi
Jq/SjVtkbc/ARrZH1aM0T3w7ENMSMXWaGorboR5T0cW9fZUosH7P/DHeMz7S05yb
AO4DMsoOeWwpeZv7HqBiwsAsAEMZ8z3DVPyvPYmAdODWPjMklHUDLu7NoZQF9wz+
uWJQ1iyNK3ajeKkG+kWh1tkNl7uUaFxtwg5CNtZMQ03z6sLSAWMSaOrEdZgO0MVI
nmJ3UN0fS7Oka8mKggWi1zY91H4ekvtfWkQG/Y3dJyeixlYOvDT0YLDpbrW67qWZ
b4EeF52Mcp3Lgaf7EnBvz65+rGuvfAA0gN7Q8aZBzVJHY780MDBHKsdg0IPTMNyo
+0AwKKPKpxIwgBoP7tXlPjJ7yRNLTnUzE3dBao34RggOMtsWN7VJ8tkLo3AlORUI
viV/bReGxdk+bS4ZNmhQ/oFjjoJZidzAAPTbTLRdfRzVEuT71yf8ZV7Jll1PIhJ3
dfXAf2fe4H1wrdk8ZRjlHHYN102sYtQ7DeKemLoCalJLUdkL3Lt5bLhCmbvgHKrU
mgsY8KQ6HS2PuGUpPg+/sHXT08QMTkYnWC65wRYoYvPadqcm9MxSxjAbaDpGBBUt
N8JtDD32tHO49C0VatIpCyOm7e3DEG82gnGbQb1VUfcbJolI9ofkSgV0wGWwDwiP
3Qmu6OT7o90/K4e19pO3frE6C1n2jtnPSTvgdOwUuTuu0WV9b4PWMxKUL/ffk1Dx
rJlK/TwtBvj+8UPjn85gI1F7wqZ8g7klZqlTIir1ibs1mkgLBFgtWiPML8fwnKVR
6SeJWKoCVLLY2OWFnyu6mwljuYNvGRI5havQbokNoOq5wAE0rXnW6ZYrv+P1GbJi
v6nriIEst/KKu7xrWzk49tV15cs+h55+l0ranTNtTvFqT56L5zg7K++e8aqvsBGg
89RQJH1yUQMs5ZpHTq/fU+JjlcmUQKO0eJdtroSZIxJhTBzgHoD3JlHsIqW+rT1g
ieSvr2THz12/noOCWu9lr2cZSwvIsHKvoSqt7gczOBEskehBzGdM7wgPed/0AU2m
p28AOnt0/I1QICCjksQIMDt08aWEavhOaTUZm12XBXOq7HdAleP5UPwVJaNfZyeJ
Lk4HCyj4oW1unyTJ8l1yndA1K377IgNKKd8GTCyIu140ATr9vt/4N6aC6CcBhPTX
WBovTNx6wvMXytVRvRetT0lJ1O5zqMOW0Xq3QWgGSX9oM6v9VN8gO8/4eMNZpiJn
nj3yXkpuu0OIqee1gOCVS9XvFj664ue5z6i0YnYC0bCkPebggyB127D9tDZkoqUK
6rNMKQTfm+8vaYTfVEr+2g/iqW4WwN8/YwN67uuLkN/1zdIPiC/ob0CPB4Sqk6Gk
8DxMUaYlLPkWDk2jffGR0lYcuw4Ewv5AjKmOrYMJgjCYLQ4Xx2U1riRArH69B0Io
Fe2dDQclByvJAm1wzm0Wd2FCeJYkRFsj7KNM1um/Jr9pBsFkPGWENmWhpkLtNBMz
+16CaSEMeipD38tA0Yof+vCgnv5U8Q2kS+sUmjvXSDLWEJG286i+IdEyL2Cyr2aZ
FQD5OoNteJ+2R2mybGn0Gs0Qc9QcH1sFIwCnrswaC/gr0p+A1D6uIz7wH1uyV8X8
oZlAEM4gH/4WIA520t5GFc6oSZOVOHiEwxekKNOBmcNLMJuh5ZmXykksFiUn9smW
3oFM5O4mlkxm4xujDEGF6vLBnLQ9p8Uq5HNrXciAnpHDGFq2bIjld5qyKrJsRcUh
SlZFZHqfRn7ly9m7s81yCNdRlP0emdldqJwpiCK/e5UpwH5jZJSVoF8nfi3/URxO
MI+puqTKqf00svhg/Eg38dTXZ/2zECPSzJf291mIO2YzOEi5A54mpNUwIeL0I7xt
1D5O09u/yHjK1uvC9CoyvPP+YLdQNemUS+dIMdYfHjP7LDrDQlqeqGYPjyQwZcjv
DzW72q3gYFI0NEk9HQFhsV8QRtKucT+hTj5a3T+NyF/s61/iyTlp55YV2F2/j0wd
HDwhcDiVjwmOZxqD0vqHnP4xIuKHGK1izJ6SBjSaz08Me+EOgX53TEG17yUk2Zrm
jlt0wDiD7j0UqZFPpWTEma0B5Z5c+8O5Nw/6ZzS6okwi1pts4ZKjQjkEMyw7AapR
Bm2Kf7nzQfTGRAddHUEBLVOqgNi05a9NIvrY70iheiY93D4zfDdYHyXhOkEGNrll
xkYI/FJ0v9H3AHAzY+dQU2LD+Q3FlZRm/GgcVoQtEKxoNAGkYiQGbNgU3eBwqdR/
yjBOT4KFumXIsdcm0FbL9IN5M8QNMLnBQfXG0AXgRxZCdlvXojdG+SSTn60+BMUV
WpUlDjpMpXsr0ipBVICJwEsOyY09SauuqswnYfmwXFbi03JvMaRGbhbffKbxBhSl
p0O7//4wvEBqa+0K+m6Y44rXTr+VZjAJRzb2lRQzK1UmMHRJz0iu9BmjpVKzlTwU
q8cyJzHrxbRjGgG6oeNN38i5l8UEPvxeIl9vo7DlsnNYW+TsnGw1lr3DiJE6U8kT
DpeAqesAOoffTqKRS2qcGo+9+X/PythpD/lZgry7bkgVuB7EhjqIxcbpq2jX92A4
QQDrTm9DIB0/ojabIRVTbYM6J1jOHpS3nYv/D2CcAX1napnWQJBZgTeqHfi625Vl
Q2lyofrpNgAovqimYJzsUrv5JUczLhG0WJB4hljzeBFHK/tesRridU2Uqz+tUG/7
w+gqUz3P7VvUseCWqhCCk6uET8C/gJF0PP4wRiqQLs2xCGAxsXGCRNz9O1mdUt/k
7jzbtixQb8jYnn2QQbXYm1/4l6rwTbEX8zjgLf8ifOdhTQoYa5+qennkKl1f8ugA
Ay4VAAJscQ1BBx+FZWmdYjXsecl/x3CnxLROkMCnG7Qw7f1X/ixLPqpe8/Ejo7zD
iMAFM10RW40BxWlWD3iz/PvymGraNeupXwIWBI9wW+ZUCipSntUzwCU9lMWZkCzL
tORSo0EOQnMyijkPmAKeYkRRQZMB/gFjFV7o+jgtNCMGjr2kQ3+uPluDRiUhdVUm
tqpVmdiM1lxR49o6Z3j3KgnOa5RyUal0Ll3M/ceNqrDDXi05afFwRNUt37ctMn+h
FnFaoBA/CrxIDNO9LR7qxDz/APd9HLEMVrf9K5rIsg42W9L9ZM1aFuy0RLnavFG2
0cev2u2//r+Jupno0QbPr6zGrKUwQ+CB4TKXCdqNEwch9otD2anmE2NVYaPc/8SC
zysVCBfd/wmZptelvDNjUk+aQnmb0xYnS0Kqm/pRiLe1yKlA0BYtEqNT6nztGWUB
+KfcKWefwG70ca7S7kPJQIvBXOyYvObKr4lXBE4/NN8lFh4ZCvHecEgPiOXoK+5Z
jBqlD+19jlHiHiYRmBEAN8HCHNaaMehkOxi9yxXQvmcWvIuF3qFuiEiXNg0iAPZs
9GvpEfjjz9clFz23MuOavs0TyT6IuDfSyV3EL7nf2FUeoAMEc+1Nok9+vTntAWnj
GLTbb+J7hcQV4zMRnWIS6nA+QU2VW7lROjzUfTyq6Nrl9sDQ9+isXAmeZ9+rpNPM
7LPODFV/NqfQvCQiPhgiy3E/CN94QG9QO7IBvPzujvFYplLNVM3XhxlYvPyN/QA0
BozzQUCTG+IoLP/xMBweTCycA9LGUAfBXkJwrG/qxIXvNXKIMUonelr3eX36Bc5b
haE4YrS1Q8anyOhVbDU64cTVBW8rHwfe4YfcoQEInATdkTSkEaR/iOYpXNkSv2Oa
sR0MegWHQoFKdFEJ7Jo0gWYXb4B26rNC8u5USFwmuFXcdAOnxmBvioUMORT6RaXm
ddhbCIfcmwEPVR3l0M8hkLZQPbNe5P8zLClKdmwwMAenRoU6otGZmXUfhUdhYQeL
/4JsFsGoCtKe/6nY5WnEjCT5+oFDPGAQ0eYJo7K2i9lDtfHcaneTRmZMHapf7GdZ
JSDxA/sBoJVLayfQCLJ4Fle3MfvbkBcKFcDYW6yHJQw3VGDRud8Wi0qaXyHzGZto
X6TdIvbHQT2kO20ep8HcIjbT/a/LlggxrL+fSk6odzzQ3l5f2Kury/YPBQPZ7bPH
TEWFgfJCCud47PRxQVoE1CZpCgdED7AWW5T09mAXKqZ3VETk4vvuMSQTivK9LW2N
zWE2p8BuSFldftKTn0IUakQPl3Z8QGiAvOTd3iKvQhi0uBc+YnbySsUcAoNhnJww
bUS2kpioFbjpdpojpEEinUh6sSC6h/MhmNxiTBlxV7GhDR2Zb2D3tpH0Dtg1rK4F
bL+p54qRVJ7s5pPhiKJAvZ3gLORKcVqI6CgeCo6TwRMLEe1M7qBZg8P4PFlWHoLu
16xkims+dZOi12w5HVZ6Vn2Ah7Mac3OmeRFsr0oN8y30K+hENX9pOG+WfTFzWcus
NcG8hFD/oJxQ1i8eGzKD82CDhj2Ox8yM/TJ7qSzk87Y0FL5QXZu71jKH2QQ7M51S
3ufpc2n0QTD2h3fRW39opUjqrtCfkAO2MYrQR+k1ddghV65+ou8Jk9W0eb9cF6ZD
TisEEeryhXiEyy9TQBwu69P73sS+X2n2dDcoOmV+3UzHdSrBbAYfgtj3B10QiVGK
J2X0o5Rj1xI49fETnTFBqmsljtvVlSxnk6sBirjvMESolbeY9yGRQN4BMJ2dEnd7
1ApEyo6OWNjDzNLx6jOB2hMH0XVrdBs5X/5m0XHLP/7b5vYSLPlBf5hd4xRKZ+OT
RnnCI9UNe39LTaZfTg82fdOfnDuIYNm0jbsOVB+lpAEdHUm1eAkIVXrlFU60t279
qeyzhqYYzPjhrvDGoZp1cEL7cjnU+SOLMfg/ccJSWOCdMHuQd3T4LU8TZK9O66Dm
FfI6n7Jw/iM9oGSoVxu76+sy/Qt+cLZ/DC9e1r2lkUM0Ahuz+2FTmT0y7V4yJ1GV
pA5JBZObfhxhnpqfboYshSGCNCopEY4wjN/O9za0sJbKjYdH2HgGHt4qCiTNIRAR
EcPUrGSdSUy5IfLO7CtBqAawamdozGdmRBmjOD+NgCUwf5LxzLy3ZvAzDSCDjF5Z
VC6iTVZEvcv4pFZTIEHmF82E5ZkZlup6N/3kzwIuMxAeD5o7VQNP2IFeP9mjvnvP
RN79Vsi17jPTgVRI5sfqlj3wpp457mDcpAl1lrxMlk/UHO/4X7REjsGZrb1VgLWv
vR0G1/osUKS0s+5wlP9RJSPo+/UnXMuzXQyg99M/p5uJGUhmFLI1MlYXOv9CpZsU
kjs12+UzeAu7v+XyJ7vcO7Tn/GkIKnCIE+k7ljku7A+l5o0xB/yciIb9+0SK3lMV
03ezLTW+PMOYhuliHMSo5P84j7RCNGaYhU0dwN5oSCZUnlw+0j/mlmZf27I8SCoT
Ls6WI84AdrUqT5WfwhDj6JQMegjsAXwJ/L1zBoQFjLsDhZIxgBN73wK8nXcA+ypt
D3rL46rPza31T13u2fTn29Ypqx6SCk03PKe4AqIJiDWexfZFIpfLWk/xKokvndIO
XgBvdbAjfL17TrBfYguPdFuFuu+G3rLja3tCT7fwXoHDhJLXtYKF/O9STLsTlVNG
FRu+LHpRSqWe0rTFCh0HsOaeRq+w4KyVVpJKWOPvvESvdL1jkeAmzfmETJ9e1szj
7AnruhukicCSGw6jV0/6mpv/R7lL9bTm05A4NYpA307BzQKiVbjcj5ncCgDptKWI
FTJ89FOjT7yhRi/eh5Oj0AE5hjj4s+SpC1MlHB03nn9NkiYhhu6CHJwyGBzE3Asu
Z9eNKRlBAP5nGpJ72AAeHN5esF93Q4ZUfxfqiHyBLvEj8iMzCGDEfHp5GhTOZJii
48F7HDj72BPTEYn6L4yPucJj8YK5Q8glqZWNwKkJDkW/uSLvoaY6UPqH8BZurAN+
YK3tfFh+vw1dlSgprZJ7AFjxykXDUn/HokxBy8hHPpDJVYLT9U+3CKeFrzCtXPyX
GegN1PDuDgTZklJQ3XR2ebf9/RVYLVLF8ycVqWbpG4aEcDoqgJ2jHptWQeSn7K3s
x1Me5O01eVlVz1E95yjbiGg04Plcpb52t8WNRiaAYWVHIEP7U2ZORRUiB5mxGbAn
fOydB5SLvs1nrHrFXKQPrXbZq576lDr/Ckq39T3ixw/t+9QjdgkN45TnoqtlR6Yg
1TxDAjbal8YoZegJTQZISdarqWgUzaV3sQWT9WabYmC+9GFZ6p5kCOc4pHAIHkDp
cqSJIf0Rql3bSpRdorJgSIWWfiUaM1fp18MF2gMsUfmAYi1jGP71gDRq3qnZEU1q
96o4+tdU/mm1d2iY8ImOMYiQN1QaOQe7V7voIThFkePlIQMsb2QHEhUdGrHy3TT4
DHWYd5ltThTsBuhZTitIqV2Zo6E1s7NnGgeJHoSmTnecRIYqlcgRU1Wb15/Pmn4x
fwHFPMsvee1E2UPOxNu4NhIcJJ6JS8H0OtBysy0HYk/E3R1ELFquqq+8okeoPoE2
269CViATaJGGBJ9WWEMHy7d2ybBvBmbD2tCPeHd2QPTVnf6lUTeZMdhJsKMggyeg
ALR3Apsjh9gJUbkvz+EeiKplbovsqbdV9blXc/H+6w2eon64w8i2wcF83EcV+yoT
j4Nl3uWo+233phXmDXgT66TX+x98/k6DPM+2pKYSegmOBfgnBQLoZ8rlLO7bW0Wh
F8R+YRe1TeGCxiQhfjvPJ2ygJF11vDxh7MEsOtATuHi0y+dfhQlbiTCqK6wlHiRK
NhkUHTkJ8QaDiRWI4kD9OJgtYvP5FJuxA5+mlkXgOojAxTLTSBw8JAWx30Q5J3wy
4vEl1ceOPh5Z6szHAFVCXwM+o4sfZ/W1C5MljU/rDfOntg7taWfkFJwqmi6mMqGd
L7VhWVERTslY0j78L9ChKDBCU4f6tusJghZVPhXn8s9Kku+IkimpE05eSpZq0NAb
bivJ0jhB5aYEN6xDfcch/Of/1EojT+WIEyNZXvje7pB9a4eKLXY9rKjhIXg59xV1
4+ljFjvV0HIhR7zKhCT7AG0yqGUCgwOKTNcxsaOHOJHioXsaKuvtzesBvpZO2OdX
FMvbu1wxMl5eYM8Rnr3HPTPvfbM3H2YnMsXji8BwqFtsSAjb5EY7YssWZy2Forhu
qMLcDlAtzGXKQMEXMTtP0FCrfkmwj3jhBzBQqc0rlnoNSPB+GJb+b74meXPJDrwa
fLAVJdTMKdO+iwRwu4JwebvIhcsZlY5qDt0P5GjMR3LU1HtDhL0tmTLKYbZMpy6t
5yAflL567/5ZCZ3u/qfvrZXQ5Itimkb0MAtdnEOHaUMuDDDsyicxAyn3Rd1FsM9r
ydufTBNQ7orZogM8bZS2Q3IX8gjJLtafxgkUJ4XDwV7BFl8J7AAgvtxgNeqb3FZv
K16pDmmiKwryfELuXbtFTdrI6AZQLM0hgIuD44ZoU3S74tlm9US/h1HvtgJOlf33
oIiHfKJBsf8SzMmDA2B28pIUbpeeA4ngYXSML4K7Ysg865+gTT7rq8dQRXU6VEmh
68di58KC3wCqR3r60hkz/1/6oe2/XX17cBvpgGs3xJvYHRkKDXa/C2cP7OliiNbN
cStpERSl2cG4rLF7Ud7kKE9l9LjXNnE2nMQC75eqk+yg5ncH7Ky6DKeKz2vMNdr9
COe/Z3YS0/zRBSOQ8lzg1rOhcfcIQ+FwHg5jZ2QYkxVvS2TwgIfi6WO/GYYcmOGD
kgd/8hQ1BSW9K8ZHFpRYEuLQu5395+NNV64jx6YZNJiI9fHCuJe4NsdeNAAJ5hly
g+XQALJ6dF4GBsn4y+UC7fprcZMKQNkUOI8mkRf/HPtNaDSW6iSOydSQv8heAqRE
CPEA60RdPC1sj/IPDTGzKe+oRFUcMHMVImyTyKwRttcsS04YiebFdaKgEB8HPpW1
6aEE9ncfqkday3gi3DQS2lPtj05RUcWkKTvGoo35fudhKGtjEJY3ebos9dlrtzew
UrOIKwtelBQ+r1HdJ4ZT3yyKajOLJdDNpmhKxrSfz9wgjK5pMfSZfxaqmlFt4MZJ
Z3ClvnaKwTHz4Qoz61sw8hYBUNbKtJm4XurVJiahcU0HHpJmjIGIueiltQt0f1oI
M524iP576GF+pzcOUCBNWljvrU8mEyFs9oLg7MmJ/TYr6RqcuiP0jFTBhYnKLCrt
MXE6Rk+ek4ChMedygPD/37bv1ydSJsbq3OvOo5hON1jJKxyFL+ucNY6+VNySbURY
zB7XKhCIGndLQN4tPYhgMi+oxWN4Esug77djod6pBfOgaWV9JrZnJbc0kLQNGP4G
M5tdIjkArIWbAvxtP2T4OvUIQXnET5EDuf+JxDFVNYl6mjYX1gFnI1E8oxlW11PU
jFv/08VW5CH4EL5W+LjzqNdDxNeGxL2t4M4hySu+IxY6ODSSvGYCE5qf1ClUwuvP
cqMpmflECC6w/iPod2QFZ4uMeRoZQx+6z+4aBYH4MsUie1scfelcND83cItj3vCu
XeGI/8wm/sv0tZtEGZFY7Q1EdDKfnDTHfJzMnciXKRWs39uqdbPGqNRV0dhrxkJ+
vjv4LqvVAc6N7CrOkquuqnIbxxIG0DnjDwzWF2KH/cpxvp2P8QwMyII/jsIRN6GS
ZgjNXLhJfrvGHfsU1WlZCpzM7RYRnReyRgYvrzmu1eqyQnnHZj3uTDtkY4Rw0dgw
4Q5aMN4lzpAfjegI8Q+lXUFiKGrkEbrufL10rfwA9jyFAU7J6c6aeUcQzknjnPjd
aFVEsNpx2lVp2KdPrB2BfEsVDG4uJtj54OzUYIgaZ7MpRxlBVC5wGXfjtsSbmJ6M
KtQdK6oj6XYmTR9T2yqE0knnzRwZK2F6GmhjSRCqwpYfaET08Bkrefcy1bBM/aHl
JnaVQirl/XpY4j4ijyNf8WL5et/scBUod3ellbGlzGiaL22vcSvvEECH0FQmI78a
9K3fywY7RfY4Nbjma9C4Mbi/gBgzmhGQcVhn+/FrpgXPZmSICFLNg8vS6UlXeyYK
UsWdMgpAtxs6zR+BKkLkA05faa4h/Qc/VtCoGPtu338NgRDI6fIRhFTc6l3mNzz0
xFMjdewNkQ7uWq+IzaBbJ1JMb0K3FmfIRS7UDRosXJ+X4vX9ToHdUxUT6wetm0Oj
PNPK9EielucNWYv8VUsa/loSFe4pdGlAMtu6oYKkRZwTJxzYaci37JxCbli0IVq1
TYb52WWWCQ4vAhB2i9AHhm1707GF7plwrWmvp5IldHmN3LRnvnxC2mhVvhvrT7Ud
e4ND2ARF802iP+3e0sFRGkaimnRxBpZz9zjPgejVFK+7POwYCT2WavngciaQsM4+
PJF/78Q72+6WbiYMf9MRD1prKg0fLuDQpTPm2FdRs2tFzUBJ1Ocf5WDTKTaOaWz6
MWhaLhLH+96nAOhVtLqmKTMhngOaxOwqWz3q6Lzf290SgZJH9WfzkK3dLJNwxN1W
kCU1md/8aScIhV4j45gP+g4hkDcjXd2gRgAFEsrVJ+9H2+Jae0uWtE0ZsQqOtwA8
pkYXr3/0sD8ISaEJfyGs9sIJfv8CDe99+rL1ALVa4GXbTlcVdk92my5DkDvFw676
UQXK5TbQnjXRBZkSrhwYGciuh85zY9lz668IYnYjNk4Im3qmLK71UzGAeGnVAcDY
dfiwQOX2nuNhDKTLN4JKu/+LSpUkTwR7Sjgn2z7jLr+7hoD+MZJSPoAvz9vUazwk
R5dXJY3G2pro+ucEjVMnAec9GLe1HL9N0FWjX2eboXMURUzG3D08zhbiecpH7985
CkyA4G3NjbOBlgC5ANXG1RDN8Eh+eb8Irb7gqBIUaNJE9jneGECPhlMK7WAqu+k1
W8bMRvPMyK5KF5kFTQIWkb6D5UbR8UZygC8em5lUh2sz3tNTepoYMxy5cUCV4u/U
6pnKobl5jmT06SqmG1uOZmQecEy6fXJPu/LTgCs9jCjWU/23scUBWOz9evG+Q7Tk
MSMlg1A4wy7D9oRD5ITdbmJZwzz8j3fJotuX9pYFXKu9h2rTruqsYXo5/5g4GaM7
JkzW5wYxwPRyko0KrY3Qs0v+vmZQwfKBSoMndFvpmNmwfbk/jCGwCaQ+pcCB55n/
Ftgn9GWQ54jxV3qEgmsJk/wIYfQL0NVwqwIVvQuY0KwMZh4WjL31N0ZBnyPh2aQt
HRtfzFNRUcjLdBAV2JM5ztuSxnkixbIMouL9uOgUQuh3Tz//GEeEfVGk17//Pl2N
iZvwttXV5eZSsatj9sVs3R0eKvVdZzNOKTXg2+joj++7NUt/blfcZKrLnIiI5wWV
qY8JbqB3DKHEHonzFuzOe6tfNhPgZah1NT2gLEzRDAVlVqAtHohAWKhBJqo0Trdi
1QDLqntzauFTMqExV2ulAvcIDt0DZGSWSMuMZsikA0SNBLUTOYhLUi3Qo9bc3d3v
SIPb8IXRDbDg6H0E3Xc7dNOUORohfUhIxxHp7rMyk9+6z3kwAEkEAbfDM5clhwkq
tZoduehuzhzMCmBEZRpl4Vfef8G4ebkKzuGNQOr+UQxUboXqhQ9VmvSrRHmbD4CM
FXUxx1q5qfV0Wdp0TGi64m8tPVhzVpt7msIAFjdRfVbm24cicPHHVGCRM0U8af8N
mlMExXvGU74Ixy6j70IDmt3K6CeJ0I2CTYcvwaLp5BJWLYIywTzmeqLuzBLlH+j5
e6DL5bp2XfIwprm0O6f0NYlliUzgIkV/76b68HkAQMR7qqMy9+U//Ptx/u+KVcPK
cu3wt+EpnMa4FHGRES5VWt67xAVpuEryIDeTJPhKzuPlWbVDuhWHH+8GzK04M2Nw
fa8p6oohCNCpxU/bbjmoljxPk39e2HOo5gy5qi1nY0WoJv9g4XVBdSzQHCPEJAwE
bu6fgHKKQ6BgBhnLADV8kIle5jOgEalVVYhBxm0yRI8wPmVkq2A6kzs3nFAVcPBJ
T5egUHX0ls15z7YX6awdm9kZf/yd7/RMcyg5rrml6SeT2PJ6zoMAMryU8ojE1c7M
qO8kDNLHLe2PZ05Y/wVQ5AfrGAgvFsDWJFxhXbYJogIrUUXyxCtzc1BGDzwz+lTw
PBLLtqWtDqMmNY+X40REu+S+2sD+sMazrKgS0O12Xhj5h87CTaEpPWadyQziQgXU
Y9Dnr1sHGtaK1yItLNy1e8nFkSF3nkAxAN7SbApYCpoF8iCzTKWKXhiQKXR/ykEr
qtqHc2FD+uiopxkVICOxsoSl2X3RulvssEjziFtjKDbO4Id2NOktIBwN2VIKXC5o
Ktp1rxJEed6FstUXu9tBlzGsMoFhE4QasNeMF5vafdoAdD0ZpepJr5bKOdSabnJf
AO3SjjinLJzJfyRqs9YeM3oEaguLujs1odcO/4QDdeTBeGbWqDJejDxdT/IXlp46
5foCnTV+kYZq0roAHsFhU3ixNuqYV3iQEjk1QCu5p9odynFcU5YFhZ7gR4JWa4W4
SfmlB6f1JIBH0mdhwTwedn37YwUS4KBClPLXgRXzHmFiLuynZSALEJo2w7xHzBG2
+tVJ3/5zYGhgG6S7K/FJuv4kp66bLNQlgFaeTvY5X9ovLYFFPfffXz+zJIdwlWPG
xoVblwICY9ZfaLrlBV3euFqtt1yh/HEviD77KfdHOeho3Vu9w95qJ3+XhWCnUX/q
p50pW36kdxO2sbR5DFf3jAwzSmQ5itctBgN3RLLQKScc3py0JZSiFOEPS9t63d90
4Vi4/A9OvX3X9rict4RAWGwnIEe0tKYVNbqZ4HasxDtmGe0/zge/GERUwLAoh6ax
XRToGVUrMBfVwlGhYBrwIgZ1RcA4Oy7CxznmXnYfVzc1N0EMfnExvJ7wjkWlpM60
VzeWECpaDHKRayqg+Z8AwYAzGv7TeyI5oamgSv6AMtdvbnbxxXS7Qm34Hk0Gc7f8
616xSJLfdcHCjMO+cw0U8MdN/RbYLbZIxzhZMXnBLo+n8kI2S0XQC6EbUWz0sOld
fdVlY+Tivu4aK3m1Cs+xxiDQUfOLsHBhePBh1kmxkPFOfQJBrBHAwi/VG59+IwIl
kc5l0OlheP+o5kQYZzCGK8VVX6et2pi+XvGYx6Nj5BZFI2H3wmYsX3/EtqNsVIYE
BTp3rTOgzX0Bo9GZJseF2r9lni/VNMsATWQfYWBxiSsu0tn9G/6BXA5eUAYeiRkl
XxMvLeIZ4NlhSOfEQGkIuG/T4IkR/D0+KzAZfQ0ntcgF+VkoSD7lysD4451kKarG
03Pcmjo/d1Mx3FegdbqD1NGMuJz+bDGv2eGs/qqSGf47mjmp0hontIw96bUM08lg
kOhbtV6DMPr35A1bsxYktc1tjtacnmfC0BnvpJKpRT7oZGxlqpMVGHjDxjF7hSu+
u1EGvdvamqsjaysHo7kON6r8k3Kvc8CKCZLltYX1++lZ3bSibH7LvjFydyEH4gZv
64AwfR1EBa5AJIDAjbe23We8+/MD0Sp9bszKxfbjaNhDv7Erd8xaxoNJMupkDDPg
vCCNmo4Ypx/gxLJF+H8kvb5LRWXaR6pqSg80Xu4oQYgPyomcImu3bGrs0LF3SjFG
njJuogv/0W+O/s4AukEwr893OGw2WXedx5P/JUBO9R6EQ6IxUvDldVDDAPUMHI0/
dDhvRJWU1Pfo42gwxgY0Il4qmhr8olFOSi13ki5mTC/0+drARoZd3TS3L81gzmCl
QotIaqrpPakTvRxycexQgjECaDN8anwp54B2dC14vIMA3hdIAbHZuPicD71lS08Y
bee5t45O818RLbeomeNCAMNbPOyso4NoXx1AGg5fOLLtko/i332rBrfJTTkLurR/
jK+yAHscMOM/82Ue8ElkIieNhpUz3YoRnskGvHJFlbyD99/dLGv79ofTkv/Q01e+
Sb8wxxdyyLbP0aZfg0z/rKWfBULLNs6LlkJblOK4CVUPtfrgq4oznaLoaMb9Lrdl
r5zHl4mrn3IOfFhtXjNPicMYDXqTKLVPSaC4MfIF2Fz5AdThqt9phudBS7brZKgk
GECXEz2jVh23aBYkGZPk8l/pBBbmwI+fgFYxqcbTZvciUtEdrYdlrpvVFmv2TDbF
kUP8H5QdAQR5NBgd3XVp1kgWA+Ph2AtY0nEpB6ZxeA8qLcBKkSS2ikhPPzZuA04f
aCN+evP/vp6DJjLIpvn/mfRh4eefUCckFIOz3Aw9eZp40ChIbcPbLIQKckxzPN33
r9l/iYKgjhNvaHdnoQhVQgR2wmYEvf8FSSsWWc3EKTA1yNHqlKjWIK/p7qcLO+oy
VuJ6EMgIGOeOGUGAKIPCu5z+0i9sXKSTZA8jp0oBwWU5siuPF/M6/tZsXKxIVTkt
11yBz3GcEB3PYq3DkOvij94eOKYWRdvlEIHfGyZrlMEuXmtSBaE0NchqspFgZxuk
8QPueH0X2q9bzTMApYBTa16BOLH3NaUSqU1Z01d10dNadHj1dMdVCvGoKvELA6n1
jjwO/b78blbVXyCurJXqw57fjDHn7/NLpXFd0agEaPLqtrrtV1v+p14vxsRf19Z9
yhtNBgLYtsXgX3wuXoU6qa3u8kuuuJt+tBJjs/k1ETR8a0tH7dDeMxygaYmnET0h
c5fGfd+YCQte6iYqJA8WTubyzZWVzFA73XKcLX4l8f9DihNjQtJyTgBCPbho67An
/cvftRNlfWM3IpiiJcDUPO0hEep64Q6ECbsyB1noqiZYMtjb+J9YXMyRkuL1JeU7
xoqNOo306tV//xgxeYHetmxv8SX4Yu2zTs7oKscU4YjWq5+4XknSKqO+EJ9KTBdS
6wkGUNavRWZHlOEYvmJ12qWWqGPkvcslCoOSal4R6aE1pfpoPEe0zIRPqg2/Isz8
4K0YBJQ35DKwIrSZ49JLsFWpzlk162ux04OASTBpL/EFKsHdk33PxKXcG2AXJ0yH
BKx6HmpRvaZCIt0ZgaC6VJVuxNVYfern0ZIcvb7L0mHHy4x+rOqVNGqchKi72seY
kk+109p+rbyv/f32ruPy6GIq5glIkb/LlAmFOK7oPljnNIm60x1qmnsXQxx9m/Ou
m/HKZT1aW6FldMEjPkh67I0owx0xphXhAjUcRTbzbiphTRdmlFYs2XshcwDVKDRd
blDr5diXan9DWoOawIBF+U9KgUR2IG9LIwU/9B2hLeHbFmQ1PPt7yznd1DVHISCk
iStbWVGbMPrc/CDRP4favuC8hG9N3qnNvaASzWJI/R3tGMR9aBlKOBUbXUm0G27/
7zAlKZaeGbml1BmnrUADu/Qf1YvNBIXfEuDABth6WsZtwx9Dwn7oEQOyCBJqArE2
ddbP/z5Vo1uvm93VVAia0L64XTYz1W2XzIMWJ1am/SS2/gtP6kO5DjtIf8xYzR7e
sNfJ820p+ybQ7lWZz+AdF5dtKjMKIWpV5ZUJ3+8rhpQ8ru/n4scjJ8GaGI1IZxnr
tQWenmS6TW8ghJvn1E586jpVmSsWcmps974ktZwRCVIWlvVFpdtW3xZQQaQzirwN
KdZ18NrgeS8RAq+DTa6I9I6SeCi/mjuL8V4IjgjxR2jpZMOaq3Tl90IGXtbA4hg9
KvP9O74Lefgjk0HFD11fePGLNQaEZusng5oRiwPGLN0DBDcGTBYsx4u0Wgx0ytLF
cLv+CHyheDu/ruKd/E/0MbCwINLsW71mcR38yFpRJM7Jrhb0M1ljAU5s1sxkPCTT
DFnlYU8NGjZdmq1rTWFSFH2YBKofs7/nL2cDZPWt/fNNOzUJxxSgUQ8Ryh9ktWRg
XMcwPb5JhbVySB0EL5wlG7aWbnjdJv4oEK4wgWViQ7egWO0DvD3dqJb33EhLtNI3
T/H6i3+WePGtcKf0B3yZF2K6YKf5x7bMQb+mqFLtJG11lIdOaUREdGD/TWIdj5rC
rEcTJK2T+gCenVIl7IB/BjgPp7OEyUT9ZnS8FibaPxMvcgzyNuzjOTXolJd1QShb
v0ag2jiqRBMedxpZiITwruyUGwG7s1GcXbd/PhkxrA3OkllPDeos5w4azJlK0u9y
CsElmOYFv8xnM7eCv6AcPIJd0Pv776w0BoMclmwcWQChVuwOcel13/ZO3CXHyJVd
B8PPQw6wBxE+QD/e8y4AlPe1vqOKheam+G3j8s/J7sF8Yw1xtC5XAM+nsVP5DlUs
/H76NHPhLUrdQWtkkkM7NfnPUqxUDmUh9U01o+0wdihN0MzVd0dt9VvheqrjAKI0
1CAF2ceizI5G+qmQnir3o601Q1nX4/uTjYOv0j8LGS6xlgo+5Lt5QxqIhRclYARb
fNWX1hk6uYn0C1xMgxYSE+VDkA49/5JxnxpX/d+Vg2WCNQXWAKPfzhEa4kYuPsc3
8j+BSc0sC+S3/JzsAFw20RQ7oVyQoLis+u7mCPdjBsV/YxPR+wu8yzxofaRCo/G5
K+slkPI3A/dG3AyILD5JuUtR0CL3MGIfI3547WekNC7jBdjS5S1FoRXg8qmjdZG5
aqokCc7c7w5RzH8xxUbY1YNbVVw/pzm8hGfM2B1hWN01pRQIlfivwj7GDKkIAF+2
7QZMiQAiViBShNNcJCr7Qe3ThYWQ2AFxv779BJXuXEnzuxVSmn6SJFfUqpeDyl1D
vepr4aKO1kjzE2kHKXZoE0vLV7g8WQXbwcy6vzJurgTDW/FGPs1nUxuCM2EfSYDa
kbp2IyGEIFybEfJodlq73kJjgKiiZlj1bJj3nTPPyD5U4ml6WRCwZWFPjDuumYJd
/jLeX+gpodw2hWQaYKLRiHdotUpFz43Aiquv0U0ylrS6T4A10AtV21xR9gBx1+2W
Q1RXle1MRKBePfWhA5zzKiwarkLDQ8wIaLyQlnmgomGFcUskvbQskC89R0jmmN9Z
Xoc2igCLvqVkafNNUyopzq+9BfIRb7aaNa4OUK7gEPaOh8JJa7X62WvjR1fOt1nO
cx8hG6cPcHzp9qgVgMonO7Dx3d2v9GsSNNhAUAv9+uUyKJ3ZxmbHDfrC7ETL26vN
4pvZ2Tyh9/kxZZ3YERzSAtVfQEO5pru6rCoBNdhzraz5JXvnxJtrZT1nz02oW2LI
wmtrDmhRRmou6CqG49A1983BGBochCQcy+EMBCmDxKNVnLvcSrvznutKAI8F+Bn6
16CkGmXcHeUuKCGOXo41HmnjZxi0Hc9XBxm3643nK5XiJlpB08mBkmFpSmxN1u18
cilF1rguz3uvKP6osJQxctkfAnDkpC9qMPZIh7cKeWvl34/8miUhzazdH+Bnnboh
4ME+5jdHzFUK4J0/zFeiI5ILwcnMuNYnno8+uUxtPnRicosaeAAx+NrVph6Fg+55
x7Z1voQLkYFZ/hevypBlyKXhrOLZ9T+AAn354cgAuED5rUKFhx4/Gg4ldr/j2ciT
UI9BHS4Ir75yaI83qVOJCd93IogYMujT6gm0pjlWR/TwBm/F8R0sCXtNu8QFfs5N
qHKTGQXIds1TVBFopCbmbYWh1JU84CuOz+NkxEw3XFCcmpYGggWPhgwTwTX0Lalc
zzjnH9eZM3UBI4OQCEcZzWq4cV33aGAohJpD1+GTEOaxIBjm/bYuntBNZGfIf7XP
y84yuKj2PF1SMuO/O7XhxmIEumJ8WB88r3zXdIig9ATndSy5JYAFeJnaDHU7RxzQ
ffN20fnQZdNBX8IJSPwZIL3MvbmTc2qEbpWp+RJNv5G8t6KN4+33chM6xeCnvwGs
OVrq3bKlGrzSXEfLRUhgl0QNd0pFxnhPue70iI9dXHRLQsKFYYJS4ciWpj7ZTcAL
xp6oA3dfzeTYE7zTsHRWIiimdw7VuROPTid+mSe69uKPdqOYH5jP2waSz36Bpd0k
T4TQ5eSyfdF75SnXqQovW5AUdQ0qcv7NLzTG2Y0qxBDjIsJyNltEQHVLc/FxoUob
F7t2t3Sma8vWq61WQyLXmOJiNMLcwopzl7I8vtPrViet9GJ5TXusjKv6u6IEGUJU
ZZMCjozXJH4iv8veKULISOUjsKZM4mz0Mfh9ng5gqwLFoFCZjAcvs7UDEMZy9cqX
a9sxl/NPSkEAu0j4UoTWhKFww70D1Z3mxRd6HzAgU9uScbh7MxkLiwlfEJLxTKAQ
UNYKsjrivDbXSWqSitUhPevt/sajLo42Jh/mop0lhALPDsza7zVzYCJ9CfTN85o3
/iInjhJiU8L8tGMMWJ7eXAko/eG4AqLAb77xQy0TJlr8mWro97za0GdonDX+yldt
G1AAqV1cfBpaHAyIMGpIarh5KNkp4srk6o54yNwfGQlrT9HX8rg8lqlE1pKnfLSC
PpLaCU0KBLG+Xz2X7Q/U9olMJljOfbnbOCfFYkiK8vkCBzIfTli0lMCyWMHkvdZI
5E5izuf18fZNfcBB8i/psuAWuijxD7OXSoSm1nGGvsNd1H771uMFYZf1gl1ir9Ph
L9bxIaaczwDi22qTwl+sXdWX4DHSEJJAeEPz/yZdA2Z3PmvwLZzKtySt2Sbuo0BI
vodmlwHSf9LYUhFUspjEOwAbg/PCi9LAZL9OdLpfE3YREmVQF00KAx0Mj6v0+9Nv
D5Y/dILAS3yNePQqoWqImPvNpjFK1XyMi1XLtH7B+DWrvAM09bqF+Ky/0FiJAJQC
jsLjNRz+1mMhlkNsoz0G/lXPatg56o+e2sDCdgfSwJ9v8Mi9ldRjjZ37tctF3YOI
9BOgfKLe152orf6QcYelwMZMVD6lcpeqopYLNT9Qr/QZUU0RcAxekyPQmRazJAdl
6EW2lc+T4LHjLL7+ZSEFQeVeEIzDmFllxxds1YMdEZdD0CxZsttTLgN2LqcxcPD9
LuAxHA3SIonvRuE7WbJZRa9mnZfTWL6wCsZU53GjFRNffhpplL+Lq5lYB6U+z/4a
bWLcQTcorshqA8jyTs4b5sxo38/hyKjPD9/vFIRwIJg55ZS5942KPYvdUCkwpLIe
ZSQvaKZhPq6Vn0KC0t8midojYYjNu77jtHCdIBM4NKj3HTGC89GNvtA6ppcqcn+h
mHpjxuR9Xc3H9v3fFE2TQ8QMsNU2/+zi89bktL7MC+7A00I75xvP1PXctbJoHO8p
Hzxg4gh6kwPC8L9c3rgXHRfOiEUgAu4x5kXkRkHOzEc9G7DsbDaZ9n6OTd5HXVVq
rhj0Wlqi0A2XpDzOu63iNSIykZPL95HP+cDoaNndCGy1j0Ashmpu8191OVfH2FcV
HhSBr/+ezZfSdQSIJqHjiqK1ZiTgJYUGwH6D3uX6XF39v6TrziBVyl/mv6Vb4N+e
AYez3+4hIXAzS8lTL0Y+eLr4dzKM6WelZa5sYY6AApd9NYaM8Exw87kr8yasx+g1
TUmJldS61ClWCJ2NIaXuKoFsyRsk65MeOFbuEiD613q9Px8jmAvaooHLChNBMkcl
oItmk96BTPXMzEApH+u+3cOy3IEPqaBBjI3EP0b8jmd214Gpb18g5i/lmTvChLdS
1HeO7J01mDcig0pYi24lFQ8tvK4RiX0Dx+JtpeZIvNPJ/Q75GRfRoQxAPgGjrBwq
ceVF3VcjRuKXPAFkUVydYymM9GJagx0r06Yet8IkNKnRQSjkiArMggjtQCts/8JE
DpQFs+hPxMJaPaMEd3l2/AwwHTTRP0Edj/VsjYDcYWLGNXNbL22fdYkZTaz0GRLh
MlYcpUVLgQC20Zdg8ShulTCiIUWZ1+f1zqFl4EvV52mGrOQNJs/Pu/R+5Tyo8IDs
oZvIBpGTOfH7dyO1vaxPhcg8aIpHIVt09PKgC0ZKVowtBmzpZHjmXRz6dugUgMms
ovYa2b+yl2ifEv8FzESD+3Cu7dUP0l9RrR52l9BoXsx8PDebVWWnmucGklHNTcRY
bKFfGvRALOcnqANg+VsMJ4lNhIl0tkGrXXeGb73EziUdF3ExrbHCJtgBQUv1GeCR
hdbi46ev767LR/A8GQjhB5EpwN5kfEUDpyJJsMAHXe2gNsBEmxrBkSjvFTrbhqJF
9l8e7YYp+JogHpnDjPYRSQ5TRpH3ZHmd0hcrJQegASg7+2OmYY7V8Z8Bh83261PF
3LPEB3IEsOLBdavNrNtEd6T4BxWhcxR6s2+aK52Uf9li3FURh5g8Ej0Ov7JGlkzJ
iGV7fdQ04ig/4SFhQvLnj7zIOvNMIjoTgT0RBFYWn2SbThio7E9pkgy6lmKIrUPw
jmm+iAnOWBAjv9sImiSanyNwYiG6zykOWwb7aPHjeuihlGda+QOMsmNeV6ksO4uL
Fw6rOJg+7iUss5bK54wZ+qWQDL3p4kO8MnBEGCLzaTDrfqMEtfVbnYBhQAFzrbba
2zgchBEK9B/lxpOozYeaS4QlHtaePut7pquZGnp5A42jAlYjAd2dCdHKLejgtWjL
ssAIdvIFhfpu5Lh043hpn3DNDo1bCeekfrrz2zedkNZ+geV1cHeHnFzTc2S/+3Tw
yusIjqP7rQ4rMb1CKm9TrjcvuAFnODPQU2tUopw1Qnb0xAC75efp1x0MjmV5w+sD
2mcUKjf1K0PEiA0D4mhuXU3BVu5giVd6GF7wSGQDSfwLgTkLE5fxOGgaUlQrNwzA
KUvmDTFV2hIsUFlRTMVF91wxe5ihE4/Sqhou2wAbdUOHtsisz3MjgQwQjxFHshNn
UI97tuKdeH6NSUImdGQBURXzDxDy23VT6I9aJya8tFmylBXBNvVKvEjL0VHXTF/8
Kv5J5GLuabL7y/Niq91XWxcj4arWF6Cc1BhUQ95ihPIvzZA/m+11uz7hL97RMwi+
dFFgbsjbuaB1GMEouUt2tN5+hpA0HfB0xTpfCYb1FPs0qIYsHjFhiBCux04qMObM
YtFKhuf5ey1NGlXB25RnCP/j4bYGol1a13l3DXpRZTJTJug6h0nayMxeIvZMl/pA
226mVj3pcA1QTRWI6OW3z+LJ4QrrBTaL3j53FNDoJ9TO6Fe4L9UnPqjPnYOY3tey
SXxzkr4F0OyoKBbsQUh8QfHaJW3V+aNqH7Zei30ak+D/0KWJe49pGbcdblwDjdNY
BT0y8x9XURTRKQnruvFLZX9/bORsJIy0u9K72eolfZENVfjwCKKXyCgSe/xA51fT
bHCh3X94yKiUKN43cuO5TO4/EgbHxsaJN1HEkU73l3QQgmPBZgSyLp7B2R/arUuc
pE5NmPxrRLmzLaUPccoZ1O6uftyi7yE6J1UCFRlPIbRh8BkaWe3aFxAJbisCwe1M
IAtm9oXjbamW7GjX7IDmFbysYvER+0x1FLB/RximjJ05Jgs4FEUeKfR7qRVBgexX
YOehATYX7n62zsMVtiOjEFXPxIHh1kP4qnud9ok0MWrk1bT2L76y81qjYeevjh/k
/jhaM0IIUVUcedlzNmhU6SUPW17dQoKHsh+jtAA/E1dlzcHq2DXOiSvjSSAgz0Q8
G41n2StKsTNuKsSYeESHrDoOxHQc1s+Cgc5svo242+wyeRRDJLcSFJBaOdPQCYBg
I6xtS+my8SQWTRqzdEmE7N4qlh+BIEnrWmi+NQhWOeVkKuYmKk61qM4jKZ5g8gXn
rn4BSAWWHjFzwWmrJWpGzbkSvF0wBd4VbBJdltpvtxSLYddm59379M+4ZNOL4GJf
caICtcCGWRGPbnIvwQIWWncYod2MGcmS3gCV7UVl9TeKKZJ6AeGeJEjB9kF1RlPw
BpIeyQRifgGPuapvikPTtzU9I3OcA53mU+xfqDlp7MflPAq18vNE7/DLghLuYDGh
e2IYxKABOYZBBt5MriT6gkCIyld2YNeGIY5+4aSmRmFy5DgwL4j+WK9L2eM1Bfuo
QdWIyYCoaTPxhzOwBJzvPNCgnVTWXzGZLrL5KQCSDaMXpVgAoAOvtFBHcCk8DvA5
a0FzJLAlp/tqbOEH7j2IY+Ye61oXlXHdWRx8fk4yTaEMkxhNXweKg+wpzyDy6D64
yoNfMna6KyGvwdctGgKm8zvxX2g6vvIpXV1qZJVqdCv9lZRsSQAJAYpZHvHrAvFj
wvi9/JHoYUwZAVkUfP6VhLs94KNxHGw9SOYLjhq5k3M+kA/+kg6Hm4V1XZijpAPI
tD+DYiKne7lMuz+nuNjO9soTEnSp+zadudOpJxk4OnOQI753afaEYVvlELWijHLy
r4SVGFbC/4Db9Hw9ZY+dDn2P/sUuEefZGIPL5CD4HoGYl6mCE5HHxGA8SmrvsoOZ
ji1tcOoQ5jBOQRJ3OrriaqFUwXum+lxtj67AKFC1MdhMNebsekLKgKuLeaG8DNUP
t9+wUBgYTUdfjKl5GS0SI4j5Yh0fQSbBgpn9S+m79I6lbsKil/XvhOMlyOLRRjCD
KzxoxTsj+xS0OEapKfVrp1jcCOCPNzDVQdNdnNjGjYHrPfQNMZybB0XhxAkJfsiY
7M7jNrPO/x8DgGI6Ptwqxtj9hX5gk1P5QGeO7UFaKHqbxXf8Q0z7jrcZSgptmPx1
+Z0U94inGktpzR6QkkuQxm5M1GCiebVK+1MShh6rCdwxJqg0t/t0yRPU1vRBgMqk
NV26BQPkbIWd9tYMQllP1TbpvF6Etf6UADCsvz/mWunD/x+ph0D3gJq7OUbyzBPN
0VXE2HauyU3E/TjlDPO+vXBriD5//+o3k0utdIy3HySx3wUtSYH+xolZRgFX5sDK
qz19Pmhsc93UbJ8zXNy42G3WxamF3O7AZmQS6vmWAG4xqEJf9CosUVSx1tSZLNr6
5QpjlmRBW6uK00WhtYbnY61Nu9VYNTKHmZAL3PoHgX4hzi7dpAv0FuEZoOYxYOqu
ys0JRpyGVY/QwG1jeNMHBulk9CPQp4eEyZ/rpR3/8IH3ryfkVy+u9NrbjbGuw4eo
r7CnHyskX/foqhCuPwnHxT1NI7vVwV8eVZjGwwSmJYhtplwyeSnyRV8Jtq4x50Ux
ILu+iPKlazRo6PgxYOex+k6O+nm3mRt7Zq6R6jMax9HUGU/0EDLE+QfipXl+P3jf
bXnfdeQ5jyEWxMWSYOKCMwlWBYxrwEfLgTMHelzUh1uOvP9cQ8Ud3x2olzxa+XYk
AKsdyNoaqJHxx9fRmD19AkkbA4wURVrztPa/2Fhqlo8rzr9b6kPCgADqbCfbIdv9
nveWWvoOmMw7csl+t2Y3nBqlrG/41/Q9Z0xtSFhNRHUoFvkOkAr6bYFYazoQfqR/
yFE8m8LXUOsFYGorCc23IPdY7LsCXuXxAizYDjeiIGCl1CT2FgMGMRz80dcQEAfr
hmQXmPW/VY9+RjOvdi6/4qqrXbtJEESSO30fgOaJ4HkWrrjmn5FwpP3uyj7gbY6r
CMhVy/6LFSW8C092V1CTPp24+OHrjnFRDUJ7eXV0qbl638XP2Vvav65f7x2kjfRT
2XB3FEMovpDKVHA5LdM4/jqMtws0VUNnCMlnltX03JFYBvrYljiQigJNMGrVvfss
+4BLluO8IHWtRXwBffkfLJEphQKzAUYiF9KyPGT4/bgQo+td5hzeKNmVP26Tk4xj
sLIgabaut0r/uZA1JzRTBOyvjpUWcS1StydrGLS/HX0bYrVW9O1/ZYI33sK1ZfPH
dgoPr5NDod1vpQzpIDfyb8VZWTjo6cd6dShlO7hy0jqgn1pJg/bXRHQK20ttKoFc
IKcQEXJJDoK1hHS+TmSrp3NV5fYBgn2ZOU8f2k/wDi1KlCo7CuyIuOJh+IDk9rsB
9HUQFPyj7R1evxV+HlM51Fis+fJvfx0+7u0sPHVjwdWecQpoo1ZwO5p5I3gtBYHC
CVRFcChvZ6empzEH0cSlYfApYy00dkSVzNVkW4qnijR8aC52UVZJMu4tBheXtxbh
xdsE9HvMTrqzqc35Jss15bhxK2SMjB5L2sV2TKlhqj9svplabiaWfHiC4n6hKwFx
NGwh8TanXF3I/yjfgMOw7cOnXCzfd93UhXI2w2xHBhAUL755E8v2xT54piJEy0ze
7eaHCUhwFseFHv+glGpSTlArybuw8VDnOh9Ow2BMHYHC8ngJL5MCBVYNQwzjy4P3
iWFfgJfi07pMHXTQai5uEoVOCNlqt1KlugQDFLG2IIFYQ8pieqQclJw3YZ5L/Ahf
zXYie2xa6LFV83HA93zvBeQaxPCWvYqP66ApyjFL0aAvTcY590QsMh6ZSOZINYn6
yHVgxE5RwM+MsHXD8dHNsChvQmLYGs1tqSLf2ddXM3Y1wlM4YqoEmKRAtXVnSlRQ
GlsULnLA5iWSfEkyxH+MliG9GAQsBjAxy5k78obCtOmbbYexnS5A3u0XQcVxQfHd
pHZPmsRAxeOCwIXl7QIgTZfK0cymYANxg5yvgmWErJhKITHTtK+afaX+ArPFGJoi
YwMBriIL8J34pS4IyJ/iUvs38mhdjlGeAjBiyJAoiYOWtgnbE5VafIPUQ5HjgpCM
JzI1pd9RGJj6BYhH4aXumFAcoDeQ16JkfEW/E4kvHIo5VzasHbdLIvN6ieQ1GoHL
kenbpfRGpkkj0n7AOqv2J3l8OHfxYo76V53CdsbJjsmTcHfl3hBf0GRfcQ6YAkfQ
zLwfxlPYktD+p2wVwml9avJ8ILQouOgQcuU9YQf9DNOs5HmMi7aOzxK/ZErSIuwb
rtsn4mTIXQ6YgK85hrp5UDi20u8P0dm/8u4SDFzx+XMzc/ePySYmkzAG3RjgGLEm
ILYrnfMCZm9j0neTAFQXfHG4t7mvRd0Em4wFEzzm/c4R/ijidDUPUtqLxFXrnuZH
mZQh3NvSbXF+oUHQc7aiobY5W22JOQNr6xk2vRk+z6HklTnO95qp5MChAtNbgP57
HbJ5s1lzBJysqX3ehZjvaVPec144OZDAql3aQgqV4b6dAEj+SgSPzYPCoIwDVaJu
htw8dAB2V3lWSoj2MRwnA1uW+8VrhIr8p9pR07RZLG4YC48j4X7bHQ3dqRIRfk+7
K1azb2lc07wnICsZrPXocQX4ZQtdW54ShWVcWf4+4MGEsMkr0/YaIQgtj0DFx2NZ
yqM8ZygulqBpYe0da7JlgC/TwCZh4BWQuYUyFk2Q2IQ7sUnJjvSPSrD6/jWIL0IA
O5h3/bYhrMoCTs42Y3rMLELVBcWuSlJB05VoVemtKGV9r2Nz97OKYwqfLeQ0Dbe4
YTf40h4F9Qn0TdsHGOfU3+rsv7nCccaD5kUTRNZwWLlU969oBVXLFz57bXKe4O9A
AKeyB2NiWwDJMOhYiknvorYLNoyMTJFXeZ8Ay9yUfO90dl7mxgahFMDDolQM4hUu
6syn+OBBbrOKam5lYsHiItNz9DpvwE5CI+8vkd2HdnBP54OtN7loigpJSCpSi5Vc
JemVeE0URCch/W6gkCeX9DfddPFAGHf6N7w2hRxO3V6lfLfvcot90Q0125v9Fz7m
ZxjIgr3mtTFhLoTBCTvb0y7IsP3cEpdr2pl+onn8VWBQiBVuuUlpqi7zRzF+CCk0
fhxKzmcGWBuWuVFzdBk9PiweT2ToGn9G/Rf4t+suqsotKRI5JeIpHeQJ5SXwgfHY
iv5u76pd8h3TypRU4n8047D5oNlHS0bG9V0m0tJ8NR2wu0kOd8qA2PXuBvzBUf2d
XgGyqNzFcMb5wKoVDMoxf14bwW8MJ7eLWck5zE1aH+P/+TmfSa8NcLyS1YdUfmCw
XYyhUwXVq1xT654UG7sfXcFfq/NexnWSsFHSuR4wbkHAIp78dts/Uy2rp4FLh/WM
BzD5NG9d7ww7arKcm7uMcLBm5mnn9yLYHoGH2GpTfV7z/w6r6oJjrhQiMQ2iQWqD
Jn/a4fMXV8dhYPoecY5nqu+pfYDK+qXo2PEDOeYoEVdDRzA9RWbHqzhTwqo+nvQM
1/mZYmtYKYqF29Q8teBwoNXpKWCD/bbnXXjV8rr2UkYxA6uPMZmZC+BnLS7aE8u8
brSkZH4K41ZiQmOpmOYsJkELOth7EZQmU8bM1aPfvC24TaURblnFt8egNWaHV6GW
qU4jbhHlZYgcS4tbN5LcWC8IqMU2kDI5q3Fy/eonZMGRJJ4nHjK9FUzFRG0sBjDT
rMhg9KOmhFRL/bZbQePi2KltFd268AbHQtFG0rlcD3PB0EXa2ga63lUJPsUfpSLw
xcwIM9NvHVVDRPE4Ui0w87mGO2FGR09/njXRovFnr3RuvB83VVk4Ly4dFACrz8JY
oFJkEHzRGNZH2CJRzSwrqO0sLziaLyiXLP6kUc3KSBQA/I5a2zcTfJ5Y9BjP3zbq
6ocs1Aq/4guiVGKdX9PNiregU5Wa1w2BF4moNkZ4IUxEb9/MhRQdhGaSn/ishjh2
8jEm5u00fgK2lKB3xQY1tKV0xkejCrk6ZbY3rD/r1ic+iqpNdk9J7IWfVwjpnnIQ
U3RfDiw5nzHm/QUiaMZMiRe7XcauBSyNtNucCbEasHcqovnKOn/0g7yDEpfkffMY
QYCK7sfJBwYUQu5IXUQk5SWNOmtvYAgvTXfXd03v0sqAneyo8PoHfepZCl0dIlzZ
+0I6LffMZGKgmG8R3z+ZP+nnFpfKNbkcujgj1HPuVaE7BRUZyrXRC4Rjj0o7+J27
iop/ACdCgMKyLbx/KS1ZSrMuUh4eyenCFVDuVYFAgyQvPYw7fZNhXTJs2nCy6ZRq
0uw2WdsHSmqxljzOjDhmm0PjJb9fNffq4me0f0gDz9/jO7+YYnzhRdpPP+7snKjx
7uhF4B6r0bKxatf542BqY7tpNFOJDZUjie9Edh4vcS6i1AUHwdccxqiiX+5XMEuG
KcTJSeg+9y8Oqh0d26mOiuZka44OGjojN3fwThwuw3yD5CnZrh9ECIJNOCzExlza
/7BRpn2/mQKpJ7UidvJpmIaMcmigXh1+uu57y0MsY6vxUR/BSKT7Zwp/aToTM39c
SeUDqHk0kqb3Eo8OOYRWt9ch7hY61MI5HOuv4DsXtPke7j5wnV6N87Zh7Lce8A0/
k3qZhPlBfEO9Sx9Vdyg9HyNMl2lvtk3ZM1QewS2xAv2MWfVwLRlQ91DVQLKOMvkn
a+A49pzEdKrlB33hbJ59zBFym84bsUbVDIInMmUWdg9n/UzocGRCA/ehYbKglSEq
Mm6Q/znR0YJQ51twxhqd0kUJvdG4/ZFjkEtFbkjrurN7KFNQP1YDVV6ACsC/1rgi
a6i6sf0adLohXp6jP8C8ckbNMf0GnnyCkRk3KPwG9y/mhAan57JXGcVAp2R36qWq
cSh7jyowCAkrqleBZA4NLro4xjhUiNVk2K8u9IfX8zDYfnNnqd1zA5fNu02GGmXf
1M7mfRkwBLaqWdeQN1yH8k8OehW7ShNP43bXC14+KA1kLuESifCBSFWsCH/0DcIa
j7d5T9v773k50ofjCUMBVP0nxZ9E+YFlBbRlbwPkf0uXM1BHpi7ofEHWhaeEkEzr
+dKBhlqQLdkn+xa4xg8wkEf4cd5BAUPXC95ar/qLpIWvp03tH6uzY8azmU9j1ZGI
e2Ojjn+iAWW63B2f32lNU1UhSP7f1sAPortrDq/2BBjxweBplRSkVyGuDYPN+Qzv
k2B3p72rOWbwWAGKQtUMyxy1MXVgVsf3sYLzbrEDqqXSjv32QFwLGF3jfdp24ZOJ
/dyB5uWrE3tOcgMvkNdMmcd/ecDF0bXJGoLmnodJaq1IkOTVB6vzW4pgRKfxciMO
w7U3VJJ1eqC9TOw+9sIFUbdpXbEVsRqUPj0UDSqj3PEfuCLRa/Iwv25E9QK/dJlm
5AMgw66fZN/qMh2VEp7XG9nmTJVXCeV1kO1f3f9eAaFubBgCT2c+MHC2j7qr+A6t
nr11cS0Ml1fhzhjLhwPp1+r+gTcmeNUq5DnOAzG+a+YDrWEADBPHCdARr1y8Zhn6
Ygo8xWScXzYXr5p9Cmv28oShWQdCyjTR/g0Of4yp1nZWuBNr+HNr/UfU8/r47m8e
8x64ezc1RU0W+npxQ4PMD+7uzkqJ/hn+cZR26okTnKHxh1Wtnb9GiGCkaeqWHvBH
Tdn2imsGw5J9M+rG7iooVmTYNCOFSR88hJR3g/7299oWUnFg2J9fIduXYWbWHdmA
3zqw/it9ATCYyRCWvQrdNAcxQvgYB2IBcZTHriqfiJs0PZoMS+1tiO2ivvpqngLe
YHA97QACYGkgThJAOwg+5+yRAuV1L4/D0+sxoTULONuXn4sBNRJeBpEMRruxZhEl
vt8WqiggYsuay80pZX7S4LH4NfwiDsl/I6qkZlI7oWOo9zc+5bLZfWl8XsQu1/xZ
zDqEG09KdzSyhQJTwzLLEqsyvpMJYWM5ie/JydkiEfehBk7AY141/q1IleQJ8JLd
uIOD2YY/+3G+45KacIWTerq9dJSQpnjfzFXv2TIbBFujD8fgo6NBvkFna8mOyGrJ
XBzBRNmXuDaNgMD6ge6uXaG0jPttzy0Q0x9c1CcNSSXFNc1ZRZ1gaEhZjPuoFvmv
HLvFC+d3TmDM1k8Vk29lmAXrE7c6er3uhzr4p6nt1stHLYiPQei376g3D0MrPBsh
sev08cksXb92jYhCgBblY13U2jztV5bNqWe80fMHiYyyXEHCiZ8+5qa/ucVeKcdX
r6uqePqh55oAvTBNbfxLr7YVzmGfFJqIt3Bpc2Z86LKDn2d3p/z/eBLDmPXLw8+z
Soefg39+2wZny8WbavOBuuehtXEG9cvjQAS/bVq7UX3kUjkqAxkWJn38RMMZ4QNe
g5HFfPIIsJbVNNJ6voV411WdbkUrItyys5hKN2klc+K7EO/jR6UCTQ98QemXFyj9
oq4g+AJpsTMM9R0Edtay6Ky/lSt0/J4wncowMu3O6u2zh6XrGsy9oxOy/2CfiE2W
3g9SDVRT8cPTkYMQpuWCfEGwufjTtldsoGRcWgdxCMYAtzwV0YAbTF6MuOIkWcpr
ge2z8lIKzwcnDWt5yvsh2yDMLa48CuVKtmUzdI+Nzx9UoJeTDmnenCSz4VQn9lbT
QvBg1SZnTVWzXYsDm5STlqaBirQRtDq01POH+Zgo9TlvMfuwZMT4t+HhbTHSgxFa
EkSE96co1MzNXnZ8LTybIN0mCod24PR3PVc+bJF+21SldNh5MBwgdr7NGmP3smQ8
qAssqiV0FmheUlnJ4ufTzkDwY4015UEqomvw9SXoHii12Rh1VQWOvPUAxKc23ry/
IPMr9FZdkqwoIb+hoAuAeewP92Te3QBNgRQjusLxjnwA7MWMxiITX+q1eZLKb9zk
1ZxggDg9Phwm+nRIWwzlR312OxjnUNlZpEOQTH7aoyYVbScFtIAscKiVM3XXz2fH
L6QLhCX7p4bloKmWcWYdIzcTQS2FordKZrpFN9VDVC5UTigW1Bd7PePWqhkLdwtD
TXVEYIJ8tIkqXvY4fxbXrpAfxIsmjEOfCtIslAmOqcP4RUr0U+4znvs5myz5d64W
5pqp6iltch6xiSe4kizmhZsgRFee0wE6bWMAaXPe/c4xaQGcTZvOkXQ5XD78rJfm
z/44YrVLm+UdpQaqAG16gggfPU5aoKjSfryq09zgbvHaPki6jYzgO+afKHA10BRV
b7Usz0jfNxe6Ht8heGDalGsoS/G3E+UJn6gcFEgW4ibydQ6gnv74/1OvhCjB2ehq
qUwIBSYjr35PA5q8Oju4Uw==
--pragma protect end_data_block
--pragma protect digest_block
MC7ggGNg4PWnyz8yTstctoonEqI=
--pragma protect end_digest_block
--pragma protect end_protected
