-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
kZDVLC/oeGAmSIdSh5Mj3zfiW1n0gBuYX46G8XWpa1VSjF/zWj1G8rXV8QgyKfZh
DnUC5VIBzYbRjW/u/K54PuK3Va+EF34pS/sSVp09HLLUV6dM2wMAP2Rtabgml/od
bvfCbmHEoghDlmwREiJF55hKCjm5J9RqVAdCPvVAwwQ=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 24052)

`protect DATA_BLOCK
JrKy3jEMtDa3uKI0a0qLzNdzIle+b16FFVt61uwJmELGZIsLvFa/JiOUKLf6UOZ6
Vtf1pOxCWmU1TFu46LiYcxJ3WAMF+CvrG4hpVwmcdci8J4SI2k7S22is2GxtzGkl
WuQucXbluMx5vp+XfUXJOiQBG52V5rT3+AUi6aPk3RwD9YxHblL1BOPuWACYpjfD
byoesmSvvi2h4pVN+wzVLBKgJGeTt9MnKKt8dn5iqwKQbS4OfXQVG6CIzk+pI9vd
WmjAFIXileO71EOR9EvPXoqOwKppCY2RvUKRk6mWN5ULEKZWgFwSB6DG/X6jMc2s
Pf4wGDhEXoK8TZmJgqqjb1tq6l8TiyyODnfCUL/PC6DH0ihzX7zK2Ej1dZ3RU1qS
TNlrTIolAMRqaNo9rcx9CxBZMxi/aT3Mm73jHqbQRL8hp0bmJH/CfQ7qPYDTxWTF
H+kzEALRfK692F8GJcqWfOHqbf2UYOK/hXOao5o7zYlB+EvWWqNpw0fUuvnPJTti
pXwoPdiIrUSZVx+QGSOk0QCJhgPsqruewb7P/PucepsqElJwJPUbXGQZW8y1Oawp
j/DEM5bAiK0swoFMXO82wVJQnjCTN/dEDv5pP9j+PtJ0442HPeY3LIn9URqpCAEz
ajxrQkHgvHJHEnhJ0DYTv1pJM+oUAM9mD1j/uOf84BkRLDVMroKTNH0e0oRoqtCA
OWfVqNNIKRY0gvirjBwPUclr3zzpSVBhtvRD+bYEuC42W6uabVlaHOCoba9dbebN
+fjtsq+MGSv68ell30z4I0WzmHwWOKU0LlUofY2FUHPhrPkKw/YBy3rDzatuCNwi
EWLC9cf1B082S+4ugiKxcLtedi2cSRzLqA4DSs/Do424XuPpxHynh5e3WTxMMUgx
xnEs6F4OCHqkqzDmua3KT+ZhgfGmZRjDG73ive7jengaCfHErNjUx80y3t4TWb9X
afJNfPzdZXaJxDWj9AHTIltBeFz7vQ2LVyl2KKdT1EISC7B7/2hfcorsf3jS0+kN
Bv1e1MenNsiBAJ0W4BWmRVAbrbWurImYof+MW4R1PlYGrzvsl8dK4DrXThvHp5pK
citwlqSePkbScMTMSqsLqM/iBK8b9tYEDHruOPZROzEMc8bWhOWMWluHm91LOvHW
9GbsEI/YtNqhx8gS8AWBju7XXp9XKosFhwum4//wZZBcNoEVnc62VgGSQcgis5ej
gem3LAy2HAEuwlwGX+pgvoRvocWzhv9S8jTzamnX6ynNP7Y5LmNMMMSDd4Mlq1bD
7J9VKXIceFmDAEjDf4sptAojtsPzFmUqcyD2741af32bLQSKHNXUSu3ll+oQNjOL
ZPAtIwjKAX/yYPoah9NXZ4o9+5LDeRiBkqbmViZxePXIU+q0FFNZaTpR2W6GlB74
BTyAbenH9KQEGREhjXFnSYovlTyolAN6uwVn6oJhMSqiDTdQeK9QcRppJzL3yBDf
MA7RyfvtolMt+4SQ7hj95l24Uywxe4PSFQH3p7lnqUiGYPOSmqsPlUg7CHd0RYhc
1yPSqjG0liU27JLeQFquH744IenzVH793XZXN61HdtH3dKaRtxW41yHNoBdSIAg8
VC8gj9dOpm97X5biwWh9Ryq+jADvVzhq3WZ2+6Vt31rxRnS44HJugvrmr/L0LcOc
rU08WijpVd6w3X4HdQc4yzPO9ZG+JFM1NtC+lwXyXivvfhn5WFJ7BDFBEFlXCFUg
dPJiU2+orm4+ePBX8lssl+IsqmLEV5QlS5/nIRPH8nvQbAWtI4fzgLPNomfMQRXV
N2d5IvBIaVqgZ64lAx/L0gytNSDfvivfc6licHTY9ckjGk9DnAisnhNSdyss2bt/
mAfS4uY1pk9ZI3YlmloGSze3QRqbwCIi5gSQzQGeUBuKnK6Q7efcLdPRlKw7gLWx
3o+xsvpYAn+Yx3OJtahNC3LITHtFWjPnSkE7AG7tHcqKVhtVh5t1b0PG5aQejx6W
h6Nk9XQNMJl+p43MlRuGU4FrtI91iV0c9NaN41mhEmxIY63Jy+oTJitbylWcK2rT
YvtJvF84qkyFZhGYYwKOSnKIfQYFeMrEK2y/wj654DyqXRwT3FEfk/6BXgq+N2mj
qwFWWUK5sDaFraIDipa9HJjQ4edRzkJI3z7m8uCqxcwI2kssmq+MtyUa/HuXGRh2
fbJAqHrWtz2cH2kUcptq4NdqR28i/+hwe1/IxohX8jOgvoTh7zAEkTYOIm5TadQV
9Xe44GhuOPVQrbZngTC9LuLU4VHQqj/RS5uN50y8wik5+LweShFH9p7ju35HTCFM
IYOG2C78ez0HCHxWgG9gJ743Ef+YIrumXeFcdga/RY0mckSAd7577quSRevM9/tG
8cGCvuLmlNvtTxdS0R6KT23853SIFqhW9ZaPMAs9/Iw429Ydc1xakvocJ/o1RbaV
wopnU7fLr6FhagVl+WwSsERZ4HjAt/M8UJHBwkOQtRugE4NjDqcLVQprS1yy71K2
pKF+8iVSf1YmkSHk7Hzu59IZoLiz608aIxINEx8+O62qi+9LUKbYILD3f5ncGEMO
+Orz8GozjgAVWG3cMo0hBc6GIdbJrb/9v+6tG0JIiH/cyllwcS3oYn9wFgUdGOLP
JIgUED7cdKu4SALwLeCDVDM9NAkzpjZRagJbO22y2qVMogV2MAQsiSVu7/3kYtrn
Ew2X/AEDaU7o1vYrpU/LTkhbHL38b1XefMlmuU+uSlKcKOYYod+waUKTV4YgbMUv
Oj3b4Gwshzql2EpOwJdXyKbv+biwV2mN1U2IaYfOMKVzlB6q3l8xTXINTeCM8f4H
Hj5XdUSWrjzrUaGKw3GJJaPdDU8kDTLm7fl03XJqA0DR6qh4pI1/jN/zFqpArz9b
Ihpcm9kufxv4izonIVbJatRB7v6GJjLIT2ZjuVMtkLcfwOPNUlva56jo6rab01Bt
+UPVHERvdgsuDWhKYjuIEG0KSiMBzCwgS7vJE4UJMW5nSQEpcSqJTf6GgqLlf0+n
F9vMvxC70SoBLI369Qa4d8GDS3nWOcYBvz1JKCe136vWPcFDvh6B6sZhGiHJdDRm
zTGfewi5MPOyuLgrfdVSTNoEeNmPmGK8+yTyYlmgEJ1IQlSvBMCX5wDchUM2VC19
akWcSmcNdd7GPTF6nS94Gf876Zo01chkEEweIC8LQyc08g4FAP3WDxElv00OlSiM
TTTeyaXGX+A3dtuLpesjHTKkUYAKvlOI3PoOpjjek/F7Hsl6v8ZMeFp5hN4KwdT6
5iOtcXYvPPU0zdJzsOrUxrCP2N+sQaAvTjcMb82m8BAacsfL02Xtwl2avY9yBxDb
f/iVpdOpiqlVHm1HWwDY34HaJXpUZtyr/eekLVFnPPKkcaa7R+clIhubDzBYCDVr
XkuLfOeTZHcJiwHOVNqOfcZLbZV4bY1LioL7TBFyEqn87MP+4vrGqJpaB+Fpm74t
rZekX487AK7WyTT+MHp60eBSCYlLH2GJ4gEcmxZShw+g6G9oKbIrkEyTR9AUlApI
GmtbNq9qcaPE+MW2MQlJMGDszqeSdwK/r2K6myerJf9KBG1WLQPeLXwqvFNpbubs
lZ3aT1CE1In4gLBgQiSc8nYlXC87LIlDGwkUftOsh3mbYFg9Fy6RtlSxj5d2WaUB
/mdBF1oNDs1SLlA11HxrGRvrEYqj8yNS4PgpBml14cLpXlTz+dmQJZ+PKDLE2Exi
YmnbsgAcEtsQNNfk+fFgtuRwcBDGo//Y6N2Y2/W33FwgbgHV5SYh+VFxyElq1lK4
xNQHxA0xu+sa7ECk4IWtg1Oqlx1YNUS2f+qy5Y9Mhkjn/mSv9RWqgQYvbzv/oelm
wPDYCSuIZ4VrjoPtaMdlFDqaOKQiiaVabxbBAM8Sequ/fH232ZeWaXckQEpiEHPk
7PkDdAp+Cczmp4KvqEREGSL7um4wJBm83JproYJOF9yROmj/x8Y2GiZ87kpDEqUr
atYfwDrru4CzlkJ0YQo9/zE2HdqHuOA7KlJh4mPXN9LspeGGHtyNdfBFh2PR0TXD
DfadS2+zX39asBBF1y82Dpw2+ao1XOmn0Sh0zoX8taeCDpe5GGirxxy5sRvX2+iG
keN83MwPlacNkaO1ats55Y38d2vVnfqvwWXu94eaiQDQGkAMzoh7f5ltbdiXjj8q
NH/jBuPqKdsrUyPZEgrUUcB69TIhaBPdPvFrBPGrQ1MYIRF+P0EoX7yN64tKg6sV
HH+1RNGiuPQZxRTAOwC+rRPbVa3+retLjA6Rsy9wxjXUf4vHBn5/rQXAke4L2pVq
fuI/yZvyppFCtxqdOVkLzO4RKOny1ZDJ/2nzQKQoQiajRBDiW3LdvxxjnYhnKD0z
AsY/kEvsG2WP2Dx/teEfAfyzFqd4ZohzB8bGaYkOaZgslHTY9c2w3Dz2dwIkZEXK
Q2r4stvg+cxkeeqouTnJ7wex72rvNSu2izhfe1l6tUm4cWnEgvmQ+HKiNkShrM6c
jufecVhlTNx4xCixRzmgvVVnyS4WDsLLxrePhLZn29O20LgArbQY83r/L+qd6sWK
nUd/qFI2KOqISGgtmGsjJS2jw8pFYIAca7k7nQOar3b2j8kVKlL+Q91AxTq7VM07
5sW268Q30Ez2oDJpQlrzqP2DPpApDesBpZ4UlNJ4nztGiQHqK94doqkAJdq+xz6G
J/y/rh6WOat4vjWRX0utqV5CWFaQf9tBLQ/h7a1e18Y4rCy3/C+z51i2U67eNbnX
0ayywQFApesDyk7ZaVNGaJtKb6skT5MjrqhbyM7LkIPv+H/F076F5+t9fUHbD3bM
42FJQdzA1M/tTZDsLosS8jaXrrCGgUWKShsMctHq9ExJ80e+XsHNOWtryoc4W2Mw
6fz12lHIzzMfXmyMB4Pc/xSdDNShNVBGhKEQzHsvzopBY1gRYLsM5PZQHs1sd/+7
8qUZx2gKJO+wH/GXZ77rKsJFCboTcCXok5ScsOhXaESdknAo5PlnHIjEqisprm4m
JlM+uGwYRy5r5I+4MmpSIME9aK3SGEme07CXXnnUyLYLqjpJfR3Q3la9URWHiwZ3
F2oy0X9YfNog1onesSpo4Q4q/To0M8IWfY6Jw3JxRAQrafdYzOC7kuo/CaIfhn9v
JIAyp73ltzatt5kNZT+XW86G58TPjrpMlQ7iQxgOjfhn9YdWYhQG0dG+/6o5sHIV
bC/Q1EECRFxCLOfstLHLlL9RWs+5lodL33SkP3PGhSWqk+ShBChg3bV2hubFrTF4
1B9n5VZm/KBwcZkffAQlzEyhosQ41h2oB4lRGGEY/9w08RFOqteY205q63AbAYxc
3lMBQaNqJXBCtJ2c1lzKd74Jd3MBu6Xi3BFLhvQGBjT+uuk2cIGcrfaMW6SuQ1vn
+9hGM7Ig8F4CIRLf5Djra2igm1Mzxql+qTUhO0pxeaTIoHrqTyrY2o5SAew9ch8y
KCCqd60sVJ/daBmRNwo7QWAFg8U00CeTckDcRjG3ECL/7ZFQqV3PDIl8qLHlaZI2
uExLmv6FEXgzeTX2aABNWebTBv8qApEhn+uqYOlXWYXZ69i1VIhoALaAxTvQkNxa
8+85FPpR9HBLYDTWoM/W0QDl02TDdZ6OtuL2oKvjXsD6swl0laLjYHei+6VxNL0z
eINkdNC9Byhycls9TXj99UQEWyRTxrEhrUbO6ZDTsfYdpclEuyUJl7kZKNNxVYwb
xjnP/M0c36zxXQNbNDTfGUjK270bqWve+h7b01tlqdI9Kyu5MZDHOWBaV0l+SKry
6+MDZ9M0gDEOMzW+s8QvJwhkAtkVerAJLrIgEpOQ7uLFfZ4mN29nhe7KRoUnXBjA
BLCQ6JbMbHySqm8mmInELRAVK7qvo8c1oBJ6wipzxIfvp+UrBIVZ9r8wNij+2gBM
bwXFMgzgRsN2/c0AkYqNmvTW9k5lb3XjTS+4gX0HRw2Mt0qCEWTJOIgCzjXdvFAA
rCs3GeOug8k10wIus7j8xtv3SQur7CXFrBnB/5es4Os0yVXG/ZYPAO1fIhjKQPH8
DAclivhf7j0LRX5QE4hYqHhcf13i9sTKdGJuC8I3yUnc+jf2PbkozP4/R72ie+eT
M/2gaZ7UXnK9zw4VWbhEFYiqtp7O/xjhgtwJQI1Ghb8gS8gNFP672BJayA9Xj1qF
B9cUZ2c5jHy0PAMXUJGrkBqdUWboJPnzpPuXLOcLLfQsNLvsJIJAiDYWioufMGet
u88KN/bv4qRnMpDDKQ77FmKLD1zhgIebmUIjyQrInbAl7HcIXAeHWHTTx1JUjOiB
81ZyPXZvA5Ux6Z6Lg4/EFEyZ5FYUpTnwl0YLl4Ar76++FeBF2rg+FiARqDKKHp4a
nDkJtK5KMIa1nKtevW4/iRsDgJXtSvyk8tzuD+H1g3TH8VttvXhFct03zBQfPrlE
Mnsd0EN6NU2Kme5G4ZCFLQgAiUL6ijsSWGzzjedZORxeH6mfjVEysGLGZv5EUwbT
UQ2yOsk8sTDORlreQ6fV/3+T/4zzbz9NLELWFoms72cGHcXRCmiDF5KCzH9H67iP
aCueOg/+N7C5lUGhUKnggBO9YgQHo/RxgNCN7E78b31vi0Om0P8ooc0plF7tzYZQ
HkYIhubCN2NVvahxvtX8iI8Aln6h9Dt+v2LclvpkllPAmcA97DrHFj3hPT3y/Obb
9u0+gsp4lVhpVAwk2xEz0DK0yOi8jsWwJMnmbppGDC8gJJiBKSDhXpheHSNkAGsc
T+Zz+TMeqwCKh3yi326+JndzLSB3yt2XKlVb2Bhr2t4tIHP9IX5uK6K0VAG2tnRy
QICUoQfdIPlTq0c8UaWkH7BborGemHiBHEmV4/894Y5GugM9YRA4K7rJPRzzroIo
BWu5uQUc9aHcWpd5hzBWHi7aF5YKzOKeilfbPTYjXCgPv7/qzGV3B2o4zLlDcpmT
YNxXcpesFMQfJD1Vyr5EjP2NWbECVSYJ7+RRis8XYpkVf8acDDwZObKTk7/Rmomr
UNDeWRZ/bQ4/aupvXJiaOpisVSt1S1QEBBkGBZLAGm/2HzR5IwuJnrVaR7a22FUm
BIZVfkuOF9moTVs33St89Qm9VsJocENsUwPwdoliJMee8WhpDX+9jj1NfAmgr1xC
lhTVc5at21Mz7Du7FmraxKCyfo59p/qMhW+AHM65hFpa16JIxvywOOCVtQ+S1BGS
Pwd1ZN7DYIng5FpMGBcVf0cHNlPXpi5TjJfF259tEBOUJgTuEjHsfRjn59BZQ5Nr
D+WSYeJ86JIFMIV9Klc+5CM4oX6lkY/h443TCdWQTnhSE1OYxPchboaY4snixaei
ZgJPedUNhPAcJfpWF89P1HlHW8lgc64pJzDzuIFwjjo4JpXFwQyMrV7k/0XiS0SR
2qgR9etHbFtRDEeN5PFL3H99MGXEYDZH/As0QhAfBxpUrLApuiEn6kE3I0tlwNae
iClrVplQlu6B3DxULG1n3Jy8M2jpAHBPydQ2wK06LN9f+yCtMtOsNMbsieQMaaB3
waRxyHs0NB9W6Y2og0RMxhQjyIALYUIFAp80JllbM0wqvp6HbfJ4EaYwPRr26i3f
JT81I4pBk8Q+7x3/g8pYEfb5jc/YY8c8jcEyhcbwMInrOghwDT1Y2g84UcvPhzIf
uqabT13t8wngJf3XVgKwfKh98XGfMdrQ1hx52bxCksg2JsjsxJuN5Y+gckQ263/m
UCEZbbianlCsZg3v0vXDYVNXV2MB729uizy/21vFiBDViv/pXv7zm1BIkWCfmW1a
PP6wum7+wouP/b904lHm4ALXRs6f6jJVKMCX5MpOM3LY+WbW3eBzJ1M31GpYPrbs
/pRHhY/64L84wup1C4gL6Xi3yMLX0lBRph7b/Z2PkmZNVxE6P9YANbenFCqmL4jj
EfJ0sK/sZG3lCCvPuKhw3R+GAsA2k75zHee21lTL7nnoBf5g0xCulwSOTcVd2Apr
G6gv+jUQvTNYgNlClMCrS0ndDyx4JCed/AcqT+vKx50Qpveh/G7h5cEChU75wmny
7EUhXSOXPKdoe5Ny8UD4JVWWW5WSutyig1izvBmPpYWMmJmmMHclSrpd2XlfY3Tw
1tkW5vPr7vGKfg2W6HtHXbyAt66aEuBvhi4E39ej5pYqeKmgAOymMGnLli06+NVh
JFHpR640/VONRc6bN21uvyqi2o8Id11X8OnmuYweWdQsNZqXZY+BUW2jWLGofP9+
yTJYJARLvCcLBiimmZK1jT4S2ni1b0idYJQ93luYYh2Tq2E4h+vOBhpk2ReYRpE3
EbRH6a5O+FiCrtHRiknMwQKEYn9rp1bcZfDSztak+5x09smbRQ0ZNzJeVu0tVioj
icXJ3ODgYfsPYfUaX/G87X1cR+GCtAOwiCQKt1RIX1EHpCshT3moze5ahrtbVfYB
Z5OR3nqup9lJvC7lAq2Qjfy63Oe1CYyQPLxxWC6BTY8O29ieADHxjAkulkwGcQJG
/McOxFWTlLaKKC0ImWG08TkI9ex/rwe0YuEzlXIi4aK8BLatGVZYGCl51641CWuY
TEgcxHUlLSXnLqDB+RfGEFPR8rvlh8WpB6G1w3y9I4DY+h6ukGAQuIQ08o7eDrbJ
sOP4vZhjKFJ1CmGyo9Lcz2PqDT//sb1S9DBBRCVyCyzIhhCUhen8IwjkqhTWqLKr
iWP9wVzxWA2QHdv2hvrhtSQCmZwU3x5/P+/cjQmaRMXukoK9oRPLJdcSJSWhUEBU
XyCFJs7DAfNQAqM/W1WzXhkLKzgZlvtvVDY0c0ihMyCmzO/xtcz/9HnaNX2PiJR9
BZEv2gwIib0TEJ5vU1fHlr0RVIUEmMLXP9NXMWbSFqDh9qnAUEmJ8ltnrn7a2Xwt
0B2aUJUqmbFMFlI8EQSIwbyG2Ftmu/oZybwf2sI63jP4xoFSAy6lNC9dyJn9yibW
YEttXtVarN1htRZ4SKHe8sZSFt0/ofSNRyd4n/hOSQ4cvRVyNz7ELZABbUoNRKrM
MvYDurZVFmjbNoq67z6wD5VwMkZ06mZqQIIGTQZ64Ikp3hikntDXLALJO3T8UCuA
j2s3dHuAt4NySa6Ure7wIkqiHbqsvcaMQXRWvx0hMJigZ4qumabjz0dwFfsI5Cko
d+rN1IzwvFLBhtc3YFRP3dPdcEr86s7U4Eqb+0UpyOzZmAyz++pBKhCoToJlDXPP
unMPJ3OFC6lcewjn9LkumC6cMUjhYHcq2gB7tMchfwhlq8geQ5yKkm048NoPtjB5
HmBDKvFHeBpmSdBAl9IsUllsE1HRGWHwMSe2hX2yBswKxaF83i+l6b9JHO/wCkOT
GHuWx68InVAhCSiPR6qxPBu+8+NN79uQ9MWQ4q09XKFP9RwgHEpLqiHwqHr0ZA6/
+fk879Ea8LXkug0kZiTnF42tHBvFkvUdHZbxbzWb7cpcAOIWrMWsz3lX9VnSLjrE
BcEm+Fjxa1OS8pogNcYyxgksqgkYWrLNiTbfQ+O50eRajHu4MHCKfUTzpuTDvk7G
or2SRezi1p3TDGrGQ1HpbvRaddElGY6O6vnZXCDevA78hEoif6eAcQg0RodLwx8H
hoIPnkAG28jAQm0i7WGGIm8LRWOeHaIj0gp2UXh33b6zlrFnonXD0KEI+67mXXQy
lybggpSk1YX0ZOWgpcL8dXVQVc0PKcz2dJasyovZ5aA5zzZsusJ1X3TyLZ2gcmu/
j4z2nUUsx+mlz0iNAhSSjGCxW0IAFayZfZWpnes08mRb8c+aMJYVtyvypvfxlMBm
E2d9/SDioB9CnBvgh8I4vICzIctE6DsIrR35ukFBSIpvLTiy61JJzz2ensNfHkO8
XI/U5J6Oy3/OKsi7qIMAvyq/QipTMRrqwVRE03Okm/aL7K1NLCJUe/zCdN5AVo11
SLfS6vtC5UgDB2BULzKCWHNWzUgedh3xsVQmYp+i1v3Hcx1V5FJWH3Im30XiPeDq
nGhQvsiIaVwtulENZaZR75CoGEv7zvcwSpXRKPvYarlgaXvEIq2JmWo3/z0aOQZT
yMZKlLzf6AngaBOWFI7kfJdgf+rXUUGyiGBAo9YSI1kuLO/ZDDY817senwALT6iV
OClMkEoLTDW/CYxTwiRTuUB+sfdz8x0antqCu25YKaNNa9kn8gwRSeQKg1Gvraqa
3C0OjlpBaRITODLQ//IJvQZttrSLAebycVVhO/u/OGdQlPyVrWBBry/hMV7Xm1hc
r/vpk3jkKfC6IOczt6b8JHLoIQDYhtMwhxUnzvcBg/yBI8Zl9FtcWGrheXrZUHQf
A1UbhASV4rTVaDnfH+1vJJ8YXj8Ne0DiV/bweBrbMWmsgHpBL5mcC2e9ExArC7JP
6cWWbeeCOM6lIeP7GZTdn+YNC9FjGOTZmLjptqAy5XIM0nUG1FZKYU+Al6Kgldd0
L3jucZH6LbA6V1LEL3xDVORREHyR6q5mls5RnM4NnX0xIYq8qh+DBN1rQp6l/HvG
h4XQKnKs5tlHoTj+vU6pvhia5AEX7u1mN9ffZSxX7lEMiFZ1X6Z1pH4gG0Gb4+7e
EctiRCruAVnlnyZXZe3oIjOcZOduv/7ZLxn/SBsvCDd52CevKtBdKmcdGAZg1S2g
f8d5VNShm1+jU9EBuTYtRsta6uqwxGZKNp9AZCp744f3kpdmxvpq5YcJNQ015Mtr
LK5reynXxZ3v5jRwwLDFwAkdhCwsYYCSGalg9OQ9NflvEpO8zlBt6E/LJx/bMECX
98ikkgqN4i5p6Ho0z9XQRezt9+Znk0SNjkt9+6bDj3nQrFUnT/vPH34wFtaRo+13
mIK1+CozKcnMKi3fRb0Gug7yGQaar1BE+x+sPZOgQsVoBoLj0OUl2O7EWD4qwAge
CmdYf4wf43q1n/MGJRS8QN5bucUd1JHoAXxGB8AlT4U0Lnj3aiDziPsov5xD6c/p
UAqw4Wp5E5qqe2bTK1WKnI+FGkv1BttDFREgKPMsXNaeAH4Ee1MW9k8ZWmclJMSx
XLu84eqlM5rM+bm5ScnOxIryPRwX8+1ZGLKHsP7/4aK7Zf5wDHQZFy0KSs9gJXN5
LPQOl7EfO6ybbOClvolekNqrXUSyzr9k060vfyWoKkZvymoVf0ga9yycP4e6t/ag
31GTdB+mqRy3dxg+U9yZFTKflgx4sK2rD+tsHNeL49vLo2LT5+oL+hMdz0ggslsC
+x9RR7LamK/iLoJvtbqzKzsnXsrNCv0kjVCODBqpzHudtxfRtQHSd1oD+MGWShLM
Hwx/p32TBvBOpfGjimaKcOs9WgbfxTlaOOZpuaGoHMVfMIl+YFJGMla9zNp73Sp8
g8CGczh5MkEYvk5u0lGGsWr2i1LxCTkXvo4dE1zwgBBaJs2xAd5fjrhGw3jX84Ku
3LLCsB8v3/WrlSmOjnvCyRLIRSy8BEtki6VCOd3gj2GcpopqXgTuQCmcVEiiBrW6
yI8cdi2a3Ok37qRPv7bk+jKmkdu/iSOzPfbmV7vK3YyckVbfs/P/L6yekf6RbyTW
ySGdQ8y6LjsCOrzrML2fOtFJl2/SgW5ysLzPdTQBDBdOekSaMiKGG6VrMbTsoe3i
GI4XdE4I7aVWf0CNcb3FBSyOLUfV5ftyq5CvCMU8T9h/ID6IsJg4YE2PM7HiLkO5
tM4I52JpUdzsXTShLLF9JmQExfS61RAL7tB8Zj8AfB5wmakyvyYHE2KscnqddSe5
ldW7hdJMQPNqMdEmcO/Oo9aBIEWxCe/D+aOcfya43oHmEPVEvJyD0n1fawDgKYiF
S8oOjbbUkb3uf0rQoeda4vTKdXBx13rUDzq7e6Cc+KGL2s35oucfS90ig0HfltDt
n7bTXyX3joGQTpCwZbEpqm4ic8bZ1bB0WwV8UEag7tSzF5latDvbZw1UBodTFwVS
LmtNnETS1yCarySkXfOYUxBWC8ZGBjguxQ1E1rO+QBRkEY3NeRbP3Z19GpofcmPA
7408a6YkP+BatB0pVE1i6DymHK0Vp+Tg/TOuEttBTdiU6G5YDTYLbVu9mSp0UnUZ
pjDkL9uAMBjoROURh5q9DN3oSxRxlkX+xHuqTSZPRzDnOHJfhopSV2omSzQTkzZf
Z7NS64CURnEG/Eo2mN4IQWUF5Oalr3H4sUuxybDcAyuRB01uD5ukWudNRHnPK9jw
3Ki0kUcFhjmZU+tzyYfQS7UQBNWn1eSfMgB6hWdBEAx6VUQ7jQTt0RYTN0aAvzfY
f9VqosnakULqnr71KmG9qxvEe62q1nUYW6I4rlDqJDe+y+uE27z1D/IqOr1hnTpo
FMeDeF+LHbJ6YlfQIwHUyafHXxHUjE4Ocl6VzCUdNcxyM6xjB2DExE/0RhqMy23x
xK1ACAA303ufYfMvCgdtxeXvG7qih3Wi7ifRYQzGhLcHylMGxZ/YIKF1NyWMIRMh
FMrrdP63UICnaocYQxpT9/SL1Dlr9wyNsDNMql3gupk37xTv6YywXEe0Eje78GxQ
L6dwcZfob0igyLHscs0PmlIVSsDOGfrjmWRoFzE+sqA3JPpjA8giJG9ffGRhyN5L
8+qKzTANKzGDnxVUE67LYHxHuFtYr4vR2CE/30W6Lrh4KCQY5leJeiJ+AivhB2p3
FrU6s2GsstyEiBpKllAV7uyMhcUo6UoJrjRsWscJ+WkDrA9t3n7jrX558hp1yfF/
SQ9wjjgT//+p7DzNphDVmvsJc6mGeaQEPT7CdVORKot8Sue7m65whmaUpkli5vFb
kSis0bvPlj4n9z46/dttAXaWpev/8oeiwrE9OkLtm3bFbFRZemEaFCHX/BmvN5Yl
OvJt9JJuWBl5XzcJq+G5fMGwCHt/WjV4elK2UgLQFCkjaiGT7DsdMNtVTmK5Yd16
c8+VObN5Z6lQKCerob11vgmiUX57ZALiCULSZinshI+H+Q/FBKAJCOlMk7sd5gne
8eqd1pX8FmwlXO7VWPQw2MJCVJoDZhNaZQWCwLNmWs37HdHKi5m0bOR9OqitGIRQ
zAogFo/H7wjJXteq2lcufjKYirGAMhprbrfTZyAWTIxAFeAwucUwsD6sQqeqTjmM
GMMcalRqqC5dkmQ5ut68esLhu7IdYCM+yyXZsJPqB7DgisIT6+ll7Z+jiiAvE7R9
jd9qO+0keeEU9n0ZM4PPqO3S53uLMaNdPH/K/f47Ufn43ZKpM4tqHNUuA/OnBjTU
aAU4lPu1UnlJAbN74KSrK2XrOTGK/gFG/GaSFFITQZ7ew/x/kqp4Gyfm7c2+4OAH
gzuzsmz4QOmoy7FeSb2Nto4S84YVytDm07OLE1OI11DrZh3UyxWWVV3vmoj2hLeV
XgoLWbonkhYVruWJPR5uH/DssctMo2iIrEPUOYRLyFU05TX/QkyP1l2g3Sm9i4ZY
BXWE6l+TQrAa7TkrB/9VRSzk2c05xPyT/sefX5lFmSs70UJE7Ae85glYd+GFllsU
ZD5pWi+49Vp4gdKuO6C+nQkUV6EQjo3qMsiohE3JXxNnXiOa8FqFe68ZCXeRQHjq
UGe04n5IekAtUafiz2Txh2k5zW6HmYDkWccBwS1xK3j/x7DNGAWhsoIz0B4oNYhe
hh1cpTb4zzR8/hbDiNzn4oG2gFB+syS+qt181JMgZ1D2gwzAhNno5i86KaCcFj4W
KQY2Fhk4QLrwq8VRWR8NZSzdLWtSbKMlnxDsKBbbEe/lvi57e6O1DtILIY/sW52S
Y0Y+AkBL+BT1KT8HLvBIhK14jA6pn6rMdlPUQ7jDrnAMjt4GVvPQRK6z80pOxZaK
Y6cnyG7k7fN/ssZ4VTe5e3p2TlxoSEJLmCrFaMP6fZjfCfP6gofTElT4MC9WmFyi
MdpajFd19Lrr2Lf6bseqY1XPzseWXBu+7DvTvq4rsI+xhf5IXdNrqQmRgzjO2n+R
J5TMsbG+HHnNlfjCvolzUcxgGwUZUcT4U8c4Taahe4WEhB+v9lqJxNBaY2QqOFxD
OEoP8nZJ/L/PTbzi3ko+L+gtVFWueiGRlMEljfUJXhawTbCpfYarjtdDTk6aTxMx
AcUMXGhB0iFh6yRbBrCDRuqG/SEcKbrRiROtLOuxvkqsGX0GFY7Hi9A1qyL7FKJF
tnvOSMqzEnMZ6/OydbDbeAD+9ljTJEArrL9yidX7KoeEAdscKwxfpzDtZcRokFqM
ZzrYkoJ5Ku1iZwoxp1D5rXh835vZ+jKtF5QKjeuPLQkpk5WyYWwiSwEgDYgz6Uwm
isahlcdVCTLbcWuDxmFuYrVyH4G00OhNbcZloK9Y+zbAEUeQWmyLk87H4kbz7NvE
fSxhkHluHm6mdjaMc7Jp/lV64INLw1l1YQ8BP9dTYpwOzuDYa9zAXmsDlpSW/Zj0
XTOzPbtSFUfKsDOhL2vI/qfT9POLH00aRmgAmaX6DEDE8INIXdJEFaQcjjUigNuK
92Umxu2SYRQr0ePFUNZGqJyjknQ1aBfr+vlzPI1tZVZmexjdDnx77I8BVH/Zegen
yu26XQ8lcTqteA8peEP87+s2byY1m8wCcBg9wNF1ujaSAAugflJ/K9iwrwbcdPTE
z00EtLwBaAYGeBpInlYx5i9bPcsPTaIr1O6cYYkLWGiMXtOeXLHyWvjGl7QiHXbV
1TnsrS/JNhMO1G3T183xU9FjOBmivjU37ZuN9HQYgv1VuCQbNAY0nmCLPQdUy3QC
WndWseA1/ctGW9chLlQGOhCOwpo8tjXq8ShOmxTD1W63A08DmeMxMSrDq5JvdIGN
WUgfCk5/uGWsawLvJqtZyNU9lx92ZaTSJJR6sCX+FbYkYzuYsi1BOuKBPdbu+SSH
RzBVbso9wdQxzmEGOmdd/DWi6hIYSggRaKSdz2G9Ry9oapUBeQZ589PCok+EnlS4
RtKwVIj28MzeG8fJzj8v1Q+jz3VSmwFbatFGWyPH1djZ6hE5Bbgk8JSfa3eTVKtL
0eFMl+VaZJCE9O/sRdZPrf44dBl33WJ0FpVyaUCglqW3rpgHJc5r6cn9zN2eD6pX
ex60QfYlJyRqpqd56si0GK2qogBmcfSLWEsOF/YKmL7mzQUwx/cS9GwzO+pjtqY8
KZCNSr8ByhrNaArA2PdN+PS75ZqJzJU0iSiIX9bnqC2K5Hk/SpD2j0Vl0rgOji22
tkSolfsZ1HcHf+mbjctAjaTnBh61ZkgSOyF6iaAh0kb3K8JkKfmyYslHNVtwaHqM
BsyIlBaGIMfLY+8fKhX/jFWAZe+6yDTNbL6Ml9ivcJL9ommQGhy493Uvwy+8r64q
l0/F+ZiZ3U51xFef009q9tsgKaX9wE2h18ceVLYAObSZDpYGmbJkAnE3+eL7hjLb
Zzrk2sZF/hJIADLYydWNZcc6w1XOENIt05ghGtlbxxkmrAziNP8zUBTc146l2Snr
o24w5MH1YSAz4Mqtz+KCiAgRV7bjW3KE/+ZlI69Ot+wxVqQqF4UCR6z6KFrJ6g3o
rvFbxXpw4ZIKKoDpLY6fddTVdHPmqPq4AvVzYmX0e4t9jo8H1qw1YvcfW9NPtdaM
SlsXY3IXrhxJ/UzfUmN5Oedi2CH9bga3tROM7rL1QGkexYl0yKe2VcakKe8eKmCZ
nxB2PkKEcztwbgH2kk3r0ASr3Tllw/6jAcAcMkG5epbRa/Am+LnGbBnt3wsQagWb
6zAx7b1yu+oAKo7HFobERutQKKDNTEini9AuCpN+/407xyTi0FN0d70Z7IhMppRy
kVajcZmq+6W0H8p3U4uvDn1EXR8ByMyptFmjse4jeHDVj4F3yF22f+cVQx2WxZaR
oxmcWQQGvrTuzRF8Vl/jA9YYFlmvdc2E45WBlZhJLz7Qy/djud0YJzI5ofk4GkPp
peAMcy0m19YnkZ4mhTDWmTJeEJLp+tcUz7KQh8BpKzMDnppFRgKMdBdVEuI5rIbU
/EwvStniG7KWBy6Mm+uN+JMayxGcUlCwY5CVBF8HX9Qj7Srt+h/ZPDdpu9vEDtdG
Vb67CG0aLxx2eCAynSj5+EOuUw/Wt6Er6xhXtOLYeDNhvcEta+eYNAZJOqaYYe+k
FNwwpXTDBjPg7eay6lSziLXPca0P8ZIRFnByiZ2OSsraStczaeS3h78E43/GLGgm
Gnu6cxkT//yDgaDiq5pR5ftcQgDJ9u/8mqcJ1+Pm0TM1KozFgyqzCP0nG8XEfTiS
HNVofw4OJ4ePW5ks5KGx0V/U++hvNGHsXr/SZXDxQUeAJki9RrZfgstywpdgPIhh
Odf9zxikYEnKC1gHOSIQ1cfEORMC1BqS4cRoYB2f6AC4IbbSdQVRsZ8lbjxLyEmA
3XUYeYWaRveUaYdZMzhT5ATTnYbWUuuktwfITkS/SkaoYEGc8PeK4n8MFOVt/lx+
ojFtVOERBkmoygt0m4Yy3tcsZ4tFXjF/AZGRsTgkLPbC++EDRYtel959EGhW8Tl0
R03ktYOSbLNdSfF/xfeQOKzqf0YgnuW5mj0mM9vjf5cLzzSgRiHELzUI9BTBNTAM
3MFv8tpmBr5taMRbUHuRfY29SUui4WofRQaQzyrab56yaER8xfH0UkxSleli9iek
nCq2a9uYr7K8L8ymNZRYuhaVnthpn+p40yGIPY53Pvp/n5y6bVKdrFHe5venQYer
ijNEU4POEcX2ForeSic63s5ECgZs1WOVYNw3MPYQlO06v48bp0XOWjCKOoEJ4ZUP
1oZp4o2KwbrJeMgdmDeWbC15Q1qTQgBgSuNnKqV+RHsMwuqDF718Y5Mi1aaytsjt
kFV6xS1fNiwOP6PiE3+dqKX+hFJkQInMWLj4fvwTfhtMhjnpsPGJjHBreA08uX2L
FMVTqUzP9ich2hdbzKVTc1lkMObfg+6nqOmfRJlAXEZiSwMzwuDmaL6O5lA+XwYC
wRYZmf8IGknBxA/LdSr5BMdMjk138WZFjPWmdiqsf3vK600dYs6gr+EwvbmxhAwc
sbHkmQLcDtxizUGYLRMxtNTbncS+IorJY95aNAR4pZoNANXx/E9cMNM5ShsmsjQM
WgoTgDyvE1MPEk+OrbUFDkDNMFLGnmUlNoVDMGVFB3/BMDC6b20rq/4i1ybeM+MX
D0a5gXX520qeMh3J3MQwYsriMW92Gf2/z+b5LjCj521ndTRbWOeKacJFEz3SvFKr
MhxFn0KIAcBpjWRnbfaODdOQTT40AfHG6ks4fOJO/qaszP2kpymuy6AdLxNOK8/y
+3D8xiDgxv84CrKrLXM6Pi8cIvCq+5DmPlGOjduOEA0zvx01XWODfrf93T3+L/lO
XwJQ+mcmBqOeEH0TkC/sg8R9QJ2Vcm6bl+p+Kx+jzE6OF0lWWrI/EDdJDSPz4zDM
ceoBlnkO4gJeFeLOwuYe5l6QviXzNCQllPh45f+6nsgF+dqfptIwaIZxP3Ijo5ON
FNXfWgQR0erpCKGDkCrds0Z7etZUrGurABq/MA0LpwhtbSTiuTarbMCm7A7icFxM
FRdrcT6PODrILblxon0LT9T3CHl3n+YBcbHD6VZ0z8B/6mY+z+7ymzNMR9dW+3hP
8GlAsC2T+HbLISPYFf/E9rCC0ghLQgG400UuCEu61fG3CNTOnmUHXpxPyaQxm66l
SCVHUkTsyf7satC2NDFR6KYEYXnpaEhLPlj95B5YSliL4xFEoM+Mh9qWqwpGpIAI
PYVhsoPQTouZ9rOgwaBN8l8Dhetra4EPLcEdxT8/ZoOUkT+DjzEkQMUxsgopkGdn
StzIjtQjInELuD2E/3oxrjqaiXO3mIPY3x2PzgyUYF2wUdvT/yd9CuFSo0dLFUR2
dv3zspxO2XaE81nuW7e3TSZAs3lKFU2GGaFDNzER4KlqDLM60rw9UXQUhNALyqOj
F9qVqiq1Kf9rxdycUH2JGd+VQETO7e5hc91TiGVKaeDqOX9uL6AoGP9vQBuhpgVH
3dhluwWdAQLr9wS1X5M3xcuPYmCAJumF7IeKSnnXzgCI5/W5SF/zOMv5beR3ezhq
0LOrYJcpOjvVdhHAvRturS+ZWHpKrE07F+wvFS0+dvYYTLGPDdvFGf1kSn/59qC4
zhOVrvxT8HYzTsXHXrFAHA86jW2ixt7hjqk7mDZmVM0goZBqQqHqrMSEhgO55lSa
PPW5f5KgdGjuI+u74UTwC9dNFpdDn/1wy0t4xPX/Bine19vsYqx1Fo9s9tDZ/MNf
ckI95hGUbCWa1cGqWMbiymAk0UlrQInsoHOgnA6w88t1nfKrmJPbKwlPnu19AZfb
td7QeaouoPT+luXkrOkFxb/HEM0T1XPWbUwaiEAIzsxOX2QvYEoOyMT5En16cKoT
+Gfdg6F0HGb0JQBIMNHs76s3zopJv1NhAplLTI05P2JjSTUFAlqnuLnDjW/a8Qm9
OTFwziMyMlYtqKXX/vmqX3Py91+6+BaKQs1pm5yEzkCFoT7zRVvKgZhYpxyuedMt
XMFwTxj1vVb3KkHxOjF6SVtsDhrgdLEgR6tPxwgSqNHozfwqL93sghKzkL2XRdRY
V0Smqri7qDQFAzcsEgOaJKVAxPYO4aMJTc93FjBP0IPoVBInBw05lXXDX2VAgi78
F02CkAlLXC9hLu2Tzl5hpGYYpXHwAkHYW2EaOinCjOBejkqE6ON42edsTGuOZ/en
hRVfWfY9SZ+pGzBjpNhB8DseVV63IHwod0QpfkoJThRzQtIOqwMWNNs1mYseH+qf
mM2owUc+n3ZeFDcmoGw4bG4TtyvcLc6Ve1JZoCcxktecpIM8QVdTJBR3a+RjpHXf
H+zcvgYmmH67k8gMkZ4ysIwTWIXprGfruQQjS+pe6e7r+o0nxjwdY6m493A6Xul+
Y4FGNRgoBTAFIOoPtASHyImCfIwsRL+v2WKPe1H6Zk/fCtgHzG9iCFJpIQrzzGa6
muc/Rf8v1hASRig48jdNsZeFmIxyol1/5JDouesXZg10SNhPtwGEFocMnYwyHrV7
W176arwbB9Uuunlvofpa0uwrw+hp6RsDk4QcPAwPboTHfthpSKzmThg5IOktkerd
nAkAPW+cssjLLCR8Ikwz2kFyYu68Q88OCi9iBSdVdscNsiLaJHuI9oMEs9fAE/aP
Ga7oKxrSFNzkO1hwda5Fov7kfM+pt5EC9VDKMhhRQXKktqo15ttJ4Z/W2/SqB4AK
Iym1nsG3KcCqDjzus4tdnO42w+XskeoADpAIsoGYDcP2z9zE0HDVd8TxlqIK8Pmp
oKhyAAytHTX+Wpyym+xKS/es0OtX2wr3rMWanJPNsEsDQftSZz/IBg/zSbUXZa/J
Yq9cEA0GIvPiPEusn/Pf494VcBA3w8lfcrpU0Ie7mEpJDoFQNF3xs8CTstd+b7Ff
phI5QBDnbxIVh5Oc61vtubXWE6C0NQVPWwdSI35DnR0jySA0qRQSkNevEeHyCiAz
kmWO+NgRFa4e9o/eRaQCCq1iMRrvEUFTcw5s4EIbvV3SrtgXWg7V2Xod93D7L3Pu
fm4yd+0HBpvOFjIDBjypOXdlOdtcbrJZ+a5OUxvL6tjW2ugp3REzCma5g2Vvmmcb
9auagZQOSgZrhPP5rT2V0PqegIB2Rrvc4Hkkk63FzC3E5JlYr9qsnhkPVpvlpMuC
PfLvPY91HM9Pc3xQdl5rSgiQL46r09WjIWSbalHvKkfTIp702Tk6Dl/4/TmTSo3v
y/ut984Sb1EVPGI0gRQ0hmRBxQfFTTNJbV5Fyfl9Lx+UShsX09tDD4PM70bfYXdR
9l881WXGzY7TYGY+Mi4LRAzUTLKnPTSaKLyU9KVw0PD4Ye7Eh1LDltWZRGyJvJDb
li83ItpzhiLUiOaniL2yuNO06oeePOGglOnW1kDoNQDJ01ci0fAqTz9lBU2xsWWE
Kzd267UHkZ4KPSYkfydCfKRwtt3IabL/8fmuGtfXvcTZz4QMec9JQiAGbhu/P9AH
0dpVytCQQDzMjNIM1i/pH1bbiOULKAThmDXdFvpOEc24pwT83vXbYa8UfTlSxsmM
ru4bcw1wZc9UzmFUZxwP2CXMXSXD+Ulj+igUJU998azKp/+56DV50NEgmLcbaCpt
h/nOG6FZ5ZLe7rDfseP4ysN4lNX3y4vbAjj67Uybpk/EJ3f8inDv0BIvSHvZBelx
18fzaOVTDxIxjlxaUTH4iStEfGtFM17EdLJCTyDyYVu10+/rp/jdhT8J7MRa12Pi
r2CsAdpNFtW0MujaFTafOXGQyfustMbyM6IQesrDdJnq6E2Vo2vawwnrfc/zLn+a
D6V5iWkwDjckIW40QJcvj8vv8aORarlHTyKAb5AaI3Bh770fiG5xz32V7C8nayHL
ewsE6yf8+6NeXBwtHTZ7jV6WHz13kEfsY3UODpehawC92npjcPeBF5FqTinvZV5n
afmqugarxvUGvCWUX5Y4Y6Mk6iCKCAs836LyrNu4X9FYLmIDw2U9iLmoPNh26Nam
9p+rFWCumCnXvCWOOPLDnKONpJM1p2g3W4l/tkzn80wSVk7EjXqcqElKzZYSXdjV
2qoNZ/pGBuOrNmo0C7AJqViYiw2GIiSRBIxYLDAhXBLn3mRDw340OydZQwfCIbgO
vus/XVKCqmfeDs8KTuC3IpoIajytT2E4ZwjwZvEHHEn8qUkPFES0i3axz9btQP9C
vbNtctFwHNOJw5M9OGZ5vihjQxT32uZBpQ7R3+7AFBMoUL9Qgns0+m0Rhb2PiR6x
QMWlgyNTvxCCFGv2Yl+Asn/KxezfuI7LluZxqAn7OutiUeAv8mGaOSTYdRXvuslk
J58sMFkAZR1H/oH7bJjNzxyqhx9JSTKLLPFGiLadg3RRaom/SFLzfnwyOXFWlUu+
o/3ca25A0ysUODRV3cb3W6lg+Te3VWhAP5ivrtH1aXQ8Ukq10BN3SdsI/guBKbCy
TxPvNfTLquSVRJX7cZ1aQhL7pvhmzQVaAl0JK5ZBuKE44QGx3davvIuYwp2KUEDE
blCJrt3kO4Ea1iTRy1UTkqosYuczrzxgJGojAbMC9sx74DHJv815x03RMVggAOGq
eHdecrZw04fmKdrevnxAFLs+l100aouMqpbtVjlhRZ/f42xkV1ML4I1JfI8ybKMK
eUOZTOxNYmN18kGaJ8c7g8NGFHhRclwtNI3pD4wl3SuzvUWwjSXLvalAd77EAE+z
//AVJ8B1S2F5KFdSV0WKsS81UYWVrQ9BT/KtibNUBbYcBBchZf50L/lQ7+ZngoRl
25dxSO64LO5Y0Pgt72Dyn0yLk6JqGq6ps5jTOR1aeYhpb0prUwtmYTc1eOGIimzd
lxDnLL8xU5H8wvLaBGjPzOZKulm6RUT1magFWyoPMvXfN1mpJNWozc1u6U1BREHn
7WJ3PB5zJortgpV9rlA5YlCMoHi4syTUFROa2O+J8tLOEVJaICsADzbd9USF5eSO
MecXOf7L0MEqU8GTt6wDyEl/llwmQ6eT+E83DPRfYOpIlP1rETA2b2E3nPlBb5qi
Rbf127BuVskKRNTj3zk5u33ZOen4bIjUZMHBm5UKSw5SUOUOzTZNQVbxYZVRJga+
KVyBUmSqvs/pyPrVhej3RueeMUNgU6Yvz7hqrp8II2HRoip3guo6nx5nhjOnv50y
Dx1FlPAjIKP8dbAvd+F2oIJb/AD+xCu1U0zfXQnqwPbsuMt1YuFGJ5ut+6N2Nbsq
4kGn0uWwxSlyeNRVJjAb6ftZqKMUjgUWvTc/GV7Y3kSl+ZYrbOGDhfvTDXGngpXk
KPNLSSDyRqXOiTk/XXhoWePzYypkuV616GIkOTE0r+D9FYAnBF/gNWySU/rlVXI5
JRq4Sic1j7rP/MDTTqKQZFcNpxZCC3Ckbhxznz19n7m2TKvGkiag2xmh6GKrt2U7
UnY4gvP6lY1oTM7RItIYtHwdh63grdVMJDze9zWZ8sLzwA9SuzTbpGBsmcpAF7lf
H3nDT8lXKXIudLyNl3v5AwEvnE/svjiVikqE7uPetzz9nnkylpZKLaJvJoAzsiyS
0ddv/ZWrMvJeSNBzatQhQ6VLVD2u5BiCh3k+0TMe3Ig/SRF7X7bDZUVcsrldtkXN
W1U7GPLa7kAV3jh8Fp0ScrpGxvEp+XT/RYrTruWzaHeEMKo1bKA3lUkVVKZuGXeb
MAaYxlTW25SW94gmGF2mvRgLZutnCLCkDJXYGV0k+pYEQ0E2hEHgFquZntDRCmec
pzkTPKa4vxqin4RnmHrWP35Owkh0Oyg2sBUUZPBaJ3B8ZIJbyh+xAgbxZdU4wfVF
3Xl8kuqQO57iPHYGLSOe05yUFWJ44l+EzSQmcVFEqTb5+1LHAQJkuFGJfxheTDvO
lznwghLVtJ6N0b90p/Kt6NiS+4+e+nwkj8K00u1LHOAYcynqFPEtPafMrcpIuNnY
iWlh8Q/glSkS1EoboznZ4O7eOZ89cRFeroUratETbuuv+tdn5nTM0QY9xAxthUN2
Ssou8g9pYL1oH37maz8y36Qi2BAL3hNFSrPxtIP7Oknw7og6Begd/QrVSPfLurwn
9pcadeuEIiAEGKLWfptZyL7SVgHiY/Or2VysDWQeZJKjn4fVRnD9VqwznUz7NjLk
5oRoM+T3Tk6hioRnsKoZPCvdzUEtEwuKDud5vkk+u+M13yyZe4QRGMkyBGEk9tet
JAS4BLTIK/2bbhVtqTW1k6hxZy61+Mnj8RKYlLf6KrdNzF/E7jTf7/F0f0oeacxT
6syhKPOE+4ftnPiE12imSU2c7N0RRdXQf/szYuAjXMYGz9Mg1mKP/QzTJOwZzJ2n
/mB5nV4VJrjZ6L0nu01T8xmOhV5n+98Xl3IlotXXD3+CFYmGf4MwtSorV7xhLDOL
kD+XnUXalnpNLWjUxKnPBOB6YmYDkaxrII2wXSLN8rpCI/2sYs0OdmogW8xGAn4q
eZZugxJE8dhYa0dGAI6AWTQlemdlaUiYLLi+Emp03RRbjdzPbcoFYQ3aHY20HpP7
LYkiMs0P4BO29kkQlpcfcx7bEHbUL4S74n1UVbwFbhxgfnynVCjL4P9ck/jDqM2P
sLZNU+hsOYzNSbUcTdUBU24NQT7fijhb66niSAqwHEB0ClpJbZmkXjNIlCZ9r7Lo
xldI5NPg/r9iNtviLcobkhssZFTvFivtkeSTTFBFk3tZG53j1J/V1fbkWMB3eVm9
EhIE8GbIIYR5QBk5NV3l0eKNSr99ZfEOy1KTvcOwRgOWmAgAwiPf32ZBr9QMqRdp
JnYjRN9J0o/fa3mDL5I6W88HC4VdpzJtL+laaK7VjdnYnhztlcCf5R5aPJbC4KY5
CrZ7HVI/iITBsg4KsWKm2jbtmvecsKO0Ad+YR3ZA2Zqd6TcdReqndyFYDVkX7xd1
58ucVHCyIk+uI86FGl96Sq84ERg0RW5Ugf33iOjCcACWPdYw0yOVDMHwcDSIhVRU
1iQZugf9HfBfFmcW/zH2efDPEysHRX1fpQ/r+0qgrQ/XkM1SgcF0CjPnUbb2ic+F
ogMoGkWkooO6y6FUZS9DWTi3UasPR96+6l/AOS4MIx7fg6JI8VMzRNorbznGheXZ
SUUTzVgiNlCBORF97C5IsR81vTmlZwmSuj2G7joD6Quqkk/6G4nXikkOlkjovQW4
ZR+PYsV95Pm9Zr1G9BQAH3aF1TqGoUoCGAQX5J/UeUMS1JMyi1BdLSQLbBhxsFUM
Rh8Y05OqZs+bxiD2AqnUuAuQ8cWCXUM4UxwowpmXDXVZFCmTbueHRe2cuqHtGCAP
/v5J428JJ0wUK2wk3hm1alPyMwiNjK1+aLkns0ukeLQZDKKNImLRCtP5aqGO3G/C
n1b209JTrVG8gIJPjfzb8Nzh4rbeCNYJcFe+wfKoeHCXkjucmLyNujHwB/FW3uo8
vMLlMjdooyKyOocmJ/6BLi+eTFcjwXa9CRIXn5Pewv9ZHzXCQBT4PCP0wILbUeVM
40SN3HZzno4Jv3/6xXAO9IGtzrMlSai4lIjUh8aNNritIwUHKJP6M6fCzSrrMOMX
mUy1CXfQ2qLKyLRYbk6wxEt+sc52JO2tveEovZkuuVG1jdCSjHnTvIJVyrx0b/kc
sMMOP9/GYY9JxPO1AknTb8Hnie+MUE+axSV2zerL3tVFCR32GW+6nJag8jP3vpFP
EIJK6mVkU3F8VaG3gGJDdcZSTKLzeSPunqiT3SdnSeFZEUtL/2z8/bkpmVnTiU7V
didZz9F/6qfV8VNI5LsY0ZuOMZ70cFjwrlsMi+TMrsowboElUXBOtLpMf5Mn2njb
gP0bzyFrLmM5wjGBbGOTgABAZ8qkUFg93/Mmb5E05KWuyMsWY1Nr8DXE8UUwamom
UqluC+aAxiBQ90XWJ+xdVyYrdLOGLi3REKz9hcRANQQSwmd5n9a0QRD8fhe4NvBM
QvqIxbCaqsB2512pO0UV19ZmNnIVSba7rSf89hSmRNR1KTDhVy3iXulrt+sBeS18
ctkyatzIOX5DIJpVZTtbLXk6YDG2/NJjMz9xs1ECzQwdn/KafRKbCJgYX+ZzWx3q
ASrNDTBNWo3F2L3bf5BzX3U6sZJV7bHckh7QWd6BF2iudDdWnzBqdeQ3NyxVFBzQ
gpcx0B3fNu1O27E4t397p234HHx7/uk4+u6J98SyHVvPSQfSGOYcomkxgi2Yydsq
BhtH7h/SK0ob/UDbHfGgVBFaMHH4LEJuc5AI0L4/xgV17zgsNK62S+22OcQW/740
BuMA35IV6k82W1oAfmzQhdv7hSQ0zOY1Ivmjq7Wfrrd6GI0dMCmXN7afIRfnk6YZ
+8z9DJ5gJreULEwNLnlUvIaSP02mo34a5JLR1rwfsbpDvhhHiJHKFzVTS8ECKo7N
amkq6THH7RZKa5KYF8S8+09wSbkvF8D/qQxI3xHLk6U4KdEB5PoWzsL6aXB8pjFJ
/IW17q5kyO+cV+g4obYWh0e3tkbRgjFPeTqAEMHoQ+UmmSH6FGb6jpz2sU5fTtXc
EOZZcMB1cj8iNn9WoYkEbUE2yL+CPApH0qK0otNCAToi/mtnbn0wZClYBwkR9I4X
TuQaZwufF4/7mCetITBESw9FIhZ4iU3KS2PycGzfa7wh55UvG2OxMUFAJ1oAhlVn
UcIHpGxQiaVbrxHJEXrkeXmBvZDyQwqibMBj0h9hIhJHRiqp7+nahUNhvMaVSeo/
slFOK5kMQGsbraLheCfaMGRH2TybgHwBokp5INKRI+4NpZM9glNpVYqmi5gNDDF6
kfK2fYwpizsAIN1T3ox3ozGYB3tuqPT+NQrZbbjhjfIqaclrY70DMSzFMwbPH/nJ
ddKEoXUNVYzMS1yuFMwPQTwrlNQhTvbA9SnBLRLMyNBW99eN1YIYzP7deA1U7Jgn
tMS3Az4PQdDDWuMPoTIJ4KGUZlSY5W8xFRsxNiCu0PYaRSGFPNjrTyvlTPFAnDdK
Q41udR3117iw88bO40emQ/GpaandGrS5xpkSC9rzzGlajZ6kY+qinO7J0p2NHRY6
sch0pZwffj/AfTiOgU+L0E8s/D+67ObUmlCjZ8Q03QTb05oQNe/y2fmfuj6LlegW
FupD55TEi8N7RWGk1las+eNvW1CTf+/YlrfQe5e7KGDhwOMk/GczzS9Xs30bNABU
uVLLVlzuzCrNyWcBahDL8mteyxy5r0uOOy/f/R9WbfC4mGogMb9Poy0l+nUFbCKk
XrqgMImzdz14v2WtRutQy1KgQlVSoSnT/eW3+LGwauD+wYikuFxq72ZRB8bUFVKx
T8xhRXZfvRXiTEAbxJul2juali+Fk7LDrL0gn2QLJfwG5yt/Lg9nAAJZ/nTTHZSf
V8+xG64MTQy9rt+rCpD04BqhIxs9lRYJnvhIC8OGMkicBofrIkj3Fhnw6QufM19s
SMLkmjrAsq+/uRN7dYRM0+YgxoCI8C7Xg8jmE0138B/eLsT+IOCbMumO4/yDeCDa
e5QGXFsUuq/IsEU8P7uqbB4exPuHRiwi6fWWWKB/IvG3eN82ikGR+f7SwxuL55oC
TYf/SgpXvNeuiAtfmVVRGAzOe0Nbey2Ya3DwaShgqsGY8OxWBAzMuml8GKOxF9CL
xQDRPu2FuXsDAFd4erMgzVVpoOGyx/QnunEg3JQEFaZOJ5J3ihksB+Qv0ahryidh
khT9lqCJI7rvBTpSjR04chkj+JN5QXP4+Aq5DkDas44WkuuaDGBTp0P8VxUOYlOd
8dALH28uTZxh6U9VRtI40UK0QmEkYaopc5xVPg3vz08XUorfCx1HhdWudRjCeOXQ
TpWaV81rhDf1x/BjSJWbGXFQxaGECllFqvMeaJRwvYwAGaBeBkRLm+dg5zmoVsTS
RpDCgW71Osmtqmm1qjCIYIpxe6YyAMkVKQ/ipUs/kNNwHN+ALbgcMhWdLmJ40Wtq
Fyn8aoSA9xBxZJhaWIewWUuPt6TSUUD1ZngSrNsX1+CGZY57u+4D32I3D9Dy9tw7
mNl1tBSkr0tXbctJ/KHBsr1OwNAid8rQepxCXXD/BR2dzB2lYKDSfIl/ew0TyTKI
Es+9SVc0x4Q1lszerQs2RLH1ONoWxvdQ7aoO1gMfZxy7JSXD/4DEOFcAL0CZVgQ3
YoKLFfxYkbud6eJP0FHPUFfBFpQmhUx5lwCy2fc6+Jh9BlN/eV08H6z5Uumeo8WL
U61a5B22mgK0j17IrhxZLsTxhzM1Mzbetq03J6BRbNFPdQPNT4c/1SF3Sj5381BF
eCJfHxid/9M6adB8yIPrh3Cs4EhQo6BhhvSc0AqxihUhkG2A7bocR502GYoYNOAK
kzfiGM+wsl8PDfX0iVr9HN9wtxg6MjhCrb5sLafySU7cS9Mu9jHEhSKEQuRurzP7
nvJAWva/pbjMg4kehcqc1u9EgeWBK1fHwn7fPWWl8mJriip2H5qhiVWYnfEPI7q9
tg6GU94yIAK3MZ/0cm4SydYCXGBVJ3hNyiaaVfZBr3ufqIM4rAQSpyi9DXh7zHaY
xktb39AZ/VntbOHxlSjQEcPH0jbDTGgZCnqoD4eGRs1q/KodbQlmCjdQXRgNRbMa
scAQyi9t1QFb5WSB/7By1aEmJUqPrfmTj9qfAHNbuRagIqBjFjgcTcRr9bQpUjhl
/GbyLUgS9pmwlcsfF1mtQ4A7lgJ4MutsEaCBtb9k+0NdSN4fuwueKdlVZADZMukg
svQiLwBm0lw7A7mdh14Bt9fbg/8XWI4KRKzUNVq9VCLhaf5qv7nAV4uxqYrlJse6
ksH56ZlYWXHDraejfwbHNbGyWc2EM/WQ6Ah8ewKFWGZkfwgOt/dJAUOZluif5/2d
KXXX417QsnixUfVgNMiozABvd3OGCViWKH6GE025gMfLmKA8OIyJBQFhN0nNdYqz
edeYGxWrFrE8+8wA5Is1GqsfWj0d4yFX0wBTRsxThp/dhkhk4adHAbuniHA53cFq
5dpHFp9hbBNpl2sVKj0BjA20FhHahjfVf2WkRjjb84rV8oisDqFAlRnOLklCuFE8
nXG9EfYA/nPN7FIymBbRnycl+vhBkv8S+Ayjgs0hrkmOUbPy0dAL3iKELZvr5F5m
b06lXzb3bPI1ILTh32EMLDPyxfVYDS08xv350jcBkXkzQ9IRSkUIvb1E69+jdOnH
UZOwbQUHEmZw+X2tmukW7nmInOGynmwHLCuoo91nsbGCx2ZvwvQIbiu/Uk6fMdmH
4MDWmge1E3NJGEfSF5/hcwQWm72Y8tazEuvdyQepLZUS5HEovqAUaDA53MhlKYIP
1NTm0Sxx78mTwhv9OaWWPssWv6PzribXWxgnS6CA0Kb90pWrJuTcV80XjyBcLQlh
Sy40o6R6qhCUViZ8rda14TLEckL9Pla401gAqqmSkfC1fyXvfEWmmtuE17vOmvFQ
POXrKPoK8iO/+DMWAub5UqUJX4F3iNjFJHtaE3uZYtSDz2AyrChPVy079cqCQbZ5
Y6wnHBAZlp0s53u897iSGxxyuVfvQU89xnobedQIO737ti+wL3uolU3TBKwqgUsf
IC15pEaDtfQQPfM+h5zKKnHJoLuHS2gqMxtEwF+u5Ur3epIAz65ryCXqk7JilTms
aGEQZAPUpzOmeVsrOr1i7tz6GiSBrfj2Hfdi0T3tQxv4Kl+Ju6G/a2wb4lMhSrOm
P5/ppOKJCscU5iQDnRJEIQc+41w5LEbwp3n5W0hiVXji7H8jtPHogp0oNYaG7lyD
n1U+Xkk1lhjPjG9Z02/DFHC9OMVbF9Yo3hZeoOLqZlJFto6GgpF0mBu2JGv2QlDf
Nrg8qknj2LOufs1gWu8ig/sLj7bKOxUO5mHJzNUI6cEflagq/90sc/+l/OLAXIwF
6sDqJGh1k4KwEuT/Q0lxO8uLnQlIuG5Iy5m3MAaPza1erJ5Dvw+k0NVliJOd5S87
aVlbkqk5NP+hnlirjeIkIUB+//HdyBCO6RAZqkHuPExgd37Kz0FTWgRHOOPN3Smp
ONMHFNwhGjGpiX27DNCMQ+7vUVb9kQIE4UzoEkaEaIRBAMeG3GuWzrG2eYhSR/zh
jifBx76es/ARFt3xHpMJ++oGHLkKZIGfujLgsCwPLElZ+/E99b+IMNSI6TtPeRuY
sj18N2Ijv/zCV94baWX0jMnhwUYr6QWGpfBeh+Mh/uOV2EE2RCdfwZOwM6VaDq5w
Z9UtlH1gqgS5LJw8S9Tmhf4suSsyrpmpNSsUv9B8XGyo7nuxjX+d4siJai3AeKkr
AJAuUxbstCXvxJmPRD2SIfvr+u9ImCiHmXEuMvZ8+9KMbNJoaTStynirBl97nPFS
bQOL+SIrY7MG9XMo3sU9pKoc/mNUibPWqVOaaZvnxKJ5E3zALehlPXo0fx7xMyUQ
vU3RD046LXz8aiWA9H2vBVcqWZtzt9DkAbs5QlBd7p2ssZ7ndiKdSu1qXEOmgvWt
/DAc8cWYIzj1lqeR2MKROZWaVtpdtOk1VQleHgBS7o+t82kSBh5wCRSHyL+ods1O
GusCVr3o4Dwvt/+2bBHbeUCEqQmid0SJYI/pDGbHq/3K3DXNMVXMQIThzHNKGmKe
cZjw9ODZm5uMHoMeq90WYIShQK+II8d6RM3q+M4w4B4fYYs4EEz+b+y2kWclEkZ6
X98cNhYzduKzZTA2y+GxA16butmgz1hCCnHUdq5qPasnnPVhDW1KA80lICW59azR
hbsxxpO3Ds/nSlT+c7tle5IGDgKBQs9POQY95Zu031uBGD2tMLrAyDyMR+Xvtb2J
Jm0hdLXwfJwGddGXx9TVBa/JDS0phb9CUgSC64+S6VA8Aq7V45z9ZnRYAoI08YPG
IllpqpYy5SU9gxAEfJ5PnNHfbwLXLaePbJ8SETRcy+HZIaj9dVqtdaVwbX1alujA
lGGHUz99Hw3YI1+9bylOBAH52V0PeOeBdZE85hVm/03b2O/e7uIFzQzTMKNMUM67
26nLYZKiNmjgTwuNEgLYPRZ2sYolg3/x99LxhMfW7RfsFySjs7YW7QikGOy5NaxS
Hr1uewjxqZRDmbTojA07XAbDkRgmxmJ+NSSAHODx4WlIfjANYDeOUfJ1SkqLo2e0
XPVqrFJXATdTtnnupk+EyJafTYeVSCIGenHUiptSjs0A4+ZbSjbZ1HR252HpfYjj
B4/9OLJEMAwD2WF+dL4esfnTJpG3oBU6a/CIsOmicBcLRasV7R57oHwFlKCBsRYb
9wAOLi5VoUqGbIt+BPRUIeExPWoGFBOjXGbkL78+tlrg80BwRBrKh7GhpF9kmtA4
Vo5jwcE1f1ABH3lblSHsJgR5UE0r0xiUu27WAEufU90l6doCZ99X1aPRr8799lCz
EF/Jk9bZqPetyp6pxPlNCt/QME7TXlU/H96AT/LLRRkYsJMRvdDpEBLDO13u7Nq5
ve+yXeIiKfOsgRwI+lNaY97Q7k7gllZCo8By5KmJTYG0Uvp2JyisGMKoBnMAkEYC
2P+MkHM9Z7Jff7GhlgF9FBiL1YvXXsoADf3DdmTCzl5y4I2C4f0ugBkk0GhUEafi
QdumoSXOKXjRZ1wNQYgNwZi/k2365LSyvWczs0twWvxxUM538Fb9yU94kUwN+vW4
wHZiJTaxB7h3sxdoa3CJWsS8yihGbqjQxSLrNFCOq0BdzzX7F9oBbpMGVowrleTT
OOj4aW0XI5P8gNmb4IzpSAgMGyStkbFUQMXD/Ex9K7jIg/URbJoMQJ0EuZSGfeD9
mO02ueHYcyjjmQFg+StLkEgXhiy2e31nJZR2TyhjDQp/RkVCWfR0CLxgY/Fbyvog
jSPmU6ogSUdy4wd4Lk62HG3iia+gRZimwQC4mdSae1CkM0v9wlaSH9+p2K3Tx6NN
83vmK9vb1+eSVPrhYkdAKSjYnS71/arNTE7zplklYAtExuWOF4UoVZyWLufvH14r
hZprz6IPCMmAVzD5cl0XIFEzwszPVBjLkQlRs8dewqloM7ey27KrxGEClBFELDBy
h7paoufOIWRzMeXNEs4V8WDrE7IgQ/aPgAeGwCqEzzPACHpDOGbU4QUVHV8j8V81
npqRWDGw+PDNaO5hIPR+0zaDMq+BNVEhOPMFUKQdvM4JLfP70f+SsAGtEcx4xCYw
5n0GA4zdeXhXU7M+4EReTiGaBTD/oCG1vSmXwIRrZ56iGrpyKlN6EWcuLRY38IHz
e6CtT3QqPYvJSuaZak/4U/eJy1KVe1UlMzXW72FUZ2iXXG3IB6/QKPZyf4Cwc+/C
lma13R7VYoEx0qYXzAsEhe5sdPkydxAhdnZAAgx9h/9d8Eysd9pDDQGKjbfGaVLr
AT9VpgZ4yFJdwObAmy69OQAnADsQ+nvXw0kZPf5rJzj1htm/6/pgNjZPlnIcL5Li
3sT2vLvtm1qB+c9AqgRxzZ2Jlshl1IGXbGndo6x94faHb7nGflSes+eVPaR00g8B
5pzUzmhIAV2zjLJo56teR2c8p/QjwyMRBYYQdADBv26POEO9NVyqAr44t8Bgptgn
oytphf4cM7E+M6sXq4+SyNMs5yLHzEhixoWyWgZwjQLIl/vtI5OPw1VqGLC1nUBz
BDaQmNkoR3n05sMqIhbboAOtg84EBzf4+tojM+Q54p/LFN7FtTOFCm+PybaSpvUz
d7PbDuShCADPqKOcUQa1haB1NzRuFM6LIpaJ5JzgRy6XBZ5cl//Xo1wm1NTFMeBl
zUKkIoD9ReTi2rXUaRWIDgk+WIkqFR4hjNSURUL299Di6RFJkY3xWBLgQVEnTF/L
5kO4ZEai0ZhvEwVMbK0IsBQCqeIGEionOdwkfDTIFm0g7ISP4qI68inp8Tl2u0jO
ckQ0in4Zxf78KFIbxqLy8O+sctu3fEd5PMIfYW/CEQ8BrLBoFns/f1t1C4EmAA94
BF27DjBWGGmB/QOZ8VqFknKjRxJjS1rT8axsEyxFdWRV1Iqz6LHAXVTpuwobB/+y
unZljdoof7xLeqOJUqxjUP3UOxK0USlFxq3lIkdjfpJCQ5AvR1XAfg/u3AcPJDc1
gogAgn69UkLlG+oLC5PYiW0VP+RoD3Ir9vPvANKRXIpbnOriCvFqJjHKc0Mc6opl
XcnOvHI73076mjIS1ZIQlbjlTfr154KLt6G1La7SbNlpO8T2211kyByiI1EJujy9
tprzMDxNfCgpTG9Hit9JRPEDpe31LzQFkCFJfYPzQaSgwe7XPCZDpSouA2Pck0TH
2jw8Wqre7iqltNGs6s0NBwwdQspIlXNc2Fw5QrITGGn/aaiGERTTextwin7wwq8O
shbR/tJeHU//1i9EK0n/ve3yru4FacmflYMGuYDbZDA28DI5MnotCyqlHuDX0nwp
pVGm6QNFJ9A9WjUD4xC8qzCguTZpG8+IRTIALEUcQWtp8cyOdXWku0Q6tzzy+FSo
9NfY95uQc4VnmTybA1mACpChYasRH0Trcmkbc3MBvMhLSaWYzjFAE4y2sovmnA2c
2hADXn1T87TVdF0v1hiSxpSGGfV7wpoxPc0TT1epTs+ZWILLPbEHTGANOtd9MDSr
oxYeb5KlsoPEQIyQSet+92uBLuK27gSn0H0XYWiq0c8Ie/XN7Mk0I5EinMhKKiCE
27qR4CBkDshNKLmhWQAPZwfgJaTd5L8WvC2EuTBFeohjMIF1sIZtsAishTUuZiBv
n2EV+6I7N6exHVhP6mAQmIWQCgx45UuDSmEvlSBQQhHAcrhRFR8PYUxv4U6wi0xB
8PHk8QsGEzMmQcOqKyw4bPEId3fJPLLU/PEXSDxicv5oeDPVxmF80ktWaUZg2nam
jnepusglwm+mfit7YxdQrylF1jHrSgKF6BhlwpyNU6GA+q/MXUiyUPunKDbNaTAr
RhCkLmb6MLjqYIFFHzNd0JynjCTY/+OCPxXN27PlzUQ=
`protect END_PROTECTED