-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
--pragma protect begin_protected
--pragma protect encrypt_agent="NCPROTECT"
--pragma protect encrypt_agent_info="Encrypted using API"
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
--pragma protect key_method=RSA
--pragma protect key_block
gJdeEfBvFS6BJA48kLPfS6pdCH/7bPQ+Nq2AoN4wfmBi1frblHd2rg3IGZ3vWUtH
DyuKcy6QoO/A0hZIkNPe2CAud+A+8U+1Ba7PhqqDq3jd6ULjWOvZnFA/tCFBWf3d
H8yi1nVRzdT7cVbAu0wTDS9yTBebpR5h4q5GaQZAbXUQEsnaM3nAy0IjdowKADns
w21tubUgF8Ugb3zS/w0zb1CBscIPTDolCGq+IoSj9mcJG7KcVKSoOR/1EkOcCk9a
jQG9TY3IHTYzNd0DuHb5jAaUVbW/38Yxru5AS8tAecorseWEXNvSNV/nQ5wht7m9
2JkQNpSz1zzFIk7Sd8wzOg==
--pragma protect end_key_block
--pragma protect digest_block
a3yKiC24FrHz9vzPNYdU2iDdvDA=
--pragma protect end_digest_block
--pragma protect data_block
efzKj2UJw7b9/BbJ3IWN4ymBiDs9p/5SSvk0FyWajGpzOOAMXXPCP3lqgNqb1RQc
mApf5ksOl90++xVGmYElV9eEuvUUb34XITqUdO34B70RclmXXeU+IM8iARy7UOXu
OMmj3CCD8h3xdVDv03pPLhYID2uusR/aeB8DfdGrlvI/ARdR2H27tQxt+krm0bkf
nv1vv63Y4bp5ufGKRBCoIwJCqrc2IbxbzOGrmUZO0AsVxi4J7RxafLdYkE1L4CHQ
M6ZqgkGsTL8L9QJi0xM2zk5gKI8/wRDag3XabM2pYuVhx3atI9MSq8p/TOf8+R5z
l9m1XKBx/tbg+s8/WDzkcd6MNZUVGL4GxdTvz0LlR/w/TfIeTl2pLmPG9+mA5KrF
uST2P0PgDQKAyVJultbRZGhVE3q+LGNel1SSGYfWeUpiVvRJ+Py447OKjmvJtXfN
7nD9OvnRG3ZV8oGi6aihlvf3XvT6FQy1UFQ2afdl4GqcGBc/2aGQB7mD1/tVCBog
0fqtKY+VYvta5w5rMWoGPsJQsqxhpOC0EsvhDnSf9hm+AcebuWhLYienbxw4g2Vn
GniFelLPOKH3jVxqmuD/Apzj+LRN/YKaUoYspT8kvtP/Oyi3O66dJy6uGWJyYztB
/slf8pT/UxvvHYgBiUsfbfHkmC6vlaZ403SXqe4Yz3h99rt6NqbUbagK4a9hlJJJ
tKttFYa0Z6I31IuOVJ3H13vLPQ7Qs7ZuZd38pDtdg4MoI5u4UL/IJOQRDjd+tQUF
Dp/ksOzmATxjJtOSyK76Vl/QszTQvMdt1i/OHB69vI48u7y2PCrjRxsFvDLpN4Kt
xrTCn9EafCbJOibAR8uyRtFivywbBcWDhITNP7lCAErv2klkbwvUZWeKdQz72mPP
rttRE9rT5IGKLH38tTI/Nf7f8BYJUDbLU9FHUpN6qEJPddNsqfAF/w1fCq89FyLL
qTb3kowD5ESI/03FlpCOzimrRfEtOmJ6e1FK6Wp0/4+cQwe4/JKH3j7b/PKf1UNm
HVSQHj0BqS3gV+P7Z2153AcmBUb+NQiHu1gFgcSNVJkLYijKwLOo11XhvTS01oG5
7SVo+L98nyRpdz+XG/ufFq/AS7PG4PFQEm9cAxoQadO7bt6u4gpUg6bvWE1cKojo
X7/xQ4QJZwx3o6Wx8iuDdlcRU5fG8aV5NHHlavBZVaSuWOYegvIOXVxD+7HL3E0P
G6HSiYxi2pEZqZHeZrJ6EJ0zcQSDv+SRr5cE7W+fMxtlAJvZpoP2C/RU9yO0wgDi
3XV1EgCtxAUPNncXSW28JtPTUIpTRwfi30dPdKYewR93ePzwJ1Ls6ZyYCLhsNn/e
qxhOWpPlQjkwbb3yZmGS9gPyP9Cl3ZPdZTK2WrHxVH/Mw3pdr58ok+EaojMpJWsa
CeH3xOIUXIbChDWXTL3Jp49DibxDlbb7fqXeNlYdkyylk6SpWZnKMPgMfro0vpMP
wPyRnD1RmKIaPZlbT1sgUk7YgNMRnVKY15lu4V0yQiPDaMxMLbgwEQH5dvsjsAfg
h1xI40ziIA+IKtW0+PXvQ7LOVMxgN/OQfBMeJVMGRU4GtSMk+b1I6v+jYlcEwZV7
izd3k4hb+0gO3V9H9cg+ci5HB1RDFFv+1FMXvbymwh5b6ZBOQ//ZVA5UKU0tWfJN
OLWEeLQ55X9UeFz5qj0EaRdJ8YZqMEpGt3fv89vw9QZPC/vgEJ7uYuqOFERCbcv3
ooaTvBw/wVcVsggpfXOJRdMFIE4pOacNgTklzmPcLys66lwSGbIoJlYkCrawYlUw
D2WGEHCVv3qOlboChOgXDq0JvAgX0B5hsUkOjY3YK+mIkms4EowNkiuRkNldA7kG
iyDhteRWJqwOrN+QDwXBydTps00HiyoUfTYX7EETBi0njXDaY45zHkYnW4pcwwaq
xKAL00jjfPiGNpEvS7fGLV8jXnWGZ5zfPX98gUO1n0Q0qpZxM01uDeM1vqKflPmU
0/cHM4l5S9Hyf7Arm9mB1qBH0HQ1uxV4FmMQVYJ0PwEP7a+FvnQC1sKVArWoan5q
7jnGU+YyfQ1gUBB8PmTsqZD/im0wbfBENwBX8PleWMS0JHYibzZbYhD1lJ46dK4D
USgEfiNoqm5MkPer//f/S/ke8iXsiRaOkJ+qPrFS1lvqgLpVt1RbqhCOCloYApgW
qmL9+YP63CEyIctFPtg9Y+xrv8cB3784h61VpElSfrYEkM99g/m38noieoDwqiPU
6roajZu41eTcR8AnzxhCkl+Hgloe1qa9ZCb9aKdAGgfF4egIq9LkRCCGlBq7kvLY
5DFdyayh9qylhlsKJXMCzAggDXXzjs0MyArfbm0Lp8BXHF/2p0XakvqDIenzEYHS
sCOncH47fCN5rN8gWpUW+lwaZRneQEU59Zz0yNIi3oVuCMies5jKWBDJ8NyVyP49
XlPOBaZzJsjUh9Dvvw0AS6bZAxwKyfKtmXGxA20pT42pLtKrE28/WatoabLeRiKC
agU516vlOsx7STqKzcKgyRtq/7J4na/RGpIMUmUSajc=
--pragma protect end_data_block
--pragma protect digest_block
T/xVFRVAv++sm8Vf0BilQ/kGqDw=
--pragma protect end_digest_block
--pragma protect end_protected
