-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
--pragma protect begin_protected
--pragma protect encrypt_agent="NCPROTECT"
--pragma protect encrypt_agent_info="Encrypted using API"
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
--pragma protect key_method=RSA
--pragma protect key_block
Z5gboyUWTHxIGSJyCB0sjT8G0jHRhEVqlAEOJtDd92ofVwgjCFGWpGqmZegMz2FJ
V/HFLlJFES/RANJEsfD+jnHj2FFNG3jPqxNDZNnORpW4LYI7VlCE8wCcmFk/Vf/1
L44O1k9s3UYJ9isnS6Npq1cPt8n8+acnAL8oU87WVzkG8QDc63T+bDbuFQ2ozRmL
2V1VMSsqwhSQWQCbViwbrbNKoNIs6bY03yxqTl70us94p/TgNE9iiiq815df6qrO
Wt1yybqOD0Z9PCpwttXF9XeOjUeJyCGn9OMNRSFygnz4XfKoWyKT8IVSrLZL+DFA
PO7wLzKMkB+DdcUn3DXSsQ==
--pragma protect end_key_block
--pragma protect digest_block
vWgH94RKpy/D/dDnag5zIBNpgWo=
--pragma protect end_digest_block
--pragma protect data_block
PIb4/vZ7hCOYCYuyfRRIpaz9J3yn1yGPf1EojLJiK9zH9YvBXOH0Dz258lLXR88Z
h1ekiPjvoR+3folIhtXPjP7uB/GG2ZvitlGhMPJxwTA9i4VVE1KhwzLliQzmuHpj
MvXf24s9hyNHIPq3Hsv6wLFZCHdhlA3TcVNSUW7iCLeAOdONwFO2Cz4Yb2rKZNWQ
52bce38oiuKqOWLX4mOCP1xtQqz6qgz0OZANYBVMfU9CMPwntDkw/Pe8mhGDBXFp
FiEswFCRVW4BZnDupAHGiIfoReVcuKc9TZ6/KyJc709nCRn0gZ+1ar8tK1iyF81K
9vqQErVl+d5ct20vNF3JMU0mMYPkhbjJu6KwYR61a1W004jYIGiGq1OHinRFwFF7
avzfQAa5PCJM+Un4GpNxgiKfDMAFTk08Gb3KZKYZZIs006pLaZW+/TXNmKp5gMkY
+xWLWh0rLS7B0NwJJqcBAcn+TPGzhAD5jGdpfpskp6KH6artfFWfIQQqRvaTsr/U
05UVfeazxApcQ8ZIZVgl5hY8QyuIvW75vciekixoIeqUYx3b/RwP8nYniqh8EX4B
0nXJ8wIaG//hYqXIBJw+If0kQv5E6P2uXWdnCu5j1xRjd84UMvSU/iVAYsazrAAO
yGGK9lD82cDywl2QzwJO5OKotcb/+7HYJp2UJs3606Ju+LjlioTeTai02EZB66Z/
KTMX9FC2lbtfG/Oq6jqKHStA7DybqtgfK2rJ8EoADyrB7JhHDmyjILxqWOpQqqDz
TgNqg6N2Zm9O9EqlGKJW1zTqi1LW4KtKzm1PBfmS9lFg8Ju3dvEPS6JVYI7yoVV2
8QegTpjoGOTy+Sdcsc8WpnRdCH8WubplAb3HpsqXtpX5jL/hkzfMs2a6vRyYZCSh
jXxgaf7DmIkXr9/SB5aw44Lw0J8EP9VJEYUIVeij3U1b5uqENs4iihQGSP66sJhX
lZRXNkK0vklVGLocNLwfyxcrtSYgewEH7vCLHRXe9HrtufIGVRGRnSaoLdduVKgW
3s8CO5Rmg4FkHv5SSLeJwEr7rySAkrUZAcFLRcYD90UhLIMcqgyKLxJ74b7sUaoE
QLIkOSOyqfHnmXtN1O7VoIEiW4kAjTweGmZTKLsAkDZZVipicfknnxxXLBsG0EBA
fWw02pbiLFoHEKe8JUUHhvhizvaFe5XojMcJ5S9jb6pb1yXidoFRrwNxZxTCKv2J
1qlEf4bLGGbDEZTvXXkqz/ivB4nmyyVGt1FNuzrqGUwEwzeBTuzodPIVlbScKI4q
qOAsdX5f3fNOzub377KKp04qqVYNnZTAgPj89AMp13R6sLNIyvB6K3RgaQOS/e3k
uOjzJ1A+OGdeAg+h4k/btl/t43vzKcuonhYSWdse00dus95UfXmoUY/c4EOCp0L1
aZBJ0DoNGLaQChgMAVWfmHr2saoexOUNyLw71ek4u/XLZy26cAC4o1aTUfO8BAEA
OlRdt4xq/Zq8rZcVP0boxWUJdK6gOpVnBz3nouqbT/fgl6+a+faKGh4IHm5fR1Br
6/VksQTkthy64lh/OP+ixdafZ5F6QzWBgkmU+9nHldep8uOFO/6NIjvHRvgmzgTX
hGKGxaA5i3av70Rm/fK0/utmV08EfLWaY6LTj5LlbAERpGYffR34h7/B2dHVA1rX
QGyLiBd2yW7ZA9Xj92NdJHkMYfH18xS/HAnWg2Chwc7n84esvwAYfnlyAFT+DDEM
Omwr01FAwNVhEu75Iqq96Hj4lRaylTw7Ayx7g3PwzlYcvUNd2hkz7bZSXf5gQwOV
m8lBPEMznqy0SV30BxY3v9f8AbPMy9C4/2f5LbNLhlVPLcdQx0smRBRmF57mC39C
L/j5MDpI3t1uWOe2M2J0nVttpbQQ975jLBzNYRibQ0Llf/BIEQhOxMKDr/uTbpn0
N3f8rs6PLKZ2QVKD5pDKzxDQogvExQ9EWj+eDnioFjQnAQnXi+5iQe+BqfiiLD0R
kYwWerxBmFCaZr+S52iSsgbTSYdXzX5aSBeQZKBsP7qn+/KSTfIu3NGI5MaZ1ZeK
WI8Iz39iqyJfrBLqvkYlg+fzxKK9slsN7gD5ljs0biPjV200xKZ29OXjzJi6tlfn
V/zsFMzFcIqNtrK2TEdCCyE+7LdZYdI6jM3yS+Ep+YMFO/6Pk7pttbmAKZ5i7nZM
UxHSr2d/XDB1zUGXRs1nNArDwB4OBUB/WeWHsTAdpBi5Dyj9fHbPc9ptIgRJZDuZ
jHIOp/QwM+XPF4jO6mHh/FEJ7chZCy8WqqklnfKtVDxd7WOh0SfYu4WjO5lqioyO
wrtyGT4C1e9ib/li5amUXJiO8HgUWinRr3MTKMiV72TTEQSzU5WQ/nbaFXwcB7sU
3+Rpxj2IoaF7YkKhivadk8CVdTiz/cq3a1CdeIKnN91Hou71dLA/0g2C0aBH2/Yt
5F5di7R1MEfyoS7WVAX4SyyOOYVFmyxHL5lacuvk9l5KCvT0vM4KpnY6YLijb0sG
S5o9X6Zy2rI6DnVFYx0zQlUMuzol4vAGx16Dc5hFlxGnsoaQTsQ127gcNAKF1Tbj
PZ6XAMrB93kL8ZbX12tGB6CHR6XDZKYEeTQl2GBsM7q1GyFR+9rjL8QVU3NPtnYl
dDJ0zvxMsmF9CarpUi2BoGqKgwlDhQ85rv4pjVQ+OctvKxn4j0giAHR7B4yy+cOO
4HHtkxBA3FBX86EdvuXKcuIOiUqw26lZyoDiP8QRjzxQ0du95yAFyMRnkExnfWBb
8l5DKlEX6XInrdvp1yOuaZgEpUtXvg9bAVU3VKc34diPjUf3zvnTKZ3DsxT6C16r
48Y825NmO0o5G3uQoJziNFjRUcqJOEZEA7jCUIHkLvBIEGFIQDW3K7yFBe5WsvVY
RFKysB3ZVpFc1rmsag6A+UGK69B4957UKACaLE/XdRhixz6NIBa3hphDAMLSHM4X
tDCZoAiPi2Tk7SNPolGUb/Cb/9t91gbTj1EuBrMszJAw9Im1HHJGItVL14L0nh8F
6CBVcybrcIN18abcfU0FLA4tGItdAjnIl06eQbrxn/LHgxOesD/NGl5yG0FTmngL
+yk2kHEEoy9wnSiSqWR+BF5iE1L8jz1GJfCxR38w7OOZ+K94N+NF4IlBajiw8Zsx
gY/lZT/xWBwn13tl33UUGZ2mqH/aG2l2kisaywjKjtx228jC6LafmK7LzyvLtBlJ
hZ1RFbGv3mbYdHEOMUn+HZ8jHk6tyMf/zVnv17qrM6rUYiA/FkBPYXreddnLqdhv
c+cNdbkpaZ9wWy7IS3zn55P83pOdvrjpwbrwSiga9mZSj7gjCvfXq3nDMkqeNJ1D
KulhFqvUMQjTLDrBpTqPIL3kEm+A0Qx5L/J0Qhzxg0HcOTn/CIYhQrK6khBwLPB7
7HO4Yh9tEYBklfrnQd6Wc3dvie3xVU5hBgSSIknH8JR+uNk7XNNEoIWY35OOBlq/
3HvexLVZ+iUhrm0utHtbozOA5DZF1WRaVBR7+bE3KsVvIo5kmzSyrpDaXND3Cm9Q
SCwxDHb1Adx9wxSo9qQONAwTHdKhfrKQ2YngjFA1GUqJZ+kAz+aR/GKp2P14R4p2
xCbMeNkHycya3UIozx2K1qkwWUOrSxseEQk2inR7HjbmU5p95rbISYTCGPTZbq3s
P2Kh0trFZnBDdz87JYUorYVCAeFklKee2phtSvgEOFrC98rdQ9E6JiJK7WexeHP6
0urmP+Z3aT4njyTasdGxAlMTwCy48KeKVxbATx2AdXBr8zrf/Jr4AUtOavdC6MXq
jREgtkYBIfItMwmfacgZmOwh9WG9PClbZOiQNiYjBZuzUEv6tVK84gb7zFN/XYVQ
eRbHJBaz8YKIpb6pE8m6q3OkkWkNx++Xw5txYnvPDXiP1virlvt9Qclaof1lEg0u
nARQdHpJngROvmeNJ+mZqYVG/t3Ysd85L0T2n5Z1yHi8wIKkJ9E0IvegTgXB/EEq
gf+gn/GTMr0qbp56vL/GuFyBcuFmiV4N3iY2IdlYqnXzfc8QOFGURRWqYIVReq91
a4f8flLXol/idbc3G2ORdKITSnpZNgwKX2NiZLyP4SXgHwtz3tvpx2GpO1pSqtlo
HSP+oEyXaS/Az9yq681RAGGLsJgfFDzAMhfb0i07UmHuVTSH6A6A/mdKZsLGDQ1V
MEjez2f2MXsC5qQXXXsJ6QofcTbl3y/npljtsz82999lseIQVCCxEdZXdCRUelk/
ms6XnekvO9vKxDzxBC5mYCUdw3X+Ra3i0B69Atuq2uNOMIBF/xN0AagfldYw5f3d
KvQuEBe5sM+bGFKs3f4S6o/uSTs0TtjhpQicWFeSTcHt5IeMkXejvtpEg/lT2J/6
sBmt0mykhiPawHZPwUKsFjhHGB7Wpp6U38BtD5LU5faiJcimhQ73Z52YX6vJlTct
DvsK/UXfdm7Tcl0DINFfobcTH7aphs/k6JmTDdeOCRtM1McJ7ucorB7FXP3RGvT0
RKPwrKkkEq1p1fxC3JdG6l+2/ZhudiLzjVazhPW8EQhioIpZbpRIezPpkp5DGlmh
Ql6lMnC+YdEbxCWeDvIaNjfweVXfSBB3HfVEtv/6cQbBL9BI4TXp77Ev7uY2G3Np
nNjXIlq7taes7I8TNILv8F0k9iK7DuoOouHeQ/1qXi2S4FR9wa+74Tbz1c1M2KAZ
HzafbPRgPZKCC4FdTDd5INGGisNeM0RfCmcBFLNNVuRV6pIgvasoV0OOuHywBwK4
zdMDsZh3wJqlNt8krlgiB7uPI87aWMi1Jr9UBsW+5P49pDSjVOknZmQMaMnAqkVX
JE3iO/3p0gkprnkkIOh21ooDwCe3c0QCLT1Y6PExsT8Sx8D+agaCB+bsS9ND6lEt
/DpH4NDzGLw3U7Fyde/HiAqVgOpA9hUZdRdG3/irq6rqynt6aC8un3Wd7nyxCIGj
qAnyNayrnEPYH0anQ2g1Bf5rPNQD19CZXzCamIBt39b6SaTCmXj5YpiXUErqED8U
/4kayTJZwAroXpeZ+klTsymJm/LTWEIPKFKV+dW8plIuwHVRZpFa54pdvXEBIkB+
9tFzkQtiDFMkB54uyEZ3IHsu0L0bfOnQMLFh76CnQcULBthvb7pDELnXjA4jIJc4
WevUvaFuyVBjOMFX+cfg7tyrdoly0a4ZMx/O5+e3NuJgRnjUCfoqktSiC8QWtlVf
ifAfvqyCwaYTXKDLHcBrFXldPg6yIU8vl6i1HoEROCz3i45aNoXoOy9UX1ShrpG5
zqDC36fQdAWJ6GpSHwj0T39YzpB/EN8wpd+fdictsb39vrT4H0/sF1vN18sPPfV2
tzgiaGxQ5sSzondGxybYQTDVpeELCuKQHnaKybcdvPbRMfTTyJyZHA+gMxy1DWWa
0Qof3FqB1bDMbMu76xqf07F6sEz0zF5PrvmLEflvbgJ/6JhFlz3SoOh89JwZLFhP
PispBgpIFoJpGVbU5iMH7J/EhXAqJY+EHDscBXcq5MeKVtuyI9mQ9OwkElK0jTN5
KrhiHjAMhk0QMvZXy/7DDLTrg9jp92CNQiOEKgesz28x4RYxJ0f4KjbUKX6lequG
DEwVjmji26Z6TAjwRlmEudE3cENvJW5kCreZlrcfWDf4ScTYIRf4VNQ9cCD1MZw7
l9q5Y04U2CfkGc/20Zgd5NiaK/FEfYKUrE0kBk4bhFyg5vHx+NkpJt+JGipi/Neq
Ecr0Q8qnjOGtGaj5zJHgTRCOltiGavQI46PfGmzIdu2SeIN4jq669jH6FS+CfoST
ZVgpFVi5t4l6vi0LhcAeq1vgwdMtHHX2l4lDm+TC0snF6DNC2g/rsgRgagn23J5A
6nbHD+7E0SeI5ost722Er7IvDSiwviOHugK0lbWKjPQ=
--pragma protect end_data_block
--pragma protect digest_block
Lw2c+OtPV3DoCGIp4yS1zNAxVAA=
--pragma protect end_digest_block
--pragma protect end_protected
