-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
W6WGwrJIG+k2U3U/vjkcB2S1bxuihHpI3dprqzWwXGXW6vvSqfEIn3076xZrtk4r
/bGSX6kUDtlHP8pHTHIoeYyV9wGV5Ixyizb6UlR+uw8AQWYd3GhpPb785qaRO6RR
ZWbJEcpG2a4MEMjinOTUjsjy4b/D65Ebupjcus+W9Jg=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 24092)

`protect DATA_BLOCK
pUd+/vFXj9yUbMerEAn0EihHGoknk9dfwAooIKAtO5bUwBJ9/gKf6QezBJzVLJLp
ydASKDFrFJ8dbNcx9mE6A5Q8kcLx9Vao6VNd5qcOQWMxHOqJbv1F99C5aS4HWIgl
gQpvCTF2WdHoF5cGTBzX0vYqa9fohjEjhd2o/FgSYxK/TL6dmZTO/XWi/C0P0q6A
etD0ZEXHlt41lR+mdOnnPXIvJUJlyigix6gvL0cmmUUbFksfbvWmB+X8WZYBsboC
kC1MkelsQLux4fP5bTw4qpugiEPI7CXiLQKc8qqzcxi2b9jzvzdGQ6gazHsJl5Gz
oTJlIUuuecp+w8jjTTFjCFYmsAlrEJuS8DXzfvf/dggpr6TXs/mqJHY2/TLs6xYd
S+mD2mDPCDsj9fe6QWjRyoWIGJbzjkjLs3hSr0qiowd6raqCIe0n3+ZzLHyvAb16
TI9zp8qbQgFp7c/rQNHxLY8SBt+qhEsMP8xaCAReIWbkaAe04m1nr7uDp/H0vkCq
4ekJfAOVKgjuc6aJwr/vU/Kf8oHn123eyviI96dqFW6LXOT1aL8PubJPEI2J883d
85LMtyfWIttpyfhpc15A/bZjfh3cy0NUR1247IGObi+AiaXPDFYSUsj5ob9cIykD
XpFWv27URAg+W/wGNKo6kAuiR2Bmhd3zcj/6R9Jr8V0O/dEINxAxh/V2LeQmmcZ9
xCrFJirrcC++PJ+T4O7+xBjzNN1Gnuc7y3CIklTS6367QatFM3JaDP0UjY01JKJb
2s2xTzdQzp3KlKL2qVXkSPT4eha3N9VU29c/p20wb7m5SQC70pMLq2YuPVoXqY1w
tXcYNlMmEkr1az2q6y8rSXtz6yVdhmLTx2g6a0AypchfGNDVZHDhUJMtsDPSTGXB
IlLR8mS34Mh0AfC8xjvuirP5qBT9h1BML0xd0BRgZ47lBV5oK2sqEEnZpi5Q4SXK
YyxTffSXkAFitkxE6ZRwxzar3h3UKXoLO7PtqYWN5s/J6neIxl6O7mqCKH8yO7s3
asVDc4jkgKbKFARuXQ5+/Mh6dbGlPqm5FuKxRcBXLq2tLDxzKuD7pn2QzBkTLVQN
faKPR2Dp05/f6Wvh/Q+yR0ke0GN4I8VLE6mBWi4KZHuqPQyOASFfnSGPfQofqpbw
gPdpASfzYPcqnvEWaWhVtGSp6emM7DQ3EGtcsf96zPzzI8jj4/C7E1jW89ULNZ8T
zOz9zSpRC8D5IyGA1HiS3CTWbB/VMN31yHrr9lWF0hYjWalDb/vKX+4gHZmXM9jX
lZMoGzJD4nNX5hC63zekt5kcVNA6nsB1gWxKC2VPibb+cuE+YNUghfeq4t+rMIAZ
nRbAuhBMrJkWs+cgFsDWgKDm1xu4wYt4oet7HZfE8pwIIDADRixDb83PFpam1iWS
8xU0SOcX7CVzMrSRSryFVIBFwqn6zuNcTkEqDWTpdZ/yiVIpJKSXaTQQOF5Z7xjE
h9HIn1Vwaxig0EF/bkAOYWizZ53Ge/ngNT1jeTR8RZ0n81+SeRmI5Sw/5jXqzRRp
LIao5WV0+m2WCoKfC7J/WkILdmw/d2V+TvIuyoQvBhgsheugBxSrU8fm7XK12hjh
S1efrzT6IGbRgey7mzCtj6ixP8Wn1hRZl8v6fbMPbWOgTJoiy7xocfR0c9g2oFEc
RJtAc1+9QXjATSqzi/gE9OACfy+9uJatcbBDATQln/S1QTxwBvsS4im/FBim5V8J
Upe/hBByrnlkcX4O0fVNkRmJk69x0Sv1TUt+Y52BqEqJLwqxXGj2nHrfP1nIFSu/
wYW9YLpQ9j6A9kTfyU3W/ZEgJhVrUJbPw/WBQYkJwmQW2aiaq7H9S2hFLGLp2Zct
6klpuOcjMBs5+WDGSToX2UEl9R/+sZudmXYx4RRbxhYqrZE6wfPkJqlhAtxc3jvR
KIdQE9M2jMf3yIVRrBlJpWRCyMbSfqTJLX/QvhgRyMCqm98qMZhHkr0KxcGxAhQD
pZKi0sYNRGWsaz9AIQdRek2aAX31xAh+/x0xRXdcnpqKuNZ71Br+VUe+e9pO8MgY
5UO05kmMbwuglSV6UtCrz+H56AwPAMK0qWo90BMqPEc9HvDnnvHU8XbdFgMDaH/0
rr7EZAzq5EbEHgh2ScV7P7dEfISMzlgmwufnvDr7NnC2FItZoJkoMiJDh9B9DOzO
wq+Zc21KpjsRSb25F8JGGHhWMKhM3BEeXjbSOYQNKIarcRVtSLl7wxYBl7UJx2ZP
jE5A6yM84yN1Bh+UxWEajoPluRvvIb/Nk0czjYjnRnAmvNPG84Pd2s2ItqLhZj9f
NyofSv19qvL78b8OPb6j1yQz1VdttxBeU1Y3XJTezlqlYC9nIhRAAowy1dfEoN8p
u8TzLQZHVDLt+472ffF/zlZVQuxI641OUKsJxfWBpMGvIe8UnEuO+jq3SlTuTMGE
J4Fy+ii9cSEr92d605v/LQOBwSKgujqoX5ZBOutSQ4s12h/hxVKRQdAVIJTSLB4f
7ic4wPIJf3my04XMYf/7BNRxCJ41hWrWURVvxSTjCa6JKRkF2RccQ8bFnqdUsNwV
UI0Vyk/3beJ1b1tUkv5LCZIz//nRz9RT3tD1HvE8PKAdetsqrIPuWDH4WNXmxaa1
2SlW2cCM/I5dqkPf/pJgG1I/rbslT0KqENWzknt5Pejlktipcqnz1z15VtEgnYtq
q9Gc0bGDgRs5sL916j7slSwOzva9ZOu1UJAInR5ES/YMN9FlZ1vbd0EgDJUXGb7j
Pm6T7AhDoyc6atoyjbR0L347O2LsnX/Bir5FT2yCsktacpY6usWatDxRAX9nT7Yq
MATDfS4qzCqIUxgxs1wKRqsZCx3PWIwtGBEE9yb1G55dZxJldglCw8dViFtenO9A
ZQ7wYtxDPEfZxlLwUr9D61HJTR/Oq3AgCJqG8vBPk/0ajzPJ+QHJd3LWahX3g8PK
d2NUFzbJ1owz4fS3NbE+bneuI5UUt+5800wGFBh/BltzsdcZFku4drKB6BQPcKvC
Us7G9ck+vY0kmfFTOyt742Rcq/konflip4x0akjhgSur5fXUfHuOvYFYvn1nblK2
6qvVOFE65KXECHIZZ51GM54oxy0v1XUa96VH2BEotMr2SqmpRaFFQu/iiXg2+4oD
NXeC0WNE88k4iRp0lq1blNfW2UUT66sxV7t+3sdnXmBrUu/4rdls2ukb9yAu/bxd
bf2txSyNd7taIQi9stJl7Wjiy2m1fJ+aOAglGpaEn4I62XSzyYpNEcwJihs5lg6O
KThpev0HWRmUo+RKBEiD30YLtQu/7dkIcXYOeAu7j9k7tP8Srzrc8viG9CYrEkt7
LXCQuVdCz8Lo6wltCPjfoFP0jx9FZ4o4BPAfKJpEKDejlwJ3CoAESTHbJlUZBOtj
s5AhB8XKT6am5N4xlmUpyGtwap54P4AoSTbK0zNy+ZYFVF4qaAWfyaHvpfBuQing
s6RBWBZwb0CIk/1Q0IYrzFkxChqjpNcr/ypuyN5cZjwpRHmJYGR76rPJGkxFTtQX
RSqhCixx+HWDNtf7qZqP0olchywc+BQtpgWi4uzB9J+MENixIhZf3Z8sCH9uDSrn
Mw87TzK6nrXAzoVxRq68GkBuD9DUFUnXdDCa/FyNQ/0uGFsTii/cTKHtG5aTHr6d
AMoyt1fmWS/1nH9F0fgEq2CNIMxZ9OI4PD+xD2vh66QUp10RMnGww8Jc2SYQOQbb
b5gatCuj+jkCSNAwu9/eiFBh8wIp+eoKt3l9rqHHmjqAbJknJHpJrqqjVNKgEGjJ
iazgReIWMpH8enkTBCOdaqjRAfdGvgcUvN1ulNOAPijaimza4ak/dkdu171iGX6g
h03kdBhnFQWCK7OSjsmEHxg2kDQuMht2CiEUtkIdQYXgMwMZbSp5EPghFJW3SXNi
bQC2ID88rjAhUJOX/bs9fP8Y8pjmhJNK/gGNXW/bH64GRzqpTL8WmpVo4oure07y
inRPt2gg7DnzZFpxHW73K8BKxr14W96F/fJ7o21qXGCk2UDvuvsg/Rek4v/ABt3F
fiLsXZfiIBPM+bzxi4sFrVJQisMNXvg4dLq+ogQXw4S7gmXK6JEy2cXf9cWGE4PC
Dd+adz0dUyBBg2xgVn90V4c/6x8jwDzTiEudoAZ2rglW5nmlegXqWbNCVtv97PdH
v9KCK0gLLWRQmWeNripCTuBF4napcPaNr/Qm7nohkoOqmPGOc02ikBjX7BNB/54/
/OV9sUp8W58NBrym0xIpNl0h5GVmE1DE0vrHppbu1MSaSuegbE0Md1yforROZW6R
ZnwKfm1PsxjtXxhiLNn6xXzfdO1OfTrWG/REB/VrItuhrtva05TaXPs74kYqjs1s
HIyAt2bPpa6+0yc5IaCTc6ky2jH0jvhLXK+cCGjwoOSvk3XtrCtZ0CpAIoyqhnwt
qfJvInIGm+OnN60lGDQUrRltXfFhA3e3VDjLZEwYfDxWqqoBzNc3SMYsT+LuDmCg
+Xcz6+khIkyqYPgBmMiJDBIS6Jq8EKh3ic9nb7UvME6mzp1bqgn4Ko9V96t6Ss9/
yJ8PJmi0sSSvsAogv6mNVc4/7wrx+Tj2GoEq3e9OxyjcD5gsSLRLRcjn4LgfkGvr
vATQEhv1beoW9Q/grcgTBe/18I7POMvAIWWQd5nJKXHoZEGvYD3Jp4tV31DEmNnu
eCFdI/QvlANZgimDuFu6miOSDZ2ujFA4MchWyTC35g30zjDFSpWs4k2h8mB2UmUs
b0QRytZ0J091Tcvd0ojNE48tiVpi6ftZcG24v4/zVxMPeD+lbfs6MWJL27ixUZG2
Wuqf52ISph19g5139qmRUCCnzjHeP9ADKY4/6C1aNgBoKNq10VY1gUa+tgrVt/m7
dRxOqGLyngSxlxRbdpxuXKDXouPC+gutq6iPuaWbtw8KjHATlNz5avE84k9O5JyS
84Lhxs3UDsjccZ5/kDndg39VltPfrEqJ1LWdNi4WiCN0TEPVekSPhiNi4d0DQxnb
p6JpXL6p2vsiKuXWL0wo7POvJ3ciX+D0csA74A5vco2wIMy5avHRErMtv/N38hn/
OskrSh5rHtbJG3OoVqg/UHYkTr4V7icaF5m5/su6lDMMsNmK6bKWhcCcSNhMbxhl
xzFx+dSTR4WZqKl1GSPB/M6s4GvYdBn/Gmoq8zRG+4sxQPHRwuPaeAelGnXcbrH6
JeL6+nrEWr3/rdZ0sDpxTRnGBy29i7JlJwi0//vpCA0jAape+28Y77d51gKwmu0G
/X0V+PQXK069i/UZ2FAknMzHSfolvpNzsS+6wDFa3WdTL8i+5qJuakX3UE6sQqlV
SmgILFk9k87CZUXAEkOVXgNg9khd/WDcX9KuyPoQGF4ofBh6FJxGtvwaVZwy/wdI
OablvVDkzzj3kua56vr8IDAjLK9SVrxAjc6+GBd6cq3P/HufeIahowoTVFEYZCoT
l3P+QZNeNVdU4R0EubHps22NDXQAbR6ikTw+s0efXOLzkytmpdq/MGLInYQNbMeA
S+yjxwKcOsX4y/zusy0+HoV3m45tJPe+l91r552OoyRmEbQp7Jdr+jOgjjdtjARR
0hli2qzFprZnbUCmH4P0f1d6t/xG/xg49MCfFjArsZtBlnAm152tl/Kuc8POpOA7
XDFR5oqBtWpcbc4JLc8ahnojTCYlvraKtO1QRcjIQjqicomtohg2O+lQceZ7VBN3
qU6HJwFWhbDVh94Gimiu+O7cF8NLzhCh4ir9UKxtCysvV6Jnxq8ssAcDF5HOlVQo
3eM4GynAB9MZRKI8u4XAkj/20eBJq3OrD2PKW7emHr7ElMeqqgC4wU9KwMzdTo9G
tKVVAFifyHtzz/MP5bLYZgFBHjIQxBAXq3otUTT9wqAgXqff7ipySUOGoD7nP0X6
t1kVtX7yJLjr0IW2PKogmlFnSEkGjVLSE94LrfWtHMbvKKgiQ3/ywGagxFUY8hwx
MZJuo2HnnglO2UU+lcXgni68siHThEOmgmruGT3MsRNmd/d7IQojq/midKeU3jEp
cDitGIKfSOquF7bZ1Bila977jIHpy6gshgGqyGWxLpOlWCR6gVBIpCU+el/OvTPP
/f8KAQJMT8fzaaW64BI6wGGeplgoK4aJX4QrHQRKer91ppZ04Ek2GNBaJ2OYR4V7
ZCvEJkwcoXSjgPonNbFYRQ0SBR+UzKWFkzWdAaffCcozvFiuuT2yoZTWjFxB+mw4
1oq8jpTh+dXIidX4ogMXlacCuRv9eFM40NkiFOz3UxKSA7r7M19n3n5q21MkuBhb
I8Ssxs6X+V643nLpsIorBdODlPtdpa8TsxJEDeUHhee7g3AF5kXpr2uzcf16Qt2w
rjaB4+3WCMrFo8eg80X1Xp/m1qtxSG5yQAEd44Lc9FDtQaaONOwXkNWc6U05eFDx
ES/IPyMiWhhFRQO0wfZRz+HkntKMi+2azQcbV4ejUe3SlcN4IVvWChrFcfKH+GGp
j3q4TLogIWX915hYvOO4ZRF6iRzw7oqzfYrvArl+dvp8kb28iP04gD8c2u7A2B+p
v7ltd4VCrDYhe7heSlC2g5FsNopEtKhGcfMf/bvdaPKtiRBRDRaatnHwdXamQ/qP
JVvuK4uH6INiMdhSckI3BT1kWFIbmzdBs8+ZiEUYvPEI/L5EeYcs1zxVTjOK19h8
qqdK0ImLzkJast+S2GSGxUMCZpb3P1T5PKlksStiX4dYs7Gson0ToGUvNu44GfGD
JKCsnaEwlXTGzrXJnMsokzmxFspCawKyZ/wr1ZWf+9pYgkrmU0WS+qOYFFfOXkbC
ATfdKqt2sLTE92UxEJnUAwKHtSRL7ZiLbLVZVYQKOpHSboGoM/+IRazuj7YtRJH6
FoGndo8aGI37fh2k5FRpJ157eg+TL6oS4UC8DXMJML9rI+lk+Q/04rMma43/Xg6W
efik3Ldgb1XRoAMSzG6tNdNURLOmwz+WDshiDq6oeIsQC1YmUFTCTI8QJ1G+r3Zn
7B7HZOWBq1uJ6LjCKJGdMAYTdNqUiqgyNN/HEs9S0JEH+JsFAuSIoelHNNfia+gW
bWwRvHRyXgiW+OfOJ0N0CnkP2pq8T8Cldhg8zxM8riQ1mp22ubU6Ha4s2+Fhv7Bj
7KkTMfy8iQgA9v3NLzuJonfLwgCiebYD/ADX2JuSHtVhHRiKb9jIOg74mZRyQVXc
VwTWanw8tbjc5o3OjTB36w8D9IdStngSLucYXU62Yc1P3Mrpbl4K2Z9tyNyoVpAK
BEJiDOeC7IlhgtadRHRfIWkm0btthHDOACHoTdHt7z6gcYFt6R61SyAgXKbWBePG
ynuvBXOGKZN7snzHydAQITLjoOfsD3q7q0vLLsO8DIZadRkAsfkK6UID6Enc2iMP
MFug+x4Xp0BRVCI+aCsix5NnibkLwv+kYj1RpONSdkvsrbs42DGOPMrUutAUrDp9
G9qkrNX9b/1Mt/9NPZ6wxS9X4OxC9JJ5w4p5dBSZkDJhysfEFDC7ZRz+h6IPwLIG
d2NFGULk2HX5fztWPLOyo8iaKsdXnMVMImK5jG1NZied+Glv2xqvZUk1PgJwZ8xd
zDEK2240NCX1j7LIBsIT+AM6XjyI/Cvg27uEFGAaWk40/d1P+csCIcxq7ntsz6+e
vHIunf2+kz36pIVeixG0279yLbyijB2vSfFv9X5/TOP6T5RPZ5t0PExCUL4uj/d9
PpyPCZdgmnAtm+E2zS9r+NZC5aB0JPZ2GsNDnDzgy3oj9KiSr1RmLw75SxysYFDf
cWem6avvqw69um9Buuj8/FwbehnSLext2pF+CalQJUBDS1nrHMLqT3VWIrs4kJr0
PR/dAe3irayPeYQK0bKmpLvZjcOW6frwxM1Yk60bcRHtW5GJ1GrAg3rzlITyzRK/
zF3djdJAbUIOSIbuwjfmTWgqrjLoaAG/INTsbZlAaHSliTs6f837iILbDv52Ugw/
W8sJcEbaziASDp9SvrfWrVFI8nwAYHS1bdX7V5wCTwRrZyKay5vi1MyAWatISrOE
sz+PvwTjNW1gPNFdPeNfFS2/Q5syrkVOGRM268FPZYRdBOzRvB2Xeo5PXjI8smcy
pvdIrN8P+gDn8IPVV2u7htOWowYkWF1LoHj78uQiyRIDK7cYB8ZEDLSgYZ7/xKPs
Xl1+5VS2jWVvGd4NEHlpOQFTgPmIBMVqzRGi4NNB0HBW8LfHUBcqztoYyRRKgU8u
e1lj50jIEUcHaxPtF7e+4XWuQKjxHEgD4DH0svIapSXSqmBNEeMjpPove0JEDwaM
6/nU8+FeKHWUGEdPeQPCXnlnDTBXKmcnLiZpyZXDQjQx0C9byd8rnZZIKZCwj7XQ
LJtcp4nTywNOPshQk8vIe3yXMLoL/47QvbB1hYlZNdxd1CcyVhHHJU5+z+zsdNTE
9Z0AUzMmDxQBtVe6oedZpqAQixGckEHkTHktmPzL4Z8iiUgYWseu44rwp8fnVLG3
V5e4A+UHqyXpfu9/V6r1NCzfyl3WIWpcan+ms4To+P5S65kVmaD6N/lyPsggm24s
EtJ9m9uF+F9X7v17S09Zfm5ziET85jrmbfsutbnKTkmCErQnKJlhSkBAGWe4HW4A
21uX7N6NSTpuVN1mm/a9TvuH0C7mXsT6AB3ms/3C6f207n07C0xaSXv4XRDhV8Kz
RKZj7GkMrEVgnRg5oDWUHC/FMF85DXNa9FaNgWeP8DwuPdAU1IDISZAogOX0V67V
Mqn+dA5CJLTrTkhA1WxsPyASRObzqpyWvvh2mLzLTPpMPHaHOlmWOMCm+TW4liUG
O4PlC8tsx/CJNI1jeYmd8wbqYJtKq0o2m6rjsN9b3Akceo3fizkY/4smT3g3MN5m
D1F4JCvkLq7uWFj+mRUVRjV7k7juTiL3knk5XCsntJ03Lvc9T1wlwqdWet2+mVG7
dcADVawPfB07JShC11+JlT+B1nIfBN5uZlyVLNjq91pZPJwPIQWBG7WYxrJdo5p1
XQSuLTEHhbosZW6+J/Mjz3TwWAcKtwdauFEJnpldFf8FSRGqaERg/NdqMhMqfJUD
fIYuD6GcJisuvDjOA5Vi27UUhnLs6f8GLERS85nDxi7aNlX3tsq8uqsLeLbSANXE
8C3whchzcOsdKg25t9joaqVADSd++YNp70K5BoDBD8xE3uiaJXM20igLQLtoF1BT
KxCP3Yp/Gt0XDNzS250852wzDv15FarulQONj1dIf2cbUFsF6t3cPrtXDdfbght5
MMNI2v1ftOkyftbteRDClQescc2JXDISkY4W+7+Rmu4U+NySvUsbfRnrs4Ao6xKT
nM+duUZX5z2aVE7IkHoeSEIDeKjeIhAV2Bc4zdH4FmIiChpkB4CorSc7EfH/3syD
pBJtQzmWXX/4/myxr5i04hYwK5thLW68cvfEboyZaVI44EYmSXp1cx+YypjzKaRv
6cpuqYd+/YmtYaOorlXLlxzxSF3/nECiFX3yaIgPc25tScq+pYIkzS2XJbz7sCZv
T+LS6seE+xaiKS6q6+YUIYVUo9RBp09B0Ub5gkgeR6znKFAUZiREDpXSvkg++Zwv
v89YqiwEYLmwoZAONZ35ZaRM/dqVklSW8FqX51OAKBevnbOe6lF7aXny+th5snNr
E6PvycIpYcI+ZagxlofpdN2RPXjlU3CGUbVKGfTp7NGsJzz5s2qXuwFkUJ9M7Wp0
50hMDvjug5fzYCoAqD29uP9O7qraop2hGcouYKIECaLO4kSnengpYprhN0pvU8qH
D7dBuvrn7vi6SxzUF1I6DgByDN/R2hjqXt8klC4yQ3H0WTUjfYdeTolVjmPqxA/v
rKH0ZixuRe6nclN7esdeRymLX83Ny3Mk2hDz+1VXHZhMcEieEw3wpgQHsre7r7v8
5RTikU/fIctG8MTAk4jejIWdVzDCZJj/jjD2gnkwFy4Q6e4ruE+D7tGrifZHMWWb
2dlatGQhfOovPSO0t1RFKG9iL3NGWE7YmIfH3aPZ70K/b7F2apmAP9Fd3B32yrW9
O25TpFGAN4lscyiqkvSqJR40Ddm5QTaVvFiNCnJrkyFtw4Q410olejrBF59H+jWk
4azJfimnFcRajtPvGI+RoswumetpyagshhWDRQMfEHmMI9zym9Fvhii6UALrM3ao
0WT3s+Ze1bZ+N4qeL9syEoWInJOwGkI0qBMlylhyIV6XIz9qxNMs312OrjLIz+yt
TjBXqpVTOPM7EeEkeoJ6Ax1yg8v1UUuPRp040+NQ5j03XnhPr4RDns+5hpHP+lQj
/ZCaujL+i6BL2yhWSJ+88gDp5OF6nBysdxJq/ZswZdh1ZXlCkAQ11btLtjirxbmD
kTvS+EJCoo7g24pyDy6kroqfYGjHnfhpxL5V8hqNjFXXeqsvogpkdmkGNGTS+xp8
G6FTfmk7XuXvNm+oigtZZcjvZgN1UqHk7tpW5mLoE4+VT3SI1UcfcbeYgFGPJfAH
qQmgbDbyh/PCOVSvpNC90EK2p+8wHHsA9SUREyvLNfcg0or7e9ynGjCnrURRKzj3
zBh6cKlMkoXAtqIeBWI72HQKpjl1lq3xomSGnoGzx1zL3OCLO5OzBQZTkeDknnEw
e/HKs3A5X36tTDgNKCgvHwTiJuE8TWOQWl2X8i++R9oFoWTAJVIP9FfYA2x0jz3J
ZyggarFRD6tM/Cm9Mds57L00MQQpRLfuNSIcrFlaUGonjZWd3RVzeA499XkLMgTN
cCjVbupMMjkKT8/i0brXzNY3+0v4Zi1EYCP7+CjxMdAXVbGcIfb737HU3o7Weh6Y
d5fF3LNXA68CSO1wx/t0BLU3SYMp3DCF15JVqvxQYHyCOzloIt3Ve2quni7rEv97
2nPDcpENBcBRhaVVTZqMMZsMY/+7PVYWMse3zOHjok9CDAxJ+/rf1A+e7/BYEjyf
g2VnWnEK077hd4BzxqaD+8BpFb2C9Q7Noc79A2PridgH7kSoJSHjOJa/SVKr1RJw
cQZ+QdT0mC8i7ZATMuMXcgeXIeOAHk/i/8QLoH3AxzI5bvP7CsIkJMWFZYSKGbqs
U0wrwy8wqdhK09OMKkzSlF97sEE0LeEjIdtn+ivj8dYEat8OtBWyptElNbKnqKbP
L4PJAyeIomwlgjlRem4OO7RWZhcE0ctIg1OfuFM1dHupqoYL0RYQtfzHOBzfcihu
mw4HLkZQYsT7TcE36rlG5/DrbGUtVZMb96d1yeJR5xlNUYxmj+aA3A+i01ZDGUIh
GSiietIuAZRWj16C68sYv8xIUxatERO5Cjdgg8AikJYCC1YvP2zc3FoavAoL+jZE
IonQ+w6Ht9/QrJlkNUcYWnC38xuYZhDMYzzCAWttntPF6c8CILbEa+WFZif5+JHg
iFsgGvY3LTPNGXWtc8VNBcfSSUl/7zixLxI8F2g9GhBUvVEu8rIueAGogetNBEs1
YXRUJpvVY6Qxst23lvfcj1myEh4LSRTrDBPkmOK+OKjMBfxGdPUZk+T6m7RXmGdQ
YZ97/NZoYHr/A6KECrjYx9tSkUiykyzoLN0in+Zt3MH1RY3gBo54T/wvGdDg2KoR
bd+l1zy7gqMu1hxLnlNiikE2U6ogoq2IcyvymuWVvVtAL5XRbLNaUwgtBOXS6oLe
eWZ7+5ikU6nAKxJBqXzpR/7SgEiY50gB2mrPcAO4tokmoe9D3PRRKaAxWyGMbRPE
b8yDWKxAcMD+uV8+j9Bwf6uMY8PVWXSvyffC7dWqENGmRU+WY2ulfGrdtBZpIdz9
fVzX7zw9E3nG4ADMY+RQ3ORXH4mBKV2p7LfGqCQphPzRDlYEdrPiRkDTDWz+8FBa
xtPPk+T8irjJaMEwGMt8xJtndug31CwPTkPsToTCMl4uPGvyC+r6F/x7gYiiFSJj
l1uLqeyIlwaf+61xt4AJqx4Zq/ARL1eO8LxoZn+8INT+SSwGZhG0elwUXVOemVw0
A/cmnjAUjvIFBoaegpb8HDRg29S10ssMsOkWkLpxIKZiILNDQv/gcSI68O+rJ194
YNUo2pfLAFqpnEaykPkFUrNvfBEhQP5YG/SORMlCmnGXPPbmS8uQCo4C0Ki+nBai
xHPYQnheO18R1yR2b/cnWN7jBTGroWNHaajB2fxCsQNlX0bGPbon80sZ5yM7FaTy
nTABzMMgmIdL6NHDw2/z6RXzdoFOMaP+9UpK/PrmYL/PZiEssihapgnWFUWjV606
DU98GK3VrjPuAkLueyeiN4nDsNqK2iJE474C+f8PvpmG4Uy4M3Yd42xd11PTWMT1
CTTlqbB29PYiWdVbNZc7WJtiJSfDw2lvQsZYqXeyqrmjVMygf4Yumk47RiGayFkd
Xv6Eqq22IQK7R7OzO8NsJSEyWlJ84xyhdQdkogbaEP19sP3AYwBwttWdMYrbYrLW
LtWFKw/ABNW2T6IzdU62bPj3ixOmesAHWNOf8LVSXnAB4fo5nz43CJtEr0DNGCvg
c27jphNHP1hC3Q+jLeWA+1iEEHoNYOYgNdm01OslH+SGZL5DEflimVxv4diB79B0
l7ZP6Y0BZhRBQE+hXxvzj3JxIuEEmqwtQO+Oa7Jqa1RxJ26va912im5dCvjv1iSp
n+JVJinJk9nzG0CH54ctrsvbK7INUfiKFIOix0bxN5rwX6IhspH8RplfS0TF1P4a
7c8beSi4rG4bL1LSgjLmajpPFCMIM6oU6I1JgBZr+86wR//9BQQbdeRW0vIB3BDd
GZAnb9SXX7exgH9y7tgtXS8R8sMbNoM+xSNjuEQaLBUYsDnaEwhF1VJ0CvZD5OOz
iiz3/OMVSeorCUxHt7frP32yXEzj/ukKfi4vWYfOy8t/9IOpp/LwaAEzsuasHIQH
7arDiKXhuynbiPh9qRuOWUWqyc83C7t+QW7wu7PPsdEug12IdM5dnnyT5yTDf2CY
WHX1XpLK9kJHcOtSySyvb22NEW9D1ICS3sCZPuXsGdNureeOJHCHRoMEsgoUxTn3
Qy8YaZ40LCBLx++/rwNasWQyr9A1cr6ulzIfTqXTmUM2+4MAZ1nTwdi7vNBICLHa
YTycz6zzCB4Eu9nAk/s7z/QoN/PbWEgYBrga+RQuulBunSjDI8A3EhAnnIqBsoQx
UKVO3qnRsgLNUc/CF9UAci/TmIbE8Q67eCcplR7XVQu7bS/KVU/pvJjsKUpk0pDu
CjjCh9nkL9HRpgZblsfm8eHFRaLS0iUewuyc8eBKkzs/dqw6WezK+yWAn2JAT61L
SWu5RD4k3/3yzjO268YdQ/p/Y99jvFe9Z8YJ3aoBIDaIU1wJFYZKruYhojKbXnXq
oKqtce4SfflBRFRSr/hvBHEa92B0FeBvj6go1HI2GpPJ1L5hrSfp1bJNpXTtVmjb
sV/LJSS3CY2YTluLKChDBLLHIhj82IKnCpJVm0KYbSNu0Qo3JKjnACzp3AP5F4qo
bkRvwpQfZSmWAQ7BUwag5huGLddDWe8EC9SQ7oJMiQRMQxTgFbrTC3t2B6Z+jTY/
q3PygwiGi/6IGPvfP97IwnQwXzkZNKokOpxqstyBg8jdCB3la08WBjHXwcZvkp8Y
4HK/OgornhsUilcBtsTECSeYQVvoyCftUNn4APfjepz3OyVMhKToeRg2AcG2D5SQ
c+PL9i0T8NDfuz9cIUd1ePUBn9fJOolGga8Ua8C52caYmlkFDKd5sP9oWg3iySke
L4ifIQsmQVnOlZNqQUah+rT8YRhM5ygzbkwJfr4be9F/BUklRBvs5+MbrLjOqqSC
t1zoMfLDUWaZeGv76qK/4RvgINLFUoVmwtaXqMdh06wbGMQDweuWj4jv7QMOJ78X
Kd3qvgL/gc3ZSB9/coxxLs6BdSQH1MgE2tdDd6Dy11qgL55ZM2cUINP7Z1KcUBeW
Cahwj25fGfSmlGynFogmKxk1M18dy8SQF4PjhYmGA9d0n8fRLVbSmevx7E4ZaJHL
TeIsA95dVbOyexaTp2wyOYJFDvZbQDsjxA3n+howLgyuaTbTV4kGdSOQEbHntJib
ONEUkReR4fnJ3XH6s7ZdIiCYcQa/6pG4rOr89nr/c1Zp8e/SjIzIZuEzhO3aV5fp
ENM38+AMDKKl9nd52p3H4ipNTw0HRe1ztTLNnE5lw3rOLy7R/vbJoR9LrnsQ0qMT
hy2p9tBmgYNiBbLtUnyZ5muidSbALD1opGjZASWWydOqJvqEnpv7nmLWuQm8kW0e
Ue3c2Py3T+Y6IDZbg5P/KhiaeLLIgnjonFZV1vOLf5MfBvwN//A/mKWrrZsselT/
lepYAjyJaZZdAs/AE3Gp3ZUa0mo1JSyhc+7iL/o3VyYsukJyIzpYyaOpXIg0wG5w
8/BX/bXiOgWj65jY5fVKqaZP3hUgQRDnhPoV55Zy5BoGiW5Q9gGyWuIzOH5Bx9Il
jrJM5fFBjJBAopB9RWLOJkZx6I6EbeHVne5ocYYi0JBMMzA22+OHgxzZPcdXqFnY
K7Sp10UGwtlsK/tmmYxjDhRufaffJBWvb0Wxai5tnPUga93wZy7juGEDioGjIsJc
ow7Mb73wqdoC/JEAE2iV0MKu6wrOy4wynvkp9UlFpdu9fsP3Y7Ht810kV582eSBg
AlVXtYXwDbq9jY8WWy1MQVNIv8XWCkH6PSrfq2EDIEKKv4DMYBZCF8PrrIYfdn9Z
Z7xOFD5De3QcW9hvH0ZW1WJ9WCvq1AZPbJUquC2Vwa/vKLBo79ww8jM9tMZzj7nQ
hbxeb/lUxv6eB/z4oYFfBks2ZbviJwz3u+ZYXSrCqIUy4xCWJh4yx6lKAv6dXERj
NeoGu+HEomH4s1BM66ItNFgiRStc4/6/p9FF/+VzVhtZVUrzoP1lwfqnIiqLEY5+
ftTevdTWPhn6xUrPhPuxvEQfJWg0vM1zixs20zA5va6qzbCYFcJ7tEAP3LIW8SSw
8HX+cfN0c1KSuRpe7TPFUaswC/wjYY/ztcOIvy18F3JMkQ/loOykFGXqt2CacRDT
psC7CzMpeIN/TJaISc0CbdlUGrQhN05KQZMbrXOIzkYtsJZdRXSkRcD/OFxD1xOx
HNj5isrISCoxmeiMxL5hzYMjeYCkmOgXjU/mPuIAdH6pK4lSCdv9jAo98BLRCwlq
6DBJSg2czjzX08O7acNbSJPrhbEfprGBlCFcGro4ibP1SmR0CwUy8oNX9bKfJGdE
oh3gNPa8r+BL4fPABremqDwf3OQMQZ4aGt3dBFgOSRUnupaZQOadFvtrZhRXK975
rEXELNKYff0kWJeQcQc9r9PCGcYRwQVh4FxHgfFn3b+GyKS7Ae44bTmqkpJKMp38
m+asBuV9HlBwCL3q8FQfpo1tekTGashcw+XvIScooP1lWfl1JH6PtOUzKDroNXGy
E633bGEW9xiF97+vvUWOZsj6zTT3LODphA01fcKQy2HTLvWqWrWMQci5KrWlxCCk
Bo6+Pm+H6gNkXWhAy3sJdBEgHAIlNQ2zSGMN/e+IiiRSKSig7dKMmkUwx5KgzLn4
P3j8D8TG2aJJesXYNKLoaklK9fOnlACJUTIiU4CQhzm515KXHsNtvc6kkG28wcfh
HdglfS/0Mpi3hmlsiciPlvBD244o/+X67cw0RTp9muSnKjyVGaha6cG4CBFW7XsO
n8KcbnHJ1qn11Q7NSnDyy78qz5ECe1wxZ6OH5uQx/J5q8T/gy8LgdjjEf5NuyEzE
JNSABHCaRHclQUkft8iy8zu0BQ4XDGm8oD5+zj/+8Q0lxqFTnW1r/DxLyIg8T92f
QcZq6KKpG5CAiqexJi98dWNMDp5HwHPaUWHpC2+bMQdvMp0N0sHE7bh15UiorWA4
85HSztqm78XpJL5nwwv8n0IpTdWWKi0fT1bJrWXPzkxm3tQUYxPFJLmx+GbnWbVG
W91sGKfqehVo0Oaj66YYuEUJlGsbJbwH/uakECDyW2ER6RjLFe6OPGglGyRyoh1E
QrtWglafS3U4Y7CT6p5gOLRjtTpCkflbXFG7ktRs9qzQUBHKXZtZqQinG3aVKDpG
mP2w6cTycJyFjXgKDbQgky/EdoapfO/NLOD6iwA5ERe9gPxF7Z6kVoRVqwph3KCg
eTV0biNDVkMAHTbjrSsjhJwfPSEG4wNwXG05o8onq+SPWdaDqNn19o55KA9R4ZjW
FRCvo2wgunGqRyzz3PvtItpkV7X5TbvQ3LXnJDag1kDtQPRPKBb0CBzbBzFVpfhf
jcoYlKl5Rzrn9zBdgjrsxpSxWDW2GANITF8lLPWCrRF+B9gpGgvN1+YW1obye8Pt
OlER34jadjFWclLOCAe+IlasGdtaHtyG+29AhAU3VJk3iEtjDG++8ytK6b8119s2
uRjEypQDHoi3hw2MaM4kK179E/QykD0to9npzq1pFvObp/iTu091Zp74l6NRUaYf
+8j2PX1AdgbBMWb84DFNdvPhF9WQ2CkQKPvHzHAsI9pIvUxG0yruRunmHjppCxYT
DRl2Q4mt379Ueh7siflmCdNl+QEPQC37RB+0wzZxDyiSyHWtAFDr5KwjY98x5X/3
cXxgKx9aaZHwGshWnNlhlBY+b0vUpcqEJ4yPD1vKPfVHyibsnZ4pl8d77xJLm9Vk
m8Q9ZaLuxQp8aanzZl3WGd/aM4N93Zck0g6smMX7QY1U6tS2atBGHqDzP2LKnJoF
8DKxfVPPXctac2hZ7G4+yC/PSUESV7NS096GE09wpablz0ucPWHp9HwJuBlkUQTu
h5OvNqfYuwuWs2vv1g5JVhf6d7bFah9lKC4FhrMSIqxWNdM+Mnh73boE6dbl6n44
Ubx764tcb62UGljSeBCqDrMf1r5y+odIWrOJLxqfYRNbZ/4IXor7D6SypohRuzt1
OB4x43OrIJV0xgQ9Cv1XqbDfiQVqlP8yK3FuM0Nkj40DJ0yGzEgQvyvP/d8UHacW
Xg5nYws+rwkvLVgWQ5yGZ+swRhn5XQgjpPnuANI+xI2yeSedzJEWk3TfIwteE8tk
uaCbamWiNple8OtruCQ3RhrIXF+p7fOxm81KH9nhXOU33WxRzhvyEQRd45bgmxnA
9SsXjPz7FZDDc/yb0fZWxyeFfiibP2use9hquxVK+qS8IhdfGn4/d6QlEKAv8ew9
EKetEY52D/k+l5FLRr8VLSAb+48kLpNqkvN1MfAnXAL0fLh74dcFMYt4I2VpcGs7
mZuEHagT2rm8l+TyCDegNIRxVR5r1kQHjZN+I25S64JPjTXK8UaEDzPShL5Uv9Sd
iptHqdVhhXTiJ9F4fhhijLHKwB0xBDW30AeuB0Aj44UnU/na8d1oKBoRWP6U6kn1
nVPk8jKQlMo6uiCRSdvvAmAdrs7mtSvBTwgYBBc/egun6zvG2A8Dwj8UPKLY5eLK
Zb410wZ4fRoPZoI1v/Uw1kkPBLB+QP1RQDYa+aYGFawEEuO601hByO23oDBDvOfc
VMaaJgEpE6oArDZBWtYT2BINO2cSGRM86EAxW9KOkwKo+tLBx43ZkGKPKGfhV5YC
bwTnx8ZznORhNXDX5CqdCwixqUdwAojRghVJlZJ9aS5uypYePudar9t2dM6XETcq
hkhAOj0t+aYHD2ruApcvVq7CQ88kyIgi7AYPYzZ6DazEboXx6ahiBlgllTvlW9dT
FWnPB7FewlmCOHa38EUrcHToFNd4SFJQLinY/znYNGdWv/jJDHWuQ/lb42yP6/e/
7inlyPNRR7SrdY85k2TYSS11QYiD56DTST1biCkU+taAS8OGCW1+sZJbSkIzib6p
NUWcBHYlk7dfWVvfhyY+1eanb68SzO43iO82ef8kUoHCZCzy+7kLqfg7MMrK+8lE
pLoBnxCQIsLz+/t8Tj6GAbSSKWx8Oug7e2dHFPOf8xH67Nr0yD3+WTjag0QrvG//
WBS+110pAzpSmsXkMPLDaYVXcy97N3aQ5XumHCrsruzau77YvCwmr24HmU/SB5tk
MDHnlxwQ/KUDc/gl2Tu/J+IJ5NLHGYWp3QFYWHQQJa4XwLoyIP4z3zRLZfyxFrPC
f+/TQoX9C7Oet9CKi0/O+p4t5nT44Yt9uMTgeWzVdDPVYoPdbZu6k3iMFwe25alM
auBXGtc5YWnu/tiME8BlXl4pwzA0Ra9vIdpLrsRkaQA9anB5jd8pGVrX5jAyCuQq
cxYSoe2an26OV3OwjO650/8CE6EwhZt8bnO2HiTmDNBQCTD/BP33RpKtPrFir0Dl
iH42dcWTtnx1YOM+U5IvBBdyon4LsQwIgUOI9Ys5EkUiLxByp1eQpKa9iWz/F1np
7oNWWwJKPh8TESlzMaSGjsWyfCGwKVINFWyR/fAGC3qH0fGqOCDmC4KJgitLpKRh
5V8N+wLxYKzgpRGfPSlQUiY3CbWhEMaTQerHJVhrrHZvhB3eDH7cRXLeY2XnV1n3
Zwtt/A+iheixa8dZQSQkWsUGw1HW5jfHbefRDevhnq2qwOCEqqAU6jX799AHV8fQ
/258PGFGq66LgWttYrM83UNHkeWL8kNuy/hX/YQenY7GHa30K+JT2JNv4oDAdat8
ftTIOdWZomGpmKDcMJYpdjfiirIGBn6zpulZSuEByhFYclMMH4gqvTOT1lXVKIZt
kzt87K7EP9sgPXVxtE+yAQRk/m2dWHwMKz1CO+HCAfXqyNiYP+V0IOAAnxiyD3vO
grWjX7mktO4I8+gVqESlprOYOR8jmaGhDnXTFxtwMdAS/oq9SNbd6RO0qIGO7CQX
vzENbZtjw9oYN5b7l032dvhSeT6YscA+c/rUe5LU63r+dIfzCKvyclRUFHxZh9HJ
WRn/9lnLjAiCmCpbEJIIGINRAQT8wjcpWTMgiJI9VA7QNyitSjgfltAp+cvG9MPp
Vq1JsYNj9OhKAwZMOagVfViMMAtSksJWbccuOHSs1O6n6VxJZntWcqBqMEDnmvvz
YlupvHUnyCNp/XV5CaItNDLP2NuH1I+nAYU0OrcaCUccUFQI/FSF2DB2D4TVRqh+
TLZ/I6wcLp1PHp5NM6xWcYiTHuv8AJFd4q0efnTrl6saZDy5eB7pLor4LOhBubuR
7pm21ME3RNA7eIsr0iBjRaLE8+vyAvGwh7JM4NZ8VjaevPquQ6GW07K6yHvLcgqM
64rmB0gpL4ue4uKRnuqzZPw6kQ8+vUpPAO7QuckcZyoPgJwd14B4za5VwBVFFhrG
ebNAddpt4wuqj+LD/IPtoMMHbQN4gSN86gKOe7bYeuHSQvbyrNX/I7Oh/tgiDaJy
5TJ7+9vtYbm2Z4Mn6rC8z4+BMyHtsX0ekKvcpjmyoUPQKkzeTXa149zutorhOdrz
MrtD6454qz4ao3LISwS5ghnJ3ngej17ru4bRiC+91U+A/poqhKtcy/rDyUQL674D
cHj0FDN6NRLBrHk9OpoP1JaQVCEu6QjZlm8MzqeJHxYiyucWjapOHVm/zH0TlV7I
1MJit0QsXWVn38Z/jbrnlFD5WHfmAcdynoW20zqqa4CaFCO6VgPuJ2+MVWQdzWfT
K8sr8GSyUVOH4t1IbT+n6EtngjsLmRrmYXpmrVsVbl0ZOpcqho1slNIS4f+OmjiJ
QYINri8UR4U25UZQslF5Ag1g5hnzaeFQ0OVE2XILHaYvYOCJsV/CcJMi3zf0/E8e
zLzYqlBkniIiltnP9Is8F0UKVpHxEYqZV9T+eQ7Ya8P79QVygTTzfgaZ+b8M5Yw2
rAs7laIHrlBswlBlf9KzeTwtiaPX/H2X67ptfEqs7FNNL/Mk9GPouIjmys+mUxMp
zeOHJHms3L8HjFvbjRQUs8bbt/0YeFVxBdc5wVxqhZi0rOH1BoX9Ls0ZWIqPCSCj
diGmLqOsKCLZt1oiKzucgRAcMgIG+0d/A9QHE4vyghTKnjoO+GIb/vvBuyAi8Ul6
YqHv8u8iGJzq1JiXPoyJYmtoJ3x89MZpFOcNGp1ZPZMes6G5Qe6iYVlmJvWIiy8g
lEUUxMSo2RjPiT2+EdiPchAtQwDQoXuNGxg7HEzClUecwyZjezF1PtRKs+uGvcUV
MDwxfgrjsFZbcGzSiw8TRtIhoNReR3nemHA3CIYVoAffNCinVNFlghpZHrBE1kTK
YyjsrIldGyg5iwYC52sV+1Srzplco8JbhQuWfStkiQigRKwe6vqqHnqUlk0az39g
AIMHN8zXfyEcssVum3wWa/HgmFQJyUBeAF+AYyZChuS+1AHD+iVv5oxxz3e3WFIr
IqTXlwgZeSF3WpZTE9/ZoSOIhQyVqb6Lt+VPUc7vz+rosQe2gcW9HfWED7gZUuRq
Ja8kafORerv6Q3wqlnJyrGSSYsk9WM2Felb39NWRY2L4mn0P3p2Gr1oCxugakCLY
FY1hrWW4xTaFBmjgAPxZ0DQsO3jzimBNUrg7nkMxC2InRLWdQBGTfjpkTvUPUWxV
tGw4IihxFRai3qLxPJH82xhmj5VboV/dKk4sau6S0E+GI1h86MyS3Cc+1u8V9eSb
ZrUPYU16UVjoKYugkxV8Hh8rVWfZJcbPR57MX8ARwxaHurpwIrZAdmE0vB5YLtvb
TOH9yN42iQF8U1fkZR1eN9Uzzd1TMcBPHa/X9UKGpVcC08q+PFpEbKeISTynxw8e
B8LrmehiQSFmLVm+2FuhMW+S1x2vzqKnDYvqHWH2ff6kwTKgSFUpML7lpquWY8IM
Mno6oFCdJsJwPZYpbrPRK0ANg/rJdyvQ69E21Q3tPGJtE+xKV77txP1//azCDj9L
Q7dSabxuaIDpVk/gohMDyv16m28kE7VVb0cdQKrHnBG2svzd42+oF7CPX6nL0ouI
P+tNVt3o3CU+YIJnWORqVIDqdVrh+hKm3vcoBPwxbptz3xvctXa4VwEUwOStF1TV
F7IffKoW3+jqgajQGctid6AMOdjp++ZcyBvjYhlq+dx/b/dwc2zyn5y4lLnbgNkh
SFaNEzUAPv9e1dTVlRz1F0AlnOpd9UsCFrwlNnALzcA9CCYEuceni8crFRCvwciq
3XsVumyFY0DbA36MYcii353W1l98zaNBDSNWAPPDLVNhb6W3kGeZcWdgfIBZYt5A
LZ5VoLTdiGPJ4W1kCHt28AxFkoLoCJTY0qcmRzwRI0y2QHYfcaHHHWcz9Pl4ZHme
mWhoTVgdkD4UVmiYD7IZzXEnoYtdHLT2zd0KUXndz5FV0ubeE8WSA/lenLDyQGjL
ejpVBQHHTTTsxLzRyiNqXMx4Nto91+NaH4vby84NyEX7Rpn6q/fv3C/hGi/l/GV9
YnsOGQQVTGW3tO2cUKrkZKuopyN0U3/71Oq6Rv3IkYZZN3ARhxBg1teodYh8zsI2
LKvEChVAZ5aFZEw21QcxyseV972kIG0vbj6797iIZjKk+snRIUbi2azNFTtfwHBU
1V4xWgLtGOue8x+zeu16siEohPmfz7nJ0YMW8MV0Z9ZGHdAV8aLtxi+QoVT6RE2t
e98U7fj82RVmhhlgO7xMIzcgFr0aTL/vnJQ9+8Yg95obqRtMULygnOiGePFH/l0s
e1fbsag5y4mVPNmmYpAOcFdg85YTPhP/PLjA3ApwTtKKVZw6UpeUSVsJWv4O/N0j
bvSm/l7ZP3pnjGkNQQX9dPcIk2fpDhfiDSq6tQ/4dHKThgiDBwWT0r6B6rAFMzEW
BY+HjaXZnSC/pjeG/qkdTkjU5CnVV07+xcz7Vx73J+ZEMuRhIfN+/0otLILo+yE5
PpzkvAUZA9PVcyeoOw/sT4VqqkZUJR1Uhc9mhTkY3p+RrQ2vHp4rGLkxy+jpriyK
DrF4pNgnvIs643udlgMCbf+gr5w5ubwUrtKg8Q6kO/opd9t4NFniohCtHkXb+xIl
5vDNS5Bu4JmJ9NBMGXb0Z0AjPJWHiN//WlQrg07nLTLHlHMxOFptwIkbl7ne8ru8
dYZrtyql4q1v5IqaqNR3uu1BZ+OMk19xdMTLtXZdTROrmXGzEjhP6kuAFmuBUu4a
oGvQvZJkWGhiB2R2Crl/boJlQIB9os0+60q4L0Q6GkmQ7OPLaiJUp0fbmvPtEMu6
ljIA3k8IPjF6S8a/3RmkQpRs7mQMHpkxtYtGka/CV+xrDL/IwUPxc2QPjYmLlK1F
ASRVcqCNnoDhJKxvwxYX7KqQHe4pPwTI2OMRg9oPgXqc4L5fMm02G+ancfUSpLWX
eh2NWMskGyHZFpf8Zrrfc+wmKXlInuwpR9qqOf1w08ytD2R9iiHiZXjEYdWJIGsN
q+6Fjl3t9/YiaWa+TsL+k7IH1SbxLh1KiVUzuXeI2KtiRt3ymmuEColYJ+6xYu99
y51VtSiG/5KfTYtrs1Qw+eQ1+V9Wyry79m+UZQFyKcv3VBDdYZV7Tof/vWRrm1BU
MWM5R6Tihszz+aD7TbOnmV1IAfzpJauB5WSN2QC/SqMlDKv7xdWGzBslFQP+Q3dY
OjfcX8ohRSdVhAXnGr/dzWuDSu153/w01pv8RRqpUZea6Zj/X78tBySJXOroP2xX
YAjRvOtJEVrp/AL+tY4py/PH0lSVCzVg4NPIhvHj4R1BPPrI3vfFloVn4oImo+p/
dNZuxyLbGNUgRl/le8wVB6PH+IvKJ7KyX/0cGluq8GswPgNPzFyInCrVaRYnPVwj
tX2W9PgVVmosrYHHzopTc3iPWFZNq7FVAAnLK1rozaZ1MFrZ92CXmBIGm7PmFA9G
JL++69IwHrRmuxMiT6PQdPSLzeo7H4JIXoESBBBvyjK9bMMisptnd5wpdxSHJZSG
OgmvOhZNBI7bPP2ueiCeLQTGde1Eg5Z4dyRyNw2KYJf7h9Nz196VtQtltUT7HHSq
rufewBbvbbPjGGwvB+1W+3mGSZ8+HeuWeCYwzfK1cgLLQqt8Z+qwXtd+Cgrd66a5
vqkQOWqABeid6S6GsrwrOeoTlprLYW/aK2JizB2Sb6OrLJEldtCYlJwhhzKqo6Gr
dRjp8JQ8fcLfb2a2T5x28gxAwHCizNx8DBosRj/8mfnJ91OL3tp0TP5CEbs8vrsH
NrNoS91jOWjeZPFaqha50K3XIeFZVnXHd1arIueGZnw5Sx9wTUqsZDXol2H2Snry
astmVmPCG1nJYrIEExnv5w1O1X/TVkdIM9My6+C+FBm1Vd9ojd+rRa5PtvVDWHsN
AMt8t5CE0UeiUY3KQuiq2luWdJi1lXTxtqC5seJ+4z5qmahGQQDgQyXELRVa5SIZ
yGY7IKsum+7HWI4PyTcAjWjZM8zWNFpAc2WZBpXP+zo1wVyNmfx9qEmWQ/kSdHtp
NN2lmLCEVSVrj/gz+E245PqcHxDeB0seNE3BEltL6ZGULtgsRxVaV6YKqj1yTJIC
VRjGBQbUcQNPhOZlcGJEl0dn7mFMFMpD4GQG5nEJU+55Jknj09pCfEo6aGNTUBu2
7QUWE3eNwCjibl/DuZsVa8NXaG9v1cvMnXxfLG+phCz819PnlDBgMSflMVr7E842
A7IxGpSwO0/Pe8WGU6v73hDxqEFm7Kdhs7DTn5NLMGFzcUUKoQkQSlEB5net/y97
L4vY6s0vPkSZU+yKSXkMwU5V/HW6m5J/up/VUfIYWGF7VU91Y03niQOtGLgKwK9Y
6KTRPgq9CymkizuK7Jb8IV7BxLJUA4yIJ/lCublj3ilXEPSHNIox6JfPyfbZXT2U
CVHnUmN25qNJCxu3bnlBD/5h+0Sqfd3sM3o5CMfu/VFY1PvpyikWpJfwBE4nE+gz
0Sx6/n3JMUuQ11KYs2qF22xQlvYtcEqUuEipROyuoyhfutMmyZSgJZ0HWTDvRUx/
NJ6qXorqdoXk61eWP/45g28Cwd86tkDZmmjt+mWGlBCJpSibugjI0g2w5PaNW4gK
yM7DYZgXCwk9eQ8VxVDdZC6PWdhaVkeIo2YznF4vkh5/MSC9C1hHvbbMq0gM9viN
k68SKkIWfrnDixpMpCiV+KSuLIqSeOT5Z5NLsijMIXU3fe9NdFBBYIdPIskhtFXu
U0EgbxjHAoTf981M02B+oTGBgdMy+dovRcCZcW2Kwb1lnrNvWbVdaAoKJZUkVzvl
9D0N3/sOve0fk3eUVPvy1Oct4ZKTDB+wSwpmXMauTVaVahLoFmFkixudz22dOzkR
1wpDnCS6nZSJQFrDarXVKn6NF5dm87WmTGGtm9YkZT1cduw1f+hYUY70BjmDdZ4i
g2gnGDKysBYS0NSSmc00QpWZOzTHXKd2GtNoOHS412iYqibqlCj9crYizaUQJFwA
L+4rtLhCbxrjP68IVVwAanxr24yvxjZN6x0mL2e3yc5oQ/Cmysan1QRdApVtkq7Z
oxGaJsP1ghY42GciXn7cf5PriApCn02Mpk9hWkARCei9ik9Y77wzIOv0vZBdClWV
RmRKcL0Q1VN6y2V2LhFOtAfDtWGpz8SCs+zOcMgoNo3Vf7cV+VERlEMjV7aYi89o
4lSc76mNSx4IyKZZLBrIvSaiHBQFMW0LAadTW8dSUxGmVEQHIFs4h79apwUkTt9c
GJJ6uWqsr4gv68atCNphbDezFQyg4o5Rzp8nQ8gVctOe0nxDS+eSIzXfOMt8M+DT
pQLXRdhyaN9+hcz8+xQbyiCwfbG+VDCAlLG/QT5x0iyq9CRGX4AHOXjCIff08B9c
85oVL3aOilEE2iBNl1n0wKjh5lLq80hwpSTtLxZZxXZa96Rz2zG7g/y/HcxcPRbk
yvSjYzQCgl51V19X3dhabtn+1SHfvgwtbOUYqhOVHxMAFCwJEwhTIDQU2UCFjxM2
11CzX/8eyZimIDlp79umdD77rWbVQJQYABWG0wpYvoHd6Oi1Tht2C5xLrU/VTk+b
skkuaznlRZBufRbakWK9yZg+Cn5+/8u1ZiYfvL2d+je2ETlqRUd+B+C5siuCK26c
CgjdpS+dsd6e60KrpsCQuI9A2LtC16EZZnek2e9CKEaoDjsvdHT6Zl9HwFJ3ITB3
LikGeqhcjdegkHiuKy2uhW2JRjyNw/VQ/XBIu8smdrME10EOlN0FITtqIOKTLPwR
17CX7nY0Y9ighOcRL9rzgSJiMc3fyxPtH7GM/2RWalWL00ILBMX+TKi6/6NrW6d+
xPUv8xmv6lTg8x/uIUG+vkCa0q1++9+7R6FeorOVqjMG2CmIVWyVuNN8gq+1QHlH
h+h4/T+iAj4oKlkIycURzIP8DKComHeKgiZiX19UD46DqnLPI+lzpcLdIX/00Wta
V5pQDbos1tqrkwlu2SFbNRksGMbhE4Ee3f+XLnJ9HeAWGwBEPLZPtxA1AC4lkbPx
kaqzvEGc6OlVDVFJOZ5i/3YG98U86GvFrdauyCdSZlcVCfisXKHyMNRTAa4FKNz2
pmulXkevato+tskChhb4YL2OnpvWL8vzlNDhSr+mGjbhAveZq6RhNhCTSoV2FpeH
sVNYl+N5PvMRon3oTCbQQbG7kSBh3FYWUMZQPBdqxW8dy53+AeZw6J0FEc5mz2Am
QBvGpz4vDfWPyx7QyPQ2myvl49hLNiL0dvOxJL1sL/06lwez8+y9t3UWdwLaKhma
D4FCViQ3F5tG+Cns4rp3mL0Q7/iD3p7sPopSSWE4kpGac3A62wKmCNxaGeP7vzDO
T2/zbPoZBX5BJo5KrEt8hwxEX0se8b8+grgOtqtyWR+3e2HOq0Rb+4yEoVA1OV6w
L7DNZPCmJWqa+GN5jOaLf+ooVB8hbpLzBLZk2qwrZ6xGhm+Shc0ei0109SJlXfik
xwN0dqkCcxkuldUqPOg3aP/przE+rl2AS3v2tSGXo3G3X0cTwRPFqAWs8u73PyOv
35IHxOPThseMBj1zHodxqd669/YesCMgDu92CTB5tp3cpdFn1IQEFpSumzL05nRx
jFfVd4397/fU2OBiXgABZQQuz+thnwxvlph1pACT6QCksGCXF1cw9zATkoJbJM7E
QcWtY44l6H0y8qlmskZUdisvr2NbiGAcT2gXjHFfJcKLABx8meztD2RB/mRKdUVP
l5TFjYEl145KyOh9eDHUoOw9h60SIUOONIZvADaDnYDwsxwGs1hbnJIdgYILP9R9
tk4UnE1lusdbAD/llq5FbtxkUUN1IyXjyihR4ny1Re+oAUxWYZCGvrCup9/T9fJy
Gc2Wp0rA7WhIdYdONZwlU2InCR8GU99Mdx4FNIsXwdy27oS+0v8KyAOwG0ieiElb
B11tAKEYcHELDeJMppSWwSNERpzL3IQLcNtA5/1qN/eMF91dFNNuofFSxE55goOH
K8Tyw/d/c4mmkm89uIPvq20NjJpWhO0RtvqrlUG/Vma4ctWuzMX5cHowK4U0S3Tj
bID8Ff653BeOulBvB6oV5CbAqXnz4sGFz/+sD5xC+Ks3SO7LYUe1rctpRx5Pyncj
pghdffSaYO+DF2rHatz4GRoE/4EPtINEmSAFadZQyOQKWz2cPwMMxXrNS3v6menU
M1lMZ37RgUL8dUWtkrXRizzgyTsKV6x9RVps5ubJQMEjbAUp0lSCTDV9UrcUGDJy
8r5iuTP0OPmrDLrg3YTCpZX/9FYBm2E0uNuiENfF0E3n4FWZd9CHpW66lJNlm1zC
B+VE8EzzwVBXM33DMJnfoUrEwBNKV0/tZjm2S84sGVB9j6vsDquqJHWv2pmYHECf
x7sICQwLpJoJMfHaTW5nrrTHBXtYOkiGXKcIzBJfCkwJ9RDgFeEd0/9NlBh5gfWH
KAfQdNrgbSdOb5lvVGkvDmPuhX4RZz0kJL31qHAe6LJPU0DF96n72bqlhlQ6aH2d
wdQpmLpIbsovvuX7N+z9nTxoRxKAD+cp/czBV+O1+ZBW00D9qnMcHlfhex/Vx14j
dx3jUYbfYxLM8jbXw/KWk8RMgKSCbJ16CfJfWO+tSyzxdtEPN07MEdDEE1YFVfOs
yDhCCx5Jnc1xs5oaB+fEvmkgXVV/CZ4MLzPK76vcqMWpeVjRObuLEcjB9Fe13Xdy
R9LVd9WzJbqXRt6RQ7p9iRLR7RPeeNnYLqGxL+KNAISEhnx6YFWisreW9wdcdHYr
iX66Jk+Ip32HAQ8m5lc6RvP4PXerqmwgMkGVLjgtSvz18FD1PwGZtGF7tVbzGdDf
X+u89psJzTzT6dA41nx7MkBa2UZsKeaMm/n4rh5mpjobUeVjGXsShOhZ3TF1ZLfy
X4q1TuZVOmVn+7h99ufTwobaWN9daIPFPEZWwGMDzUiwg4G9+2vmaF3i37tu0nEU
hLRI+q8YcSjsjlojdWiaqZfmRSmzUhwOr8sU2EJiYfvWdF3g4qz1GEzc2h9/OveA
Z6XLvyDyC6IOfH7o+Q8X7dgituwrlNlcAMYtBPapFp0XxqBHrncAftD8rxsEMowT
iNBzyWdecxredoew4+e5IUYBRTCoF7E4CuJtOKo5l8fmTZXHfMEv4GQxOEsTunuF
x9VOGI058tXPH1QXHnNIfPs62FB+mlRa6qLzJ5GvVMxceIYueiUvLj1V4UYho20y
+iz4pFaCGbsNFY7zaBo+TO6I2FzUxHNBUvWXmTpTNoySkKdX5HjXiWJ46TpmIcAt
6OHOd6J2b53dLBzrB5rcNPVZ6trd6Hi8WiXJWBP6HJKlHFwu66z+Cscgde4SI8oy
GzrtvFxs4nEZbnqqoBeDnzNcYnKUIxePA8tRzhXqELZjnwnzv/Fm4Sg4BkmHxXgY
e2+yWqBJrK840ymFu8cXqC3x9B0QvLnTJqq3mRhd/qnyIwYxc8KsD4hWx6onkwY7
wgEHdXkJOy0OCT+FiSQJpzvkwA+0Eld8ynOtym1imCN+VHnaFaFXpCaV5l69YHqF
EC7tY8sjsVBuNEH0b+3mcalsoYscmUMSXNSmRhGyj0ZsIZM224dBh4NlIFYEHiFz
yPWdEmHjvEBLJzydCT+xEGRK8lIjznd/qZe7TnIjgHyRJ7rLwQrChUjJdCQIL9oT
CSWnMmvq68VRCSMQd6uIWVDwvWJbnDgi7NQBhP2DO23w3kYBAAVCRt/cpNO3xNcp
z+NU3MqAyTbpqK6JVtY5X55xIlXoJlwOTr/bcUmcUuj/aRkDXOQ93jyVrb2U9KeP
sv5KK3qR+eIhRTrPdSaOQe3bw4amnM3yaDRSranrfb7PBX1mhuCobErofDu8Wuud
ay1JcSYBPzaSL8QA2IghrwKg7wgeCJqKffDLdjS99GHFKhFbX9KFTTbWHGSb4ZlQ
BmPUEz1UHuCr9T8dUZjcC3WxO6uoKcGMgKb1B+bgO239RvhPfNK0uZ+Rqa/IV+mW
eLBc3KrWZHjo4lNMxS1fig9d90hY6PrHRRsx4t7QhntHEu2QpRrBLspDYTU9DSk2
kvgMSjw1CFC5V5uDzHU1JtpXWmZAi1rwCU3UNqKV6yKmtLbvCCT/aoFOrYnRM//K
XyIePyFXt4vjc9aQJ5hhULfTvBPOUHZZI6Pr1jBXt4dV7CkZKzc3y0jBOE04dq76
DMgVmorGkIlvr00xNZdiWZghNYN/nblCyb9UYG5BielezAyrCVZgsVnOOAVhHUQE
tIQe0/Ip1tZDWf8yx0PAA7/RwnsLGl+/M5aFq96D2l1elW4qPiCMMZKeqs5haKUh
SpdkqcQE8OIp8MEAMyJwFSYTX+rTRQ6goaArXT4wcujEy7Mtb09Aox/U6QTVVC3U
6B/++jVogVHajNadZK+vcS/maAN/sr4vWIL32hASUTQVQlZlt5nqmmUJ0IrPzePp
dSIOVJlzu1LIYQTOM+WX7F2EuPJoYlLzzArs7JP7tmXcxDj9Wof0Ho/kHbvZm6xC
Sb2WcQPruFmw3F/rJFqxwaZv6X1l6zZZdfXsFWnno/w6Z6HfLBBQwarf1dJiqHEs
mB8o98/lDez0TOfPXVhzc4tCY6zN6DCJAf8jz7Dh1UM2TWsOkuOS4xp5BT6ER1js
iGF9Ow3oF1zIAL+NFec88G/7L38hIDIXA6RSjX06ltt2lX8xk3owA8qzlPskeCbY
PIY1lWzwIFYd5/QQfXxoptkc4auOmJ5byFqi2xWVbD31vZbQB/EDws5NVrO9d0u8
7s853+2ceaT1qBav/nOeKCUAhOy6mWiYOSkO4jGxS3wIfNMFIMQrJeDO14TOsBr8
vhFuub9TAai9p5+9+p7ebFVvVCsJD5j4HBhfD76HehvBIuh2NcC30M52bI75kIGb
m51OHNdllAcAGGtrabIQWaTsncFn8JSd+N1ekt25tXduv+ghuA0PH2WxoTbWqV/u
t8BhTgf2iUVJO0ry7PYhRIVVA5QJXc2QS7EqGfMMTYXcvnxStgZSa2BBAESmp8Eb
Oa99XNawfz7OL7FPmmGcmVI956jdE+cSFtCTqPk4o7E23NWEgqHweha7Jo0mTKO2
uHV7nTP04t9nbGiiutmGdSAlJw0rA0syFoYnTL1DXBujJ/IlqVnFCOQXGTr6Yxn4
E1X4TNc2fG/E6UF+IiTUVWp9mzK50RvKLPIdLVVIQlVel9OkWVdpxural2FP79vs
eTsTTCvcXE+QNyRQ5fUwZZaLrngv+Brww2C66Pp1DM66nH1yyEpAaQDfbEKRgPcD
/1bXcfyucZSCs7PbYDTOOuPftqc573Ld3HarvR/qryd7nfdOF0PIy7F86jaMIyRS
MP/62ivTtuRPodEeVbehRXhlfAUD9h3ktR/1C76sTETlEbAKDFk5K4NgXvIjTeRm
B79LYGWQJDSS2iHY56lo7HX1GvoueT5Lv3N7bqbkNGXQjLOhp3jCmdm26ILaoOo5
m7Hjq6ChO9rZXnyezCnJdgxx9eYRDoLhkd+x/X0HIC0wj1tpT9euwKuazcS3XtgY
nMxblLpvlzoM3E463EgyH1gm9EyPDczGfRuio9RhmQgqmlc1DL7Hre6BvyDxE+uW
mnXmv6wXtxqzZ9hErXvnbqXTgiW5nk1W/pUo61C/sWaGtKzJ0NC/oAUtxkjRV2pq
jSHcIt/Dfinn/sT4Uf6INfY43XzXraIKZkO5osTXMC6yfRq2HYKyxWqHxk2iQdqb
UxdONMDLxkeHR54gw/ilDXrYDD8E0zXviV+0wb9SHF4nRn5d5E1SCVwPXnZNBL0o
8bq1erjAMFBUQahsqyQozq9b9f+Ivi+UiNQb/RWV1YCc3m5sqwDmREgMr+QmdfHU
nqpxxYdlmXnzxlWNHvAJed2dLHBaqUbXZdrmYS42T2ulerwuIu+A2dNwIxdtbesg
f4L7VYWnyKfXfrRS+pz76EHexN1v///EkbbZk7mSokElMq6XD3kLTlwN6rZk61K2
REjc6fw13ZdPabk11brdf1jIgukCeKyoBU8TxZwvcYHT3jHKS5mJE31iNo8+JjVV
3eVsafV7LXv3f9UxQju7jZqJR3dfemxvUHlDaQLzBhh6smulnXQNGJw0/ko2ie2o
xWbl/l4+a9Fi+I09ylmivPyy5O/d6hmu2UA0kNO2XNST7wm1emr3CTyNFq7OKDK0
3tmVuJq4X2WBtobJc75NJfpHCRgpFNark9BtRNiY5kwqYotR1AnwcPlSKI1JNCVj
4cNhW7t2U4WFvhOEuyI8ydA4zzTIknEFJYKyC18zP3iwi/ye7ulM0nRtW6y/UOLQ
YyxupfGyEDZ3oPCUafseJsfNeQQp0Zsgd4tqx1sJQjog1b986Bwe5ZSXvZr67npb
Ro1pkEwr7hVGVlgBrwUeRdiZemte4c4mXpi9+vLKZ5HgA9v5fJS3ykgjL73ipRk8
DvlyYGkzCeRSn12Pc4VJqc0P0p5KyJaZOZUqgHxpSiLu5xRy8/f6wMZT+Haf2Kg4
7sk8U4iKPkuXwtpiS3GNc6eiIxgfEheshdTfroNafEz6sYHjWxf4HXXBJJsYGc7C
7MFIx7JtieVw7nqgKgC+LrxFTNBoc0e91ITyjm4Ug6BnLf3qaUEPKFKsCUpL4KFa
TGFrJHoA3kz1qmehxNp3eTMzaBizdDtVKJATj767YTPtBt5UVMkcPVdiKO0IM2Ce
1B/75ecMo0Sn/2D0jw21KnEpiZhglxA6lXGzJuqzhtXSee6KZJXuel+30o/KY13v
nnnTCJGPV/VE74TBAv8EqAYqzyJCkIoAJ0cC1bqmSHktbiceAikGawBGkw5uflMd
cu16B/GC93Xre6DlNdkPiVLGb6f2D0YscnWYD8f88sT3rTXH6EisZprXfOKb4VsE
X2HOpMUXDLdV3JKMsjJRURBtaUsWY06IlJ5dd2Cq1cr8SfKQjzMozQnFZH00hS03
d1W+Qjet6fxX61TjQ6MZBZYzMHC67Gij3eqCgeFPmh0vSm9L8HDJ9WquaS5tPwqJ
2wowuGM7z3ahDwgnx67yyVsUMSRDb3lPpXLmVnWJ1IounjMdGEYioTx+T7TICHIR
qJR91BRdxHl5ztVoFuAk5HartMbDNpj/ptt5r+iX6kgYO2RoA5YeBzfNPOwduJ5h
QoAU7WEyGYM0HkozB6gJQkfp1Qus55wWk0uSTOPNayoCwjs9cI/SQlsojCsow0jx
fmULSxWUUPhycYnobnrwQlvz1+F2FMsHBP2c704BL0gIbmZJ486elkVPVAEPOEZx
XZI92Yy7hUd+MJIJ4vCVJHMXz09AOAXRhY57kNIFt8aqceTErFgeuTeCmHEt8abJ
NQrmFIi2LbGilDCiYYCpGRWCDc1uE73xHt8exIb2gT6KDmaj482qdgMQ93oPAPS6
5EPIQjkF8mQeQOwZ27gtlx1rpB5DwzeVHfeVlheJBQlmIJ094YpgQnjNtXtD+geG
cG7P7Seo8X+AYiDTzLvC3PbGvuKKpaIdiFmQkAjZjqcCiow5odoKVNt0rIJnTOh8
3y0Euv2ay3Vrwd9u/6mIEXnVcW3HGCsDfMvU9U1Xal5WB6nmUbZUpMcT4gwLQxUH
Pf55egWP8Yf1er+w9tjpWwTEbjKHBhCohMaOACXGx2Ziq87jisMV9aUACU1xQ5xV
iaRBwpU5t7pXMU5+iE5MZFYeJRTkDqg5+zDK2yP2qIp0H1j72CYkZ0Xtk2U9azfT
lwKjlerLO9r/hbtfttU9yPHQzegarudBivzUGBiA4sVH02kl1k/UffwedC6GqgIO
IVnJdsRrM157E7968HUgqSA0GkVj0tpJav1/0xBgjs+z6bhIlpqqZu72WM4R32DR
BsRGTnwacZW7gHCNzmobDMAN477MyMCfkvGo8B3BECOoel3774mMvFm50StjQ0sa
RfK4JdGtc1b88ZDJf/+b99j3vmzgB64pCDmDEpNB7owmFbPg7RvX1e6GpYTdtezC
DW294C/s0pcjQLtfCW4C8fPWu41TldS7KOzI8sK1CpOFTCJyMDMoE7lc6tg5keF9
8RxV4nRl1WR9bvlcQX50bTAdNPn56g9o0OYa8myDHOkGNrwcL7b4y5PxX8Pc4NLb
h+ogi3PQ2TFuFaSIwsKDpg==
`protect END_PROTECTED