-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
io7+X0AjIydcwOmPh0Tkkdn8yFrjTq9dHGHyMt/Us1nenDyMLhlm1y9B7hBS6l4yT2LmMPYThrJw
BjiFPhIlsa4QvGodx+gS3FEFUcjwhQyAQWP6V8JI+eWUfzH8ooEFE4nDtAoDPHbFMGbJVOrT0ZB3
doriAkXMt8HB7XeT+3q3fCbLC1KyDqY44adqmgznFJty9bs+xZ1PzGNBRjAnMHvHEiUoJflbTvfU
WOFXHJCXae33vJReIn5V002MLfftuZ0KzKbW9wvihrdaSTIIiDzLb2wEUAdiiHCSyX3V04/+WCye
GABWKfvA3MSE+YfuvZiVoWEaScowfIx202u+gA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 23392)
`protect data_block
PZMeBkrdCnt4icc6YJAflZuxa9dywfNjCrjJdpPRPrjlE5oH7LkEK0DhM3/12ytCsS2ejtzdaS0Y
fJ82jpfGtaaq6P7QTTuWkaDZnSnnb/VBv7Aenfx8GgUJC9oW3x1wuKzIF4VQ7x/1EWHkkdvZfYhM
yJNM6tkSwtZuIMjwQQn7l8mCmq3WqD8sgjxRvM+zacf6pFQKEw6EZTcXjqAfZf2O/bbEl50m50wV
ggrW8G/xX8E8FUCR6czu0eshp/I6zUkA33P8ASG1sRI8gelZW4sVUTP40mExuArSaFAL0soLtGAT
lHHxwnzijDn9RfIBRCt4HPnVAKXwwvZmp6CSPlH71GDFgU763kCJvDzt3M3b4FsKA3uWZBYdF9XC
8PQnnwlJXQ6ZcNrXjymZOwdymv0VvFEEZR4TJ32nPq3HFvdkvZq8pGuFOUQl2HIEublNVQSrMqQv
DVbSBKjk3tNHC6KPLrom6KAJ+wvp+rxnZGNrhyQVXDCPnfyhC8UoTf96/ptvpOyPIZPvAc82YsrO
uStu3s9w2zWCeaXBcyl3o68Xnm0wDhaY7IpLMCBeGtLSeGBmF4ARETXaqzg597Y7IVWaM5n9WR5K
1pO4coE0C1Dfm1Fc/oa8tVJFQVZaxPKaFs/aG/u1j/3ti4BAk3Zxd9U/yfpyS+hJr/+cQh5oQ+s3
TbUGBP77zXQecam/eiks2Vx6VXb70rALO/fOaOe95PupmIGp/eEN6lp4oIM0RBuaduiTGpTPOWhQ
AQsX35DHo3gCya7xiVZSsizERMd4LWijtkbZgq2k5BhKcTWbdllUe8D2m1xwJ/uoG/0Ph/WlK6nw
5/oZToteAX+dgrgRiCVzUypWXEQO5OvIrw+Z5iHcy3Ra8g91WBJ24wHXJOElEv9elraDbcKWKchD
YwH90FUkSBQ50T/isma+mWD1coecuqESeaZlCI+UB3Jf25xUSI9It962NEnb31aTkaqJYuqTAnHi
zvW4ymhT659ONNFQBAXLmMN6nIlcS72kPSzHe2vM72MNytzq4wp539kVco2L6Tf9dAw58KC0nypP
zSlrg2MfqSDr6a3pYrytthu1exXZXbz9r2E3cy9Qq4OzLr4aPTXYxzvgM9RxMN+Q6K3Jjm1HQbdU
zhxWO5bB1j/oPL16syCFHoUK4iY4VmSdrpcPEmum891y1vhME3BgZy7UHnt0mNGYvUbM7D9wnUMJ
eKc16OLVHm3ohwpnBoIuIUqIZPs4KICw+hCKcVmPPm6zuj5Lm7gPFw7scgsYB74FqSHw6nsAdOLL
D9rSd4zP+owv4ZVVI/tKO/qWQHm7beD4yWHoe6OQ161Dg0mhuW5rxQObFe/zZqrZ6PDJHHw9qoCw
eTu3t8H0GgcHlSeWYpT4ftBrbtYC+PmyWD6bCdsfjZf+87U+t5ZublOOaCnglCuzQIfKOYdNxYEj
LoWbrlNIiAZ2wW02NOkyZuEREIDBcwBR5SDPC8fFdA64UoOdXk/vtYTyusO1S+5Pb7q5Ut9XOcpV
Fq+MQICTbTu1fGwCPfkZcPWOLSiXfctIQ2Tgia0/lFZTs4a414LZwHuLd70kFRFm7CA3KWlBvrb9
/mbbp+GPO5kUMzMJ+Sa5qCIzEzIHXzRmdtCM2mS+UpcW8sryffWAK0XjlcWFlXw0uCZjgSX6dsW8
TSxI5TKNEB3x2tk2ep6jXGeHNelUjy9ZfPee6JHfNeV/JzlS1y7f/NKdbSLx1AWedTUx2a7SyXY/
K+r/3MR3PNRwVRMixbkmVYaKlUf+d4wgyOF3mgUxz4arKstd0JtxP+iBBFdmMdhPZYIewtuz67GT
6VKLraEkzdERBu3Qb1FQg3RIhekFCUeu2N5fqQ61PgQiJbtw6QwOy3v2ZET2eGJEOwfpgTQ7+UNL
bkyYeoPN52NfF/rxK6pVA/AZC5fMfQ+vKCHHkZ5b1OPGR3Q5aOMFyjrPjp0kjYc4Vv2OpuA8TKd7
OWXTseR4WYerTsckgaWjVH5WGXDjeP8II66drE8kQ/lKe8c/kqQjIkFl1YZLY6/nu5T6A4XHswsB
klwQbNKA1F7T/yOuyKJqHdzqgQ2fqViTSp+ewovoiQpHUUr78PYO8jls4hQTRP5kDssiWR+zGDKf
z4YY6hW9v6H8ZkLNWtMsQTiL2+i48wU88Ywh2In9E3fe85Jpi2z61FpA49wrITiwLCI4UJ6nxsK3
9XJFhcXweuQW+GopgS7L3xPgWcWnKKdvG8Pnw9qXFOFJXKDd+72NAdgjjqhL1QMz2siRJes0W+BA
+TZ+igTZdPEFZkIhVN9czfXyArp1/SxXBqvM6qvBodFMu4HbbThpVUy9DKBkG6klsr7kZ4zGFQR4
99dih1XEyzlJhtScsIwKxdY2FHJLFB5Mkk7gd47cBsxj5ohlxZQW/Zy1LKsmYTTSmHbKGs0nfjHc
biiYEVogKgZct+tXR6VjSIT+zVZemM6UQXtkcgKIjs4v22ahArcuGkxgou0bz0ljDFymkZgqwBaL
W6+o37DtxnafQrlstWkVb9CxaBYewYRx4Wjo7O4jcQp2YL64n2lGz9XH+C1oxXcEkpwJJ4jZAEyE
oHGnDTZLBRdHgh5rJb/jAd8pRQsGSPDdHydHsI4rp8nYlOm+pU4RWRBPOYUjBOkCtv11yjvtJJyu
tvsgaogKfCOTmn3EmDmnN4nMwINDQ2j9zDN9RkDfY3gDrYOvShzBFP0IvWfZbxhxv3o4xvFdOTy0
glN7qlxZI27EvleOQ5DGBPy33d1u06USBHA0Lv491sBSfcls97cUgoLcWQ44Ou+5xLioC/ull+ef
Fg6Pbwe/0ow6kPVTZFGEb5SC3HGnU7bJ7YRph0NAPCRTkIEcubCDUrWMQad3WExvKo1VNy8lcuBB
nZ4wlTtmf/W/enrKYhwU0Md4hJmInhx6zE5iQ7vF+bwZBlXMUvK68WpBhH91owIQYnvv3E65GVlc
Vz3w+8VQ1/zajKWLWk/QNshXsyKjR+FRyhU1Z5MDKni2TtrcDwl1LwV2Pavg/XycJSb6kD+hEWAH
qOiu1tAZEpkAVGO1ym2MWoFtE5I2I//bzQYPG7gIVRqLj5j+KBD5skzTudBrbGofeDUDd6phpODJ
aZ/5QfC1UclMERnIEEt2qf88oZa3ZyeK0zj1A7rJ9K84S4EPmWDJJkwVnZHYm27Cdowxa0NLSc0h
PW7is0IRJV5eGj/pxNTRRUrqHLtIteVrNiCUn3RPa7G9O+9QIwTvY11J/3T+oZ+TLq224nzUtXbv
prEGI/n85kx2qT0CC37oZZl6ZbnqyWAQSrdoeAkEztUR4g9d9DwicuiJVczFzD7So6+iOnDegEkE
fAvjt3YhWQYxXckx29u3JuYK0+g5FFkxSEKkxC4eXh2AoMq+4QNr8RqjmiOXJdZHFJJz9HI09aKR
8jrbuRGgQuy9WsVD2CCLP8M1GY/0XYCPBmuhEB6wAkCi0aB0n9XX08cRHU7ra9DuzN644CHa4+7v
fE93gwsbV79gTltcLKmR+gsJGwbBhG/PE2gbSf5eJyYccDwss62BkUI/7kykUxurW20QtU0a7eeG
Jn0YiqV8ZnX1L/Wii923dHVQn0qS9oJ0w5SPavp6V6+6liNqm3SLG10uzA2mUCWXK+I64jBWj/B/
XbF+qng+8P7+roOnD5STF35OU22tNOJEHcJsdp+QB0tRRXsfGXoElNxj3yK7fZ2hJcnkYZ5tPkH3
v/Zql2VyhEDEcufuPcMdU9Vrz8Mwo5h/wZAjMMWMKBeQUXPLblZWBwBoxgI0X+ESWBEqRpDkYc2y
6TPv8jnmagESKznM1loGZsKYMmAkjJwzvT+XTGQ4wR+a63/qOgpx4H6xbe5mVIibuGyCQ4cW8vqN
3nynKhBcKPuJCMyluntHhhRSRwroUBxretoTw18RTAdYTGkMax4bdMVHZz0XOApcNUd35oPy5fNb
G6wj7M0Pyz84vVS2Y2+w/JzSh+v8IyrI2QnpTF3wVEFZhd6ERtRkZ2ORyMwg8XeZqEfWGfkr798I
nfgkfKBx/wynHiWivURwrx8pqwlYC5eGP856rbPT+zeZpc1XszFnfLa1a3dreXFjW4EtJDuudzBY
9KlTomNDrdMe9kkTn0hxviChjKOoLnOcCTG2uu6cyI04SSMvzzxrnD3LpCt9Z6L+vr6tG2YHhrNQ
CtLkcEymWL17xElrADB0csZsNhJkp4hN6oQ40bWtACpri79KGb2dsRB4NmcITqRwDpmKbAKKdSks
x4YJV9bP6J4HlZUQX6Pf/yd74P/iuFDfZIVXzFF9Mx3+YWu3ViiHv4mefh5CBlsen3NldxMM/cTh
vEWSMIsZu62I7cSkJahxBnIS1oAK/AuTo6BPomM1bNX5AIt7DYr6DxFHCgbxMfNm3IYGxytgjyAE
KWVhXF5+HX1zwafZRtYtrMvHJGaAEO39MjKJtCcyaYFIG1GkOO+vFW864PNyhzc8DeGudsxRBKib
79Bc6Wt5+ZBnghzdLcBlGgxjpW182ZCF70QTQ3i6sYXLrPcpzpV+CMlls7TxPa9V6TmJYAu3hsQz
qrlxgy04ezfr5y1yzHa0w7B//Z2K41BK+idhKaML5m93X2Nb0M+S8k0rpJnxThRV6vn7pv9H93uo
CVLtHKJ9hrzC0HIA1AtvkWlLbnztl5fss6OK6qwgeKbaUDIG2sUWA0dRiNBrcj/zfyBl3reOkmEA
CQiLs4Ge3A4U/KQMK/bDUXLb/YB0YmdOYcL4Cwuc+imlRxkuBr6ce/Y0nBzaOGWbQi4p+hxlyHiJ
3XJOC+qXt5n04zixIz+m0VLkUvujviJLa331ZA5DPNSgJDruJA573gCVyfWqOajLSYAVzkTqvTFr
hWK5YUWXUlwAsr+d4htsBC0AsSDpVUgyVE46LDN6G7Siu8RyOm0gjsKcjocikoch/z4tIGJulHSt
1UCGbktY7U/2LTCzfmG/vK6YKmEkGqlQrMol72DpeokfuCTws7LSOf3VFYj9VxsmkUEY/vCegNMd
oyrTDWyHfcX4uFpqAfq7yW3BZxiVH7OIwN0bQ0FuGtdkQxxvleIAwXkWlSrosf6yo0J8t67uV6vS
/X/7QFZQwy9al47XOyiZQi0gGZWWV5ai3MjVcGwcDcITwurVF9+1iYuGYmQBuWg2Q4N7ivzxpsUe
wai2sVjfu77L3ewyXBcZE1VzaIrrCpk1wev1y3FDq7bXGdONylcBtDP5ktlgbEFLmzIF+bHZpUEi
NlOsJW9NAc6lJNZD+4TT75eOTAXqygMfGoWqLn+gCZFWvD0d5CHe0sqEU0SwE5icC+jo3hnDey8/
yiyAntqlIvgAML7L2BO9zonyK5B5aw9+dE3rHUJtcE8gFyj99vOowPtMPyxuJoV0d9bDf97WxwBx
F0KsP+0U3QSbNwGQGwpkkNMFzA7wadhgQnfuwZbfkJgFOuCTf43bHHIQUMvPeRU5d3R4dbDqM3nY
xAELodqcHUbTwHTkVPUqjyT2ZPXGBwqFuLiqEX4fV+x1KKtTEcwI979+R8kE4UiVjycNy249lfuh
dmoWl6MoIjnJ/EcHylP5jmesPVCTICTV0x5bqydC3ed4Yk3gpOkpSPRQr9NC6Q4iWGfFDc/TqEFB
aAPD5BAEAhQj7C1Jw/MYQZTrn/AfeZeBvZytIE68j+fGrF9WIp4TMvKpLSjW0Sp5tJ2MGbnc6mzQ
84fnyicpKaZOFDw+6o48zr3+DBLifBuwtG2mIRmqKXn3/NCo0NKzN59rFkFs60/MQ9DAG88pbsPl
GWFae+iKIfG5BwFnJOCP1zpnQvNl4fIAT5ztl3SVSKLPk6xj3OI3TLnaBBmvZ9pTQenpB/6wWaTX
JLLeIKebMk88V5cCRuhwoZrkfY26aNL+p6S1K/xnX+Qzo0pEiH5+ZeVMSUkeMBHLPKQohn+CVws9
hyA5gE/k/3SmZ1YMD6wVMjWMalqoTs2ZUGnEy+Q5EWPyHyCl6s8T3SYCK8SmrX5PzmvLgTL0EzY2
FDK1mVrONpR2Kogetth256k5Jy4/TYKdbGkl6CxRRy0rWvQlN7U6i2TNMA3AE/aVWpI/X/etw1Vv
ChuQh+Xb6ir8Jav1JNmhLhc3cfKQfTfy36CFsMBYc6R6c8yx+sFOzblpv+rEpd2JC9I0phURXrJa
gyOVvbdgcsnec7fawe8p0ksr9VWLo65SjoFWyC0jteLJWZzFIZZ8q9qOdHYDnMSynskvlwOgPQUH
iAJYjcGumMpPEik4YmEB6E+ULT2+9WFyGgZREdn9pfaomYNv3E8LnycUBJW95zccV32m7EDzDou6
ZbDBQAaFFDMnmuzFEeIJWVzVdOxsqennH+3sF3ixZO3ldCQKtSrycbrOYRQwAWxOvUBfMtcB11CT
LBg4sEPqg/8N30H6mqm37UY4QR9+fwn1HgucrbxX7IdICvpxRpzp8Av/Ux3LW1yteWbBi1NnTEmq
QKW90mQP9lshzFXDlXD6IU9ZObDGHyQG4aWUAhlKbmKdTxtE1Wey1Gl1pMPbGAgNx3qVTq6UjWUB
d5JVQExswa/6c68ehWKBDg+HR8BMEfYt+ldaGs+jhTEvR1ykk9hapihK/xY7np+GDmjZzgA+Or39
il5bfTo9MVq0tBCeKAfT13lDDJBlMagXqmivnYi8UdDQhHJB/0KMY4+ZnPRfriT/2MdhEhauqMeW
O7L4V/LURs2v305ykH0NKjcMglRLvKhykioLTtZEiOwJMkzvptKNz6VNP1jQ9Na2fbyLotUEF8VH
m0Fv7jjVw6qVRZkvmSBl0ZiNDfXNhc2JPN/ftfdP+Z0mRHeU26+IQcC+MMFIFspFJ62pqZm0OVcH
BdhfdII35C4sfQRZBa8/lDI5nFdBJLrHPOttNQNGcj5fgnIq6qrhTNBaJJ2eaUBG77nqN34XImEe
7aslkdVijT4f2zM1ipKGroIqwdqcL54Vqqd7AOXlwpHS++fu9kpGTAlhYPskl6goqFKp0JAlRX5Z
h0DLfmBJBfnkoR9V68zI4SvGhOswWg2DiPFiCoOxdwQn2vrKZ9dQ/NMFT8fDFYlf72YM1HsgWOJU
YbN1VwTsA5Y+GGyDVoKLCqOP2BMQN0+IDLQyeNmAwNJGRhT5PzLv+u8jt9CIGOe+Mo6bjvzP2ZlG
NzdO6a7dsPdKAA4rHdENMcMB2ESC0EloBuTH389lJv35Ki+NyaJu+yb7glUQ5D6IcP8ffLhVFTVA
5W674YWaj8rDSbocAibfgiBrLGtl6In82moy9JMe/TVa3VZcGxRBHHIVk5Kv/hLPyp+1Huu04Dws
NbbN2IRnAHUocgztkV+Txk6YHAMq+imqL19S2vCKquSL9VgSyilmQYk6pDeVFq8V7NoAWZGGKV9N
oh1T4P3vYTDVjo7yRQ3K0whpQGtQaRyXRD5jwfm8/TbcQcaRANm0hg5HKLB9+1BtFFtFkORghzvP
M5/fon53uO//x8iD8w1FOHaLnhZVwPnHWUyN8k4uffOK9BxHkmhzCR0f5ZsViVIp9wb1afLYsKml
RQi9FEYLY2JcLcOJZpEjmXYb0e4OgNh3YKKInv2c4h5AlcGdeJ75AIVXnqyubWZKvjax0ktgqua3
X5cnujV7huQH2w13yc5/Xh2hI90wNHEZqix5myqQbdHrf2zlbBFtZG5K8DLAV76c1d9V2PYj5847
999tqF4JxuP6nkVOtncJMg2FuqeDHldMizEPVwh93noxFE3TeUXY4HmE0CLoPa0irkpC3tpZjzyu
UbLtoivxzGot85WvOnMxHrIeGx49aGFJfdnPjyh4W0eTnxuHzocRC2+JDG8OSr9W2V+5KXjJOv/R
JYijExrIyJWc1/4z/T7MJYESZnmMZiBZyLhvgPjqGpeo0k9oBcs9WrBKwfwylQ8Ff0WqXMX5km5T
fcsa2xnXUK13jc+OkEJuGhG+gLrF5ODmzpRfJ+Z4vz2+f/eGV+0pfTU2km71XjGK9t9iDKspLSNE
sBjvwIkhJeyFODjperxixydVNJBBI33VbyXM1Y97ncbi+siW0euSToYQx8dfJAqhIJGbFWL60Yl+
3Qp80IMN06ztU9yosNWXb3x184cy4MKB3kyZxnFJ3esStxoNZ9nJIPtmn+46SueMnIDH1YGBjKuT
cFPjuTjk5WICJTtKa2oD3YJjXhVt0KiBy9McrnRZnms00Nw5PJ4NS1CJNCDFg4tLTK1BXHCP1dOH
qBMsY+l57wH0vi1h1OCCSSYpEt3YYpDh0RJVjFEtq97yMFOXPMXa7JiRcbDgnUcDfbaPWEapowJn
t65esTLkYXXZLnRkO8VS/lro5h7oVyP7ewpwTaNv1xj5kfY4OyHgX5PFexwuxqqqD1dIYb06vfjk
QEeC/ga7Ys6TUrKldNZzkowWHAuEP0+RL5KFE3It3pNqXZvHr++nUvMjninz0/ngXsn/tH5Yocs+
LqfZAa150QOHzlk1+8MolMl1wg7pIe7vNC5zKk4Da9p27lYEq/JD8DU64S2dhqV7TCQ3ck/s+s50
h3Est4+SyzpcKG9po852xOQhOyUeqBReF1Mgg43se093tkH+KGHyFTJ8RXlYWSo9ZgWE1PH993kb
4DvUG4IqWiBR6aRjkUb4GWzDQGfSfkCueUQUKV27ajcx732BdNLxxqQwQBKKv2FIGAjr5htOvt0E
szmmlo96+0J1dKxVJ8LFnrKEAE/TdHw/3WVLZlK1OHJ74Dyf+OnVBAUWgYs+aCE5Z3y5uK4uBtft
XPHGVGpdhP+FRk9S2MsUdCVYVtKfdomNm9Ngqn03Uk6w9HM+CWB8RYROOTPLcvVsa3/Fx2n4fbaU
K1j2x9djfOIxJ41DdkSp9oHKeJqNoXgt7Ev4QFYMmfb2w+QLs41jNF0yu0/lPNyeYCozs+t4XgF5
zZkVCbspU6hdi/LQsx68pgNy8xGj9VT3+6DpMNIjv6bHIJl/0KFO6r3YyKGrTyEKGiu5jbtipVqT
hfteqkTUUszeGji23E5sIKuncQgXhl60WPf7PhWs3jbyktUphobaAoPP4H0EbXr9jF47D5iyRIDE
3LpBnKtESh6uOePQpG2ERZJPDwOyOg0CMS4MxRFkI+EPIP/cI3zCvbf19wTPCgIGszBGdQA4/Zqf
fqYbc0xvsGbAEXmv9EdiZgiAnydl7wXxjiQcn7O4qJi/i1gWI3HmsuNO6SvFVzU/OBvRd9g4i501
p9krryNrkQjol1fqHeH1BUFsIZTJjYuzaFhLcCI8B75y+mdXRC00cNn0iTJJVwc/lNCkADsqnb30
YSUM2iH9YYJ88Haf44AAgL8BXkZD0bOn72mC20I1atkj7yqp11TW8GqvMiTD9Dl/+Adzo4/3Rauo
qRFh0qSMELCnJGfSurw4QcmvpkYKLTrPCwkDN81mtByq10oRN7gaKzQp1hDWCxas/6eFiKj5XagE
KRVp0VM7pPgZHU9hCKXltVV0Q9Cbuk8wm7lonNLvfnRsttD+YJKPB/5kd38ziwMt+GGwSiMmgMXl
znRNky8WMzYXadMV6uSE2sGLRjNSxxfSzwWpXtHTnZkJjjm+LFO7VlkRFxmzCxDL8LqrGyVLKBKQ
AAf+H2Z1bSWG3+8nnUHjDw5TMSzIqh55Ajl2cLTdOSONcbtWupRhvqp8IZB4QpuDx8595AYxKKnW
7oeaOCq6GQqFvp9ukLpeABf41eNMP9gtk0NlMt/uqDjKO+h+JPOna8eytAYdiuW3Ap5bMgj9Cfos
R/REuSKdDkMYcekliW2V3NClFdggiikbIztBc1Tufe5xjdizPars8K/V2TenBLW8LT6T9+xaJ70H
YDKcDVe7q8R8yNMoci5COfq+Bdb8Gt/FLC8t6zz20Pe/oNtKHb/KkamnqaiZvYvJajCfc7KTikbc
qIpNG/I4CRaGu2tT3yKByfvsmdtY+Cah9o3mQGBU9JGqIw7aSBLO02Ts37WvD2CmhX1m2usAJN9y
xC6XNO7Q2NMRftA75Mm0Mp8CEjEU8Ox7ugRnyBUWQj536zMRElZvCry1OxEBt+Kq5ddoww8r/bwK
E5xsZNeF5tOrpMBN5H3FdQaVkyxsWoCxy0pkJC24baSCjk8ZIOksye19/4D7aESr+FTQOCxWgT8G
nEihTDBm47NnfSC0dvtsI6h3dh0Hx95xn2x1UOGZcMr4hZhlh4M8AApy/H9EKdFTTAxosgPGVI0/
Tpov9UJHtPRe3cN+UgSZhph7AIL1ETBSDgPwy/eIJmTaXas14fDW2Gy5mPErkSMixDtcGIcnUzQE
2DxEJqCG+MvSsdw4J/zKov/fFhdBJA7BXzeLMMlfAjtHeJHOTRHq9+M8Iu1HO0jN0YAutask+Dmo
nbKic08996aXhHk+Y103OVn2kDQvZgem5N7+l6BQQSIyC5j/M8RLka/TWKnpQh785l6vZiwmlaFS
9G9kdQgesYPOSy7RygXd5O5hWmYxLVx/eaVOxlOs9wqU0Mf355VRaF7mwpcO1S9JXLZl6kAgZ7MH
7zmuurRKyeuKdI5an02q6f1ed0241q1FDy99Sp+7crM38vUjnBfIZgpdgbyNwCuqPX2eDosQ4DeF
YAQj4n3OGY6JbjJjzS+jSm8c93ArG4hQFDMrLWtPKxlJDMSgCmKHPn/86w1GQA6De2El6PgkiRLR
A8iKwlj6OU/rY/EnWHTwhNAZK2VvhjfaksS0CZHdOoqN5d6bxs40WMYywrP94Cfhg/2p3PJ/eftF
DVX5D1Li8dxYAKAMq6U3OVv6Uxe0GMYDSboyEVinvn+So1GMNVIGLaa2eP5T2MwZ8AE7NbMwcEU+
h2aCdCIdJhm8ma0BWcr+hJpMoGkIIcAYI2L35AXcWcn2GT3oeGQhHC4w3nZx79NIeIVbQ/wA/7yA
ky1eeGy8JYgYSWkMed7RmFP16skg8HlIm34f+0GaEctdDUB/ko2XxeCBdNhIqXCtsciSOoiyMjjA
msPEJeLKhfB/NPhd+bNwUggRYYDQL7SeqN04QmMh3KPVBfWTywDoXImmMF+rNFzuQvKwAwiMM8Cw
b+eld2HH4zcZhF8Cq2+AcWx4Jkowrf3GlYfqZBftbP3pfD4xyo0GtXUHx9ZdXn8aksNRc1p9QY29
I1IPYueW5hNEci8g/UEBAbaLRsGcu/cHxGX/WN8rqsgT0Iab502EFWDo29/X52fnQV+rxNPBYX5/
uiZRZixyWL+NsnSNMbTQ6vJ3ojqL1SLl00B5AXUftfRhSOXyQhyZQdZeuwRVjAn0SYlMQ3KDJE3B
B9pozpigPjSKPkotIgLLSp4prV2hA2VQk2Omaemd3a6DG+3jWXV84l8pgLhXrUXV4C+zx2ceu2H7
KcAKB1cVIexJmiGkgK/HZLyfBifJRlGTeCzkOAEkVZ7vFL8p5MVlh6BqxvJv/TBeW478TuvSKl4R
pGAqy6tcfA5oHcGfRp6IEHuyaQ/xKlHR3aPsmZY4dDHzN6tHsztel4MOToY0D4P3qfLWupnzV6Ki
FSscdrzIT5ezQ76UlQofhNSCceMvnCCb8xZEQpXfI/UuFGif+Dfknu3leAfPrt56gagqWgRmeWpb
eDlXSOFptYRJvrpKHs2ZDudZy6fxmERhBtYVyeggLjluGJzONvlidiVIlRcDaTDV2DozOa19XbqJ
xJjkwUgPUlh7zSPHNZ/Yj3IcaQo8nIX9gUo3yKzNEDtZxvqEedPS4c8vAf6X2fi7tG6U37eeY6pZ
XNuDZCZ9l8hRWWopX02vPxt6ulrhS2R9UjZc+cQ6WUlRXqHo2Oxx3Hq8s7rKtgHTGh93khaSfVw5
2+yv7zSOllDz/BasvfIb2XmYcAS6kVHKDMFQFNCaZd9hbaMZb4zZ2VJgDq4HV6wh+FPnmCW72DUS
XgDq9356qnFEwMz0sjeRvbaurTEllpt5AtBVHXGdQaMW0/k8VIEUeNZJbywqH6HSg6vL2PvGn4mI
ZXXh662Hv/6fmHviDnmczjo2nEqthHtPZUKBeLxSZ+t/vBlvZ3AlAQLf/l30H3tO53qnnblIN7ah
mgZ4z+WJG22pGjNx3MMB5ZDyKUdrJtp24AQOz+cYzs3G/YY3dWSh5Ri9B8aiCbKzB/chkPQcSlyP
j/57t3FFTHB1+U4In8SjDzixpz3nfsCca0l1HV50HNyS6UBinSP0dAXM9kTfssE+7ALAjOZ2d7So
3TfK9xNVsSjcm9NhGtfGX0XNFkWDwcSWRuD82wa4BRoat6/ySvJ5moEFWA/L0KIPXXLjzxrlm6vB
kqYdFnpXHzuDhkpOhmjRhb81e+wxsaqZeC7UwK6Cay3ejHbNol/npPcElV9Q4LI9QhHLhI6KDK85
oILcCvKDb/K6LOnQu3j/ZCFs0wSAHeFZnz43/ccOnDz+NrR2JVkzk5ojxArWJ9s+6UkUD97VYekN
cQGnbP1b3CTplnx1puQn9w2wsstjTQiyBv7nIlFGF22aiCgt+6GmmS3aCTJuC/Z4GylJe/Rzl6SE
6BxM9qaRPhJxYYYjemm7wUMV7mWSytu6sHYU0/z7FmzXY/TFadtd80nAGw5D50953FSz91CPnyzL
ARGX888naJ1DEJTtJwDMw+gOanpg0aVc6SAKU1nfWNDBshf1+wGxEhN44XcG7LQ5d0kTpXlm6XOe
2IrJqxKZbdywiXylA+0usU77UX+xLSIBYnlfL0k5W6tGiIHroDBzC2bg+yryhWdx8kzEnXMPvnqP
rhBdw83z2OHNq5wOT11n94t9utwFzZuGxbzm6b00QtcYLpqlBpUGETDpYjjaxjS0waNQFYorguvb
6S8dbHlUc7fefsdiQN2iq5ALRpj+CQV3Y4OiXLYUh67rAGG9xk/7x9qzyIwfgQYLgmoKa7mua+jO
wt/3qMRSIfEelQrC4WtjueOITOUHSsOW38+/V6MIqlDc8UjW2p3hlO5axpA8qbw9tKRlc7mvHER8
8+7+QfJV0ya7178lL+rj2Me8nKTLihZs/trb31hlGXTjruf361I29rn1dq6l4drt6X1Rb2y/GgjE
CMfOFVVUiTQuYeO+qyHreBRsYBfk3gsM9/DpcB0MPkwP6IM0wnpMP1mTIiyaq1bUbQAflR8z/djp
/b1oLmw/ELZV4XXu5ZKcvdAFxJypatRPHetfX5qeTplksRfhLKVWkaU8O4ftavAAl4UOquRtqiKh
ArBwqpxlrULo+kfjo7Dmyz1EMXuibgwkYAba5jjFhwcRSIzdGe7EZShmxJ2YbLsj05zOMaZgOd4N
cB4KbPLjjFf7Ys2nYHZk63mIqW4qbJD8mhzFMyYuvNFVdTU8vPPTJ3yNZPG5x0KDL8VByu9Pb72S
3HmzZNsoEJ/8JTQ65VnTfm73SsijYF5xcbJ15K/ZYUhYhuuedzshMnkkll+o5iYQma3hjVenAqnD
PG4VNgDD64DPt0/7jDIimNDrFeBdxfEOdwEbWfi7IX2mufQEzPQbDb1EZC8Nwt1uins+CL4RsJLM
8FHYXkXK7BZaGR62XaBdar+fvekDhcosgIB6G7FmRk4p+ruFqizYpsuRiz8NjolQohubeXKIlIb2
b/IIocmCsB/EZsh6ujcj9aIiyfn/ZcXFQm/9KHgCyfbyah0at+S5C1blZPiqR7V7yK3obea7do/d
Wa4vS1j53PguAih0GeLc/jrhlNMCsovLARLB8uicZZmLKE7/y19dODRqiY/5jTdIeCjvNKVVUzpW
Wksg8OIOp2fsqZj62JDEHgWFMdtXnJ7F3hechDQoMvix81xRrl5PTiSnt+tWHTmT8vZLfxoxdCGm
7HMktpukRdh2SC2yr7aME3aYDrYNLN1kWyr4Vg3EIM0OMtR0ENujhz2hKHwsW4oiuLCF2xEvWieR
jCx9CB6Zn6vW0YijeAKry2E52rBa0jKRYwVBJrShVXoKahuy0QM39HlBD79+bTuJU+BvEwEYCvlb
+MkSrLvq0WHTqzUeow99+jrGzmvIiDerJbu/RlL1No6Kdt2MuXZQPrIDHJv4bZrXYbcc61Q59IWi
+qgN+3f9c1BznqSJWq05Pg+fge1kMpc1HzQRXhJvsaCsBZvvmlLUNu/2AAMkAHZeg8FuVh+ziVb9
1NbDpEfwlTigW3sXwzSVMlnCCxO8+90R/pWzvmgxLUfk1+ot784A/FWObH3Xn6a8KaiYnXPJ//vN
9xMMCt/sWoiBbSRvWFbgg1DwSGnyqh+DcrJXZ8lwwoXotYFpALIHhkNvr++BQCjuQKS1f9+P/hvH
7oYDJXoDxyUJEMQkPfd4QGNW98mEcUN8/mLVIATY/NX7TITDCcdsUqbRY+5hbHhGqS+nEL2IPkZr
Ii21oETaJD07f15h5/z1nCBZlCdPajOTl6yjshHrKF0VVjxjHL4IQANfS7Se/B05W9tiEjMAxjr2
6pDpWUiqhh/uwhniZTUuJOGnxE7nh9ThTV3ngD90tMNpcMfwsHEOB27bkMqsbgbTj+CAqK20QvEB
tC/It1PzI5e2Whd3uLoTVZFszO6coZI1jP104rpZct3n02KKhpTsVBx48+Duffi42PFPQ34rcCph
nHJYeukDzRbQKYPnOrs+RLcR6nFj0zGRVSVFo+lOiTHNNvmc+/mlrUBBZKt9O8P/9TELxFjAgUL7
RZhRYdarcsORhV/R64uzcAia+PXEc0Us70JGlula/U6AuIeNXfpZGHOHcx7R47XChCSi1qy6bjva
24XeoyZwBYjt1gFAa0SA1d8r+ROmu4NuaFYVJGaUidgWWpl08N2ybzraSW3RMGiHmSpJjjMpN259
f0pX5cGwkGDf+sRY2CLyu/GkNRgKecdYOqwPmebzWFligJbs35X1e0OCyZZKp4XVYhdPwTMCknf2
VaUqc8uUzBlVN5sd1v5hLNuQkmv6UrRoKEsIMI7usc495YsVPNTCgllETeGKykaUz6abpfRzfnb4
uPNBYNHb9zq6WXmDpBJMOf3ErbTdt+fgrw7RoB4E5as+thkNP5kMp/alCOrYH3tJETFmuKpoUKKa
O3/ty9liZMXyB4MjSDVPqnUcxrtN8jgpq9eFjG6oyvE4eE7Ii3X2TyPxlK/FyvxwtWn1whpjEwvh
zPwQqyDtII7lIIq4htklInPM5hc2DUN7wYQ4znLaLPLEmxLWBW85dtq/geMJhP0rBNTOJAVsUb0G
o6fJuSaYaYDf1i8XS7p4yyAYsUDiHQeu3gcKHz0Iu7eooPM1jOgHcRA1wdjZ1aSj3Z/cNMA0sQaQ
Y6PcJpJDU5RXAoli8xTmBKulaMlzsa6/rdRduY7eG8KGjxtgmGdPnisryiCcT8TalDVqh8p15Uy1
RcFz6jSqqH3qFYRdyWzmXxL4hOrq+8Kg+Af+Tc7JVjDRDTLIgoRdb87xFMSQne7J/52qJyG4FM8N
9yIFErky/8ExJzHpHgzkZbUI02d+n+TCbsWQSnhTgVzFhBcLaXIhwK5Gn8s5YqWc423Ue1e0jDGo
mswbLYTi6IytyBV9+xMgmTq51bE8dbDg9wHcphojOmCl+h32EO6+cvnSTCO4j5t/BXHn9jW7kyUI
p/bxkiJrMtJCnOVe3j2zaeObtJujVYtajez8yGTBqiozxk9J+8ogieQMc6sQLBHxAUHzQkzwNX2b
11D+FOiPBX3DfccSQfggP1bHTSTWrlg4ao8Lviw9XZNl21RALZzGejOGYlHq7qj9qK39w5jPq1eI
VNYYODn91HuwP7I39KJL8DN7NaA3ktv80F9O3EKxRrV2Eb7VsEoFpoK7SwT+F9RRs5YqH2m00s39
1U/zUy55EkrmLku3m3AnVLnvRbSobhft0MctJsfEEAA5UOinhx0p5B8aHdaq3X36M6RE+wBcDpFi
PR1Ys92OOvCxnX/WeeKjxRvmprkNucGxBNuPe1s1iqxpPPx/SV/kBM/KBkekmYQ8uss7Ie4MA7Hl
qtP3Xf4HGbMlRoNWNmQrWEDJFHaeBUJLkSddcpIn1h53mY4Qnmr72wvpP9sg2y81KUBv9vIbXxTH
HJjmI98Ckgq4V3stVWzhzdug8TURGPl8geggnpoCaF5XzZp44Bw3BNz0oz6ohYRmwrKzP308TjJt
trqDhEAAtOq/mKzOJ9jcdjK5GIObvprQfFUSqcbuDPdw2TCUZVShkHc/vSdMKSqLwmJMu+7zEkel
+H1MavugS905wjzncQliAr8hM3b29rfQxXvhMlkx0Vz1CiZm1ybCe/fn8KNhFIUBJliKJ6+Dz8GG
UET56c8A4A6JezQOO+uel+cNfmnwsk/KeDWxjs7bRklyV7d2b+imjErbFqYIdHBFeMZK84udH2Zk
U3RajIgxnqxkIbSiOvs0CZuI51aQOVTRWvEKWoYvBKPK4BfxNja48qug5gnvkFNsavmt+we6jR1q
NSr3PbxLfTX6LqUD7bqlgURtJ9BAOpm5+q1Gca9V+Gxqwtiq3giIbQlaCxy5opvXM+7NBDQIiQkW
TB2pS1HfksRlsaIqJb4UIMtpNmSt8+yeZ0oExE8Per311sqPRYX7znq0nKIQypzpYbauughelngW
7xNEd0AoZzJLjp48cSjk297Q5ERmTVmzTItdIr6wtVpPJNyM54SCRUx4jGoz+lRq8rJxmSGrmAK/
+B+VFQTcE8NDks0XN4T+UH8y60jqcTU8e00d1dNIOpfuawyv9evNQj1UphCcsW/aLcc6GnRkotg6
kjCHBkj3E4mmC4U33AbcsFD6+8hs+DPx1VqWnHTWFNTpSEYkg3raYHyGEylIAy+TZDkj2Df4UGwP
PbPmSD8oS1VRrcMrsJz1Riy+u1YkcsUZnoaq0moTGv7keyMafLWxaJ0YZBrrjmx1wrNwVmb9OZGj
lcdMexO23GelrJz2jtQHn9b9RbYjim6NAybAye0y3IfzuRA+0JNXXQMgyLMisi49AHqCZVGcvB7j
xwKYI78ibfcjFAqJhpImebcN8+p4PhaelNjMx3JR81E2rUWgS1nQs0MG9GCJjYP6PKHO2UynEeE1
AHtgH5QTLronP7RC87QXt03Nv0Wrl7KAPj4Q/EMIzzvXUZHQqfDVBdqYBvKCzM8KRJhTql2I/59y
8hDWkW22vAnOOYief22AAS7+ApEUXDuZGYbcCYP+Hl06ZQM2nn0MUglrr3fJR9JcdlUiMRYm1fYG
Yi0E3rQy0kOyTySUnzRlfJ5XHJkH2noFILSOQaOhFOl9EdVAqkDSu+Q8TrtGd0TKqH4st/lERKZ5
jdUR9g7Ekb5J13pTD1BP1/UemsItomqpoLj99kUkejgPSa6+FpH0MIvPmHn8oWLC2iKTWVrztayL
ki2pOqXmfGFqL8W/9cn2z13nAtQmdW94W+9p5SIizncmwaNpmEirpQE1jrr4IsFUTOqXr1zgFE2h
gYGUt9ba+99UPxLbo4f9vUjhitG2wQS3tD6H1D38auQcgIcJVFleY/AMriC124L+hYLVtQ4oYkys
kYhU3nD1qgOe5XM3vBxDV11hyG5zKIYKrzZZp2Y1CqL5dxQ+I3a0c8ET5O2YoGZSvi0EFN44qfw+
Enyspkh2ukazWmN5rwc8rX7XsRXhOIeq7rNwvXqg7U5wgjeLynjme2psLlknir+YVmsC5SqMHBeZ
myU6MNMQjdk3jER/+6NK9fIPJglAVW+lZJtCsyYwiiL5TQQlqj91lLT2AWnc1MHy1QZkdPMDYQ5X
hJMsEDg4Z4lT0VHkmvpZxOKYeySZBwfYXzxHQQNYTrdgybuSzky6qdoRZ4FR8dGGChxERdJttIQF
GtoDQlpyBrDo43M2SSC5Ct4TFph+L4+11xBRbRSVXE2+YLSmC9KFZ34QMRlmhHzyF9sHPY8dLPmb
1sddUitbVKTacU3bStHAV4DUTnRsJochBafdEg3z1UAPUePP9DHgqAv8I2K3zNdrR36g/lcDqZ9z
emtWvkoBj2wMMF63+G70VN1OSVf4c4zB02Xad5EksNW3D0jFRJfL/sYHybC4Avn2Dd9vegIb4CWe
wxchYkn3eeT6p5xmEoAYzfGZaVNoqmgYA6v75M1c+gpOtCC0Aa61D1mM2jgYjtqV1et15BglCCle
qrViWtOh9b3Oq9I+I6Z9K4n6VWNzOd1u5C1+G15t/opjK1n2LNmouLSrKxRKwU8JL8vwJnKIair3
gtZXS5luZTHH41QpSk9w931UzD2YOroDVlk98Ljw5UQBgaZZBQG2YxscvDHgudTmq29+LQFpj9hM
lhO+eWU7djrNmGoIBOE4BI61tvNM4pg4OKYCu0QQkVRJgsfx7lbQUQ3nnyQfhj1vaBxcPTl2CTgu
8gzDn3HdBqcGcnN8AnA5XwE3SzyVT1KEaBItshlcEZmCHqVmqe1W2pzPR91GOBkW5LJVoqPaYVuz
1FnnKr4Ag3To0GHIQGOsyqlZ/QBToc2JRRS03itbCFWr7ewKAKibJGpuzc+rEOeczdqULdSn01Na
+CmaMQ/+9LyOF5vo3BvXJ6vK6pzMeKsjzQ2CNetGOac7OVpUuVnru+7ObTeNUwJTSPfEgE+2/O62
XTYOR7N7bf6old58aLnmgaQnEiKgXdvapZrr9d2BumlutGHVrCL2I+oObkytTbN2srXRyZZIEUuL
yCIkXWW4ZTz4zJaJYLDzPNICmA82+yrwWS1GrxMsqu7xnGk3lvF4NrtO7F6IhjGjkJfNcm1FNFxC
8k1ey32O1HHPoJJPJe6ZBnrNs/Nox3kyD7Nsg0O++USA3aXe3Wft41ccMY+YL6IHFi3r4nDhwHhT
dLAG3OI7A5fKT7INtEtABJuZcpheCJB8CStsXpKkugs3VhuqjBEH6F07+bQsllY2qL1PmxobWHl5
weu8GaRCE4aN2UbPsJqLOctI2q2ZzD9bUaUjMCpO4Od8i+sEZ+34XyXCjbJhkBLyKXqP03ivwT7H
40nFgtLbWanQjiXljnbkzW1PUNhYCkHedE1KWPcrpBoARHAFOA1DzOqgKAP/BGcKLMEKX18Qk9LM
HGniYGDv/siKV8Q+/IsUQA6Nom+l9nmXiPi7NITSmwcYTtuMYXcjd7WXjS65+1nw1lkYuVOrnlGZ
WMKPoRNiH9xSs7T7Kwya6nj7c17i8p9D4J3YHL0is4LT7iewXR8Xd5k/AxXV5Oh6kNcvCEItUgbt
TEwIUE6XZz6m5Nyk4FefSWJw95djPWazO75hWuXu7l6YHFm+wToMwxqAkJ8XRWDPp4QpzoAPjbWD
0ME1uhZvcgjqjXz3woP39O05LUnGQ7ndefZeb8qN4Fgo/6xaDSkbwcoLvw9ybnsaWYlNHKH2PzLx
jFIqutam7VgnMagLwL/uYfl51HmrlAoq3J3pNZ9MTq9SeMxmkRlDmzucQDexb6Wq3yMF2emx4PU8
mWwVPk+f81z4J4RnXDEF7qHPn/lhbleerLhfIeia+XmnLWP8Og8kwUd2hyGaQOwS8u7sMobve9L5
1MiZW7qGX52s1sTg2rZvoSOyMWs2m5ragn192qJBv3//FciiswkAFORPFi9NQJqjKT+oFPsQ2Llm
H2/04FNd2K+eq2boZXvRMX4MabUxnRLNJlv0SQG9QJGLbObpRMqb/K4GTkG06H/tgfzH4BnYOKhs
FdVTE+W3gIA0YXqRo6GIjidIDIoiKYTdNxqGmC5SRfFE59cV8P1Vy6Rj4UgoGIOgUzsfr2/Ux1nf
FS0dvZ3HYj/pf0X9cFUqhnlpcROXjj7tPzcbi8B20Vs+NFlfuxLcZeTVo7IAmLrgfVnPqmuZlw7h
15nFK2AYKOZNfACFVb7n9lPqgsP7vY/9Mwh432jRVWamq2TR/PJ6Z0Hggs67ZVK803cRYPswvF4v
j73pZJusBZrliLbcmmavw13DHrH1v6G8pgQP7I285EhXgAw+f3O4PgpuqHlsID3YQp5P4tMsEJ9U
f8vxne5Rv1nM1uTwwmC/NxCgMrFFzOi9fAZzDQGCs7TSyEP5SE/N5Z7XSBR8cnqka/V5A3osk+Bd
nP8+QXeJX9xbGxJl2KCIuiXJ+8275kme41CuJRRspKPkHmNtnSIQQSc8cUX0DZtQlnSSOO5b/VZU
tQ9uer1fNG8JegdydeXenhoUGC2TWNNGnWIzg5VSSZxVBSpcicXs1nB+/iwXOdfWwj87H6Tsvw1O
6tIDq82scw+RSpHM3RcI7MuHMwC+h27Jqv3y3hmu5+KH0SfXqfzW78djCadQGtkPerl8JGab6igQ
en0IOFZTTpg+1jqTzZEiTLTtIgjUw9/2PmJxZRHLWY3aY5QFIdJoDZXGsF1WBdYlWINVVjB9CpCU
bAfM6fnp+dCH+B/bWI45fAWiVW7vRiRLpzVyXHiJIuyoAWZ3e8OS3sc91FJh5UeB/GfWvg9S5O2O
ZJRgc7aTV8AdsQPkyNITD2hwUUuVKS9mhSW6b4WaiPjs4NWERahqhqNrw55lJ9cjrQSX12+/5Tqe
39oUzMTPU4E/kcNBIUq0mH2JE19psbW3MYMfVziTpY+L+ieH8D3QA2hLgwky98YHkAPhyGkLx5tU
aIj4wZ6+Vqy0jx9Zv6F2tAKPDX7+lTthzUUiC3IWK8bED5paVWlkkl1EWoBYQc5UT2Rl/KsTTxrG
rXMK9VyisZu9FSrVJBIKDBu8U8Xly1YU0dNFtDkCCLlg/Mv1xVis//UUDdsA4T+FvJkIEkd9O0By
CzihUEaPfem7cVbqWO1/JxsC2O0ss8hKNj7/YQ4dzlTnY2ZmFzNhWM5TfWO7DUlgobzb7d7ahcW5
rRGfmuN9bzU5eTSjEdQcoMkQf3mb0Mdc6vVNpOR7hOOlx/W5tB8v1RO4v/bBFpmXR5YUqo/wIJmJ
LqWyw/McNqy4cGIGbdWZzck35nfkOeEzhlVuKoaoau6Ladg3Y6tBAUegx6jHYlHCCWsnyo4MxHvr
wl42g6Ohb5D7fznqpcdrEADS22gctVVhDD/g6+2hLF1L5UD921SqGdTTIsrQn7xJtpID7dgPBu9+
INtRorQyDf1s/cIuRjeMH18oQxrtfN8Th9NVEG8BlwFwrRJREIbWGvSAp0c6o0SGht76fNwmNWk+
H3r/KeTL4RD0WmVdEbK5Qmdwa/npUsKHouJ10DKNLWt4K2elz2LpR+97ZWWzW9COYsK+dwTdD84D
kMyW+/LN0/pe5HQpw6BAa47903Liq1hfzikrTjJxmvc0D7pC9VRfgFeUq/fgs+A7c0ag88/e1vd4
W6X/WSWG4rIzdKVMQ9FkAdxAMRLdrWseaftiI+5yYN1FrZ6HmdBpFuPkNOfzE5o4zgEYNP/pc0OZ
qtzuNeANavisNK8KQsOdwmFhJheu8zKDi05xJNrjbkqij/goe/JlqPZvkqIUbH1OFIN1ILzmYk8F
HMrtDlCAcs4eobqIvHxdfa6rYTBeCO8Tz7WtpRxGHGhY6d8y+2cQMz+x5yZTBA6UqnDYl9EAjwyh
tebR1G1ZTRnIorGANVZ1CY4AKKgt6iLeZiGIazXI+xs+pNwVYiI/HKh0Csn6tPkGkEqvR+/JJbb1
kewkBywiNphjQmFZ5g9n/IleEfTPIg8Eq3CasZV7WqF6jPsJ88Un5fxXrkJDM3t8Zm7FYxD6WxD+
e6QFtMD/OKDhKzYtIUrjfF2UQyn4gSBzRLm2Yps5fhZ0i46C2TYr40YW7jCPfmLr15zKTUYYNdMe
Un5J/KLK7xmEokqela5R3N2sGoggezbPRRTD//J0cT/oO29KpCFnR4DS0UPhnP5JYlldkIl863r9
rJ5PWi6jBLpmmiQwkhmd0tCkU4LpUKeiJsQYmfXZhiFoX96JuVOFGRwnxTo97/lXDjPldOKMQLd6
e94IBCXgtcWziq5PLQc1JNud2edZ+VYRlidzHn2Id3CWLvSNOPi6IW9wMF0U5uQRKr6Xgavuu44F
yZFkyD2dBo4m5SZTczEeesX5hk1FqCstjkc4JjpICzwq6ItICvmOuwDkl9y6c6k7N5GTYtk59bn8
jPKNGp8ukWZ7oLiLzjTN8v39/cQLXZmg5vpPZNBDF40TLMnuI6xjS14rydV0Z6SXQF10S5WE1r63
nHx3PdEfEVhJ5EBxhy7ON552PaiBkWDlKR0HaeLTzyecbJa/YprS/I2B4q2+PsAGOQJ4OomhYpqO
C3lXnASUHOs2DmN1l2K3sSw+CJXE4n+Mx0Kxgd25lMLAfVOhWVy9U9RARE48dJkCY7bu0kBTa4it
QDpKc41nLihSQNccEs9BiujSGtJYj5CzHL2i6rIP1RCVYw6iJdp6oR9sB+LGgLbGNIMYWAzc0STv
r+E5+mpmM0mZe//fm7041LqrFgykrjgdd+Rsw+xHeWzOitOW9n3d2peaO0TU+1ClOSJWAl85vjkI
WqQ4KavezqRxNDsHf/Zgnnb5UWttMg0KcnJETEmpRgfMttWALW60KtLAm/nAsF+P1JqpfomJ6P8S
9WX2HZVEdapi4I7hPOWdHAqtmkF3hJlprnURrsOFcvMKiRfKN7aHhIxD3+m21WV1ePH5e5fjU4Yn
nAlB6F4jeQAUn/ADG2LmFu63/kJIPJNeeNucoSTLG4otzJORxJwuIBeJQz7FWv2wlXimROukgSn6
mo84XUkI4HjXWDp8ups1VVZB0RL1Nj8o2PCTotub6o+2cDJDo2+Kww+RdVJQTUcl/evsj+H+CH5o
FUHmqmLs7c+e0ZJV4xWHJA36qO5k9E/Bc2HLUBgZh9kxszX2Hna+jc74bmwTeX7pm2jmkRyebXSC
MiTF4DdyGVCj3STas1ry8gf6AL4bBl5g0AFcxlmqTY2DVpT4PNi1W3E3gaG5s3DRvefQtlQ0Dz9L
Ge0dzByK8Xei0QCe9+zFln7bqEKHJFoMLgC6qFJdUdFUYS0+zcZPLjERhC1+0FFhsnBgDdQYeLHj
rpaDaWWpfgguupFg+OIC9szxY009UFNtKqLvImmdCS8kKcndQbrHqmoCGeUYiiFOBvGe28Edwzj5
ar1eBLfL9Qnj9AdeQA5OAkn2JyumbeoGarWHciRnNENS/JS43ktw/nbre6B12Q6F1ZnJaGwJCDcd
QfBgbKwXddiJQ6zozrGStN+bh2WUqujn3R1kSrUAPpFT4XbplV8UPYwhniim6HFMmdAqKvk3LOPv
8oFmOmwKUDDugySuYb8mxt484voAucJ6qtWDDM4fO8G5/s0mFQAu5g77kLBTau3D7i9pxKl+BhDV
YPFExUuPeGCHtKgP64wWJcEeixTgYbHxZbJt4ZFVgHnQMOOS/sGbLHqwami2qSyQxbrKC7TFNF5J
hvRxversVXCCDquyVnroDdoWl+wVkL5JjTHRcJZ01zxkb/UVdwg7j7dVZc/1jzsqtvSI5eiBYZpt
epGqK4E6ZamtuD+6H5gYl8N+C4ftnMkuQc6BI/2Sw/aTyanRRkHxob7p3ZYbWhFxPsjVRzRWTB+s
FjPIVurQ2cWORjgdvo8SdwpBQCckjWi5BdPZF98iOPM2SmrtlqoTF/cgq1TpoCQn+2BVTwD3h0hE
d8UojMq3sM07rpJ1j8Uu25/mDgO/foxhDrD81hA0JcfpjjO925R5G0Fu9OHfCfNGoJx8SZXE0J78
hp5be7lXNdB0dZG5LaBRrN02A8oMc1aC17qix07UUMPK1JqBqvLt0D9keMHgaIPkrS/asdUOqHgd
xMWI/q/T5KvB0zQJfibc3wAbeerXHDGQPCV8GU3muwJ47JLxtK9dFiAwjEUmXN9TgFRxVWON8BkR
kEudDyP3gvFYgkFI68SowvWdAesIeTuvbX0XaQyNK0Yv0FXahelbGnaK9DX3+scwv4AV+xL7puXA
pxe+QiRPP5gzl4dtQhj5kjcsjrTe7pEJ8Itq34dKHzNd7r4AWGy0nwxwCqZw6+apVqGcnDGArCQy
fMhN7Le7PJrQOkO1wqx4fxtmbHCeilYeu9DjvBAixpttIG7DzWIMHX8TecoNp2CvV8kl6tYp0Mb7
DN5PO/A1jBhUpjh7YbCbj8oqO6K67a17iXiguSrpMAYjbnixZA8IBeameOC806qf7En95cd277y/
h6VJaMu3GqyUURMmNKj8/+QpANwGIjzZp75a4HI5Kxv00lx6vo3G2eQWs9L2Un8HPwulLRtqUnQX
V28iRLmX551T8KTsQeZXnQ5vGlDeHHAI0cEvGZ5+mqSg4IR1taPgdOtiG+unr3jRfMdXYC8YyFhV
D2jJfkGYZAm+CjF58+cP3li+KmCK0Qgr3a87rHW6soXsqbSF34bQo4VHRs/xjfbFmJvVnu80Iey/
JlJlLOzceHiFKmstCC+AwUPyXBDB4e3daxTcwlh+hkUTKek/hB0u/MYr+Vqb4cvvPIKjzmHDXquh
c0rAxFxNCCdkzet1di80ADpCSuy+PzYxUi/kz54pitPp7XvA1pX2n+gq9Iq6Lkewn253A4JIeOz/
frLvxAQuVDE+6CBwvyqYyggRA6lJibfwmE2r8gNsd5HNa674G8+/EjqE6hXItWNcLwfw9lb8jLb6
1mSdKe3UjxbNtp+hO0J4W+xi94/pn2vNtL7d1UxD8BxyO3NH/43amxRv68sq0ALH14LIz1dIpcOV
RUcbcRh4uGZyKkInlwKl2ekpEG4R5qg56LTUkaB1WF3wNC6OuqrLw6tUGbvUt1ru+Zq7zN1/OdFV
kNgQDRjDuiLMJvo8gd6T4MKiANXpO2CRA7d0JAeww4rnNv1+UVMJvEgVPk1eU7kofU6HbaJkFgg/
F/KIXXfl5T9e3tjWhQvLR8wlU2V6r/OPPXrc4rXSxVQMXLbA1JIN6yscM/EhHekP2B15ERveorc9
4k1CsiV7iSDekh5oS+lqqKAhYzqCWdMvfa9T15j7fmtwLxOyZtgRMwnH5+bfp70Zc5kSIoHYq4pH
0EUCW4Z6NqGrWlk/pBVGXdr+16zxdQXHWm+OjyGBjwTypfktUu/szTVkqfqY5Zt5rlI8iZ53APaW
fur0JAVIQPxHVpPwL+nfsj4Gsxiizp+SulJtPii8VBzjIqDtzb22zYt3QSp9CMXyfYlyTGP2tyH+
+JS14Y6HBuLnCCM30Ohm4RNalnB4KS8Blgh8rNEMH71Kjy2heIHFC/rS86Mjj5h6yQy9fCpRuPWZ
DQcFC0xIT9vq8HWqRulVk4iBaCalZhLG3ciMbNaG7wxgsxsgEPjlakMkFM2z9iThKqqJ6Ry/XE1u
I6g/GYhspKnOeWoIy7xS8zExjeRa0Y+qMAKhOXKdlSjUaT4sveBJM5uk9x184UcE/BUDg2ohR0gf
UCXRPKMgEvOKkEM5VbA6hR3iv2e4ldQMOgHqZkQJUkDLCiuvVKToICeVi94cFUHk3QwxruYNfSkB
x4AprZPRiBpzerwHuOoaU/x9cZCB1wKKlIPtRoqYQR168wz8Pu9b4bqoa5gxY/LTNo58tQOPHCCo
l/lDAuP2EdW4M3w4KXKon5wkfVL+Xsqv4mLTopudw7zfUnJ36NFpexTq40zNiuGL5YOcTOfCrKvy
CXd/QBpTBhyECOcotB65phhOPhJoJlcNDQb8YT9WT/ib6byAIdcQPTWTzsSn/RxN+aueOoirMftW
La1vjUE00LUH10X8I5S9TuzMJvn/8Z9Api4kkhUFxpEMM5Qb8EjP1wuCnqVmqJYss5FPosrQLE7q
BqApMxnySh3sIbpnymDM+LOpMKnCchGp1b5vI0U5oFNZOlu9hlbJH9x/AXjseWHKIybvTYST/TdA
YTcgEIkWh1EGLN2S+FQMN7BpSlBM/iEhD3tpBofvmdvb4ELzSaqfa80qeCuUUtvjRqh7R6DIKQmA
2mndD9Djtz5cGb/yLBdPu8y3p+SSsjVgR4NDNFpyQFlJbdmvsp/X+jPU47SdxsoV9Jv9uO9pEsG4
B/GGIBGK6K5aiFVmZDlKW8twQgjY1or47F0GJZPmBK15koj+EjtmR/BGJOy20cOrX+izUz6An842
UhlpH8VFGVn6mKOdjmjSvLhXkCE+kbvx/LUAE24M7mJr+/aDXJOSqOZzvtLXOx4RT/9CMCO3EgSn
QMKbZN8ncnWKrOWSH9sHx/cpC9cRYC49iZbv+rgOgp9DNURR61OeNBAXfejLurlaWP5J7EVa0gFC
/m19gK0FqU08VSUrKCk80nowm+7uO02lelpFVOxWzH+ySUhLzNdSb/bQUM+hcjEadTaCKcLrz8NL
DEyWy69Wa/ip7FRJqyDgyzKA/Y8pd9rj9t0Xg5x+7J7879UfmMKTK9l6rIOozqVBdSeLQdpU9Ruz
G22TsfzEVmglM9oS17ABKccBfj/JXuzDylo0XFLywHFRmB5RYErVZyV1zLdhYqimrrY0MNcNyspz
C1lfUIK7bAZ+DdyYbdDA/eA7AH0zgeybpAW00VLud9DRiBhBvrUtAc/8B/FBoRDt6faUwcCJW8tX
pMsWG5P84bg7oucQGfTYh+6jHRAFH9AlNBxiOA984+nYtRi3Kvq3GJMbnO20S/3Lk/O5sGOBJA6L
quV2piB8+VBazpjfnFwOxnGhYxueGpSa3p7VgK0orylr9KophX2TFVBe2y5rsDGDgLI4t7moD8JB
ZKWmHqD13ZBp/Ezdsb4YXSxv+ImUJ7Z52wsO6ryXz0V8b99vr3Dgmk/OBJrdK6sAJBE8vUwLEGrx
/wbxCcjRCvS43V7JvK33N+OAT9GQJf7FTlRaMRi0Hcvwvw5ez76wuiRFv135z6YWrKiDr/hM0JS8
xOvNu7a/N7/S5K1qcPeH6sypcIgvQ14DbWBmO3erf9F+AS2qElG7R5OVD781DvlXMY4A57zthuzP
P3ANzp3BxPDHL1rIfVQoIYUliNmOPnE1R9CTrhDpmLI1SBZj9PF1yaSHouYv0h2Ttf69m87A7213
oN8zizhcXh7pVCEEnjn2vOxhG3sScxFR0qxU4GBbERE1OtmHOkzObyG8+bL51RmTK08nFkQmDMsr
OY+isRCw/CJpXjjwBSwQtlUHakUptu+/v8N2IF3VgScJurQF1lb8OLW4Sv2F93E0SKbNqAH6RVE6
3F/0AwEqKSWbL3/OKKel8kiHZ2Hgwkn033rbWy2yw/3Fp0I+kppI6SYN5hXGYcBV3kb4jM/8vze1
rix+gDn90QCtzfUDo6LT6Ohpmvo5fyKkXZ+VDSMWa7pRw2j0ohANknb1SDs/Nuy/ioHLLkEL6zYP
SPs7MbL5/yPR+It6IwOw8QFzYDJ78OVjKAevaUZKVaXONEtJcUJe2ETRA4lQPxI255IpHOZEOWE8
VXIQIS4w4NNQoa/D3TKeI/uSET6IkENQ318323FNtec9PXMpxRJZvFUzXapw7sFn1q7pg+H9DtFB
B098PjUOD38bTdFAh5/1JEMWESu2/64dI23PVBfc0Y1LnbqVQ65boWuJpf/ea1tkdwc7EQxOfSGZ
hsmKcOcFDA1/xXVdfUSPKSEZzhQoYIWNJ6jsoIGrvd0CxiZh3opJJNA6Z+qSC0DKZtHspuXJwZ25
tMnO1pg5negDpp74SBip02OiGvq2WVd7eqMVeGeSJkgnlydw4WMWkOIqwfrMyz58GD344k+0+k2p
f+9KASzeItMv1UEHQZE7hDEh5AJEvA4ZudKRzVhP4wRi6P3G4bduUoImIB8g+vVo3rX6AXqUx+t2
O5+kwOn2CMx9V84262fRNdar0/V46/tYEvmDWFV3cNMc/JwcqrhJs401aNxi+pq7/39/lL22/aGo
2XRANRP3K6hk4zMu2PXQk5lpFg46P/MT02eoxWoeWf4AObm5Uz1YHFWq0OHKR6SWg18DqOUti/xA
UpdyECKENi8ery7r0SmrY3j/U8vUjJHt3SsnbOM7crINi24OaHNmU4b2LWvak08o1QWYD7heHoUn
SbHjjJhODYi58Ce+u09ImQj7GpPtE9EHTLGyJW7RNt3xodnwXdMDVngJEoBn+3ttXyHIJCf6l5Hc
5IMgKOG9y7Ijw48k04R68/s/L17DO2zoL5QP4TFvvYa9Iafw3cqmqH0ub3ih2wtoSL91xoF1k/lh
K5OKabDj939VqbJG8q3U/ApYA6fxzEG2osrFbozsrZrNSegNX/f9FvthywJbo7i/ULYDEvLFDKU8
Kmjqvu2eUYfQRdK33lZwFRXXGdRbFG9B6OsZvAfo9rnE9n8V1E6/9EteqX/KO6ZM+nnQkTrXZQ6w
Oftg80qUQhwB+O71uY61hD7qVqYrsY+Q+NXz0Q+ZVQQZut18QIMB8XkXyiWBK/1ta/s8hartgwl2
1TxHL4JCPabbnVbQgYn0oDzKqErCBqHS8isoBlTL/m2kc+G0rOiBG5FaEe/Bk637TLsg0B6hrBur
E0OyBeTE86F/1pkz3nS/uvCtFR2ndrktNym3DbOOqh3XsIsIxBpjp7R/mH1BGdEMd18iyTzPArt7
sjj5Z4BoAoev8WBKorhMXNllQso7ryPwBTZ0URsi5Cc2IH4CwPonfAQPLEG89EbvkvlEUJDM5385
LlsiHvCGrbtdvOAcvYvEkcU+6CWBhqVsm18mMpenIiq5zkzWcFOz32f4uWXjn96GPpGlNyAnOCV0
KTHAsTscH5H/Bp/Knb6GpPMP824HuVTFnFq+FLVPl+N0VoTVml1p24Bhpe77erFYPlpfvJiRXrAa
hvr0O8e2ulLemtHbYjQWAuirNYpi0MIabJ3zXoDO7UNNDuFvw0z8wu5NCPM5Cup2YUGZarNSy+Mu
D4wAIg3W+bRL64cEAzRTGFStQ81jgNk0tZdJniZuSQfNZ8X9u82mPMt6dcdxH6AOwaSvp2vmKiwG
lSA0dBUGGvjiY5FpUyhbqygwC3FjKoUtDGhouYpRu/jks9Hm900Om9WH3rp1YpDFtH7eW3NItgwC
UW/QpV9iLbLfvf2+hXrTeSACqwOKehbMI++YEcVNBbdaAzBcGPn+6cINOsCQlqukCMq3WNL1YA2u
WEnlcGfnMZDozEbSrB4RneBXHEgye261y7hcNcrrs+2Fl2Zg+fYxVGSuCikFc4uo5VqiWeKDixl9
zBwu+8u/fynth/BYMw9oTd/X8IiU+ZR9v5W4GMdi2AMg7wRzhkiUVDxd823lgY9HqHS7JDbsIjms
ybXbQiosOsSjQO9Qh/0ux0Jf5gd391oUvfmKgkE9xMBv9qDQWYQO2WOz/Y/fEIYcjSm2IJJJoDLW
3EWdVrvd+B2oQbZjERnpWPiNytxIYzWtBTw+vS2OCFjLVdaJx4Wtx2Eg7SdcGxxaifhz8uz9wV5J
hG2/diyidUKSxoR5JXOfyRmSuTV3z6ap1iHLiYwfuNnfJWf0QMugu5YaRT1UR3IPnsc6BuLkeVsC
/CHfYggC7UKkQCXrkrfG+MD47OEwIXkXOZtC92JLCqPKkRRM/qkNjpO6/W28lRgOMmILaoIFgbW8
v9SxnrtGIy3CIUD0pXWuTR9OoPSX53YVvK3nvGko+b4/xVtTn+z0k1nUyfbDA2qghixlN3K5pLhH
4A9GJzPYHjB93k925JzTBRNRRzDyIBsQtb11IfcqbWW3wjpo2Qj1dW5ejpCJRiNM5t8qhP9C7PB8
W8I3I5coD5BgPJYRoGnbYNnf+QIDBxC6+T1h7LXIOqd4GxYppWS+v/NVxSSLI1DXJmCNHv2dpncl
NGc9Owt5kLgyaI1xWO8T3qah+8oQa7wKMTSTfOb1AmFzPQ2iBnO0qkyT+p7M8zeiCDRapdaGLbCt
952+DfiQ8mC2NDPBRCqCSiwjYKgjoeLBqcHjBQG3DZ6oWdUVYdcIeEnR4GAHevbpZpwO59V6eYTi
3ZMiAVXSUsnLAW4/nEze/jTSxUBCzeGjBJuleBSCcAnW3k2Wj+NMSy15xgsLVq3W0RX5vSOT+CvQ
keD4/EhCVHPg3QDfPskNSdW1e7/io72FEk8bhnKaXcZaAydag5YPjKMjwaT1hPhFOPtZDJonXSJo
ElIm65/480WCVOFhuSz1ZaxK/oRTBBKZb7zbPDtygslZYu4R5MwkdKNEiYVzWSLaw614BDPiQiDD
sfQuh+zeO+pMpZR6Exj5NyYP/8azYsU9xC57kyEEscOA0xZJG23lGsaMCpWxPtM15TfIs6+vrRSm
nbYdzH4y7Sj6Z7Wj4QtKVHim4fZMUVqjtfRjLi9plOyNB/VTZ7euWrGa3IQNpxzbUPVQidkMcXnJ
Do2IZ9qOgVw3bKyPHKAS7rJGVUetyaNttDwmiK4b5mVtFc2XQBKaLZHBb/WVyzQs5aygt8/BG7UV
fNWlU6elRG5Id5EgUwhLf+IoQzjTy1tH6PiNMefw8hFOLTJ2yWB7o1OciEC0F67jvf1xR+Rlcm+a
bPOKsNht5AMWd5groqZM6znXstPrYlbv9SD3DZwXOGbAf9w6GTpdWR5EoTya/J4R+zjjrMhyMdZg
hEnVzQpkYSlcgj1xOXDa1IUaTc3YSHqKA9nxmb5Fd9VqxSn9D0qZFFSI7/YCamYLJEDEHcUReGSD
+Ye2SJecoSw9lC25b43ztQR8HQeDQr9PLiTjhrYUAckZPuFe98o55alxob4YeGjc4jBNb1koCGnq
Iiz7goOAm1vQN/mHVthnRxmAyzU9yo540bTFDD2QNsjAkCRhjjgrjWqt9UN5xa00ej2yrOSNArTc
mvnRmeMAJfOV/vh3Y15hxLedXE/T7FbamSgMAteFdwk50UMx5viDMeErdC3TzOc8glYc/XIs+yFh
CdPcGs6kzLivvVvaxODeP8sw0/C+025eTxHmtZfPtrgJ3cGE4hPjCMp1h34bjrH0mDTBmfUlszNp
ZvyGV9IJ2gEWpEJ/6vRhuGmuQTidvIlwleIjLo2cqGfsxQRTX7h21ca3PskMPsiYZGrEdBkS+Ozv
bdrLtO3T3JYV9A6H9e5uLoVHmSBXOhaKMzvBOW1s7kFtZN8voOdyWXwFqrhwtT7MzBtHyYWlJrhe
Csy0A0XkKhV6VnrtHkw521F3pPq1HCvwnMKQs0BkdDWzfCVE0FrrihK7JnfXVbv7u+pOin+jF7VJ
pl2DWpk7ONP9hPsIIMNDJOSJBT4Cg0WDEBpF2n3eLgJh4v1NCV/NRMucVWRNJBOaImZcFb6cuIjd
54UXOVXTBOktQq2E+1soh/H0pX09WLT2Bh5QP9ydt1G8gX6SwTfH2RTdSwtUQGDUTX2WFG6NzA47
PQVHi/TgRE1FYsr740baJxxYYxSiNxlmpnntdMKssSB+cVBNEhnBo3vHJLdKCDtmC3MFAlISGGbn
Z+0Ms2pZHf9HhkeramCs5r6JPngZ99h26N6BW3riHO2DHkeyGz6GvCodIxh51dU0iRnhv/upfMn9
v5SwXDvWSh7qAR7Bc7rNzBf46zlf7w==
`protect end_protected
