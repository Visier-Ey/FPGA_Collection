-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
V29SnZsTxGLkHtRYC2FSam4ZwW9DkC5+TstvZTQ42VFxG8MOPaikcdfXmEwkPLzCh0TtP2NXq90C
icnwa6hR+EWrQCmkZ2XhhifqSFFBbQvktDL2gApL/0r99uBj4+t+nOjKZ1Myh+XshUWF0Oa3MQWS
HB4B8zixLCSgMVjhd7qWWV2ZR0I5gaFatOzmdIiASTW7aib9KKsZ3JVkrVTZMYdBy9adSdv8LqBB
Q5l2UEmGajRndDxoJOPV8fwrGVafYHT61jP8JWhvmFHLIr6e34el+shYCO5Ad/y9lv624ATskpy1
FNaPtJiakcKYqxs6VtV38FwyTUXEfIzRs+rhGQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7984)
`protect data_block
1WEoLwM4k9YFuT8qG/flTBFejABsCrHQq5k4u5kNSW9ND594kXrjuAsowxQKMBeH3xD8Hov4+r3/
vd+kVNLHefCJCBq85BMxdScq1lWXLjZvBj/Wv5xbGJhmfmbodI2IjH84GzzxdALrRE7hiw+pF0LA
qP3klrLXg8sTjcgsLHiU1Wer5vkKXCsnntRSgskjBCkF8pYw0geyw+wthPgz5xgy8YYawxHQyJYb
l3FpaebDFQ/qJskaRQvVtwSk0fcB7GqGk8kKghrlZ4ctpNWNwEK+QpAgwRCMYhXstIdDMxVRjm+W
HSFgsWTSloV6d1KVTxif/gOSMFlLlJkuFRCu77yxdPf4obCL52UgcwNzEHuFyoDiOVl5pQ5bWTzJ
w823JsG0NaMCO9hDv6fJAbHWRd9mwp1CuxShqJaVuOugLwMiXamq2cIOActWOMeA3wvAiCB54VF7
abcW/3B9oKlPNV28NeGJhTPm8ErVNrvuKkO8rbD0VOt0aGnwCrkLo45xJEOnNDDi02mvLNhArPDy
HeeYJJXi3uAwlCYt61ayPPwZ29Nwh9+u6+SabfPyIT6KFZlKehJR/GUD9SzBQkCpldSrwHgXXSLD
Wz9AMxaeaxa5vjSeQRyQZy8plM3WqRA6WypAHg+R9G+ORyY0ocDUzzQE5XD3UIKL/YyXhSkp7ycQ
6qzZ/wqJXra2J3KACb3WWZ8clKT7TMcLpgA5G89Y1YlnNa8sXtJ5yV0sruvMv1az+bgiLDm2USgt
1/eIF4JO0HudBbq9fMR6YdamzCOihQeE7thAHYuxkVRGHA1qjyRDL9CjS9XkIE5ckRf/KEb1ZKBK
ozezbNT+kPPO4vqXur6oIOnLEmc0aip0fB8UVkzK72L9hSioS2l4bT4yn+sV1Np5+rJKOyI1O6GN
jg8bSt3feqV3e0Q+JaRdGieKaubHDHEYCm4/OzRGqWHS+7LArbKbUHW5fJLb/dT4bd6RpPIZMTkc
bxBAPjPab2UFkFLA4+iqsUw8+rpoFzHRvDbhOSQDyLa61YA4wZEdeMEschXTa7yBdX2FCEBkLYEm
ErOL4PFN0pYUnTF+EXNTYG12kyS3KSbxj/2mTzTpZDRofzLQbLqlNz/JO5glsg6W5UBFtEaC1wRa
6BdldI05wMPb9btuw1gdQOqbDJqouZFA3FaF/vcZNKtrCQ4/IarAazW4nv2wEzdQRqYfdovOerVf
0ETbmswU0/s3r7EEc3Vb52vKpG1zG55y1lFtHG/3pyfu8hg0hD7vYG8Ff6C3DT/Sr6+TrNu3dN4+
a8FUpdQx2TBhIr5UchQgPY1ziPHaWzkHdN2wiZ4nfmjSA1j9xm/y91s3a6bU9YeRk8aMSnPaYwzH
lZ0axub/cy5yxdvuidyHykxIjC7G49VT+xPiKmVXvKIBunkihErqW263KBtZJEt8hKSmblaRolHe
4a4b9wnNrWSmi/3KdZrho4XUGtQFYd6tfKUyABKFGxAwv5K+dw6ronsW1oRCwHHTnz5ui8shftIC
NnIahS8ITmEsUq57J7iOzr4CObP2p3fbhA4vaj3CQ9+K0lb49j5l/3O3/KARxwf8hm25xEXnDbfJ
GazGpY0LAT+6N+0Q/bS5IPHok4Lfl8FQeKQ0xj+jyIDzX1C0Djpo3jiO4sbefOYSTtNeCYI3okps
5NjvO9mvykCYGa4q6JfmZcznXrxS+pZHT8l96I55c67pkCkEgoi1v1ARUc6SJYr/w4RoDaMhFemr
s0YOgYMRBFLWBNW2LntEp704s/op6Zf6/wqlCwNaG+hqAieHVKDg4tduu98KhW7YFNPWFzGR8Jpe
0hFywO1/errBk8FsRgBtA6qx20k+awdduMpOlmmz8cnWI6NkdfnnxDxcRJ26iaTUub4dH+nuDw07
nXWOi6rReVXYJVsZ5Cn2NVE1TKIcPo7Um4Oh+53jlOiu4VBH+D/bg7l1Q/wZ3o8SmO10IMW5ivmh
I2kLPYD/NZUxzqnfCiAe4n5EMgeF+KclPAmx/KWqSBrtupHLwNL9iaVTEp9LWkVKLYQ71gJgW8uH
gZAS7PhhW22sDSGnlbb/dkyozA98FwDsonuVxA+xfUoLZ5cdPqnFjI5w0HqfCIWtmo8jpXPqEeNs
MGOjXw89k9O3MS8FwSc0GvKLs0kR4Mi/GKRJ0reIJpRTPzZ+bvC+YpAw6dZXop3Iu0vArRq8cX6r
b2nlP4vEjBEjkv2G9VLtTO6GW8zqulox8OOBWfaSv+//lPorF2aJp6nhuCHghWnpBjPBR/Bv3NpA
6aXedRgWmF1zBCidg7pXHfHKsQ6ZbFT8BU7BQgUfsXn0oobTI5QY3i2rUJoBTMtGE7G5Js+2aaFc
xuwkE5DIphV4dOd/xYkP3DN2CgDIGxlyb0yly/o41C8uLmwK9HqbFRkZx8Ra0eWItKtBkud0qnS/
aUyxgagIWwhnDzt0c/fXzQqa4wvolIUd2PjgzRyJs/XQHd7Tdu29+Y4V69pc0WA9/wsYBpQb1i5H
QPZ5iaPR1Hhbk1GskglS8J+HA1m9dRghFMQV2yxL/O2rPvflHtD2pwNeElwdMMgYOfDj8DT/AEvn
Jh8oHmYgyJX/I60Bck1vWqPcPl1z5SmlPzYuOFJYFM0Cb5tMPtt/dvBoXpHy+mu228H9ltSC8tFM
WLixBIe9gzOixFV5IHeUcfj6XcMo8z1zKbp1CD5BSNHxYEk/SkgkwDBw8pqEES+XT7RIwQ7zSWXk
oscDgyiKYmMcedU6uTk4n2CpEs/XM5BZoHHQEGBdr+DDfAtJNSEY65x1LbJnLUybQgI+2EnEXoU3
j/DnqP2kF5LzCQDJmynq4jewGRLVKeyaCaKP7Vb1mOrmOeUBysxrWBDseI+2yjRYbSeuso3PjK7U
ROorEqYu7lmXIXm0mmhpKEX5rkwBU10NptpJemB/MQdw00YQHReW1muoA+SByBWCrLYggXTTTrTP
x1vAcZNRGQWtnyjLq07mRI/IELZnSfmwHW47ky74g+wC1RpRSAzCNq91DdVMjRdBu/M2+gIP/tDh
owiaavk6DHbTdR5B17/fht69TCcVLGB8/rMvifkUaHdM4mfbTasBQtQd+D2JBO5NFCybdBgbTIvB
cqz5+saDvqUnOgdrzdE9J6aVVWU3eVYb6OBTNj1ZbCdI4M+JW2h+dR0+uy61vx8OZTiHDcP5TWIt
VrmR4TvIXUjwAqPRpi/PsGzRSqPLafem5qKebrMjJ+rLinfr/2GSpyZtCFGIWjzgm8d/PF2ABlth
61e0rvKOuJaLdvuYdkB3lh1B/ibz+7sd11LyIi8QTxo3i9LcZItBiL/ihz+zjGlJDSTQKmEZLjZj
osJALGiKgkejBelNntgC3/Nsx1ueIkTaIfUo1Wzh0LM2bWYjE4/TyP3df+yAPT8NKVcvVYQIahvC
famP9MrMXfbvrV0y6GoilGXE2dmDrmMRhpnMkzmNFUdMAQ//SAZA5YCb9Ha8DJflnJo04bk9KofE
aHE5yx7VIACtCvivE76NLYo4PDKIwvJl2Z1wUn/NL14cr7jm1TsbMaTDWYVbkIQcnuBQIhEs4W7o
WYHK9V9hLMvdpb7PKjyYfxbNwHpFI8VYOdU5U9D1cxti6Jd9nzQH8CDNeqv1yulVUPREc3NVS8P4
+2qpVyNjh4HehR1Y9kK8jVaNk4Tc4VU5L/PioLbMsGNI1pdYyA6jf6IK7Tqc60cfGb5cbIGRSMZs
DZ6RJqHp/ARMTOBzVVtFVRiznfcnG2QzZvtITLEeVuqobJR1VJIkWHSdsdnHMPuaT9U4GpF1er3h
T2JyClEto+75494yNDhRStazHPuvkJ/7tvnmkZx/tYscHuZzG2NzODr4CceKyjIXSVPeugBB053+
PyQEyZsWxZouZU5XqFegnZsY3I45X2tegRSIzBDy6NofbhsBDVaJRfp5Kt61bfTPgWjFUXKjdfBZ
9azVReR1XTQLtpj9SD5qD46lNejRiquvjzE58vSKmGaHpRDdd02fhV/+kbkEMKYXOVix+8AZti5s
X9Nvz2aJDGHKprKyPHWnyaGCFPhYzaItU0lkrgbCjnmfKyc/cEiTTptPLhKs/Q8AyqrgyHZYbIs0
2ZdlOzKptawCXimRRDO9f8o/9cay29Pp0vOfYSioqpeMda07ZN2N/kl8/fvA/NCzaNxsmaz4daqk
TTnWaRWc///c2e4QNoCOskaYAqz2MKkuRPuJL4VwJ0ZAuEbIApbSutKLd6tPfjYWrt+NrumnQU/O
WMgmq1A/V7yisd2MoDPjT55htBGHEyEc+az9gChfLrRLxQT8gCUvA3ie7yT+UEOKDIaod5CDq6IL
U87HqkH7Up3xzQkZYnPXdtlYcg8xTgStgtQv4SRGGKQORAgmBJ0Dw6Np95g0rGMy9JK6HVDxJCuZ
nQXxp2MyFkFWBH29gOOhUlN+msgnfON7afwAVF5bYUXPX0HjYk/F44lWr9CT9fHn/mmGYgpLTYyt
68rRKxmc/kSgh5bfCkkgV6XUOfvTST6/Xq3wBGD2tMvoDfEvfEePF3+T878y7h/AEi/Ao1yF/niw
e2jVzIOVmpSxU1EaultU7inMbL9iewuon4hUirf8Zps45GP5vdZlNuxBci6dIMBjatAlV6whjmT7
+zQ1UHhESjdRR/nzwd6oWPn2t1SBua/bGBzO91OtkZk4izXFAgC2imBDtxReLy4HPBEK0cQuBjvw
ZBegczhnBhVobMYgESEv+YX9fdmBH+LtnyIkvIfmZP7iQQh82ISjDUcNDOz3AxWNQOLFNFWxTlQ8
FuPlZZvB/M3HDpgIgjonv2RSn6LqmxpjfkGFNmgr2kJPtBDVAQFmsTXxb9m6mws69R4ef6f3NHQH
WzZ8Jj2QU3IKF7Ap8p/se8NlfVMBeX5sMUXsB2NW/jg1G0C1LvNu2RjVqdH48CHL1Yc37tLF8dzo
3L9hIZtyJxFva7bgGRWetC9LbXblD5VnAEpUnnx/Ueta5wbTz8+pWko4xgDsK+33DniN8Xm7f2W7
JJNiqtj0z1VSh5Qo1ffKeUDwrvcXZTpesWekKqxXZSyqd4EtxozSaZrdWP3zSjlUlnu1ixpoa1TL
RFQ1QF4I8qUkOFbYDivRBYXCRzwYNv8GRODKreCAT/+dszcGEMCkS5ujnE8p5Y3/Y/UtRyRrStWC
QgGUjZSHEF2pS/6B57SMYQRt/lv29Y1w31wR74FAgxI4GnlSOSqpB/0ZM10hlWF6N5bOvVrlGM/C
P+xPc/bRZXc0MvE7pdR5jK3YNuVdYVRcRnJ0acpCGFSVXzZQZ7a2tEYpc1/bC0zBMtz6irJaJyGQ
ZxuqC7LBpGiVAWTWdPZpeVS3QA98hRSnMxO22fIV+7BrftSsPaRuefeV/NVBj/2OKc6J19ewxn8P
ov8MXLBE6KcMdaLKnQ0tnFjgw+F3gF63u41YTYxw5tEjRAxTOQmTkJqGD1EJ9nvzLht/xlypsYaf
rpv/DqiGOhpFuJYtVNeeGECdUALmUwLLn9HInQ+OsEaprHsFkNlUNKrf5V0wt3wiM6qzZ9nvURXt
qFkIo7nfY8YhQvjW2KIwTgrz82aOWfej9WipP+7dJoH/2lj3RHmLUwDaKaaVwZM+YOMNbFv7AYM1
fOn7mNluTqpnn9WLHJADdVVSojrUbO8Zjv/m+K3fX47MFdalgGbTisFKMuEKbp2UOOBDPOnpvtLl
JgZ32QKqLtOGBl/Jan4+KJbH4LR2fsWlw/r+mWJQSFrrwCC83p7jCHvYhjnGyasNb/ziVge2+0oo
4iTdbljMLJqnm5+SoAalKh+FPBgiYYqojOyurwSxBDxO43XGVG6uDm3TTKI1/cuX09bZ3qRCsFNg
KfN6KP9Z73HS00EVBroggKyWElvaHekYAn5LsR3TK12IxH8Jft+gwIsyASQAjloJOHjEJEdupqXi
xeh6r1xtqnEhe24hT0RLwpnwL+h3Dp74KO37CtdlaaCi4262ZxY3InroD0ZXNSZMQXS7Up+8FxLl
ts1fbDKoTBerMLgAja5c2pcCPTMj7GihosC3wk3ngqZ8YW+g2SiYbRUAMk7lZRo/9myJGGcaYRqi
zGockoOwM/0Uqlr0h4yl5MgVa2Z+d9ppKyHkF2V/H1igos5Lq6ZobfLI5LlnYwd+D/TClcagBi5a
mg/UL0IkNdrA2grA1foOqGWxJW2+tLkXtR/m9iCTV40x6Qgce383fsvpwPfXdQNVHO3DQJs5okFN
kFexLvLPvJ0dg25zNwDtzYIK2jZswh7WXZLBZ8YyZ+lbwZGWGJB99Avp8eLq+xwOjxKLzyz+F8nd
CiMubNqaVzyobtlznwTnmLvKCchUKL02VXJ+1u8OUP0u6E2C8UA2DQ4/zIbSkGAVgff3zvA3x8VH
Abq8ekJY7gktqm8OkSCgY/LTDQT38whfCKk/yxOwAaRJ8iS2yGzD6Sqt8tOKXKOrRKf+VpyJQXRt
UoSXaIxW/j8RtP36oefYWsHU0IQkn2kSDleJxauHJ+OMnfegjh5oATLfj7MEN027fOtWefTX9TWZ
iI8ySRl2YNI5BczqB16EweHllkyzVcNJj12EvbQYSn6/hofD+bpnF7rPespTCBrKDgtcsrDp0iD2
gA/wzASiRBN/1t0+UOvSmJPqO5aC0A1EFttC74RzvoNd6PSn3rlE+wJVaPeSqy7N7QJrhHhZrI3b
TfMELn0JYmzi96dVrsG30WbHhjOufRdgPoi0cM16HdnHCnsV7GZSsr9AVEAb8NEcP+zcXQE+CHiJ
L6Xc+z/xZJJD66rqd60rp1/OFK62aGPzXrnCZKSEwk9x7Ninfk+o0Tm70WpC7Du7aw0TERTENrJf
yg06NsbSTZqwmhQnXSquuTWu4m+85slkJW3RsuRhLFfZ5UKEhrSKG71r507+T4nCHBLU8RlyG6w9
qVLko3ggEvKuyDIiCllMAy2LkLe+XW6zfcSZbpTjjdM7zxviDybSe0YlwiUI0U729e0f8bh2Z1zH
cLHcwowoL/o7OBBuApgzAQ8e846NXPLjBaERq6tAZOeRApUSq+bNTgFmP02KhqDHYKg0yA1pkA2U
7gFaf7frmdDA+mWzW966xsrwTxIA0+RkTne7hWz+yWclvQK6YNUywFKOMazt9CZ/kpXdoKJ9ABCg
iGgDWpQFQH+kf5+llVtYyjlDJDMtr1jDy742inajcSBWVh7yOLy3yBMSe0yWGxoUctAiyInItS4t
oHSedLwbmCUEBHPMyt+t+pgpjtJEUNpZlEefvvlLN0PRZFMI2KZwPMSzzXVP16dBWSRG8fIUGmcf
ffjhxxuvMahhHDfIO22V0uU8FZPpSs+U5MupGUAmlf4be7xix2oQnQuh/SyJz6dnp48iOEMH2NCT
EJYqpjKWv12jqTCR48rc1zwLZsI+dBSp96iITWgK9m7Q/jtif69sH2fu+WwTL2FgeeV0Q2svPcBr
QVBZY2EKkoGrhaojbMPyy7PG7h1BWok97hCebTPYnC6hzAaBgMmS3urDuS05dzYSJe/VUghotqgz
Q6yJmpR4/lyLqwm8vQ2b3odAhXeBYviKr2YHmv6RhpxvSHVhSaj/4o7ZfX3uaqzpNYfFsA+zUd4p
HzlZlle3l05uEcLPYorz8eJHasj1H2KnP4VoRwFpaXEBm2Ai+QM4DwRcGLzVSvTd1VxqxEuj7S03
o+NuMq7IC8Jgy+Hdf45iK970OrfiThAvJ3UGnm3TrooJTXCIva8b+R6K/QO7UdUwSc7axcAXjjEK
2qiUSR89AABkxVaQKRpKgJ9WkWWeI96WwBxReEm57vXkysIRM7HrUBV1VrkC0Fdr+WiSTNT3Eo4p
yDTAKtWVWGyMZKWjVrXA/qHXhy88L6XQ+8DC1fVBVme2H8J4RAg9da9EGMkjC8CYxbz2ucxFYJT9
Gd9XpjNoHcXRW2f7OpklsgL1A4Tx3lhnG9hhyMqagm8CA4HQ+CKSQVBXneZ9no+apIEUBg0K38f2
NNSvnTY+9PwpgaPjQOkwvYrPxWmXz6enXoxAnxzhUkPVybiFP1ekbFtr8dXLhgSW3z3vo4B9ThgK
sJ0W3YVPSZ0QHgRg1FAXUMfj7fo/7txr1+B/CIwCxVA28rLxqNYvJITZE4kP+6UqcaFIX8oaixmo
4ghsMFzJsTnGrVvqor9t/RbnzDzX76I93l9x0uWa4m7Wy3tpeBIipDH9owcbGierCFhsglfYx3ta
rTnBauRKKRWL+BklViMXZHEpB+RVifTUN1UXqq1jWJqF9bGLAy5jA81c04Sf3e+NATuIbnhlPmtc
REdCZ65v+qky07Ji1wn3cCTDWdAAeTit05bi13CZHFFUcMGeWCRM62sPvf4G5OC1Ouc7L7lY7wMs
4iWM7vP5MUWD4NX0KJCaL0BX+Z04eto+vmzfieOhS1aqGHMDnCC0asIjvHanGo0cwjsHiiedrDcW
C2rhO4owch4r8QtC0Jk8ddoKlofs2WNVNW0IEFNFlbaHdSCDRGJai7+AUggN1g1ULuQDQ9hw5czh
KTINU1nuZQT+CeIuYFs34deDScv4NC+5YAgxk4pXJi4RHRULxyWMWAmag8n+q/BzE4G/5O+KcS4O
jgCr52q2qUJiYXhOv02DUw5BBHDMg7YlHFo12CmdPt5Mden1QNiPboyxBYfr4gXd3maoh2jn5l1R
XxUmnBtpgUZa8owDyejKoF6yb36rb7vmHtmMuqZkwLZ3zScGnyOuoXlTIHB36OrdVKi1HcgyAT2y
rWouTx4nchIG7AUZ7UeNkllAhKUELw9oBDg0yQjQRwRHaGFXty1avlUlFvx8wlhBA7pCtLQQWk4Z
fikke7qad8wGwc/51Fc5aogdDfu/GxHqOLODaFH15RmjIOlW9x9XndhAbiNem/QbNkjvcfFW0x5I
TBd1cEwpN2+W9VJ2Aj20RyN3WtT/B0x08O24ReuTl2SLt4vEFzAz9aW1CViIHVS6dFt2fIcAh9hj
e78ua2xjOFjcbe2JfjaKNB3DPpIQ4t3CF+22aFP6n6SQOl1/l/hnxQszDwTOEpkh2Da0CgmMW9XQ
GR3hqB18ycouwKtGJkAo6S25RxHOvERpF2Jd45xfqVz0ThFkyG5vT8ma1LzxU9Snqf+guEOvqYwm
hosfEQ8T5lZcG+iFZEMIclaFfBJEqHyx+AhAMOwGw/MALuwBw4DoeHLGGnVv8Ifh8UQCCIfcLWTn
5d4yj40YDanJgXgX9Mb2VLJlrOlhgATYPiMMzHkLNwDv1/9AQ8ra2ogMrVqPF/NSLEgxvf1V9YXu
p6r/sUfiKDQrlEatZ0/QJloDMRu15rlzKN48GEs9E7/GAHELT1G9Psydm3fdjtCb7UozFSn2ov49
FqIHYgrARdOegSUSm1klOxBzN+OEeyq2CXIC17KwB/L1aqcJFYYp9sgFqd2LxmQnLIpDbhKwdkaN
HCHrl3XtgBMplHTQrN8uIIT41zIyNlk7FV/yEyVIo+M8/US/dmLeIOLDDxXJPyA+DhpW809tKyix
wZU+w4pWTwx7wJtMUlgjx3oaFPPxho6y0QIJeaCk0XxjK5/WF3JzLRXcy9wx1WYKWu6mnmzEmO1z
yMrNaQ36us1z8zo2RRURJuBWrCYp7OT+aiCESukhoGSaurxlri+TzCwJzIxRAPlLpuey44fcbbEQ
enxyuLLitptzr34+0mkVl2Yq63gs8U6uJPMXkN1hFzD7PFgNO3ND37f8B+m+yAQAAK3SnXdN3hRT
n92JVpXi6PBsi9M0eAvdWaTixYjANCefrWDdofO2TvX743KYAq0OOQwZMdEGzEmDlrSD0/0m1++1
F+IYXOV44KqRuW9O0YILWDmPfmuA1SUYHBFQSYPT16K2qdurmzEdvHP2Jar110EOmj4jS4P8u7Z8
DcCQmCvKsQ5PsHyoiCBf3CAvfMBsLDlssiWdf6LRI6VAKUyo1YoO9dF5A+B8t8GStQljHkaeiPg1
8liadlf3Xdp5rlMNT0EjE1x6JxoJx5jQ9x8pgXMicmmGBHIrg5b0CD3qBOzzn7lLajAaIDl/H/z1
tcCP+8PgK9ZNzPEATrEmhoeLkMp2XSysaUFEmC5W5COzy22Rder9DnOZTaSXekRms0U4/yGA+R+0
ADSRpSqY+Vy+MYTVb3z/uTU06w025FNlvZ67La7J+kE7nKZURyLehbrjzc7pdu8qXPTdEE4l4vt7
JcksYCEAtlQZ62h22cEi+VtchxinalCo+Q6Gj+2N7uusuHacEXpGEZCwOgNrV8YOAu17b05PkZCZ
XNvieSVgj6JZUEuEgOYcMkmJKO2ZkAeRrIg865mq32hzb5Hy0hs54lxwfqCwe4qnsohUTWnPsqVZ
v7mg+W9EevmalWxq/swKEM/ODw2/HisgCAp/Rsg1XjgVZyIk9CX8T3KMWiuTkzY+GbHdXEmjgKlJ
mJCvpJ5DAzsTEEZqSm8/h4d1iPoKBBuR81g/bt1ZiHeJiFzw0UoUtn+M4/0XS4ozIhc0/u1UjIhB
I0xss7+ai44pmgEq/iJMDxkVIM+RZTVYIeeGwqtmbYjHtnVF1skNB8g1hckB3sTS+hNamocO5T2f
z6L5iz+y8jUvS1S6xa6cD5qSt/ijVIzz9UEQ8h17p3vMd+6Bgo7ZU1rCcPw2qmFAr3s9QzbOc8Nd
/+zc2A==
`protect end_protected
