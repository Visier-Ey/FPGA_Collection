-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "N-2017.12-SP2-4 -- Oct 23, 2018"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
BvajlZdGQbMyN1uEv0W2z9rUgL/+yiIclIIcqtfMIxCM1FHoHOYIA578LNAGF+ao
1IPEnPPWGEPOpOrLy3vmT/QcjURBxb+rw4dcDbZRFO1a6CNRdTOCuEnz2poMw+rU
l8ZZZ4RrHzSe9b0QVz6J4S6oxiEEEncDqPyNTe/IOos=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 24704)
`protect data_block
nfKREVa7Xe/Lingo3N6KtO37UgTZmckto1u9RU2IYS4Z2bPAkmOKSYbzZ4Zn0Hpe
mE6NGt72DCY+jR6/Dm7hhob4xV+TxhXqNGOgR5xO59y1fpJsouNXccClvwgz4ivn
+w2VQKY/z3LfPlTGV3xSVoY7uToikRjuJijt9wBKvnIQTuJP+VI832i5CDxdwkdx
Kd6WYORD5wdMicu1A7Zc5ow2W2SfeUD9LYjJHeEuUTCvljdVbVuD2R61LzQdHNkn
+tycCHi8nFmIofcAD7rlw5PGFiAzgiBFk1tGDOqgLq4d+n8FCNSl8jhC1Szg2ocS
Gk5gDhE+GoOAs6WLMHq/NwBNXNfSMMaLdIsM7Vp738nq8oUQbx0501fdcKayl7Gh
nKz1/p6nrf96+paw3M7lZnDoEPmDV+uuonh+1afdjz1HDk+stPHqXFetASALqnlX
WerqTVCXUbmyZqXlHed+3oCjWrxpyFmJpHRseDpkbw8VmsOWQbjy50ZFK0Taha/5
AzqUGWhEgnxspNwlbo2bsM7hCMNaSRVX0K2Hz895mFn7xcAztSzLUDyAlvcCXQkU
SxoG+OIv81n8R6EPryaMURfRD+bsa3Sk3ZPHjQwITA2AI02ho1CTRowyuQCjfL7p
KZX83mcqHwciJibP2nv3gThamJLlYciJo86G1HzTMZPe3SR6jpFmVk+H7IuEk5XQ
7c4BOhwY31z4zh4FgnjN+Nn+mYoVDGSB2EWCZeitgtFYmuhLO4/dvLVdegyKHoSe
lRS688+oX/NW3dSzJNOqHPylMXEuLbTdqg4rZwYxQ990iy8cl9l5sg38lrYgoPIF
RIpq2jbp6oI5IGs/Jee0oxZFUjanfzRm4oYdnLsONUjT22oc8NRHGuDJGYmZ8Pqg
T7zEyZzM5GrVUaamvq1o8QKt0NKsLSXUW+BAoABGiblE16tjgab5GQqRf8URyaWI
UdabK4oSRbsgRVieO8HWFztJV3pzfalSinlQvz9XnaEI1lFUq0oHkRLao0FHLf3c
b9XGBNEntUlrYTqH6zMYpXEczA4Wx62Rn6Y0Qm8dsntrNpg4uHq37fUGBuWL9f/Q
PbBrW4oTyqIwZaL9IN9Tjyl4b+AthEeJtzz+eUY4lOtR81oVno/D7GIEtRTeACKg
FqWn/1hTWjnWQKsrAmw1Mlr1Yd1L5hNH6sSEv/apd9Amdzmp/sj4cqvsXySm3n9O
A1xyrVIoaIFl+WGpW1C/caBe9dOFctsRN8+F6WSYCQNTNcXr+3elJ4DL3spC/QHy
r0v8VifXJZRNUGSr9UFzqYPlnd5td6zfoPv0shVP3gPJBe6XbishYATOOzCL+Now
NtOxxg37Wa5a+51OO7N6kk41suQEWugCj5jm4WLvidlnLz6LNVkRSPuQL8apPQCM
FaM3ZwLu2sAO9dxvMInkH88T0azvIl5/g7w9Kn0UDC8dEsgojcJgohqu7zzQo6ZI
N5Jnf93dPpMK86TRam23ydTL7uvXXOe39wE3RmLdQ9J/DAbRzLnQ8EohMgj0gcYz
hiyqjyzxQyzPNoe8OoDsz0jUrgMcWggCczbq9/3ZBpcFW/4YoExm04eelUHORiL7
v43e58Oxbgsi2lWPn7iRd2yNBgVKXm7IpNObKV5N4zA/1FS+TIybEptfQs4jMk9a
4jdP5rza7SZuOzHN1WdwAQzFJPKCVyPX+oyF/B5PfHuZOmEpK14Lwu0yT5BXpO7q
kHYubJJtmBNpbTht7s19Y6oUimNGHO1NqrS57MQbbW/dVEjifcpavjj1N7FEf6eI
5T24LPEFt3Jy4tCcAqwSMZZWl9SYWprrLz6VyJxvgrRsC2I8NDjzvnhkkZkU3CgG
hiLV5FGuiw4QPEfYNMciyisyOKGPKIxUGQlBGHDTryYBI85G4zqUX12knxSl7mZK
TzNnDKETFOHG12G5wZPIvyn9Od6uB6Q+oE3i2yRZ70Q13IgpGmyJ+sRzpUmP0RVq
6lOE4D7S3YpGbR3uDhIq1uqZXg7YiNeg8of1VnOWp2uHDda7hUgblYewkTaF/qOG
uX4GFcBcORM7Cr2LL8aK0tE70/q3m7BFwW48bEaiebeiFb3OlGhHTVsyklKtr/iE
TivJ159A6Iadt6pS0fwzHf9kZYOCsat2vNy4mJPiRBrDj9R2MtGfq7KQMIPN6wFR
s9uDj3DHXEjU8uO0c2gb5CBZcxj2mpKXViJ3soOjEtL+6y96bVzst90HvtqK2rFR
EKwmg8IhSILqN9EY/fqXfChW0V0blkBx2JB4bsjpgax0gDcWGdENVzvD8FC2t1Et
poqEixL/SXiAM1hc8QrJLGw/fheo8Ieb0HcswEY7X3Hogla44hZ5dIgxVFFkgNfC
YHtS7YqKbRYVPeGAYx30ziCAjSVdA89H7Behm8e8q7q71IS8SWOJRzN2/bvuNQlP
iwxL6s2fDBfkM/n9zw3AgJf5XJiWAUUmcApDKD15IIyhZzEDekxlMGb6Crxdr159
zNeLQ7Sa//sxLhJfylRG00evEsSs/5/tOix7U+xrUpBP8xuKua3kGvsByJ8dypHq
jvEF8NPN3QADg3BSYAKJnRb4DjxNT37xAWJZqhZsmFVDG3Hf8/vgLzx+bu02Wd+3
AdBcPaMxnTdXYgI3I2lUkcRLLIe4nvBXZBfZ3mLpd0lyQvHQt6ZkXCjYl4Bb0Z0+
W3NXIs1/l9ddIQ7XGF3XUrrsbnx2Yr/veY+o6PA2HvSp3QN6Xszy+3vCz1HpKaLD
+RUtMAQCzNz1P2KphILbxG/08DiVWsTUbqSLAF+y7kglH58Bt55yQTB85LdAVq9h
gZgsFyyU3qejTZwxx6zBpNtn/3rjFitE0KwbWmZL1h8R5RYLDidvuZbLa7Ls7x1C
9wdWE0mLVCNOGE9+WL/ND2z6HNDknzJ6mq5oqp7R1kejnx5WdMdnmGRsENAJFemk
Ru9QL/iU4LcfKCcV2FzL0OjVCfGiW23MaDrezTapkTX7sk7XwASeTY3kqrd0J4y4
p8b61xwQYL0aCX0MhH/3rv9WvHC8gFTaqdrQbJEU2vjJyg0OyAfxudpmGplr24T4
l6GVQeYUja36jpOF5ChX5QckuyK3+t9S93rR3/xLFG69wtBZOU+uJ0417tQ+PRan
miX2Q7mZCqGmOf5mYzL7de/A/c5+ncOHYG7ca9yizlTdPiwZsWqsr/U+iF/Nz/Wv
REDXePCwiQiHyCCfYI+uF49G1NcQNwSkb61P0a1843v3v2blKxp/BNJEdg0heAx2
GmLK3Y5frZGEkRxG5UAxoaDGyEA7Em8THm0fflwf0APvryri6RoftwF1DVp7ir9G
YCM6mZSu5+BWovKxQulCXFEIcBMKJx4U8XLOUWgeDCBKzBkxPjn/A9CsfTxsSGwm
w+5PehpP7xxrk1vWUm/G+/s2JfZFDXjhO6D+JPaUePluM5p3dWw3BhIIErLi0TBL
nNftOduz2j/PT0ExhGbty54iximGdcAkVkvK1aySnAHnbs4nfoHZA5qV6UxFHxFv
sIwgUsf4V+d+iEZllgz2pCdOt79V8RwDJCAsUfY810ThhrVkaGT67/RzQzanN4t4
xvn6ORZCBvRqXPHGU6MDToVayC6yqxlXW94wpqmwKZTmt7tOv1m/rjaRIJlGdhVm
YoeWRqJUIko3zjhPs+sMT8VSO4ord0Yrax1ap2KKtNciHnm8DEeKE0QagzBgVEqp
2v7Fi47A0Ofsu6isdtioOgvwEo6TfeBQUDMy25LybxJ0nPa+bTEG44qbcBmdzGKF
fa1gQpuYgs09wNnfFAyp5wf/jNnDQWsIx5YPt7LYDtDmz55b3K1gDYZWF6NtJ80B
T7shMsG5N6jBYeo5LZ3xiG2G4FJWuq5klBOzUw0vxJ43Cr1gEdAbmS3ePxM1iJNZ
plBOuF3GQaQGoHfMxd7MTtaUZpzIygurc5oK9JYSAcs9v1aJO6sr1pGVlF+PQpb4
uPgX19OxWXjpdu/9gTmNjOz11N3aB/GX3Ys9zoNKa4RiwK3PgjgaOpuO/ohRAA8A
sUDwePZG7aV49ahu+4KfqnR3ISwC55M30tcsb0BmQQ+p9tjokPT/qb4LQRN+f1I2
IUBIDVgjil6SJigM/Z6cMtKL8UtYpeX9pHsaiZLHRyHH3Ej3wnAGwNtChjgPwrUj
ia1RAi9TL+CT945gDAqm6OiiANWVrhoKEAf/p/trYPJrUP+OotCfc+8lmvrkrY16
4adsgK3dezUCo6087g0qc8Oyn/Vw5PTVtZuRSIHo6cciIuOiWA8n5+dzomjnnX42
CUOTY9eYlt2Q8EbDOYiOcm1+Qdzwu/1sbhLx8qTUgikndTJtzIePMis3p1n0w0k3
5+Z+Yx+Y1K+bGpFQ1CLSilhYpkLwBBNnNDHvG9eDVGyniLGu8xYAF76IP9MBe0gD
ASl+OPkWGmeXrCPYB0ALgN3F6M4PUMDCDX5e4tsi4Y/cBXV0niGYmM2IA+yucsRD
sg0j+sxAY8uWQyXb54hYzbMG+a+10gEmv6oXEjUpj3TXa4CfPwWqMBUcbg6w7Ke/
18fi0hQI3Qm7NvvnQnG8ojWKBUYxSmsu/hhFDnIGvBcQVqahLngHQM7/W5Q2PKb6
Z1/+i/P9Kuts1bPaOF5vKVoGecFqTfvC9oHu6Dq8gS3ZIXskeXCfei4R0lLfMelo
wAKIKjONhKtEOGBUrBpFjoMKlAG2jklg8CG05utCw1Z8Lqc1qTSJb9ihGgiPrF65
wVKBLURXjF3dcyijurc1WoiPyZrPkA8Yf686wRx/b/nkcl2II2V5pfiOkdKwQQoo
061nwAojtvTIrn1d+Mojmt+Elh1N7x2un3YQE4RKq15vqlk9ZSP22tawZAvLF9IE
rudnM5WwePN1QfZq+5Z0i/H401GYt7U0VZCL6i7FYtbSAOoSQsfN02OqAoClELtG
5v9S1qKLZe8wMy4lxGkGEse/L45lj9UjY06ZZe3sHQu5MCiba+3nhkj1YlcxEs0D
f7n7MVq39Az3XeJe8T1kNztK+Hb0ymQTFFxA3FPJyFLqtVGGmnb8yJfrM0tiO489
JolVY/989Ecfl1SnGIv9V8bEZrpEpgapaLBr4P4MaeAiNCpqjmnOkZbjRy5EXIVO
Bpzb8i/ug/5EZixrgQm3QA9YIVP+iXJI0vE0Dwnp8pfO16jf5ja0nSDVYLJDHmti
boFAvak0yMRRjFlPxgwgrIaeV73HKc4EqtTlKBE7leB2XegTwwfCW6NA0K/QaQr2
CEpdiSJV1TBymluuTAGaPMPkFT3yOP8QvXN4WF4qXWnv+fKXdIs8S12zmmpxlUq0
9t2pty2+Sv7UUl9xZL/fz3Et3fySMVGg5KK50qyUa00QCJIRjAI9/LRCNO6vymDi
IwnNwPBv9UHQRs/iyEI5n/wERB+barKNVpfxnTKLWbKaVClmJ0SG5cgwF7QFCj05
jhE4foS5RX1CSyIpeOGuKjQaWXpuzsysvFcfPuIyHLMDGFQ+wIZAtNUEXWmgVyn3
ZW1GUNcL/21aWkVJi7f4gD7WBfqbGR8bXHjQZYHJSIc5rFMPTCGLbwHznsUjgFm7
XvvnADiRZ4/h19EamR/VN9fzwoA2I7/V9VnVOCwSAWnRgSAf9CEltAXmMal0M3eD
IDof9QmmJ1K67J91dLdOP1KfdN7YnB5Pg4V6fE+VOCydYf1aipJ+155heg8T2Tds
XpBEXrQGd+bWy2p9mRbppvaugpGRHS+n6BbF9yim+NS+FOlT1EkKIvbxs+uG6Hy9
YDcTmAsBm+TEov059jMAKnjNpx1IqmHZKRF/3EV1X1VU9v3Tx9Yhf5pCCY3KGS2m
U6Cfo9RBJshKWgibiYjMQZhmp8xmaVGP4x4bK+1zNvzgpFr1Pni5OaHZexKc3s6t
BrdDOVJxFvIOcrLthK0Lfj+aMPbpe7AxCvLQeCZaXuhSesp5SDEMfDfEK/tCUBxb
UdteOhYWvCfKkqUWWzFrQX9sjtzNc3FVj2vwftSvD+oT3HReSx29MlRpISQzju7f
2ye8mXZL6+5r1F2IT7RDo09XZBM2+23AAXJCXNGMjNX3sy1TMbG77+hXyCnZ7pqg
QvqON+u1h2aH1zEE6I2BZWNxXbBMLWy1MxQFTGw+NK9hQRPyz7D/LGvfdWIGasjB
ZDQBCEd6fip/xAe5HI1P/ZR2ekOScCPfFtoD72S5veC+Z8k9GxLFf7yyt1Goj0eF
JnMObSE//6+mCt2seRQ/f0Dk6mneU6LhFqj6SMEWTFRzhMi5Tun0WUBCpan3b2ap
M1FQWdjtALrFkp/1H9dfOz3ltKY35OWcbsBPL6LA7L+MRPp/BBBMYr6piv10Hqfu
PMlkPhY2hY+ss3n3gVufOp0vmmNNyEJf7JiU4hMrNeXK8Ey2rEJI6fkcAyERQujI
+9etFIDXPQDfCbHN4UhoNRuLigQrfd+6UWXIXkeaCUE+9XOJCe05MI6G7drykldB
WdZ+rZaUq5xWhW3225ih/KfIByi6MCKSO8UJk2rrZk5LssBAHdkEeRrqqL0eUcSK
8LuW+C+49XVl2/6rbknpXIxdWEFTbqO9YyJQaBMu7+gqqgSfZKMqHCkD8ORAGem7
X2RFzu8gQWNoYzAR1VDajQrGvyUR/djr7hCTJL2YbFKreWzFRCAkI9w1Outa2lDp
CjzG6HYJja8i6PJKd9r4e/5TGqXZTi78DJPSod/K3Y9qOv10jiu7EOVu/eRKVMGQ
dRZN9nwcOiUto14owKub7aA12Crue6jYRYXSj3sx8X0mwzeZYWBm6rPUr1QRWBo3
FrJx/MKYzoOjfLe8CvtOO8RwSxvR5c8QfNk/hC50+Wzv6goRivSx+gzI5xg9wHRm
Nr8/Tg60NUJvOIpGU7z0F04h+VEN+2ld9qahhXKmu3JIYU+mNZQtQpaPOmRf0FI2
IwXkDMH1QKBIVdxzRsyNZDXGIy9v8Y5J2n/7RxwWpHer750PNN171TJ/3eDAvaCh
O90S1oPqqlSaAvQiE4HVHoXrFOr/Jaxru+dYPDP4OrEoeVxxo6WYvL9qKK/o+Wrv
XP9Ut25rgpl1Lauso9AxqLniqOjJlcK7TXGuhQVMGUoVgKk3QwqTIHC5uyXvtqxO
cH7m/b2RBUTL3AGzUw11mj8XkxzC/lF56U1iaR68v0+aoqmumvB68woahJnzj4No
hzKs+WPISpWU7pesmvo9txDXpr5BmIFInkZmckbbshaxDpkvNl9pXJE7wEAXjp1A
xKxSvr5oNbkj/2E5ar2mv7ip1b8LiqmZQGc0Wy14zjceZuf3zXVBdLnnVGmrjFsR
mSWZImDsrBMsIxmo+e4hzkFBJJ2flzCSR7RV87iTTSIE1/l9w2NMMfQhdk3ia2TJ
KtoltsQ127sy2q2ieFhtVrg8KnEWHBGy35wlaIhu70OK7ZtVMPpEMPA14pRYjUVZ
3BuoXjWaTnZbsK62Niixv5pywRXGruptrIugxcD7Lj6iB47I2d9qDShQrlzyu/Qc
FX87Cvh8q8/wkQvtDtN3T1PLb5fZVc8O0iHUDZseoAKJkFSLHQX0wbz6+3tGH2bv
GaYjejl+Ifm+dibkGrd9GEPkKfiGHk6PuaS5iJbGfOrxWU4fOQvCOZ6n0XK5MGm7
/jDwBw2+c6n3xK3mh+w4phjD441KXApoEqVt1Cbf2eWQy2PnxcNuvXDZsmLNxvLf
YC+JjM0XMOVDM7FgRs7i0C7JWLj7KuIEx2iij0awr/VJLDxNqOxD7GXO9FFMvISN
iFYeZZtCezr49dCN0ZLQR0MbGW26XdJqOJ+OKJIe+zuzqXZ+xHliY0B0eHqmTRXo
6TrMXNMWmSQ1cKKmxlqe4VbrT+ZPQYVhPnN1L00ClC0xFry0r3Q59CxNc1V6futE
jEuVGb1TaHjgxi6/Vjxh+xpBTOBsR4PGo9VEjzmn1NpQmj5b6rswf8kDVT782mvg
orOlGcqHs41jbU0N/NxkfMwaHFdBFNfrPZi1/hjc3HQO0dHb9+aXGazvcygZa4KT
MeT6hobKvLXaENY4neTIkE0nGXE91lFUPjO6AEiINTkFRfUlrULdOYiK3dzCFxVh
vAwH9yJKa0JBV2rfyY6RbZgd3qWIEdZQ7LwBF9pxmtCf/IJbreAdIWwBr4MQ83qu
D9sbxZzqzmN+Ere6zsfwoYqkLJy3bJJrBk0uc7mm7+KmbDnG+yJF9hi9b0fUKxPf
inE9QB+/1W+ZiPL9FRrn0YSB43TX3H9lIDjT9isVtapBOqMMSm0IVmf2s3kKoc+q
17AofrfL+lm++bOFzAvFjYxqDQxaBqzhjy06ZpebG497SAmwTZjwcXhx/WdgLb6A
+Dl1eafLo0nMU3xPfs7Ms5Pi9c/un6aaBaEt55MHb2PCeUS8UZmALjv+hRma5g/o
vf4JZ3VWmUZwYYmVMYXpA8IeSf17xBB+ck8zOiIHXL9Lu2yFEe+cd8ryy+h9rcPx
Dl4CN0/t+++aoEmEFJ5pNhBNtR5AXfmneDj+zN9AmznNo+IKRNljjMOj6M2S0hV+
jo0JHCAA5MTKVd9Fdb3JRUvMUjjaP7DuZttV9dQuqTIQZKajXjnOy3vPhLa1BVIp
9WRjFa6i5F+gdQ2fCRq06glgGXheYN2goqe1o/5fUM4fYW/DrYbZ0k1ivQRU79tq
NC4Z93CCsJg2hIP4ItTQWlsTguNuIfbTN96xfD4FL/rrCOwD+LVlBNn7KV4F1XTo
qlkum/vwJB1VXbliWT9b2StHRITrBP2mAZRvWm8OC4asav5ZwAxXOSDTmisu/ngG
8yvzm9EL5m+CRVyBodzi9+3vfmwVC3dHM0rQR8Ny+Idd1Co/OMeATxFwfkngX/EG
7GM38/pM8Tzq/tDfO1mxpD6eA2ugqNykCQImz8H4BXxdpvtJoKxHJZpYd5MOrPxv
i1aMizzqOkzhfmiA/sKS+XkHZGmEyQXaQyS5gHP+eCtmGpPFSJLUyWNzNmm0QF8/
r9b81zyd9t87mJwFA7fVyMrN/5VHpNB4M2DvBWVpW9FNRT6bMjtBfpOIxwuc3fuh
NPRQKG51yQfLgYQOL8JjxXMQIXUgAPzYpzQjl0HaIMhv0o+eKT4ntOWS4dhhG1qe
cWlQyL3DWhdweX+ldw+ZqCu2gS5TVMb9fj49o+TjdyGHKF5r4GvuBqtbi3khtnD8
jUlz9ksVKGcLNUZzwo6lQSPtzi3M5UppL7bl1zEcKH0LNbTukgh4sILf0aH1N3Eh
m7PEqw9b37/Et5Z5jfFzdba/X+wUqot9Y4Q0ztAFHWxgwB2MbAG/FdhJAsiheA9I
egtJaNPbkG9xVraFSzJaT/077fu9T13elJdZF5KmCZGCRbaYNiGJMDN3bf/GPdqY
DeAaTpfbHqLNkGX9ufIxrJd8GJvcyX4zpIORTUPM5AVv5+pmRW8kBlMPZ8GbY0o7
WOw3lJiznvYTZxMiBiWe1xXBYugeSLeaKttBIMV16zlb1ZpkPXmafLY0kjiz+2BQ
eMi0erQ9B6CVNTut51MqwtxJnMGgQ0HE20IgS5cFFZ+tcMHR5AwqkCE6adIJj/OA
zNnV3Xxz87MQwRx6pDXWlOX/JPguHD71hHs+3xSc6zxyy/ILiyfNRfxdZcZ4RIrK
zhDYqa+R/pe8v4+jrQ3DuH0wgdnveT8dNzffZDfEJhdIGFp+p48u66J96OkOmH91
jb6Mw3WM+l9CfQGR1Ya4GqRLKuovxYV7+F46zUyXK+ANyx2gzusLMRGjcJAzH2jf
EmCetGdwQTbjM1UbrJObm3ReonN1ahIro1jWaUzL3V/URjpvpz5hiOVKF1bGeFy3
w4pre5N7pgmEM4kpufE0Hv35kzaPSmmLEPfJEyT7cH9heqhgV0cNi9oyKPYgoXoO
8R4neYnTG1sbPtHMS0nyNJFmLVPKRDnrksEOPBUnp2rblp//KEGDbiGxuCa54rdB
Kevw9nNy7/pdPMYOUMH3vHWVoXITsbCmQ3vvpxYszJfwSaLKUgQCecIHKdqTpPMK
Fz0KwEvrUwAPP84IVZgzh9x1Sbh8aMa4H1rIFLlPnoUNkrIUVumEW1s7S/6Tipms
djKXjtVyoaysGzCiKoYDxUUdYjcDmb2kjiKqR1jWl1LUYjHqEE+T/xg0p4MAbN3J
qT3FUJNZm2ZsQRS0FxxHGPXh7g6ivMGTLbJk/1RLHBmD6RuyJ40USdq4NtegOThd
QTvj2rXg06Mb0DiSiKT59Z+9xQMm26ogLQRO8af9PD15LOPMvJaccJrDrdUV+PuA
zcwNF16G4GwA+e4z+JcJ9Uz9Gvu4eMlZ1DRDnOLD7MRQrTGUQIOxrdhhU/8xEcs6
whLQ+uyfifO1mDNh3YNOqH51x/RGTXxHs7bGBGY56darAQv18ri6jeHKxz0blcvm
65oFwyf84kui5e+sTe8+LPNU6HCIEGgpg1d9Nx2hDbwQwkhns32FEWWZEVziQI5w
M5D39JGtNQjCt3Hzp9NjcR8DefxxWteiakQoopkYn/kkxqeNEpSNyA5buSA7fj2R
/DOB4onyvr3LqvTTYymr1LACFiApvUCLiRp0o/I6KUQjfkjZrLOBishflvKUl8bN
LLYU7WSImOQgd86InQh0p8dX03Uww11sivQ1bHIeX7Qrd+n2g3s2YRWgprGxmL6p
/sBzYGyHM/+1KJaH4MFgrSF88xtl6F/Kwr66i15fS239JVl+DsmJ0+ByJUKXqOc5
LLmkY68hQbvsVtNFSPuQjlYixWTJDYJbnhAHadvFmKVGCNRJbtvfZbR71ON1fO6Y
rx50LpzwNO+GgmgmKWsOs3UyOKkLc9GQExH4Ey571h2paWPTDXsxNsUIqD4HZKLU
7wKD1ghuAOl2B3lpvR6m/vJ7Wxt5u1cqeR0ZJ6HVrOv67s7nH/Fy7Tck+a+YSRUf
5yvVb+bdn8mjuE+nzpP1ZQ9/snYRxN8cY7vvM9hWj/a6hVhtXuDCFMBrT/5r8brM
oDKoEY/eZat3RtUAKT/CR5RvvOJfbaexmG2RBVoKRlPPU9mkKyaJCNOfakNiKjsN
nV5B/u4R3y2y0xwhmH7uQeib+AzfZ3/VmBZUem5HvEF2pqUu5Sc/XVPhaA5dDH7l
se0/DPYQgPpacQb9TUSvm42iIROTOcYxyW2VlmKss86A/PelUxofBWqT3Z2HkYhE
lqoTMd09MLU79jz3Igz9I+9jDFNFA6mYSOoAy/p7fhmdQfFCfIuslLY04WS8l+Ux
PtYLwowMrqJ64sdA7lSBLSUeaq37tRFA77q2+hK6HriteUx0fj5lKRQSq6Utt/3o
auqX29pIwNWdY8ZVVvivemhC/TbfAoj26+Xvf9ltqFmXZsl93idNOtQ6QY40pZqa
bmDz1EvrlkezsFZyzWgdyGHCsZIs6NMMCPxP/rfdjkY3HN81KsbOEV+6vuKIPzZ/
A5NGOzAZOqwgbukijX0LeRDxHL946HkJ686b1duDcxb8TdbELrMi3pVDX0WJkVdg
X/byQoYrR3lc24uXuTktqUltFiawBWhgnjrHSvShGO1fYtSAYQgLC+MSlw0HM8i9
cqRZO1qmVfSFuoylyX4ryHmKggEv8uyUIucFpLaU02zZTo2MzT2YafpvfMH9kNvl
x0gbXyyN9N/VVLzkmrHw63Oy1krBFBlEANnbgHCdl5yNZyqaDJy7/eIGJ8VrFv7E
gS7ZbEVq+8qtvSloe+fScdO7f9nV+2+ackn3pfmPSaP2AmDoaMR/0huh02a9FlFq
kdr/s9X2ILW6LdimB+aTOsKpGZbGD74RJdtwMZrs6sIGxsHw5TbmGGH1C0quHkMw
9ZRITbBAs6InItelz5qYJxmnMQeIspWTnSyw9l5BmIhGPjUkAXgnWf4oLRX5+R8/
KT1jgWBYxetNKX+j/d+FG8xUVhMb6bXO43hbltO5OxIsJ5/2igd7CXCeUUaUUZZk
TNwCoVRu0zjsywtZ9f8Axc6UtRKvRMbjs/ooo0PS7HGst5Qh6P2uP2BfTuoimqZk
PAUNTaKWZcTz8E5jEZWAzI2vfIySjDIrURYS5/nAkf0veN4NGXXzeKgn5qEo2crt
o+pLTpmZuplOj3BSuZHeX+dd15kLvVtyskwuq5hfNQ2q+9yX7if2WDQqWUnFAm7h
XlPKIgAIDeJEPpDDTrHaS6txDAvmQtlBsk1UB1t1MgXrJLp5qJXmxvQbKT2CBb9C
pC/az3TWl+AQbY+tsiOHQQdHRLggaARWYSBVoee/2wDWmKdiirk3853neNOwGUSV
WFE7/3LgsJ/raUoDJFKJesfTowrPRrx5Sb/M57JiGJ8N5j5ceTw5vuxDTBCPJtfw
mWMEXsYjMqey4wzSlPZUXEaJYOxLn0Z29lQKKxdYm2LEMEcHW7ZAm3xNjXRxnWm5
IEhxHAVCJ+coy1LxQb8jX3ltzb1UqAzZRVOl2cYh3aUDFLoQzN4zM020H5lQremW
ypsqkUG3Z7F1ddMHOlnGpD+plyhSzdE6vMOYpRzIWbvKe+4iJQTGEvPpr4MKMhL7
QL490EbASI9mEEsf1kbf6HuHS9jHq9W5p5ISN+EzmON1dvrMHLvUxCGX4bSiO8gv
p1xtIC9th0dJ+szyo1oOLsDpqGSIEsWk43nEvj9Nw3ifvWkEZ3l9v3LWzcOgTsbo
lYOIRs1Infw+wjWJ3hWCiX53zAXASGrIpdKujpDtwGldnMhRTq7Jitf4Fx6eBvF6
RvQ+F726lVoe8lloqmLGdS3LPpgp73OCP8Qh68e8UdbtRALVuVxVA65Cnc7EW5Dh
c11pdr6dKl3GtQv8gtZa83zlHM8Eczm0x21L/ANbX+D02z8j3OfqB+jARBxdXb/z
IsWwjkOYH84MYc8ZoRiVOyiZ7rgSm92gp4HMaOiUki26UF4BCNY+rAlrDK0qDRgk
UQK7kQm/W4DvVq5pXz6gPGNIwd1NKld7MN9sxHXHzQVBKeoPo1t98gQCqYvtndp7
ny9++0bMYFiSkrdJVbm3JMCWoFjjFVYs5ZrsYVN8Gy41SuL8Q9rBlM1wS1i3mM1N
e1ia+xwonWkMhcgCXSkGv3f3kkxKsOExgzHFK7pjfxE1g0FniXhLax8VctqoZ75N
wfws77oCOa8Q2Epj2yOvFaoc0g493G6eNNCJGk852QyyeKw1K9/ivcyZjvf0BwK7
p+e2IFS5d0WXCtcrlXubyQL5x9jjeJRE0bXkfTCRVVLOxUuC7Uo50rX0pX7aDCRf
eULMumzhhVQNgxlZR/5Lgw6Swf91Yj6IbL2gi8mcu7ZmnancKyjjtfaixmgnz/XL
7qOMNQAKt66dNMtdMhC4pvNgSZhy0ThfkrU4GmoKtZHAgeXIOuOGDgW2sklkbBHs
iXprc/j4cgx23n43kF2HFU8eEreDJNwnWFvDvToEe9Elc7u/MVmTzKpOgpnkZ/+q
wX4ko7Qbbs8pS797EtyeXduuwltXduEwwt7UtIAujmY9CS0iH4H7Qr8Y5NXtaMgD
xLE61d1As11QNFsa4PtiUG2XsNRHTaerrd5v328OAI4hgmc2xeqgMRDXihjO9drj
chFNJHxvvPlCMmJLO88A7sYVs5Lvh30n0lxz5lc4F/G4tzBk1YeYMwp+Bk/m21nR
jYCF49jWAg4bWgFhJvQbEtrS1UPdMx41GB8Zl7WsUmrUtnMs0/f2aW/Ju/Pp3BXA
IgNkzxdkGoEj7pPflQXlgLQXVr3V5xkA3slnMEFuMrQWMbu/b/nN0zcxDQ/l1E4m
ihPxTWIKF9YUFLlIb9kl4usjMfa8ErfKFSoc4NdGXbQ6Hxys32fnHGx5cjaX4mBe
nflwzSoFNC3hDrZjkwdMuTr7fOmwmukIMGzaTnr0seDrjnBt9IAfUxXFv2FaNDU9
7KwkVuLNr8RMG1Fz/t2/3LDpM5rZ1QC9TolFuzBaqm48emq5BmMyviBvku59KeMV
8DYclHzDgdUr5Bn7N8Pw3R2zsuAVnfrnPOAtnnjxmn547wwuSNuZhj4mmmrHbLyx
0Np/vtC4lP6FcNTUUi48lS70j1ZikW3O734CAgi96s1hvpfjx8LBQyfkjyxx0M46
CEg/7KXleb4Rmo5clNX73SztbmsScaL+MoJ3mwwqKStKCCzxz1QoJYuhL1jI5HVj
J1+7ml3Liu+6MEgG/PsCF9+JmyiaerIYCZ273yYJPF5Ow+i/VSdgFQJ1pTveAyD2
4Wkji/1HfedWjI5aeO7FsZRdpprrFjxKdJYLv43L4MbcaxRUbJLSgWapcIX2JHot
LenBklcdRzfBu07pqgPNYZlwTLCSJ8j4JhgEVi7Ft5Oo7B+OtpiuWd0vfosw20x8
Wjosrz3/16cwHnGEzjgZM1MZ5WXzXSa0GPxuHfR4KfFheM1hKQw8zz4nk/6iORO6
gZ77TRCo8gifOFsT0M0gxzzZQpsHBYVWYvIIlHi/WWpxEASEZqXC59f0yreYmhfs
bI1Re4b3En76hrYR6nxav2mCsmsMIvLen8mIe9/IU2mVFvJ1BBjNs1HA4qzZ7jzd
bcrtZxVJHguy5p0Cif9CdBOUCCAncSKTCL4JyjLgYvNjxjZNN/i+QUx40sy59/ku
HEj2zq87i1WIPjVSkyTc2trmV2cNmHOqsbDAzPklzgsZXBgoGbFX+px2bB4U3N2G
t/zIeEzsS6TyJKatNFwsEl9PquyjWAYfHzcuoWftXu0tUrE9e8qcoiqJxfnEkV+v
XnWoHoG6rUhOLly7qYgitfTGv/UlhD9jEeY3x5akHKgkhHJt3sptLrD3kQjwujiW
Nrhbvx6yh/cyLm+QX4zVr6XTwMqXmUYP6sKYyq9M4LrV5Z5N9W8SM3ldDwCEvPUi
7QZzRYqBFfN3oHvBlO9jDdlxOCPpkuSmIC8IVoPcKJf3CBHNKtdZ/VmZMvPC5TVZ
RFp9rBoxqNzHFIxoFUXY0Ds+lwB/77o8JHyCws1pcIqr4hCnf/w6qxmU3uDbDMdP
oMnViYrvPEZmzTo4frTJa5jbSQDTQakY7/5DBCAwoivI9qRZ+kexPAkZ3PqyGPmO
x4hXd7JFT6Ff7dVKUMPb5cXrJvo0MyEguA3myX8zTgD2p2BoZfg9+YKWn7TeG7GM
TZYVGmgnnOqBDAXpWpXYPP8gUyDI6Ac2uRq06G7M+0BF89atURFUxeCFwOfX8Wkz
mwwlpL3ugGg6fJqK494OSrETMPvOagMsMyBMDukmQLz9M3wSOznzo4RuodX9OZ52
KhRMFcyKYJoS+CSP46KZUEtnjM/1XW3etD0kHU48KvovkX0GqL+iSBrIZWhE6aTX
td0V8Kdu3yie/jv792FCme/RoKVE0087VoTCAhtO3MqanvMfi1ZbiCnVos21MclF
I0JBapsVnOQPTe3HP1T7ItU14uxHEti+fIuEs1cgi05WUl5RnKH+3nznPN0ceTnN
VqRFQnnRnXLxSbNTD6iZFT5TSgas88ajyCgHmFshNKuwfyLEHScQsiKTAn6inuA9
eTuPsyinjs4yrBqnFtFyhpUj0M6hhNRfYyRhNv0TUZ76NZoLCKoLaEap1oCJzmGB
gmStVdBcCuf+KOvpM4SmG2D6V8TFszzPvCxNUXFJeiRbH1RYncesmEocQq5ZWig7
RH9+HM4WmMHIyybd2FVLHfTpRRfunqRe2EwYGfXC6uNpDpHUa6pZHClu6jvbV0iC
4y6ku4Z2ancIKUN2Mkt+Vc9iw7hGYekO5jQxziD2SSzHrHOBW7JRhFxz2L4MgXpV
JwGYC85DvsawDHhu1x0lzGqdo986dGVl8S3VwN7imqu3QftrEEiQxCWeZBybcC1X
4eIxhzeLbj67Z98D21GUwDhKY344dUaF7TTZvi7A5/zmi9cMsY+FJ/Ma7PsenzeS
dG5THOOt4e7FPWUDk8Vhkn/FyEfo8RnI867nViPikxDHNG+He2O3rYuyJL1pO3oH
pmnV05p374GyhPuTvMEC/0dOkNhjebM8wn3XFZ3HagTWmZA2qAe08VsxR+wEieU5
xJGu44bJZ0UCv3LAB5otWqQzrMbmqq0At6cQURwme6FL8miLYkjDJNzbzCYmqc3H
fuCEeGL93PMUVPTXUMjLhRYTIgS3c7Fqnyakhnegi1q8Ls+ScaOSoO43rUSXrdkZ
ek92bkA2BHmsW4tZk8ph9DhdiqAqW/9aUJU95WqhV9/NGNHUynYyoMg3gNIqo1IP
aXht687rUZ6trcUzHenXV5TV+SIwjxSq2+We5H8T+1nuU7KI6SejXSSwGOqqctQZ
Xof3QXMlc3JvWXNrJoGgwcbMwkgSD8aqpRaRdbs5meyh9lP3O0tiPnqJsLUDkOJ9
9Vl689SKEJbseYGD0p/tStQteyKMAGr4g6cGclhBLdEuh46pXH+PMdptcy5xXZst
vvKeP+LhASVzb5Fa2IgUQU9fr1XhbyFn7IOteo8NHnGDQeDbvPy0m9pslpDhtMbo
AQGxjJI9rttPDuxgQNX5cH6UV21/7VKoYZhsrJlPWs/LXF0RQdU3dbG/oT4dYW8n
NsLdnT1g7jpv2/7a3mtgKNJn32kgEQNdc6zvmIXr44uWFU6mZ7X92TWKvHvI20IT
GtIB/vDPKBCrhdnlG16LlsR1+d1zgoJCxBPhe5xDz+1oqPFGjOmoHS29Y2zq/Sid
ac9yELBAOa1zuVCf9oIBnSAVDBqil6BXeaPRTmRVRnwyQ2YQyG6kk8kQ86AYWy+V
LkNzm8lmhYym/ZnRJOhSeExHnio66yi/kGHg36r8EmTchSrLGfEhlKg+/CYNBKgB
MNN4tGc+qjDBALmCOc4a19SUyCDxpk5SerQxjyCC/CWLygjmZZvVtGh+aW0jPT90
iNZsqNnNAFaeCJG6FHe8sqFoCU4RTCcoX2h9FhB5kE2oxVYz88b6ZDRu/B4qYq80
4j6OHYpgnExohrAPKub3IE9Exv3Yq59AOtDuqMP2PMZruFilLh67IEGEiry5h7d6
E7Xp6x80I3ssxfrrMxNKctCaABhxXppiBZLirTXv9OMp9ojmFBmRzLC8spr+q3zP
0ZleYzhfVVbA2+uzLo1IWVvyZMU4AZq5Ig6Zqyue4n7zQb4X/H4vl/k4mRjXRh8a
jYdWaqdoEqTOK4cYCFW9XqTKJXqI1xGtdo5W3ZP2T3lxmvSb6HCRqBU4qISz58Rw
jfN4eVQr+YyO0JMlcYjl42lJxO8zmjYZhVoSKptS3Wgo287xWh/ABFl+Rz1dUOrR
8JP2KHsM2uVN9KIWMGHIxPDS1IUxx56cEaZL2vx4gMFLsZOJN0wYaiguyNJpeTFm
Uiiq4QdlVb1qDw3JRGedV3fftTL+BIKDKKJigeXM1o7RqoI4vqKYLh8FvyAZy4SW
yTyAxxB429WAL/lRzrha90B1mztI44Di97GKDrAISO0oBdK2fjQR/2lGc+RDdmvR
83eI0Vao1r5RSoM6I1PyiXXzQhtUDJsFbn8K995gVPKaeiwBygL8affabI4CFTwW
5MFZyG72ap1t1cXGbCrNEpicpvvQ9vVzyJBGeyJfw9lS1uuPpUgDgjsXvL60KKr0
CktzsdWrPaJ0olb1yVMf50peK15Ea/VhEFHlfQwMmsi3ag6KfGBYDGolx7ChOu+G
Vgs6RIXkEMJWZKHKvBPHDj4r6o6n0H+4P/NEHtl+l5xNIheyG+7lOYtL7sL7qRBC
ZBQNsF1mWk32FGv8UdInRmZN5pF+cfudwkhNKatSuPUFsk57J0CMwwYq/ldtm98e
k3SsIpnAiE2eCPHTEzVUhMw0qL/KfMzLvPJHrzMy92CsE1CJNxwRFqcptACMCs88
EB1PzNWJKrlyT05v9kCSOOhz3jyya0L8ROViuyhzsWIdsR+T59qzDbMJanL0slAi
/8pMdJCZQDG2/PtDADD+JxvYhkrZ+HIPr5ul2Nciuy2+hL/X5rmyerpTYNZvhZf9
qHyXr8w992wGhWZFt10dolfX2jO8LULOHtjzJtEjqfdZRBL52QAq6BT7AStzGnw1
T+2zYXQ5xxDZVLEsZCb065p9o5tiqwFtKQfFRHyhZ8hRtH1Ddx5+3uqASSArPUAQ
OlvqTTRIXKurKlg6UVNW2Z7CqibKP43sRtMOsyTvEd5V1cGKZT58tCV3Ui+TMydR
4OS7pIR9EVqCQgisHl7SCgMDV4Ohui6sYW0k2Nk7xfkHbyoqeY0kPKEmGIt2lpBf
0UPLv2mWK4PCYeto9nOtXbHmlK0sJ1s5YIV+lmxGfL8puJAy5ONGs+4ONlwjp2nq
2pa/HrX7FDnrD5YYjsKZ8ZbYLvvKhzqf7vfUqQH/Z7kqcV8EsGYUEF4m0TcP0uWJ
pL57uDeVEqQU/vnD5uDR7xzNoUKnJTekHVtg+9mxjlXh7KC9DjG5qo4rNnnFp4Tw
X80bJdOHweXyznBCwwVEUCJRm3F4sQ/BzQDS4FxPJ40FREoqiu1S4rItRmq5OG+G
70tZpiCF89Vf6sNUJIWYl9JACcg8XUPVitjv+viB3/dmfFcCDWNURQGDiffgMxRD
fV/XmltorNu8cKubsD3ao+TUGkZ+yzPI7yaOMq5vwRIfJzi5MsssYiqWVB5gebpT
3WmO8Nr0VZMBYNkZI+krECgg2RHXmy26OOPtGBsgvMRtCv5E03qDO5ZdfhN7xI7a
tj1dqob0J+lmDEM9RkJD5jQhgUZbYjjP1rWk6Cn071139X2H2MFp7tTszKlYVM21
1+xY5p4OZ7RcxZ4/q2uqbO70pVJMwpH5hcM3okJOVl8TQS7/HgEh0DOVquj8MX/D
SKtr/PGhCNo9cYQOLP7yl2RpfdoCQROJbKQwpOrx/OjI4ENt8NsNzGwZuaLPTXXh
ETgVdQyWz41Zr9sd1dCoAm+c4ZqSSdcWCuA6vQwj+o1iFzZ4kA6VApCtrzbGn9TY
XM+Ttw5Bs3q1FYBxj9wlMpf38pWwzP6ljny3EaCb/PUEWjidOgYYQ3wvxnTDHuP4
bAEe+QkxlIya9ZOVatr2ScZ/4iIL5Lv8Hun+hw8GXh3AGEqgyjMhcgS6jn4tNSqV
4nTvfWgy6AuArfcjQAkqpx+axowJ9CXFHAokiiW32YxqydDyzFnlXKgZUyPVTopH
NNsYcz2wz66m+LtAv5iKqsnIIsfvL+khpTxcESexNfsbViz7oDvoczeeO83dvT9P
P3x9kUUzWCesTnwDHc0PLP/WeSJN/A4e6lB7kkD9WzglCbi0XQ1icRqK5lGxKuti
WndWSSpKbJV9MX5VaeE/buqNOF9NbkHeEUoKhP3ryeTAwmJr3Y7K7PP3FU7GKdlR
OT9KdeMZ339HZfBdrO8/WXI4hs5Mq+nWRDvcz0mi2HhfS9MEqczkrOj6S/7ruwWH
/tRZVMJ9YngzWzHDJCZLHou9SlMgwTUerZ3DabOTR3wdN67Rvgxf9FZxUQZmA4dP
Ne/BEPIenhHMOwfJoNcXEuur5XJjWTXAryB0fIIx3y4ojSfIM21jTDz9SEmgzpmg
AqJjN5MiMrkB9YIfB9N2PNTuVFF9/pZkndfpzodhOnNzJo8S2Roi/5t+2Z+sTTmZ
lE8WWsUe6bkROhR0YKt7WsktwuyuHkhUY6nUhSTjUbcmvHA9XTBEo7Vr6VW4kQlA
JLXR2+K0aSFMotmY+ADmassRfkYRbxrV4V9IhKUHPrOs0ZdgQi3AuJzJWet9noGi
AuvACj5uldNUQb0NYDKRNUkyaRBNmk4f95lkLeSzYSoWOKvgeb2npO73O2Fq8cG9
khtIQR/8+l8eLbiCljKImtyebjKc93Ss0kDKgk0q9TaWJQkVTvU9zjb1TCFoqCb9
V63b7xLZ7Oy8bivmUdVza6xonFIfLp7wfFSQ9kMe+TxNgb9u+/9g3ESl8bjU74fv
ZV8WiHrFvShuN3KSyGVLEvHOPF5mHRNzcvjWhN/ld5IfdQrEUCzClZdzPexUhkCD
IyDj3FUNDZn74FC4phX+9euV1TjJ/Sy8l7F/bebV21pKT04Md0AAshdJMdV38KIg
fgwU/BjqBfw2aUkrj4J5m5BDxBA9zLbd+w1HiIcHqcjkRsW/l0R/ivexOfm5ItQq
W4ergmOeGUQfaYZf1FIYJFrKMG3gOg1wy5ocuY6ZXL+bWIdgHjsL+vl1pg+5/4wE
8znh4mqyvWy0w56zo8RAVDPlt/xzk2pyBolMZPEBzAAYZSuPKsonN3wViOGM4YP2
KcVD/X7srud/PY7AT/KJKym4+M0e6CWQ9y49eHTGCRRR7RTzCCaApzpqMtkBWnzs
kHZxexCmH1AkY04xp4VUPCbYH9TFEawPQ2mioycgw6H2pUUQKr7uURo4A9D5Sy/0
QOhUBXp2pp0yA1ikNayigJjCsuoO1dSsfcwfX5LwkXqWgsLzcNprpdwoDqS+GMEX
/vxvKZOxEVfP8KoOmed6AD5eQxvhUJKId78eB0xCLLapBONK2pIdckhqA/TF6mKC
VPyT/uJmrfBVDr1V0iqvEHWjY4dTqocSdOKbW+eYteH2JJ2NuXn3QveuoPJ4AKK5
T4QL66BN8EEjaPBIm99DT5DCeVY4zczSjUPRe0cd4YDnIY5TBCXShIIyEQgcI2Bp
2NqKHP8/vXZ5PaEEVdBdNPC1XychRDpSBoNb4XVPFZvZGY01neGx0zSBToQJMh5c
76m6tCgNCHRo9qIrsSlwiAPP7XxshswHxoQ/OREIbNHzOZcRtEXTUcIWoRSkQrox
E8EPuEOwFYQr5fRId9OHHgiEs/eU4aozu46rQPh9ejEtqkzqGfjAKDmPnLLCnFOL
XXDplTYpzgZKm87kxrDlJ+ZkuRuJIsEm1ESYeIPjoCWi8UiABD4z2fq5q6ygGjD7
bbrIW6NR4iTW8fyWXNZOniNfpUk/FbEUCNOV4m+oSaf08cWG6a1eD3AlrhpAjF2+
kARRVx8JXnuhsMJ4as15Lliroegk0yt768Kdhhu/g50NH6sUi5fA598lJIgzN8D2
P7EfQVvK9+aUDotIErJA0TfW4q7zL+XRoCkNCZrTBPIgxUZlbktsMamz+DoLdn5A
OyWnAdKC5STHHmL02FEUZc0+QiMwl2Wg/tbV6gk6vh1YKL1MZRE1pdvbicSHMskp
iWvFns46tHQtnG9Z/P38I/TrRfae8UZXeza+hxtX7yw7NK99uarLSs5Dk3tP5L2H
w/36rf7f9J36hGl28z8wJMunP9Z2MpXyLVD1ZzfgXyiJ4fX14RSOo6V2MzldeGok
Se/mY+yT8E0NqGELG7Q1jQNPnThPWJCBaAMUMpx6otHcyTBCf5z+wYsSr4j9hMXr
0fTou01zFV6CICeu9oM5+maBqcT2daOaNNAMRp4BEN6pMu1e3DWqSuUnGkG+aGjl
9xS+uxVtdeAU24nHzCZmHziJUXQ/sKeXYFReeoUt/HIiS7cQL8LqTyTo/wsl73sU
BzFCPOrujNIy3+JqCbT5aAVQxcEeXcSJiWE+mBjlziJZ9CZX/thp8DckmIZ+9JeF
g4TqLOTu+JgdHXE5Ck9eKW1n0V962YV4vqWEVcxZZWsL+r+sfeDgxVv4/gXPJ9qy
RGWyWnl2Kdl/kUKgvhr1E8N8eaAGHq+PV0cbnfZFA/28oM6FhPozU10iyWBfSkLE
1m/y1O91zNYpQ4jiDbwsVlWQrbMaZMOa1CVTLtetYujR4XbnibTVljw42xq22EKf
yjMkiFGWF5z71C4sY+UcvXGsHxVe7/IGQ9IvNwp9CvwwEavFOLaaD0eN21FvoZ9t
BvoTEqGa8sleuJmxBQhLL8kqRL7DcBkdrhu52hfXP4LvB1CAD1EaO9C7o5/jw1yK
9biswifHLibLmiWnyDm9Mv3Y6/dOdPXERWjit9SuYjzeZklzMrrehpCirXMAnngK
clTcf3CitfSV1sjjihdQ/8lFQxWIA8L4liZbHxwnYkJ6fGAugVBq1femcwIAY3Wi
y+mer0Vl9LpkKMtca8cZk8Gh13aKZ+2N+SBXA/+EMIu0fgR+WvZ9kSdNBIa/MABc
clCZdBuhonHaD8S5BoljlZEkb7F1mVtG43Iif05ePUCQz1qu+YngHXIg6IWMN/9C
r4WVDpl1ffM70sXiMRknuOXkOtmaq5gXbYXeyDslwP+ZHZrOHNjMbxKrXy+7hZsj
vL7ySilZ/vty+XSrJ1yOSjUERJ2tnQXY0bIIebMa4VVwq3l3RwOAdrvuIoknQWJ/
dmhV0iUN0blpiFIadF/pwM7foKFRwgD7nOQYMBMf5W+JufWJvsPIK5EKowGXytRu
pfY6tOfiDToO+WWyMsMYKRBd2HYjow/+WryeyrAuKRWEF1bP2erJj7RnAedIRtWK
KI2dhuDFH0aCRQwXEkbJyO3EtBbwm1l4oCuIJWZ7/HdVd63fsd+eUYnybzbbezpN
FXk3SCh+46ceG+cjDk/+7D1/JXFKKu9X43UvPjW8d2sl7Urjll1wlHr0RfM1BuLD
j6eZlGBDo6esyHZjxBI4sE8ozMFiJ/A4SHAjLVrt6oxsTNWu9erTgL66g6GFW1fD
6W7J6JSBwGJfq/xVDu4x1Z22wyuctn7J+wM+zLdiTBTJgYdGDTeGoUfjdBqI346r
JwGe//BWcuJG67LiiD7sNkYVwyqKIl1TNpC3HPDlkzr14lC922d+RfMGMBbxm8YU
hx5E08nWWahRxC7TG/mLd1StLE6Y39UCeGvGZc8MNTOh1SKi6YZ2Ael9Y6MKviDK
JDHtYOrHlq4CeY1Db3pr2ZJfb4cqEPtWnC+nY4xoV62EmHgoz1B3pn4NjsqrVnPT
ZFKzp8g62gxvyQPuoBPzYnUXBBoFrGu4Iqua81xe01/sp4FbgB+krDd8D1jdMdJR
Qa3NzyZ80bZ1lCE8QWPbAOHM/X+SQlYXlARi47xeG5AZhhullQHT0+MF/dc3OOq9
0k7sky8b8ZdkUmDHcWDU0duRPmz7WDHYtGyKK3SHr5vWzj0e9gAqBkQmp0i7eDm4
YTeTGdZSei/lqMSduJ4PG51yMlWg6RoZ1e6zFA5nyMy5DXiSkH7GYuAiAPIqlC/T
yNrS0STrViWEus/yyAJijPK0uIQkQUNZiFi+bU4PACy5pkZdbvhU8jFmh5HR/6k5
cagzmDPirzuP7zIWptL26p3kB0rhdr/FWDdq8MT+slHlQywu+KIu4D0joDZHhGhg
V14y/aXOu2LyUTr1fV210SWLCsHr/51v643TrpRg06/0ppYhx98dxFhFaFacYpbD
nBXRQUcjj0u/sWp0sOV/aOb04Cc7B7W6jg65VxmqTPfiLHdT/GEoSDCIT+DThTZE
rpwsILnzqH/kmqdZPaXvAZ1o8P4rkmG1EVK9zE9ixCWCeapm9gqlMCpE5aX3SRx+
pjxDvklOfmGO0uu9LKqJaKTlhWuEluV2b5F4urk9hcPEhtr49Wp3NjglfYrmJQgq
yEmqZIirelilueM0d5C2haJoB/gbw5M9FHp9xMxrBIwHOatzOM+AjQ9Nma0FkDiR
xrAi8lnJ32A9KJQqGYGcRUHBW6B3w8XkQKCtikRoemaMsfKzl7ho/Bji1frSC9wr
ZWIj4J6IF5Ubae9hyDC0/gxhb66feK/+Hn2pfnyp/u1yv2lbTdoQzfNavkQmkiVM
Iq0h5eojgtOnGxyNSV0G8v0qvwnBIhQ4rEqT1WykrXqTqqLnzS3vTci906NT7Pwj
h91NKV/8UawZ0GrCXEwLbV7FvDiuIDjv7p5vnomGpOurMy9oC9UrYzefqOLADh1Z
dkD+90EjsuJg6orXm3yvJ24gB9TnA7R5Z1WV7Vdw+KKdVYB3HhMxNvkjb8Qy+EVQ
Jrb+RQIbQbWN6FQEBnmKcxb8hi46VA1gDN4Qf8Msd18qovS4yS3bPekxEKhNtW2e
0AW61fljcuLEeIVHDUCMcMCtDtcioZydsEWT/cODeSGmEVlqZVOPKqe9iq79ZdLI
I+vvM6Tgi24XcQ9x1wtXLd9OSgLFEinpa5qAIdXVW1pkEwY+4Abzta7mC2FMY5xb
MIx8Pj4XzGMeBKhEY4zxzQoSAFpGIa9joOtijCxno4Mp28XxTHdaUCu/13kEfurj
UHy4JZnUqjjrpUdu9xOkEoPVce5WelJAWXZGgw5M+GEtb0SMtre/cz9PSn1ojjjU
n98JC6K4xLuuIbX71JDCCwYEKyXTPs1Ql+rTu2ko6hqPeAUCEwrssxqHk7V6+qYw
UWuI946fjuo1EYgx+bu6w1nPQfmEIAnkr9OyAF+LypRRNV1wgq2u7nCoFGEh4AFq
W3bBwcWtCTr5+O27ZQNF8va+qn7hsbyftL2bk1HxUPNLNA2x45j4d78Iodw35ZPZ
sNUmubaW1N1XjBfLC7+0vGzJgrD6K2E1jMvK6U5vd4vLFM9cgcIcqTuKdwpovbdZ
PZM04Y4BiUx9Mm7SadiVlmAyHEnfRGBzRXYz3H/RCoFOghRAPAx/VW6+Cs9Z79y/
nznHnvY31lvE2Ke0/ikO3f6OcUtgv38cF42t/2cfB65da+vVDk37KmSIBuYqmerp
KnS/S4L4ynQuNmSwQWR9tnxNxHRfTVCObMzTB7eEq29g+QQc8UUZhdcKl4mPef7B
EMZEaURSmjUp6P1G5uHPsejDOt9O5wLgsZQt76LDhgHS0imIVD0zwXI4Il/4Ea0j
lqeBfj/HPxucxoR599bF5Ie9wLImVQo0JAjs9KICgsq00zdzcj2VS0X9mUm7EnWK
rlIC7KlzgadKEjxmRFVvKc9l7/yB2qSSImpmxFibLE2qAq2jK55Eo3iO2zNTU8Ps
3c1tqVJOVpRWps+wsDXl61J9M0UBUMHC5O6ZDxvd0iJ0lDEcwRGmg5UD78Cvk838
kd4H84IsXJkfl7sOgvCSaCWnqMeXocp7heS8sz+hegvQMvf7Ne0zzoiVNawFwgMo
gKdNNdkPY3ozew/ZG3ZqMbejLWq2DoIThfe5mV+/KT0KGOkOdbq/FXmNFgR/yoWo
5ApV+3Y1/J0m7O3F2sHglmxPuGKIM0fGUtFqtxLuXlBfyLV5WsEI9f0GsPISPZve
FBNN1FCGdvf+ra9VhfGvFC1rRiWg49+O9W2vt/VJiXnb6WYevtGGnRYc1+FK7Elx
EravQshQTU2FMiHc/kL9Sx3SYYvlBHdCbr8fDNWdbCCGBWuJh6L4f74fBH4+wuPR
nD4Z2bi/6b6ou/XBfz/UEXR127y1yrV7lJUWJCLn/3f7Ocw4Yj726Do8lxLpjixI
BdEFckNF2wYxi+An6qyE2/Jw9JrHFqVvxFKYHmob3lRtIlEyhX5Qc2E5VL9bCplD
vmYEVoKPHcv3z4eTALgeTYJiVTjvZ19UYi0mwLLi37EQBpVd1qbexrQbtuuExrdP
PEWof8x+oxTk2zplV86k5M0O+fnvLsFk0j2K4Xwj0y8WoYJF55rIGiQeEO7GfzX/
pL1J6YUZ2LVuT504zKNdL4hN5v78dNV3qB3POW+S6NlcHPc0LUKfRMyBTaiZIqxb
dNtsbJJbVynBPOf9OA9D5dcgN5srmCsCTneK6Rw7vBwsnixcFduJJAobXl4DTqKm
smKh9y0bDsiJUUWGSQYdyfZeWgEcIPkLvWBHEfLgGGrS2YGavjTKbFNhSv554DSZ
bgdzfInVLzy7aA+64TFKpKPm+X4L52VkixPMdj8goXtpjlnU/2awhPrNoCc/hDzg
BPHXojHILj20EFsnZS+LER+hwvPaicMyH3LQULZrR8juj+0kWnMduuAOqIrM2zlh
3ChyrwmXiJd08vbsj7HXoGnjYKPmv8n5RiwNzC9veJ03Wr6dwtKZInwC68aGB+mS
dV+LzDu8oM7uifbnTaNPeVgTQrcon214dXKvu4NxKMNkCR6rJNvZOqcg+dUG8g7E
aga9KIqpvgoEfRzQad3m9FILk/Q0GZas4lS0s5MXoNZOgs2r4aatm4mWinT63usq
dwrxIhDErbUPq/qi+zgwpcG7ceDxNTuBI7KB4j9e+XSSn3XW47VZQmfnV1kEjQs7
Uw1+JEIUPQSVa+kGGMemuzJQ3m71U8KDR2PaL92fQeYtLORuqmiH4eZQnXdr42xZ
XAETlKbOXRHktzHMXG9PndKpBjdsBZPeQ42apinaG46uNGHFq2sqVsX1VGwwdf6k
6FPOGe4YkFjSUBNlEChRRJF3B4RnPpBPEHcP8VPVvyO9AZUpKICzl2IveFce41wz
byYFmKPjr2FBDsZSShu+nu4eT+6dl2vprjDX3Ukynm7SSdXLwPmB5pqztr42UYq1
bSiICPRoakVVzVBvVuE3+vkY59XPsO2omc+5h6v7QyZPwufLlwqN/Qy0uif+qjVh
S9AZ+lboxpR0Ws22V59537OvWkeEkQkIASrNO08K9wKzr/sMuST+lEmRsi8Iiiux
yCaTZEhwpcvSiGcGlxHTtt7dY0pPPQ+/aivtijuwbyztEQPuCIvtQf+F4J/SuA+F
UaBxgH2gndd6Wt8UHvv/Dghk5jy8Xs0kMz9uG9BOkp/AzjnYdQm41HtrDJwvwxhs
WPpUd3hCs0Ynafscl48rwc4R6HeL9ZyB1IHxIMg+3X6y/xKBu5fOlD5lalgQZZnu
/okFczKO+UlOsO26QoopluZqxSrBfe4LdxsTWsqhkkWpMtHuUu75U5pHHwoMWnVB
KT+cm0qGs4wT58/Iyvd1dBXPD9y1FVnDUd22Ds2LFq4afQnjdF2KpkOGysX8FIDJ
SRqXi0fJdUOSFnGtwh2yTRaFaUVVr2Vl2aKcbS3xeJKfC6NEkZM3dFH8Pf5ajCUo
PJYv2WJpnvVKbsInnyKcz5nc8XGbQWxANdsf9LuNWAheEI4qZ18+Hs5swoPO/AQ+
CFTxpdjLzDXZf53+2nDCEmQ6YmJGGVlEKOn4S3dLyK6Lh9AdMEWfQLXMqo+cMOGQ
fE5ZmOUNU9N+Br7rf3XpzPiV+rpK0pdZ2rt6PgMP2X72EmOumaLe4jGJuAHuC3An
h8EZG3C43VVY68zWVpSTdiV7P4dvoK8jREmSKE5i4G/enk40vuT3DH+PSkHJ5kCF
jlcSkOjTYmmeaA5E9SEcOoZehxjYJbjN+tCKlaUdrssCXFu5J6gfAlcNITY0Xp3d
HvRAxlms49w0lJEyk8Vu9l4hEqjM6kyBhUThJvRLHF0QCmqOzz14NcsL5ZCJDv7x
v7I1vi0bEUrhKDXXkTjsn7+TMOlJTQUID1KF92G83qKGd2FutAQxr/5oy27HcXRf
KHcx66OtJ57ebV5JSeCpNt4BWjYPmXZGQhSCpmjoDkyOb6fucC/AmBv9GxjfY4FJ
BuX2DyMGEpeB40/qkDqLn7JhNsEKTvlfHPuH8vuYV3u1pt08iKn+pa82VOvaE5qO
jk70f0NKa9brx3/N60Si5kd+yZnSSlDooPMl4hmjVpaDpNOUhuXfj+g8qJIfot9c
0IMQtmD8PI4a8ZrJGYwypbz45vJFrDbGnew1jxsVHur65IpvmkRkASESmO/gUDkA
yciM/7vsyKx1eMmvPqlQAzj+Y0VjbinNBhhWXPxs4cKGJsqdAPvQMwVBns1/PsgF
u49+VL1blVbYMmjBW/olPRcvLx6M7WkY2BBoqKeMSFWwrDALychyWkBaARgBRz3J
TGlL7h5hvMyfRbxc3Juxd9VLslK/T7u82BSVnCbEhZsqStEEP58Pt6DF2R6SmD2j
nDZZQ6k2G5kUnZi6rHUJ2UIDazA921tHcWM13DerNW5OjH0VyE13/YT6RobjFnJ7
iORknX9NM/Sbp7bbEtZwIq7DTMMRRTcPrEAqsjZJDBOjZs76TorMRIuSQBYgeygF
oHeDLWyPpvihTXYC64pWkLCMLE8Sc7f889Mnmg/m/VOa+QsNC7t55fKZMM15wlJ1
Gx5Ulu/Twq1kviuSVnGHtS36SvpF7LJWpXayVPXiSJlA+TTAEvLWIibjbjl1UZyu
EvRRODsGru0XnLaLYQxf9OmNVe1mKY0hSMVXd8y1n4vBBNHNXNSSEpOgXH1p+m6J
79RYSYAzxp3H6e2uv08uebwiAACAsc306OMTJ+NOBT6C4diN+vjDdDmUYrCWI9dH
l7YUs96BuMH1k1OQhmGTmTUDSo/yMNECFfCZkgWKmU253VNBiAEf/WkDcL9f9Uub
crKSvA0IqXG5aGSFUhLRQAmveibd0ZG8nUkHvX9rDlzwMXr1L3CmDXY1qdQMxagT
Swd0xsFQ1XemiJRgbXUZo/dlzi1wa1h8MePOsKp9fAxp4J55YrFuB/4d+j9S1EtG
GR1Z++0Chngy0K9s/78Frz2kphYL5QvKXrn3QtMstAn7Vg0GAy6tMErX3dLYAbeS
JeyiiycqKsShqtijQWodnLGOfCqb/SEjNB8jsxj90ReX1ySmEQbc7OIH3zYn1c5E
Cb0PtNeP4hkBRgakoRclbHy9laOsGQ/7b2QqHyhEvkKo0ssJ6s1omVBs9gK+dtXQ
0eYsleBLb6YAjp4fGW1jSXTjjXeyb3fc4UPr9Acf4Lsf3G5R5Y9rG4of/vGjdIqi
JSF7ID8olBLlkXyBaPa9RG+dXgBdlgw/4xj9dLYIfWWWwSOIA7ZXcucT0+Vsm/dR
FLYCOtpNHqgaj9x4hr1XBVcus1OtHt6cHom31cT40fvL4MCUyxAG381cVjGXoSwO
FCGiYRzH64DHppiZk7ckfvws/HMoc0ygZB0cRNf7lv65J+PgGj5PJacgD+W4PFE6
dbK6TX1ig3NNiAvGBiuhLL8YI8EIEx0R/qjGuN45dEmZ76w0uY5gewrsXmxZiUb4
faKNRcMKDrNIy3L2qjeMizxjVC2MK5KsZmYwqTTZrsIyDVxWoONJnJJTkfYm9wIS
ZxLhkJHjByGnXEXN49ZbNH3EVr62fcb8ofUC3dVJh/PWJPVJzzQdq413NVgnnVdK
llQ7kV2CRfSt9Gj4ffgAA1ybfFOMwMm1fuCe9dO8LM2H+5ufAZcfCAHEyhBDTZ/o
6SOCPBwUJ5T/CwWBjs/QI6hpMqJmhMqMEmUd2gcuwguq18ACZIaUkSPuQJpVBify
jyG0uypQhSY2W3PcYOCgH5aA9wweNOQhcv2XPgRG9YQOYrfjU3EoVZUpNHaxJMvi
i+Bc9L6w0HoXhV1cfbefZ/L1qHVDUihCuO0h9O1DV6aGbz0voqkzQ52SEkPOmSRR
ce2Ee7y+DjsiQG/mMtwo6Bo+nP5c+QK/HJb18fvmvx8lnsZLASBox52Is5wWvL9Z
PVbD58TC43UFSsC3MhGwqfblfLVCa/l6jr1Tm8OxkcER1S9Q1wqetNNV4gUjgec4
O+k3nWp7jDah70q7Da5c9mIj+NvXSEBqRlPNLHvfCHmEjOil4+UYJt3HkwsNPOW9
MYv2jjahpuBf8/VG007E9eauRpBztYi1HJ0VSlG75L5n7Hu+gidPQ9jozlviq21n
DO4sdWmcBBeGGXWCw2sAHsSlc1iRXIzF5uigGUL6jtHM4haRq1jRuKFrY4oVwc8g
Zk8YdTJ0G+GWz7f6gc6NGfgeU+4K4wRSuOb9apaqM6VprjPzfQK1tPODr3sDSakQ
JWXStQwVVSMsWm4EPORqmbQrDoDtJOGleT7LDFN+Ut238h4b5kzm+YEcl6raRSnX
lJJ9kvztJfQAssUAlSCIGfxtFLsGRlRLeWr6BNO7kB0+7qT/aUJ57vzoM6fqijK9
nsqN2QVObpcYAaVD0wdxLVPvrdxUolkDDJrNmc5yUWmu0RO/N/14iAu54EEyjszg
T5dOJX9XRTDbQY+oYoB4Ph573zGPTjDFU8Syy8qm6rgjUDBuyZVXd5LbfQ+MV0uc
8Yjzugwg8M2djsb1ZDfif1R8Rko/3Ey0r0WkjSpRqvF95ySEQmQLjJghD3Nh3+GC
IpwwOM9Q5Zn1ErMzyBp8q9zMmhULkNnrGf35ky/L5UpS3eoNoYPY2+EYII4JodvB
iSL/ozWV7YFimxw/HgZL6S7dukyBcLzBZFmvXEaEBxjwfGXi9TL6DiYKzWrxeck8
JUXbEUrX9u8uFetaQgAil3thq5NMnk7CoUuxCk0POlqaPDa08Eu0NkzH8AQ03yZb
dbxW/p32cUvsM253wFGiGnbpD34I7YL+tFdf1PSDdCV7Vg3ZfFIiIZjkP/yqXPYx
Zb7t0gUqxHJ+YAALhIgurLZWxugNPEOlMfDM6yubeZfEdXQ5/3rTXMopIQDIyzFT
VE7C+IYvlc0hGAcaEbPb/JmGNha6w7iGdw7kZWya+4SAiA8Ok5vGUKFBIZYKN/7M
VIvoc8gt34Ze2TN3QAsR615sRIe8EjR5jHYzCfD26CoUD2CgZKRjNziQIiS29kAF
H/Iz6TjWYXCiiDus9c3yMlrnYRYK864qvDpRa8EoKONafQQDANeVEAjuwfrbqva/
2vxTVJgU/DJYAeqSmt3PTZ98RipNrJzA32dvGvXiG+GWkePc5zEuxavSr0ntSKoS
QWMXX+UwYE2DLvuELzBOl9Wzu7RxlOvlOkypDjbHWMORIrfyRZry2pGukOe45Gi2
u05+f+33wBB57grRjWOAP3xH+bI4eZ4ro/w5+o7IMaOC9KW1e6m1sxihAMPe/VkL
rc+7cqNJAO80ge0idxADZJakgoZFhAR/2rW/FtaLkpRXPKs7dwJW8mFajr4l9JJR
95YwrcO0HZIdmdJCrSxJaeMvtMlJZioNuvDzZ2h8Xesrly3O9n/R8DOGU5Y6+N+G
6oos+eYn4HMTXrYhF6XCTqyubaZhQo0SloYVuV0ZSggDJrxHf6RJKaCYyeTkwK3c
0lsk2+vFuggAUiHECzdJQFcujSrPFxgCh0mdhHgOfLvVoT2ogBvlNmzJ0OneM178
0aRKN9DyYqykdBMOTG7F0sseK8zJiiGxJxHw1nUZr5jb2kpMlmO/2egmKweDT2BQ
1nmlwpJOYm1r7mJNzI2++OOUAYgHtiJ9T313EebVhYV8DTd5V4aF8x0iXten3E30
u6q8JeHfJKF1MBO+opbBSruxjnfD46xpvUcYWB+ZuIOa9InT0v9N0/JS1PbMgqQp
dWb0AWeP4NiKxk6DxTYKfs+6OCVjA/KguO8Nnylr74LiMcaDhXaLEPKjU2a8P48O
Q9bv5pxZVesSKQZiyLoeV6yNvlAJNq4bvpAo22AHeK6b4CoM4tKrVftMHmSS7KCq
dE/ZkhdE5EIk/ZoJe+Wq8AdU+NUvfBL8pcXiUs+Kmh6QIvX9MMGO3FdiN3d0/Wju
Q20O445cZLv4X6fsfFuqEzesGb5A8/tNKChiyC7Aa2Dg8Ee22PR1FUQ7Q2gfirPr
M8R9pV3rNZtXu5QfILjA6Oh5LERX3D+mJHs66l+NX5oi/UPd4j/PN5YlWzPRHCQ1
RjqOX/y2GEa503Ma8AnyWcYDnBs5sZ1H6y4Rlx24cVhFBZ+7iOTubtBQwxNpCRg2
V96HtCS9cnhjnIOsIAhLd+QIY/sMSMjiXN3Zr8PcsTe51gK/GlIRh1nGenr+JRdK
xJkr1v0CtJzjmHyXxxlQiRH6xTVix3aVzIiy1bfSepgovDVmgSczSaOJCDArOdnn
Vqz5zuXf8dLI+eGKhXrTmC8KPgpVS/xELlq2vbFNX0X1+MgtEk8spZUv8vX1D+fo
XBzWANqM9kpdyGDCJbge/X1W35MbHum65OR0WAMggtRGmilMZHDE5zwHd0amynbt
j1lWBwT7kriC6GBuLKsnG6ShbNk0RFWsOoEWBaM+uEIlJjeYasosQuKTMYbVa1WM
HoEYX4J/KBQeIV+sy8Qc5xqejkSgtBHd0jXhka/AFwR7OjjW0NwhYsfPZY34wCXg
kikSkMXLEXjki6Hcqjd7MTKLBOk7fXWYfFFhoZMTlvWswa/VaFa+yCqVuap+iDb3
MRMkLvLSoWePeVV45Pci2ycvnxgrixK0KFXTK/Ug62luEm5uDSSAEfO++tGomRVg
QdSDwDx/sJi4GfsJnGSr4yI5H/BQ8fwud4AqmGUYbxoYV6OIVQ84QjgF1t6LMiEE
IQbMOn9M54eZvC4M5Ui5FE53vAFU/tinahmt9uTKm0NqBYmm6HB2LU/s3ncPj97e
KbqVu2FGwhWqCUr6J7ILH/qqKPMuEihdBXM8sgJs9JtMgUHvd3JCxahRxiC+mDrT
6ANeMsd99mBS6FjeFNWAGIuyt+KDu6b4aRCyq0aah3eMEOMuVnULBImhWmOVDOff
j6kI30JKNI8NjrgxjndPAxwllOXQHPg/5BwdsMZUO78As91riycabYlLqXwiUKTs
V6utXKn406A1KRVYgkx9PupLr0QOdTj+crqiLGVwH2fWNxrE7SnbsHZ+xUdsgRsO
evm6yd9V3cYHPWOW7/ffldcEIR/Ioc5Tg65l4P6gI7Cc2H70U+uarp61tBJquzdx
PI5++VvsUVHIEp6j7fVMH5COObJn9yD/dxSwe/xFR06uP8ZXDqBvjyFJuUN36JBl
F7h9CgenN9heFHCZ46rIdPYBN67CkhBnRxyOWz3WbHSWYwQxwFEitxfz6aTYohC9
AXxbxMSuj+NyUbbgrwGx4sUNA8E/3oQKApAPEi05PltfMNODIqUnGL8YtLLaZwku
dX1BTZ2NZJGhG/rfnm84oVEi5KN6HQcUf/Qcy08MSA5xUfevOfWy9fBNfhMYI9Hc
cjycP4f2lS0hl1CCUIntpEHMJqMlLMqkdb6yqevWHCePj6NEsadr2yhY9VWVfP/N
+uvTZ4IPFaFbpeK5TE2xO8Kk9l5CEWl18pNbp2s0UeN+BIcJY/oanbnWWKDtlxFK
a/QKyT7u4JAr81JxvHpk7auBYcg4y30U2gLCb6zHAcd7nDBnr7BWAx+8I6xuUqQG
cOX3yr10KSwoZz0Ci/mKPy1aQMpjkOaJaZ8GwdGc1bQ+/dhugZMakwnIwXm150dP
xdbfd9/W9j0KXMr8+uBmt+z9FXA8f5P7Ablv8nDfRk9FjEDoY8HMgwPHEGy/Tg72
5zGlGc852oHl5qCGAT6tG0wYA6gMRXe9IIqkbrDN9Wf9fqYSGXczuo0U0nwdTb92
9lL9agLmH8P00iihRSE4/HdERYT3joqzUD7j4IYihITWq9xMfGm5T0KtdpWSWKHK
srMcJeMuEOoupjW0/tkOHzM6/v2rbQ88/HQCcgfxkog=
`protect end_protected
