-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
bhaY/LuqPFGxNMyau9LU+zEtHgNZs7GhRvTQJrF2mA5UlPnAByD3N8jYP7qFznH5
MHa7l6atzx+330VNQDFfwseL5iUqdgtgc4etEUg8VhTULlbfpFd08v4dKFsVdYiV
qDZZIjGM8qgXBX0QjmNwUMgeuO2BXeXVuciGTU+ms+I=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 6063)

`protect DATA_BLOCK
3GEVtzZmdT+G7s/a539SX2wLmrmO+hI6ojGQI6rvGtc0IawybvE/px9L0xE/RNc7
QBvkmH3LHPmHjuK3niQpHvaqm+TC9Avi7inbtKYt+W36cCEwa3itPdE38mUmYBFr
YR9o9kGdFNsG9uVbKyo1JWHyBqEX/uv76eONfzjG6987ibAw3eOESxF/HSjwBGhn
baBd3YGy9UwZLvNBIB8DD2sJlmHhdq6yJGONl/ao8EmNc8twYfGFsXbI5z4nJCyu
2cEbuOzkIdKp7X6sNCZ0kbaFBZAsa8ozwNlQAlYQhAfg6Z6c55FSpWNhKKUq17EE
q0R1sQyU3eEdG0X7CJx2o6NOQUCb62coYcp/nHTUajLzd4Pwd5vWSLYKRyFh7dBJ
d9Vy2W6lUseiCbWo8gomQwoOH8F/9RvNHAXsVMkZ3w7W/Fs9mgeJszRPji2EtGhu
m/AFY2IYL8HF/D2L6FYvfQL401R95iPwNfeE9tb0UhZJ4lZkKMrPLlXw5h6ed4XA
798pcqahhrFfyYhv0CaOycOBEUSiGGKWDuH5ccW+FexRoqLgUr41eMLYAtTIu8oT
oJXG9RKi8QO8is8NEpnOwTMgWOAclFDHa30/1PMaf2lNKGrn4wRc7Kr6ZR1jrf5Y
biDfv19VznGE+47kPXcuJKAH3mxNfspLxYSsSh2BJiy8BpwEeK3Bcwox9nsZLVwS
sHCtDBAs8ohtAgg7ulAQmDb/NJbbHlFuVrloc8oL7COHMrSzXpuYACih5MNU5FRm
qGvtRKCXTcwkLHJe11J4c0B/SDfKFcVlIOGAEA55J9cTQgWBmap0m7IYA4vjr7Yg
qCf7h+NEka6tXm8Mq2AWLCtyqX7xub4+AwQhIdYKDVi6CrP+LqtJifk+AX7kuK+o
2MhICK7wqKhR0UwIRBeL/NOUI6POmAmlQCNM8f85cuaNKUqfih3Nup1VB1O+/0E5
x52UEED4NqZbW+qqnwsVNRC5bDsjd03g1mumYk27ROBn2NDxvKvpVTHPbawReDo8
tkLJaOJDzPUGpzPu8HqRcUy550xDls8TIzu0Yd/dTusSty9EKK8HXmWqtoptNiQK
AVf2mUojepgAjAhn2prFRCh0s+f7YniniQJOSjio2MdZPcvGJmxyLWS4wQ5K0GOL
4nd0Fr3ShPV7BDsIudjIsKF7U89Z6WKxQAQhX1RpgMeG/uv0tna9vvso4GKZb7it
dHLph4aLgvcIJjqhaDYUwyBZ0P2tVwpQyJS097OButRX+GwAVT3wBgUNudJfW5fz
iXOyk5Kv+Uwx12nhFvQ1DOLKN0f+ae6nzK+Q3HXlysau2MOOu7mcNLUU4+JlHkFd
m1wzz6W+EOFFkMRwZDknU3ehd0obqHL4Sktt6E3zZCRPHPls1WJXpJZeqg031iMF
9cpFMdkvCtiz9/9sikwQvz42p+3ldtgPj3bMhIKgXEi4wSX5Kibxkn7dpw0t6Ffy
nHHa6IfK9N/JlBZZtx5rWDn4JNIDP5ZAkv5M+7mWB1YZMHCAJNowxQ6X7WvxQEvN
9al6FGL/5FnttH7lOkNFWhb8rhGQKzOODPbowPR4Vfq5rpO404vQclLeZSCM8RlW
P/fgs3Y9VV33ogi8LGY2z9Vj9VKdYq9b9EKHuDOXMYphPLSXTnd32FVsMRyFHVqb
290LyUSuJHYmqYOJsMk0kqaXhwk3oex9sbevRPiIye+fEPUEbeTKEMQmtasJVXFz
t5uDng1ea63cfpKNsKHC0GW6G8d7EKq7OS509oCExXvrmibsLz5cIXSxdNWNp4HQ
sJ6eJFGNaIasXia+u17l45tsSs4MbR4KMGjUCDwLHFGDcSIrR5jwfb8ajH6IvnDh
lEqo3pPWctNSITib9a8irbNv45pKp3jd2IX6RAqXelAEmljZOePm2HEavWor4e6u
dnUkoYReODjhM5gYycmyYhlbLl3hux8wapRUSZ/Tktqa1Yjkdb8EvPEjED+24z78
Z6pDgeRCvZhdak5fhPLinSBYU2qKQuAPy4esDi4SKdb+V9TFfson1AQ51pUR+0ER
rQ4+QN3cqsa3hmVanPiVDA8xUyv00x6rodbd1RbVBANQ7/jFhIlQft065zGnqUIb
Eae7OkfV0Hr3EIvC/SVnW40DUZ0BCyqt3VfYsmAMtiXemr/zpG/S+lzwo6Z4f4ho
dDFKOVmtX8NK/TWpirWJ7wiBXNzt9Hxd0A21+yaeUifSIyx8q+iGH4peH2O30Ctv
KOW5SCqPiDjdsG0OSEbwFmXzdfR4IBdBpYu9ijHrJ0QoZDrpRV7T36VG9ujjc3Lk
7ewY63YNmKeRi+CIjZfm6aks30lJvJUCY00P53BO1G7PkvbCNLnLFYP1SKA8T6Ju
ZknEHHN9iQ8r9qAlKbTxvwkL5FhODbIdr80o+jQXAtvSw9eKnZ4tqsE+TprQ93WM
xXjrcxEk7fNbhxQntVHTA9pyiVLCuhtswKpt1JQvYiZUFDugF2VhIRVBQEdnpOs/
JF7iwxqq2LyUM/hm1LeJxOeRnwx/NtOI2nBL5K6bhx+X83auLNzb+70kNnM7zEtB
B4lYmcwULI9wPo85s+95+JHL+RUm7KXzuRBRxrNrpj0JcEFMezqLOSv7t6P88fat
57DoU+gjMlE+wqhVx93zliGt+pHMmylq1NeGRBweC7lwCzzc4hfUHlr1ymfocgl4
QIPm0ZDvtW2MCPg1bXXcSGxzopgl8DhNeX7oiS6riIwZStlTQVVYAux7xZb/R54u
kvrJz4e4zh8vWO50z9eFdZ/ElfpE80+7a0Qxhj+/frKjvmNgBViyD7AzSPfslV2p
rZHglFLV+ZWHSv6qLv0FLG2e14R+j35GQn0CdoAei2RztCdZhNtmhG5F2l3p5oJS
m2xspvpwkgbEf/zv7/qxcakw7pP3Bi/Hd+kF6OjuphNko1qeNgLYoi9oLqzfVQ9h
sI9vCxVOO0c1r1lAlGxT4LHW8owfeK9JTWzj87Cxg2kbBgaXpPU0NvVihHGVzSCD
6TTAL/0FOGuRDyFb3qqXVBXmtfpd51TrcsMV5OBxndCBDuJTkWrne1/GwnIFZS+e
Q5/7I3uzVUyRljvNBPhiaxF7BhGHmxsfJ/U/dMa2/nbJBCEktriG3EqxFH+LO17+
DKDpdW+730EOoKoVxiaFUT3ZNLnqjduBg+/eJljIIiRDkQAu4zGhFsJ0BtbdQ5qD
uYISo5MkHd2PETvyudK+TaaS7g/jpuZxJgyZ+fXuufrzPvmM9ESq/wdcWL1sfF0u
JL1JqGvQo08k/4DsEH7aPKZEdNxxCOu9hl2QYRPVpGcJsKF5BVUkImfizNg6SQjI
nzIGSyymvuOd/iSNt4rqRrLJorfmG3nX4kNE/DEtGiGTAOqyqqjpr5MNG6Hh0wF9
enJaqpGb55ej0NQFVh/WiN00dRectWJh+Nft0b8RYcpyESSjnDJYQQHOfBS5jFds
FGD4j3MwGBGGP/0hwxWHkhb0HYU5tiaNeElx48SLSxmDHsHmm8ex117vxE84GZhM
PvPP1kAuepnUHEpF2g61+3QFS5pnj6jHYDovmiVpqpnvtAIei5ygpuj1scoaY8qV
wrekxzQma0prH/D0DhQEDjh67hssSDjLEXGaP+kb+x66tm+QBaiYq4WT+NJsVAZ3
892DqrzlqxB2gi1OldS9ygXVb5Qeu2hfxAXWYC+15Acna81q8LI6BTdS/M0m1rPn
xPy0x8KoZTV5QL86bFzbWbbBCAHVtdUKCsPiP/URglsNtI204P+ZKFglz0dqOysS
13sfOL6mWpvUD+NTaoLAOnVRnccNXlpHPBFlU5KA7M2JZimqmDsHOwOj34VXPHsj
36iB7LYb1Ie3yMPz3YPXpwbwcmcfVyqUeLM45dShyqty7696IBgQ5PRMEdDvAESr
E+22USEPztGPgqXNx6k87XnqZlIJfW+UBqt8Ld2smACUNq6LT7QuAk0Ll19nwBy3
HzqT+kkgM6ECx2U01YCbuUfUDLR9QAoMyy20BBU7hHlWSVYI3n+BHafd6rolqYVV
1l74NeiMZQTtNwPppIRwNz2Ozcm4bJytrzZXVh4JrC1cL9gknbVqzmk1SHpH+wUQ
DDYEHMek3+WWSXkOTNGzHSW7thGl9ksRYvtjjfp+V1b1SSTeOd5yqV92GkHl/eAg
DRl7igLzlGQUpWywFJEWnW6/EcNtl/SDxGy6ppKKSMIAshMoL7TIsKSWnZ3xVi3w
Q03pCsyrTx3Vf79w+1pCEijo2IpGRpA6WRPEhy2+PR4WPLI3fGYlX2rzFfdsPl7q
OIhKNVjLjBThaGkmdMClqXgVhMA3bR6x/G0OxjB44foUgGaz/TBw6lcyY9LUtLPs
09XuBLGvHPv+qNpR6i//gGno9phqiPWGDRtAwKM2bLLHirgpmOBSb58bnXI974Jh
KcwKB166kBlYqU/o1A0BoGpf08Bg84ZIclonhnagt6F87wdlolci5f6dSo1KqRKh
qi03zFu6pNg6iBBJHH7lm3F6aA6NQb8x0dKqaxAdwJovEywWLWcI4/B2PO1G+5nX
UUE6e2i4PoXakZCmTwPdJksGPPknllhIZMzqFnjmNjrZ4WfF8MVGjJGQXBV4KzaG
L+r2FEUhqx4cQo11K772l33ETUlYGeRFsc0D6JFD6QKh+yzKuYIYN3QmeoXOmcpP
9qbscY4cELI7Y0lU2k4DtUK8xyQ2mjor6yPHdP4lwlv3WdhjdoIgqnH7EtWzNvop
SuQ59ehOXCTPwxTFJ01VauPpsxX3yHp4jtOBU30nUrWPPw0dtCdGTYtYy+NvaqqO
myD8RT91qiy5j5OMmKCdFzddUfd1oPk/ph5f6utNe4N1xrlDAlsrWk9kSGRM2Rqw
oIyJTahQG+IUoE5Wsj47XrNkkWvS4g/tAwMq+Xx8l/T6ZMg7pgji05tmMCJqu5rz
oe0x8abH409ZTBJ6/qTMWkehwxhQoESIAx8qPElLm4DekQMgg/71CQeS4P2vsGH7
1/+ZRhznyHcONymXguNBO3frrNNSZl0Y2GkudwLnLhTaN5s6BNCQMZXcQ5XoXZ4N
/nN4iT2P0mcRC8A4zdIAtmco3/dbdZf2WXkAV4VSeJGOjeOjjgJysrxVp6QVFoHs
Mf7W4cxUTdbbKtp+KXYgD+89YxxXe6WL04RlpPPeAEGPlV8fklDUakXguyK6HrO9
66h5VjvW8pG1px8v7jyy1jn99+OU9lQMHKM/dZa7ftgb7hHhcpttmEnWON6Kp7tK
nYvc1waHyAqPpdfrcuB4h/F+nhY299vgxjpu52hhwAuft5MJsxq4K3sBsNSgVzzr
ZgtGJapC2WcOtKcViGNN/tirJkW2g9UpTJ2Z+iHSsqaAYBFYz2YLo3GB7h5koSja
L5uF0To3SMkFhSM6F/oDogho1QLsM3eqWEIZ7tdb49LlHx7sijWFB9I+T1Jzcn/L
EC1zlldiArCQ0onecXUJCq8Y3HVD1bPlR+rzL3FAkxwvSvcFI7XI7u6PqDgKENoa
ebJl7ApoZckoAOC60Sn9TfDpNxxLqJQli1LJmdV/uJaRotxyTM5cVRkLoHLSWSas
zXYdALnye0VLLEcmoz3uTTL1Doi2xZWsuwrPDm2U5tNg4s/WcxBZRWMA8K8WJUdW
KYLWg4c+oEIoCt2Qx1CvDQkItBCw81mhtG5iDVnxhEJI67l3hfKfzU2AvjeyxEOq
VLYKOb6sYPfjXd7nCmPm9529RaR0kyTt8Ol3OdSDld5D5WmSGThr6/7AhrY6Ntj8
qdkQvQrfy2DbJgVZT5n7cV3DvBFnJK+0Y3jhOH+dP/lFQ+gR/e4QXCwCXq6ev3Ls
GAtGCCwG6gVhKkjCcBv3JiGWS2xqE+eVtyMEbmbqRSfqysiQFATagQL8J8eeoVPM
fIZfIbqVnCZ7yPSYDEXwznA+ZDcCVS87ZIc615ovpm0xKgKo+bFP8PktC6jmBnGq
LLegMIy5hkJWqlHjdnBzOuhLIEsXjI69PrFegK5VpVqQkTvPXyW/rVUZyk5+/Iku
TSTsZ/BftgOCoNaUTIl9Z6PUQElUkiPtLJ5Kow7l36xogTS8+NzodGIbKeS+5LMc
y0TWa7Z5VBv18ArKMLdSmoyMvP+iVNVlU4ebr8vbcKBQsDVGH4V40RtiGaGtWNMu
HOxcLFRMrOcGxNDVoDceLy21G2eqDn2FHm04tcA96FZj4WePgMDFgcP0pJIm5cd0
o9Q4CUZaFN5W25lazycIiG4pFyrsVlCgHvfqu5MCjBT0LYBT6LJnw053ysWyifb7
JYYi32Qc+ZEXZIzFaTMLNL33T1J0Rh6xbDpgLdHqe2ZtbITKSS0dHQiJewY/3d8h
aaq185BvE7alNMR/B1Ma6X/RSK7gEo5CLUtLMlVHgZCOPNzrM1Wkcd2/MVxPX+Qt
E0tuWTzF3kzneCu2kX/w5ujDuh5+z+Z100dRtNpTYDvbaWsTk94hrTRtPIyCCzl6
4Ci91v6hjVwRytACFJuKQaBTaUEsneJsy8ldaXb5/2AAhOtEoTIve9T2nyXYUQXx
odER3JvtTt4iEyKRb4rsrQb+7AvKDbs/2wD4Yx7+eoloOA6t3E2HVUzref3m6wBF
QH7Z6WV/nclrNH5l4U6RJPrst4ifJOF3qJ2UMriCG5D/kEVzoWPRkftPeBLL1c07
yyrGtlyFSHR/kXWm3MzNjXvKsi9n6Gk2xy+VLl3LPU6TlDKOxG6oknTZQJzv99rO
BmN2F7Fp4HfTM8SK1rH+GNdjvyscvIukzh7gH3mw0JCPBKz9PW8ZFFMr2U9All/Y
x6RRWL8PiFgxyrxUHGa+4qyxnNdWtNoy9/55h2nMeB46CTUFCvmn8DGGNovIiFnZ
q0g0YqBfTdCjJkSbbOY1YxJWj6Bt7gjLVdvGvqEJgHZSbsqc92B9+qg8m4YUvUia
hbhQA3MakFNiz/SlxYIiIVqsqI+NRoBXE7zlLYH1BWUV9vaGXl5atxA73PQTYTlE
jMvmsHh1NwykUrfS5qh/01Pc0hW8XJ0/cLDxllx9j2NNO5Pazp+MqVoPaaffeFcb
+vBmsD1GqPH38pSKwjff3LnmKjvhRp3WcBXOfXeWBNKtLqAKPgbYqNDrecOv0bDn
X2GlSO7ntNxdIWp4biMZHKlyTQcypWcCGBzcFE8tpw6DXUVZl3H+R6geRLr3IIGb
y8vfWW+AdT8PeFtIgaWyJt3KZSSLGKfCv1SJhIE5mA0/TaWoKKMJvQttac26GsnO
o8QTQJx8XcQdqVNmIOWaGUxWZnBI2mHZcHGIszC/kkXWDXqyj+59u5SBi/MTUYea
uH1UO9/roBuzSXdl9oXbCC60qdna9+1NvQ2lBy/eQwB4mskn3nDCTyoZL/QYTo39
PJ0cHICZ5kWsYUcFArCZFB9CeTHgYpmDbXR2GPm2gKBeGOO9qEkRxXp7kkQfqd/5
/Tx5oBdZpmafEAopPWcl5Fv1TVNdoUwRG9ijIcdoCzUZ1S6EnyOSu0rZpvAB+JDO
vqGppbBG28+tw1QNQcRFk2SPAa0URrnwFiiFvkyWdRgtvTTs+jDc2xxmJRk7gFnE
3PVEWkpee0wQrLp+WUMYi/GcowLa2usjP1e0OQHhokjGxIWM6UOU6ov788j/8skC
PtYrYAnmCYzuHvfiDhhhlTkmDI1ZsCHXM0MjT42Qhehdp0okoFUFWIV4uB9WU1nH
SHusZJHoxvxFxtAlMy1JLzXiScT+6XhgCLz4URkO1FpJlzdbUeOCP9m3cagRUzOW
fOZeQ7hR2aNhs2Z4tSz08S+eJ1GwXeHZXGmTHJ9ctLGi9RLkZr17QHZ30LY06kLs
xe1PvgqeoPmZ9yq633f6NpQ1VNd+bg15E86fdFVNklaVZyw8d4lWRF8QnyV9V7s/
085KQVEZQzTQfUV9X2Y706IlLJ/ixrvZW72MAd4/LFJtHLilgIGMshTZ5vxkYToR
TcGB4P0NtT7lIcHrNU//8e3/cr9eWVng223xRvJhKvPzpqS/B/YlFNWtVwbFYqwv
VQ3IkFLSr4gSNwC/6Pox0EnsuYnwc5hd06WDR5idxGhK2g64wC6tA41MFMdaetmq
rFBEYt2ojfY4pfTSJtWqFoaiORB5sosTyJ1vZMOq75w=
`protect END_PROTECTED