-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "N-2017.12-SP2-4 -- Oct 23, 2018"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
GwwECGwtZ55KLZo8hwWHUeZgi94eEM0G5yKuBEY6B21jjq61DPT28hrNsrJX6cVs
Gf0jwQ606C8cX9p5EVckoSb8uwHiJxuM3y5BQG+Ls8t8vWVC/d0HV2IMd1hcmG+9
YuCAr3C5C3+2Szxh/YK/WUBBr++VUorheIIQnMQgcC0=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 111872)
`protect data_block
o0TOghvcVSJx3WtRqhfQ/L4vKa5gEKjZN50v5syfOhq2c51tQIa9C9IPGCmfgPw3
bBWWA9e6LQdjOYSdxl/ZnfxtluCD8jocdQqgqvC74ntuE1Jno/vqN9OEqV9hQKs2
kCMOwQ07aSmpAAnoUvgt1VovHi8EFhubAil7/4e9o+ZceMEfsrA/SaU2YDqDyHGC
gQ6bC8boMfQVapzBIPSJB8hmYoSetI6GJnsEnlo4PUWD+Cjx7trcEtQpW0ego51M
S2GMyRlp6RO415IGAyoH3dRJqvFtCK1JNFQW/1FxfIdV2jBVIv6Yfr/jctE6MQeg
dUcPe+lIWLk1XlZvXpECO2MtA1cX63FuL9HI6zJyontdYlO0X0h9POoXIzUENNZg
c6nbTqtf1DfItsvOMkwXFRazE+WQ5gNGTmIZi2XHSSa8dm2SXDVClStRm4MinIo2
5iorLdOB8TrF2QuMunGofSEAk/xqscKMXoLVn+jkxrGIg6HyqR5Lg+b5SDGifjmR
2DSWF4UJKiFXElYOFtDSUWtJDnAtKmKE0zpAqJEPes94b5o0GSPoxFUjBfwztH5U
kuzVZJLXmADEkSMZ7SYex3o+msTQNnRGqch+ZnVpJYL3S9XTojuxToLJoU9DUKCM
A45owNWR4+ViScu9jsCnx4AY/lN/BPfL2hkA09Zw6DiiSf6Ac0D2gBcHbvmXcEjU
7LNBrDcfTQVI2cegMEFvQW78k9uvrvCREhBCduGRtdPrwEmVfApyJ3fHD4Iqs2Pv
14ICguarlVGdCQbo1Ty40+nockUE1DpYV67FS7EPIdAIB49OikPEMVuldgJGg0if
NwyYQXSxH5VhGNBpw/PQJAvSExigcqHnwLTxjp7JGt4o9RNuE0dbvf1GpuCG17dO
gXJOn2oKxMUY93OzQJw3A655voLxBu3xbJqVng5jke1xEcJCGIxntn48tFz98CE/
SH9IszOFQ+DStjTRgoVCWLxl3VnpKm39GdzWWwyr1l6MwSWyOcVRxmYu4phBfK04
H+d2Rf0cMoG8aWRnPSnjCM+ZibtsYyANiNYk79D7GChPgVKYKm8rwnsqBXtxgou1
RkeRpSwIrZ6bEdzp8TtTpdoYNpZdTz/c0TUGrc1WX7OBpgZM4Fk00XQqVmwbgtjf
MP7rUaDOz91pfgCoF4Vfr/jwjm7bIF3dHqm7MVx2SDrLbscT9E9VXobPwl+TnF5X
XlyDKiXKet/lcPdKEbG3S0RZRa9j9nR7vJLJntL6ZNBDsI1y7tI91uJbMgpx2ymu
I2oCuwePxW/SIS1XLlZDi5kLqzzvxQljt6BZkgQHkHkD6jD8OVOKAetYQjF0RS18
uInqtLDCcAjI9/EqgCLqSZmlzmmunQYyHodBSjyTeyZqu6KBLDiauBNo6ExW02zw
+0UDI39r8f9rtpFPhcqY8BdT/oZVeFv/yFEPptB4msIij4tTyOHXVxgh89DVmgry
TsgRf0/eIdvXYvxxMe2wdl4KHHRiKm9fQ4zVZOg+6Qkbh58ytLn8/e6hyoveegmv
1B8qq396+dtSxq/xvDsFfmBZUVhawsFRX5Nn6oJtcUPAUK/SPGQyfcZ/Pv1xNaYI
73N+6Q5C6m7mRoNjgO5D2tGsHCF+yOJOZWwveuJSuoyt1iEipMjxsmxcP/Z3cdob
qA5/AqyJpNa68/AFzTYiKLa4ancSCp9nrnY4K8VTPThuWQN8zNXCdBMke3Xhi6Ym
YuF3w/rcH2grPpQeWsLGrewo8KWwwSWdp/hP2yQDNW3880XGDp3++Lmu/qM4z5jx
wg88/DDs6T5YT9oG+FeeOtKITtiyJ2RgP4eMUMgF2mcJMpmPwYUdisGLqGCxnLDo
5JWlSBLGoVYnoxwoLQTIHg4iI9T9HQ1YZqIRqCMt6E1OdDkP0DdsdtcrbF0ute/Y
4HQhCzYO1zxbtaQwu4jVlqQIsetEl8BZuHLDi4XDw2997fJbGWzGF/mSroacpkkg
gZSDfKLb22I7ibDjZ9qq0fR0N/Rak0NmZc2ja7Z9FAc2+9MAbTyZtkXWaP2ryeTu
vvQlLUcmxJyPhFyHBPeadUhbVyVXghAkyPOMnbe/qNNWA8mU0ZG5TVIw+IYJCb8g
0J/REsn+M4SJCOA48wbSHQpB/4R/vVw0m/xLgcy8VA4uyyR/w+KAiYnvoPx1Ji92
z5Mad+TCdzYFmbJLEMo3p8mpM6ySw/ixXPgo66wevzas4fuoDrdvESLubYuHneez
VyW0CZPFcqkgvdJQyVThPIuDypu8UVkMMIETVeGafIVNxC39+IY8w3UvFmhJUuAH
gHQ5leE/heuatSx+0Z/30N04Sk0fGaMa3orzT/vCTSkJP0mW7Vck6qGO0Wq1QNOq
z59Mzi55SYh9wvmGOfivgKlDmLqHP8za8l6XYhjMhW+yLema7vCGnYaAl66VcrZO
YT5i4BwtTcb/mAP0/dNKuKrHd+5TV5CkqERUemOVoHDViHRSlYJbTDJSiH3uivrH
CrE7MZ4m+PsEXNZmhxRZRbUthF7Vll9HaSceFtS//PVGxmhMudiTplLc1QINk7/m
MGSqZ0s5bQFNG6fnLyHrHe0X7wL8VT1Bj+52/r3m6AZ/pjxhG5ldEwkgkKd/4JvP
fLLA4C5Wuzbos1cWJGJayDNPGljaoP2WwabFk+Uee1mJ5z7BMoyTxWm5xscDvWUD
d77yIXsLN8CVvFGhAvcBSOyxGAUNZxSURtKaJWIcxekU43xoRiuSDZ3osvAZToex
ZCm+/8G3nKZVr8ZLiBLg0pv/rKpXxFaYrhkuxQEhTIqxLlNlG6GzvU6gLuykulYr
bHf4SPpZsI5E96iJgCUdZlvsVEfM5+jqzRMM2YjseuebZKHcYeY7/SoikXQmeNI2
RWxXyYhbF9ksk+f3z9TSPPe3ifQloCFA2mUP9LIMwhB5flb30GAsAPFZHZwK2Gwo
ZexSstf/83/Rk6EwiAL4E4NBkzTuc55M5YNzPOhL2MP0MvWbGR9cDP1J4wY8fazc
WuTyDwwzK5aY2yFG/X84cFoeLujjYxNwDNlZwPpSVadj1v6ZERJPjUVfAukroP86
JluDNM98B6LHBKNVpn9667N67bw30iKI4NGPiP3UisPgK30gRso6ulqcYZkGiZ6G
BSswQdTUUbOgoRWWCEV9OaF3j+eow/Agpn9paRrFtzCRtRorTWyVuq3hqEkRsF3E
NAhbfilW4P7ShQuNX18B9y27Ojof0hluI07Aj55xeGO7JiQSoxeV5GuB6/6eW9iP
Nnj7XrUXF8Qi7wJubOVYJtJRTJATaZvyxTIcGEeIah5bqCYtSthTQ19furLGWoki
Q3h39lta+i6OY9X6DHeXSdHh7OiNs/Ai16s7aZn2ZCZ/NZng910cZEw8u+HPIbUl
OBKxo2aQecOEeHoSpl8ybORh4Si01R3iPG/pCEtsjyDRvQnELk9zV1ZJffWR+Yrl
1vh6GUAFB4au84pIG35N/mFWLxZrSd28o0+GwBRQLtnAS5HAPWW90E/GEOjsjvWR
j6sMEj9e8DLcAg3u7IvqCtxPoj//X3/EwtF/zLFdb0UrBFci7y/bDyXVl18CU/wl
hSiuIZ8I0mZz2GLvCkp8BJiQYoCYFHWv5PTVFPLzv71KuCEH0E6HkGTnFA704x3l
btLuN8I0mb9yrYFXTIYXPHj+x4TKknlA8YCYKW4K5EzCIFhSYz9rB79ebJxMPKwr
Df4f6t+zC5QdlISpNBZlENNUCSMm4r11suFJU9Pdz2OWy6RRyTFMwPEv5iC9b+I6
dVBDkkrqqYy56pyACJKc77NZHB4y52jBCQuz/9WXLuoQFa46qfp54T3J9LqMxP6k
f7Yt0GTCKiXy1seAKR3EEnWnWi5dIoKVpTvGCPQaok2smTYfA1v5lmZ2D2KXQBRY
rtIGA4Pe4ksB/+pHHrxcva+nHLszVBAbMQ+h5u7TBLjNY/lREdcgp3Q1Xs+UOY7t
x57YwZ9tx7+TdDQlICh5RxrEl0Cn6uT2qXfINuoC1+Fu9XzzKWNmCtJWH1CcRJCb
b9iDO25dOk72iC0eVrLZBXLXzUBHOz1xPCFOCwdHJvtHIpEr3faPqEAqbTaQdoCZ
kPjK/gOgQPu9LaUF8yxts6P07yv7fxzXATMJegXtIfZf9ycfU/XfpVIZgpl9a2bQ
6bZyB4BWDlbsOicgj8DUjNDvMrmq5n6dhKQSi/hJS4pwVRw1r4q+qvHZxXl6GwhE
f/+r/ZsYdi2INkImzP0DnIvtuzUrf77wnn8EX9IxYy15PmVI9wz42nQUh7/Tnm/S
fYpwxaa1tbgM3q4nArQmWGiQgCS4MivRVJCiMhlNxPMkO64AV8G2tuJVWhS1CTKk
mGBbPn4Ak+AN0/MIipnI+fjj8NzZVJn3U5QSwXq6r9rEXE8ggsapyIenc/wh+GJ/
60bSkLfHLPQXyYmJ1XtHmpRzKeO/ge4MUgJuiOzbUpCeoSkMbj8KWgedFHt/cvde
ZqocKaU/b9fMLlybN5utb54tvX0Lryed82Tz2TQKWryHjqSqZhbjwMvlFE/b63s2
pQrB5dWmVTx5vFOTaNSqKvodp94IJyD+GOARiLstdqokdcOq8F9vvc+YHASodQgY
2lkGUHZxUSrwUcUnrwIo4GRignNG0d3wT/3qzPPmohWMuUrZye1ZBd4HLrSgUqt1
P05onBDyPCp4qwSx5sUQW3AnB8/0tpMCtpaevQKMDq20ovFQhvRx+PwzWd3NuaiP
h7D4arPHwDyk6TD1JztE16hSDOI34vHRYghsoPS5aDknoT5ZAB8YsEUkBrCYM37p
qn/SWp/EMetjPAaHJDXH724tmIFx6LZ0BnJIxJC8sqhJL6m3sMYtSBnwUxXhXGuu
fpP0ltdP8BMSkimBXCjiIEOgZNKZMMY17cJDQF1Df8+dRtpHM8a/YRKu7EsXl4Ej
jPc1u7GYicCdNybg9PrmD+SRUbSoN7JUzXUQ4GtR2D1VNbdtTom5G938BBT+QS8K
odn1PO463ZXLSj1wMLuUc810dTg3hX02GVBb33J6IBnNEk7a9/evy/R1Se1pZlfm
UcLJcI+QjbhcaBb3YYmDI3Nx2Wj92nTPYI4r84I4QD0RSAgTeSJioXE7hdgfqLCY
iLUgNc+VvPs/yU15ooiJXnQPfEhhDJ0/nkIACKKATkFkv1hW1qyln4fCrDe072uy
Ja362kbyFztI3wZfcyEVWGKlMtrsPcGnhV4BvK7PlDxPxP7wg8BVyKRqiKwiPvKt
NKeK0U5IzJjkrx2qHLiUBu4jY+3I+RYl6vNBHOuVGlsWWorZ8RdLs1T/WJvnsmpP
wXwLeCl1Ek2hPFhjocSUrLavNGioIT+JbkEo/P2hoC98Kdrkbp/NxPMLgUOwGbPU
KL6HQ2kEcdiYtH6qx6vsV7TUMECbPm4Vg3Q7I4aPp/wefRVZRreye4UDaNtjzbCQ
dbmwGhg0Yme7LytThDhZgU81vz/4fD923rGWvrsliQgG5Ji8PytXJkRmxEvkR+BY
y53QTgPLfdCCqwQOiTZuCmBRPXoEaDZI3VfC7Fl8MtYvbIDqBhceb0Yy0UtrBCyD
YiC/RpdVHiTJMEgVW3PLweP1MUf0/Xv3UZe0Tr7Vn24w5A+tXhM96sIjV4hP9O27
0so5i+CK4b0eCt7Aqm+ysz9xgrO1kbM5542NzwSzyOXFylKXoqjPTPIs5HimKTOO
f3Qaiy9X60gCU9M5scWVSPs3Zv0FCrrSxf8n0Le9cIlWNDCifnA24sJDYalRMsoa
VD7UgZB3gIiuDyVgrVPM76xKnayUx2GERfg6H1E9a2oll/sniXMu7tv7EYC4Diyz
kmNegrzvxzc+wsQAmsGgkPPaMAir6LF8YSTBp2frXd1USOIhoiN6lvd+OkSXjhNt
1uFcEOOBsZObwDZr1OLUmEFct0d1e+QEd+hLBncdKaDYyfoFZVuP9ACi5xikn/pX
3p3lX4NsS7IuhMrXo3MN0qqepyIgaFkKwECq03MYT7IGhzr3CfN2dCnyLxGDKGvZ
cFcNKm687PehSXWd0fjtqsJ1PdMQCLjWnqxIlZPrZHXOaiAfPvfVPQStz9/EN73K
OlvNuTec+aSt2T9+jEGtQ7TeqGugNiAC7c0+osoaX0HpsxYZ6NHRQ5jzLxrKmBxx
EpMOBljIDaoaI1KWWp5tW+WOB3Eb5ttEzxa6obSggy9OUEmdJx9TiAaiDa3XY74T
wPAbgQRRq5xtYfWVO26TwamtQm6OoigtlilVTUpWOQdSrXUiRQXN55Tedq4WxvK1
2zytHXdnoLLIAen6VrsVA3Fsor7HknLB2tfCqhr3r0UXpATTNLTLGPfAWa2ub3nA
R0cZmEGfSgmCqBu11QkyAG/nY1uoV8hESGPYu38RN94P1oqHSmlpabHVfcXUqRq0
PBC365GOc3wYxZxGAUUjWHpxS/W7exMfHYc8urjQRld7f/Uj7rfSI2ewoClptLzY
P+TCMBZO7S3DjJIjQT9MJ5bG67Dl6YOHP2QXy0W3Qfri2WHjN2jCf0kqM9AhF7DJ
HxkwFU2cXtJJ+FYuIoC+i6DZkqk8gfrhpYM8I5nKj+e+1aPHEgnq5NpP2IsxT8/0
dd2j1pOZUeLu56kBoabnYnynRG3Zn/hoMZJoHZst76LBHd094FG4gvo17LIESC/v
urc/vzjx/YYl47HEQjlL7a2QF0AVqGb9rNxaxebq2iluiYCFYNlmfWd///4HL46m
BmBbmc/fiyVxp9Bq8zCV52P11VX9iyDfA5x16VdhxQDtB7NZx+i4yksOu1oy6c2D
XPaKUaP+G3NaF67NDuypMMHLdiyYGUfr/RVSVDR3cX+KxoAzWCKFaDvgK4OHgsBn
ubILz/q8OPO9RKBmZ5Uh9QYCuh2Vs9uc1WuroCTY+5a/FKrUQB8BMveQyEI7mOHu
HTu/bgY57wADgX+0Oava3zPtlm98CvNOqMD+7JspfHnUrAC/HFwD0NRR7WPQAt50
vjBYd1lO92D2rk5jzKeeJqqiOO0S1a4Uk9DnfW68zbK+ywX6ZDoiWVdf9erXCMQI
xJlomDq7HTGN2LAZ6e/LKMG9B5w7RfB2v+2i47/aoEwA38wtj9m3ysF7S2wfAX9O
wY8oWLVL34k0V/YFcyROLjeiqs3vrxACeDaRSz8zowoekQMZx9kMKTnf/P+ko6FX
oUbLN4ts6SsxpzutczUU8IJELo3P812XoqVqFi76RnIT7C/GfkcGeC8MEzJWNG4U
NUK0O0e3IoTqPsTnakpe9uiHlTXB50J1id0Mk0CrHZCEwPq1ASlGsZntWHBByLFT
VY4M0M5Qxft5QokOlUZrKefhvEf7ehYUhw9e0qnldv7xa8GIsub50UDHFhq/2Zse
mn9f72jRbYWl3AuIIQJ7ML2V28IDbhmhqCKWHCA4b6cAsxyzqVdgSeQRjVjqDrLl
+FlcSok/cFzrHsWThCtKY7SrnUpQch9mNyn7wEUNHBeqg+p9u/vC7mYzaZHYQtRO
XpcNNFXeDvJfB+05SXKwMRx5IVtRZStjDxKxkAsf+qdR0VOcG7UOj2yQEXmd+tyW
MLtCuX6FpjQZBYp7IFMjCM1Ljya7HeW7BZgfpLIJ2zpW1ZFyglCTF39hgtAoT3fB
2NuldES0g79RtN2Ins8U4BEPVJjQAJFi4HbFZXt2+sv6ey82e4iRi7MrYKhVoVI0
FEL15NMblNS3kqOjI1iI67c/Iu1TVLhLAf6R/vemy6cAt2arNvymDRB/D/v19LsI
uwZx2EmHPt1xE1C5xKqM3eWsKD7pYQjt4EHCkpBcwdZPy4+Gk5b8CJ5d+opPWb5D
RUikPH30vChY7f9VhGo9jsJgMNeiMmz9Wq9BhLhnEx56+lkU8kBxN2dwd9RXJ9DZ
GYkZUKiOr4Jm03Nf1HmXUGJfhR9yaA+nZxPIIjD0F3gsqb6VmXT7VRKVGtnaa7Zk
9AJW+HaPRqpokO1BSv+cwEgMrDbRAHGPmB+fYOBxQ+MYj3FFlnA0qikP07kDxplC
JiDSQvW46LmSstF4aLeV812iN9ag9x1fa6WRksuggpYd2jMdKadb+PWawxs9Iqej
tP9qcKwoDVmx7CsuxHDGgQXc6q2T/8JhR4IfDxmNbVFr70LatlmB8UUW1FvDAIOU
9goCaSEToCBW7xr7gFLt1eW/V7CxxPUMROKt3F+kFT27ImbdLdyedwMFRWpSqKTf
6XGLmCTOU2eoEzhQOuOlWQG9Q5VsqLoYbqaFoOaTVXKJu2f1b5WZZQ9+b56qPzMW
W9b7WjnAr3AtgUPr1JuUj1XzHUXBvfe7iwnNsS33Aexg2JOJQm9N3LLvv4rjgK7a
gCsm2JDgvNJF33GorYRPaC4IHRC+PeuqpIcVzIjAIf2hBytIKf6A3IRuHSSZijiE
DUHp3fRtmr7vnGJlYg5z1fq8A5jQro0NKqs+OV2LwneUtq2Xz59QB8iv6ptUpyHM
l8oBSoqMoe0hpDZNYr9bTtE36Zpm92bqxaE+S7xu7mZVDORzVkY7ntMNext/9Msx
Z4SDIqs3HoICfpAyRZfb0XWw0SWyiNmYfeWmEsPSdK6YBDWz4eI6mD5xrcAcmext
ggEo1M2uj9ScGiQZCpRHpOwlGL1m3o6a1+hZOVD3EJfDWOSqK+s5okuAuNwhc+xt
iLBfj8WVQXFpRNfOeseXE6hWpr6dhiPGctjacDYXSaPz/5NGkS+l7SpYyIj8bSiG
9Gl/oRsUUxdIebHGm2GXz4kErqQ76d4U5I0vqJqetdzbAF1REwJPpwfeM5P95DY4
bdwx/XoXO605ApGMdzsc0Vi3i/YZ4LTgYB1pg0XCxvExS5S56bpEaWQJflHHw0rx
5cTYUSJzUY+kajA59kZ1ddgWzw7sRpwV1T/NMJOYFLrj5UXa9sqq7txkVNi1jeYh
afKyFWGxJ1tgzV9lGm8oaZUFFW1CRfOGHk3snxofIbdvgDTUvvCv0kIzpRYFdSyR
7XsYYsbZgVMBbUhiKmiGzkYVajOFBRGoRuu2H3kTz8QwhLgD4wlDjUIHPLAGMoKt
Prjmg9dyueUK5RzunxYzee6We4VQmDriSVqcKZyyD2DwlCJA3nudyxCMAblb8Xdj
0bKJlRnybghPYw95XDAUj7zXHsKki1akKdUJMDyAaFywScE9Hex15tCp6znY+0bh
kFRbYU41PuqYbQ0/4tbXPY+ugz7NVcjXJ7u/eT6XPWd0YCVxG+cQKQNCHGbU5P2v
RhrjIUY413acsSd5B2kSrBugAYR11xGbxJFxGya4bz6g0W2oZblndCpITAbiCDBL
3hyMiU0q8yBhryavToFKE3qX2MB8E58yT7YWNPK6DlbGZucbkpDob97tfy1lbvr+
Pxgny9Ue0BalzNYoTNPwpY7X+FboMJmUesLteuR+yRQhpoccjaXEq0meIfBLfn53
3nu2rDELPVGYFJomi4MCIjKS1UEI5JS3jmvEbF6ViFFR6cYkYZpN3mnQNzMmtiGy
mziWfd8u5jolJEUxJOhm3W61R9qH1m0lcqYfqE/CzKk7NKxzJyP2h7XKnygrosv9
rZ918NyPPkE37MP3h1wLVVnfmloSC3+iSJJAaHGvj/Hy3hSGa6hgEKL/VIHolqdR
YZ2Dy3mF0wiD2HzDoiywbNXgWq/KIU6xgPjGHMx085wIRH+T/Urud8696XZ5hUq5
6RcibV12xCnLosE5/k41nBF/R3IwygoAfFvpR+JdkeUIuooMk5WObJ4cH+nRaWF3
Q4rstE792XkJmaytlFG1eM5WvpTQmxn06iVIiKMyu7bY0nes2nDook/kj2+GCQaG
gbMYt+yeB0a3tZ7K0p7hNXokoesGFOS+lZXqGlsV39GI7u4swXCCN0w+7kjB4spJ
C+j9y/Qek/TE9ymlWtJqcAG6SLdHOVQJu4GWkLpSotVjLemWPzZ5dbNyOtjmRTRW
nUHNJhksIQdf//xHUJzbAuu2vBuHz1OOWMr3qvLJ7kKJvfJEkcKzeakfaHTVhImp
/tryaeZgT0MBxxZ0OVDdGIQnpKTtZAB6M5Yru4DTlJzATHnl3I9VAOiTaZAban7k
gLGaVZz0FEF5p8Za5B7GkUS1yJL/CKMqzZCjmRrhtHQH5KPqNAqT8OgtBCd+QGtb
jLr+dNBe1HB4snJpNBOafwshDwB1edlgcV6/wY2nLF69sjCRzkkHjt2T9GCQ34xW
RUmUkuYkG9l2v3irCUDKjOhGidaDkQuOkRxDELPnJvnDamtE3XzBD0/9czrv8E49
S0hoeHt5IGPh/h4AJ+3U1bAXPaJTnLYehP/Dj7s5stdQhbqTk/XO1IcFSDue6CI2
J1kBAy0nSKWiwyAiuVYUCK1p85AUkPMWp9C2OOOSPKSYyrnCP13DgHIfAUVqOvmd
1dqTnDp1SeEDTpPC1T49QkVWmGX7XzDpcPk9+mNU9896q9ZE2Yjyf80k4M3x1yue
FdFx5UElEmT8VdOwvtLyIy+mbhzb08yCxk/GJyqmECfBy9i0guFZOiRu72OTdCgV
t60CHvo4At4bpuvzHyP18Ww/YC5FiRsN5tqmlKfryT1SuDq1OiKbw0Ntt9zjuVO+
M8ovlaNF0riq5glfY9qeI0RBfKGHxW11hR3BhFqF7obgVT2HqlxjNQEojOBkF/4c
PWjF/rDj4qUnsKF9qqJRFUgvXth/icWZq38OjinpphsPMGZUmY8lYTv0+Dkn8tvj
mhmsRubIvc4Td2hD3LBZ14c+P6BsSI9stOTwH6p4+DgWl03hIEp9m038u7gpfkOf
KemQgjPwm2028i4+QJc68KBbYSHauVOGlzLXJ2pwRxBbswNpGei/F+nRlYgURQPs
crq6NX1ppzTT34aTkUE0dSBk1c7IH+IyYuCY5yWzdfwq7L16VEmLBZYS7JQ6d7JZ
74m6vDdxs1GCcqsj/1+yeoSI5sAj85OxiF3PqWHp6eJGEkOaYxmshYnXg04i4KH6
t+P6GDvjvwrMj3FyF4zCTCQ5bLsZlzjZZp1kLM3Dz+D0lGL+zYIoYeV5B/FrQv+0
xFEf/lYkpCOTdvAoQ9STCM6dME0fUMSgwNLrG1ZFWmy5hFIhO2d99kJC5LEpg9Vj
395XmORF1Al9duxk2cHmBoBoUjZ3rsLZfj2cl+D1wAa6AkBgoNibTg0oAunUM3s5
PceuaCyE9aZCOkR346MUDXRTN0/OPksYSzkdeYARpIruCjw2KEpm5l8wDC2jXU/8
Dd16ZqzXPGZjGVptyGYSJiqpf165BAzqqhYCKYzMF3zqVjteiEg8rfArpgexZSX/
x7ehDkn0STgSAAyUqTtJ3XCUVbMbwHSyaIeIlvuvzfqYw4SQkSdMYuodSl5xmw2c
IYgRPV18RQY4+60RSFFE+xRTo+pLe0QoTI0Wx5x8vz5+ZQ98JaLgCLVI9cZgVtH9
jc8NnpgsVy2CxDZPepN+ey5R4dZVMt2JaV/jDMMrDFiC1qTkM8qepUKUJY4Xfy/S
MMCFWwrLdFLK3HvDakWDjx4Mk5QkC4I+Vax4p1RUFJoGHA7b0XEojdPqxquF+pOG
sKtgoIqxgRZWVLkv1h71mTTI+vVFss6TDCWvjsir9AOQ/Sa1x3jcCp01vGdP/OZw
/ZM68ulx/RfmtwJ+et/I6fgScssZLkrWazuiuQfCN6DJQjESM7Fi3/9TDMEflnuw
VZ8YRr0DT+Qeo1lSCDwQ7o7EjQ44YYWIPjTQFIxazuR/KeqvJvEhWnUE+f/2fIzO
rlZkoWkn6t8Z7yiCMa/z26D6Ij50seFGrYMPDlj7SQfGwM+H5yX/kXM+VVanMRsh
PzkRT2Np7QcVLO12o0NNhy7zMfy3+CarKPzIMNLWA8U3oA92KpNgRyJ8Bn0QU1lL
374QADtn152JDZ1Ke5v+HPVSxo9g35luzYjWmuk7aqiKeFgvrR6Bsp1WApA52j5P
6oDzDvbTBykEIgtglYjXDrvGHrENLA3aCJmYlbAuELLWSPg4JQUdNbuebfvjyEL7
CliR6n15gW/ffMoEIZS1/7lKbNIlj7eWsV0bLlxdyCzkEjCYIQQuPxtP4nrE1T6+
5kFI0tCJDvht2uQu6Wnw/G0vvunun5lwO6y0uQDkg9Ro6THdQci3MUp8QWwaDx7U
/bGHrgfT4SAuT/MEW97n4TLxxE6TW1r9cEBcp4tj1XK2QRd0MSoSqGkGxVvKFy+C
Euly2hHTZI1byp4JUR2xv6fg3VuhzLb54hiTG7JlVMc7SUMNMjiuAejz0Xs4iL72
UhrRXhkY7jGwefI5Vlh3y/fbUjtvZvQagJ8WSIpCY/pjYi9kqynYxitMsgGFFmH9
5+bpbBaY5WgY+q3FlbeN7wzvFTiEujKphQatsomQr+iOg4K7xQmizkXNJ1gx5Rep
gNIYBCoHr8pYt/lZat9Ca5UwyKxe2VFT4YJlDbXqGXK/XfTf5HQrMNBIYEsD9qm9
WJ1ykj9h9TrK8hfsCKY5i9FOZ2GBf0lJoeuEdaQB/cD3lk4ypnXiTZCbTaCwny7p
qxpr3jO4dclXTGP0VXP/Ew/bI0ae5xVbGMZEiC7hrmuVwQXSJUZsLGiQy3+PEjt3
bEoeqBIGUUsnPokXgeUa6/1aJAm6MHsaHepKZ59PYqseSVo0bwnDRMEK0KcyFpfj
1rzhQcLh+YYb5v+T8l3u9QqURAzRnrGQBOMtzDxfRZdv9rP6U08Yr/b9EH5Dajoj
0dg6NLlXThKCX78FMQIsyKBF9cbKL2l0WjTePh1+u2f5sMb4mA83lg0hb+NLRUVw
YJ9feu49O9tcFCjMXN9Mb61LT0kAhIRJROKAKnd6GhS4GFVUmNR1zuCs9xT5q2Q7
yEGFaL+tkHtBemqCi1FVPfQve7wZLVRB+hGZevomrP9Ffw4JQlI2HIJeo062BEoL
w3Lo/gUoAlm3a0T8RbwKj4tUVgBV1mv3hXWoAQqeCfwSJqs0rtdfVr2K7CjdEIby
MjddnKHXPFXs7OZF1S0GP8jRllrbZBmnQIP+DCm2489hfeX7UiUUtjWsiBR7QlZH
qEFTvp4zznjdN1zWQaTuET65bX+TTtr43s7QWhmAVHyYBkAMZtOGIzIRpZOnDzP3
GAc21Nfzqhs6uEOHAIYoGTwpx9lPNA+rXRGMYL5bPxBkrOYspXWFfoARvQXjrPdi
ZiJj/WP2FxSsH18KX08P4baXNBevigVlQAGh8SKiMy6iP9RsJMppAeyzCpZ+2vgJ
nuf3RR16cztDDCBJZWQDRcYD+xPjPWxlpvuryeJ/G21ABonRqDA0YdHm1XtESHZ5
GuDMSQaCcb9sfLwA8hkSalizFjeqmyhIwinZaVP4KruH/Gmy1JIZOb0qyyo1X3F+
+bpHdxR37pq/kot+e/n8L3xQoQR9mBtR9LuO2XZGZ8cZsk9Poal0v+RYmZrvohE1
HF/HTNMIpjzpITpyuyGyGiQPGwKsezKPvVTuT92X1oe80F005/sAlgovTVe3kqFi
Hl5thjZuwpDEJ6+mtNOV4tZHG/Aac252JvwGKwRWsoglEWasI41c85uDgSsI5ve2
4ZaRkmP5yGWGJkFNRRG6lcdg47APEfHe5cwfKeJwX3b7Z/gLV5Q8fZAoFpOPTwcu
ijQ27yzZDOezry+JFalgfSDYLSef7UH1ZBdahprpXBoGQPe28BO1XWrlWh9kN0qd
SojPO724OWfPi6+aqTT3otZwQOPJtdw770XiJnFEdCLgbeVAlSSraHKAtj7DoAkO
Lme589uxTp5acAMQC+6dAs8vQ3dLXk/ozE9EZVU0nTQ96g6z+8HpdYR3IakMfRk9
EJgn9/dGiObV6sQUNu5UiH+wVmLnxAwJnhavLhtpOmhfsXhC2E7MBGQAh2H5hDN3
DtqqAEoxxmOexeiF2SoHSoel8T1e7c/owBDJ4ASEtFEHlQLGUhkhXF5Xj1imvOBr
P7inmWhbrb+JA7yeET/BFmi3M7P1EeBN2UNuFULXTmdEDrvmW0ZGxK1aGSgLQBnF
Nye2qpzHU6acWAtYPNZpHBmv/2Ulc5eD87AfEAjgBm6AEhoQz1buOeaBc5QcZTv5
/zeD4zlD1KA3bR+mWE5jYufcEckL0qUne1ycgF1Bt+OhoRm+YvC/Tu6bBmD3LZOD
QegMnkufqX9JYpEsGnaDQh8SQNtA50cTa4LOc02JTDHcWw21EwVD7ejfztMUy2N6
EHhO3bBg64XkNV6z/kKxlxpKFBkjE5FCAx5a2nu2x8uY8BcaAwxbYz/xFchTcVJ+
ilrDTBzxVrQjKpUSpnu+MwTHAbnaiUu5I18w6nNImcG+Ihg0iQfX/ud3ffohFOWr
FpeRNW70mSdwX9cHtEFnnRt2SjDo+7rl6jNQvK0ATyo/bWhQnRSKmWBkIRFoJu+h
RGHZEq7PXQwyf2n5UqFjibcFKD3cJZbjNtGwRJjOoIij/AuNKG7BaZlDGUnOCH51
AOf7xAuJ73cqsWelXPt3iorpn5+sofw40Ly7/46ysKlk+4W1uuGHbuMaoea0Qk/T
6uSKEHXMZ3yG3/8SQTqAmoPd5IG7tFVQIRBXkOnPuXow89y/4oE4fLYdx5QfI8X9
4Og3p76HYMit/1tKljzUT+c6TMnLmL2Sf2LlNZ302Tux/tZhpdpxaqE9/0tupE4u
ZYMxtk3yXLRxFF9f5T5vAC1xYJGIOa8N7bS3N0M9bMk5Q7JV+/9iBpmB0rM/2tcL
EfRneGBei3+AJ3gpnQt2zrYxs9tgMaA6cihmkVPaVmp1uofH0kwJpAGCa4qU1JP4
MFvq+GrMT+gttYoZFpxI66cqbbJ7HpMuCtnuEA93PPglM08ZDLI/DvxweDEwWJUU
aU/OdwIs3fRM07l9JWpgZQgACSBvRrRaVFSfWGdeLeTyLRj8vQmMVBdg2wXWCa89
FBzNR55actkDvF/WG4CG6SD+mn1GDnROY7e4C4aR4rAzhkFiM1HSsYkI+wKrQzAv
6YBpnWJrFafdDcUsNhvLD6SOa6ZsSHDLtEoUZlVLLRrNH9YVAJv3QhsGQDpO3rEw
D44eOps8BpWl+JGdT6h/HRLKf/E5N7O3dEHrIMMny/5G4rQgRUk1kLtd52EXyCPt
PA/f5YsPv5hMaXZaCfrkrg/VGVp1XAem3UYBM8gQH5exnZRSL64PQ7F2xvHO/++8
LRDIzOyjjEamMhgNQ2yLXD2KnG7RViOQhXweGXqIXvIBCBVp1xsKc7W71Fx7uM25
3+QAZcoBnnqqidXkmjUZfF7w7kivdoZ7H01RWtNfdXlV4Nt8U0uHxq/G3pSBapKo
sAgpD96P5YxRlergqRoomFXrSqEPGO1fRRcRq+3aguDpt+pcY7YJJkLtpzhMu/gw
lI9QQ2GNFZLJXAEVnbeleSd2F9m604UwERRgAwieXqTENm9nqxWgolIMOY815qLv
uD847Dvp1WN1QJjzurwBNPoqAdnuILyuORcJeZqTqFQx+mTEBadJ0lvX/dQenQ1o
ZTRafqAzyTlBGAJ8Fb1uhBmjOvVMq/ketvB98rRBwnEWUedjgcgtx9uZPDDwe1LP
HnS4eYSsl65t2UwPp2VszKBK+P86vNGen5XQcfu232EZIVdwPee9gZ8Us2EdRJxD
t5Z2I5vCt+dPywtp/Ir49WkDLyXRtx12+T1c1IqKriv8EZQWC/lnPTedSu2/MD+t
AsI5tZ/w9rPHIiwIUZv/tt9S8CHMUr2uyNqUMT9ldVHWj5gNctnMmL6dwhP1oh5D
U1jKzJdDlDfQhooHv0Vo0jEx4IjPtuKCEcF6KzOpII2RdCnAV5hcSoQJhBsQrl0S
dC0RklKQWmEDNPw0ZZfACdqT7tRrEEYCWNn6DrShpHDSMJXYWZPU0PPTHqheO9XO
bVk9augp+zpgh4/Nm8wR+qfnUPeJAAX0QhdpmC0UQmHvYK5gWr5n1dIYiRUwwaQ3
qLBKxmgFwLl/ist6H38GHI89+bBgTksQuIjQAlaVR20pS8RR4C2lCoJpdC0l5m2l
eghMgzYi+fchmuBhqGG2wv8zPNK3APunEtherH33oV3Mm9o9WZpKvB3wIkzbtHsa
MJTyUErkTu1TL1FgRBnOwr+/xQqTzWjHsZEkqBm+U9cWr0eNSV6awCgVj/N2q83X
3dh85C2pHws6d+0bYq7xqaBFZuz0n6FGpDOiJBhB2R4Hr3DJArmg4YypZ1kfZ+VA
F5VV8gcGQLjwVXE/xcmcglB/vPzzsOnb/i9MBUpFcRt/UmAYneY8wqxDEtmX82P+
wrouVCO5wev+SdKtt6kamRAJeVsywjYCU2mDZga6wrab5E8217b4pVELBxlBYNfc
ngNVWfbOcd3HeMqbBnGFlEvBAo8PnC3V8QA4gybiQIN6PalFC4C5vpkak80vELgY
2LehrDBVtB43hODYQhN/jh11APBcT0J39Fjs9HDtD1s+Kp90xaCRo93ovOdmmDmZ
7kLSegrwebqkyiRlybA3jrhFLP9iUfH8s9ZJgS/KYSXt+CQ0DWL2aC1vFcpo4yPc
+j+wNKplEffuHt3AzL07OqF2419vkdhkZ5CMPulsZ6NvNnG/9XC3Ze7i8w3IAK+6
GYOTZZP03jltKQXzaXHVWICCZu8pI2x2L0mInEzbPW3K+U6K/UBlc8pxvML9nvqu
9CLUCtcl4dFhNAoBC8hoWH8uplhP5WMgcWiSTtbfDNEsUiUfPWSWBao9bCTWThct
xNjgZjI0ljVdr7iRJtXQeC1tAkjW/31jepW+RUjR9lSGEDyTZBHTCwgdmrv00jo0
vV/EoTlJ4twkTbJRAfC1+FcoBHfPij+35G/+f9QDD07YMurC9fBumY6mUYBR/5Jm
4yqH9M/KbvGPQ3piLCQhIC4qKPHW+lAU3UjcErDAL9dIvFKNOdvcD5elRE6vQPqt
QXjXTGtWqHsSXAdN2VSL2ht7CiMIRTT7K96jcYky+W2ALAz7oiYyUgv0VdZpJ6SA
CX+FF8PnNXoSji1F49OE8rVGV/F9JPcFkafxvAWUszhw5TauwigotnU8+O6buHos
uFnVvRIKn8XTVSlu66Np9Tus6ag231oFsNS7B3wGpk/1whg5d+42IsqXYxWOR+rY
55G3RL0f4twgsnmWt4BHklQI0P04tDamT3+S1hbgMWeDw89io9E0hbRj/eXhqjh+
HfMdUYIStpP9aTR/cfPaZ9uCrgRgcbD1pbYDSFSUdOWPe4ZiqlSOCXlRWw0WXXeM
hqI92PmP7/EnZLGk1dDdW1/IiTBR2OF8BEJe/2MJBitjbnlI6KhFGIAMKJ6p92MI
vmwk9CjkGDo6Y/onfpwEQ87894mJ6Ml6HMR01DO+gwITW6BXlXphhbasVODCFhXi
vB/j4Yr6z3ZlaSTL7u0iqIeJS5bWgPuD3IcBMg6k46nXxU8my3679G3bcdESg1BQ
2wdSr+dO8+OwyIABYmwG64VqA9q/CfRT9qM/ZFVCdV9KjyA+zOfv9pHKb0034WFf
tKi9C775Zqg6gDDvhZ1DjNR6/8kjTLqEZ2dzdb5C58ZzgUb+4rlLcJghpd2fsEkM
RtygjnIhHVnSnH5VUvZwGBu2rDSMZsGVwh8EV6/lN5I+OitsHOOQ2ccs4If2J+8j
2TMgop756DVbH7/T8zriNEq/JmDG8IZEE4dKY03pwfE4aSLBB/Vcz3SWQYLfc0vK
2bUuuxaYcwB7POZKuB4UUbQudT3Q4twrWGoc/rC6VOZoQ7qamnXngdYLve4FzFzv
kkssk9O6AXKwPZrq9W4V+FWozUNgdNj/GinMI0M+PAIMwwad5LajzoAQfgeZ4vfh
Ulnz2Qwg/S7OnAEbKCifJBwOpGjIVSZjZoHOOlA1MbT39xNSMHfj5LFawWTqbjEo
i5CZW5sZgQb2EhrsBTv4X9prcgSLBWI6KbWmwYyjwtshLJT6yaj0Ohe4bjLxmUgI
wOMO1MujM3AoYTgmdi5HNGJmRccrWXb0F91CRalDonqT7tR5LrBWDMbdSkmg8iAX
rePHBTMUI3NuG/tAS9Ai2EXIGq5uZYjRVci5sVZtFkB/hphuMkRMo91z0NhcB8Sg
BZ+hfDbrCQvz12YWQOoUqCbsWaS3r6D6VoeVxQxj88MWz4ZsVqEmY41N2njaxdW/
eBrD3PBwo3G5Mr2Hzgv+XbLDzn+agzD74KGaM2s3rPCBRYvZmDpGrQ7mOz+pHmOq
mDfnZBdo4WqL02H+ANHyH0XyKIp8QLzjlBQbN6CNyHzukACC/mltImIYBmk80wRl
FQGcF//+nx+1SZJHD24w64AhZFkEBuFQTCVuADQ0XkR6u0lKslcAIrFLohLmkMSb
jTM+9qf7t+e1rMpzdFwCwrvISwuFMlFgPNXXWcIxtMouLvoYb043aK+wMgKsFWdj
9V8t5O19jUpV30bhN0IKhLrczNdt619ZF2YrXMr+aJ2CzI5VU2nouMhpkhdVbeVP
ZqtGtYdP8m8sq2pntxQjSBkFmLQ+3i4B1p8+R5Y2CDVZ/DQWczW4PE1Ny+EWpb/a
wBuoKt3GhMkK+XWzVqMbJTwlJnF/qtjMovW2z4wS7axCBrigHcSViMh9PRCCr3Z1
pqS8aKkwnjXcQ6eklOaR+LCIVLX2ktG4Sw9z/5DQI+eP5K0v7xJ2OwWRnz+vBWqC
Y2eeCrCvhrwpMlg5p4zu4ggd3ZdQnMImg1xyAocnSUpmvg1eWGjORfpsqaucHftJ
y1IqU5lMJVVGPpTfhRqdpNbhGTbFKWdcXrORcI8MALjHAYRBkN928SKkbChg/6xI
UH+2sHPF9UWbFd98j4Y1Wnt2I8CUQzDlMAZwzdRRMIJkbVOjPB+lVm6OlJR81Uuk
XFwV00YwrwvqxtNPezf5Y80BtEBpk3JTHsBnIkTp1g59MFPHJzeajuz+b6jEoknk
apUkBL9f8oTO2nVhqTimSOO5ySh49z3+P96MwgfL4/Y5jeYyhPSsH5cC+P4qce1i
6mkq5adRFbIBKJ9Uu0ToUlSLCgSPOvrY3ZjSpxPsx5mmT+XbQKljLbbcLpx2o3r+
wjH0L/hTww6n7VDypGQpa0B3Gx9xWACb1dU1dyZWbvj1dbI5nLYxsCI7Qi1ab4xm
Kswxpi5teCMKtqXMCURHUEoRlHmdnEuwOieWKLds0UXmEPcfK5+fup5f2B5FI9ah
xocrf3N7niepuoApeAS6n6UkbRO0IVWlidF8tlaMv9GbOe+vNkpq+qN9YH9hiAdC
co9GwsBgvKxqTcQNCHCohrzAMEYWatTaTld7Fe1mXYplwSmyeDt+awQjt4nUCeu7
2rqu5K+scPUJmHPxged95FufQ3KUeLpP7Gw9/9/7eeGIvx+R6pkDMu3Prz0nWMTD
7B1/nAC+slRoqyXX6/4h6V97Tx1V30iyeN7IJ2MS3BtxPbgBgeu9DshMrqWVnIcY
UqXZ799TYUL7EeXpsvBq/Yk0iKeTCLkUQT1hNJxUZ/uX75NST/+flyj064i9ydJm
lPHObZDaKgQkW3ZItkESpPoCWHLr8gXFBZXQKaVvW2qBsaIQ9mnOO2mroMFPrbFE
PAyt97vZgzD3+JDKrkE6l/lULgvpVpFnzE+GmOdnKnn386M9PDnmqj+PJnt+ww8D
ZlL7uf0PmZKL5UUrE8QAfVFl9VPsZiOEkpwcx5qD9ZM2nRn1Cb5Kqp/NvHnbkV/C
K8KucdNf94HACScwL2Ly4KSyM5ed3vSwcoIcJLNoz5tGJq2jgKbJda2ysThig4Cr
VsDbQvdZBfPwnQax7K7EJ2pgX5JFS6oBWAnov7JwO0ZZSxUYeGzHMTSwMmqretWv
Ml89Hh8Vp3ciVHS2COtqm9Ja8uv1uD3J7yck4/fqo371R50pFQqu1KQsyHahU0i9
7Q1G1tyDHFrAnIZohtqM2sM898lny7j9N9St23dxxD7oMr0YffWov988Tg9vteRG
tCH/qnAH3qCND6aPRsVhspIqlQUn+nKXdsmIbHaWxSgPtK4+VgxIMa2JiySG+5gZ
5l2TX7FbwRnvRC2xElcEJ3nVbO7RiqNhLWGvzu8ldyh1kQ0SutJwM+1S9yaI6OFO
bOmSmPt7KoCwe1cRC0F2exAW499zsuUZFOuT73omz8tgIm3N8jr1sXVRDZi3rKaP
P94Pxz5dRFE2XEmAM38MVDgaxSPOPanJi8kdtKF2Lm10HIyJsWUBAvw48XjShyhe
XMUjJO0+/gUyXHxS3VyH1RcRkAB47y69MB3mAYVI9FOUtLPnWIdabT7C2sx+yjxO
eC9SVuUg9cRY61mzUqpOomb2LdKHX7MCbba9nIz9xGVceGQ/KF0Tu1P30L1gcc78
ScII/XipF3Rb2CfArtSSYtQjbj1UrXsiWeg30Np4Ym9eW0jHUZAfXvBW4elM74Lr
xlUuBqt2xerdtCpAFH+B3IBjIkAANZ/HYMSpMWkf2+X5ORhu1A/neiaGu9TmbZg3
43U9peK7yjJLAuwOsLGw//6thsOsYBOXd3rHwkMA9XP89mTX6t83BSh5NUkIPUdR
Ja3FfJSMfi+1sNYHnOxx2bVBjwQ+kgyfjJRBxXi29pvai2ZeXHgY2d/6tSnLOGWe
whByYMsKUXQWkYku8GjTNtnsA1+61tIJp59l5V1O7Y7axC7eqoAWcssMRwun33KW
o9pU2CfgUqxk9IihJ+ip6ci3QmhsgIy75ASvs1xl9USbzflXyhuhbz4n2udzuX8a
0ORHj4HADVRvHfDPkQluBlN5cF41ZtLCEARgYW0VYPEuIVDxvoVnXYXxq4FYTU0+
X67N7XiF1W8m+r4i2DZitkthtMKhUSTaX1cgkfvgrYaUyo1EO7aBj/PXvEcCwIBP
d5obYVnOpcTWL5USHkRyZXAzxrSVsCg2YvIO60j35KfGBkdmMxBKtviiyekVudo9
zeWx0S1yypb16WVblCUtDaLOJ1AjwvluHTNa45ManlVa7/5IglzfH6eHyBp7/xFu
oxaAq0xvhKWGtXXbRy9IdjP1HKi57Q0Ui9Ug3BYlh5JrjaOESuTczuYd3yEx7pNe
bcmGNyijuk30jDKfrk3UEpR9bbL0znTyG3t6BObbo4StYBu2dMFO3VY9bLvXduEG
s74Dj5mYGv7mglvxW63HP6OQkgCO/zYkPTtjoOrcgFYT2JKG6L+R1w2bGEfZSnpJ
CEdM076r3su/9ewa/TPhk+NVcid0+FIwKACKhncQcy0dLgTtxI8a8vrdeji4YxjT
Vn7x9tXYxqN33RaGrVgTKwXaTC9Kr4QOEKC8Dpu7kXHOwV4ZqHFxnpMpAwqp5ZBd
0sUD0Il9yn+MiZf09neCIbaRKcBWLFPM8gEIGsSlNWAfkPJzK0GUlH68MegMsl/X
guDHNNIBn9QmfHSgJ2G01oujcXk384qOrTyzR5Wp+5HFBY4qije/MRRDlhygOe+Q
Bz28mmt78C4VWfxiAJGMczqwcKILlXDf+c+Xmug4JYyBGRwHbDyM9n5sE7I7ACkx
DkwCugh7MsSi/McpBDltGYh17HEXhDfx14AEVmvCKE0GRdDVLAqJPHcEvQ9s4Wxq
hzmi2230DBvragu4MAMHawuw3+H0jXJ7FPHwfhxEgnboWu1yNqFMOoTTHyb0Ts6n
fj3doWkuX+Jkh1GHRst2qEMVICm6kjG0mVLeugbKNtpJ+3/jifNn1hgVxhyuioK8
eYBEgSk9NXDkVTaoVtJBzH3rP8nHJmjuYsGCTX5+t5D9igruPlysJKEg84OiTZQw
ebDgM6SS3RWEzre76bDPVW1WyYcqXuSEpSSzscfQsP3o5IBoCUpZpfOr68ZilswB
Nw5+2tf80I7Mp8km/Q1UXBNcmXFeGRRVQOo3DKyYz1Sglz1sJpNAOe3mS1jaJVga
H6s46GRD4Ny2PUJeyKH4aEciK8+0CQ6iYr1a+kSNanPH6VQqvMOrYHGrNbvgmZFi
I0S/sWVXFW5xomHn+5LPgEJ4omMpe4jY5P/si+oCCsww6vS+FlANxcToCrkHg+mO
5N3PcMbZ39veH4XHv9Sqqj75H7VwtMCqFJSGT3uUp5JAjrnzrRe1hkaRcrefEcuY
z46H0Q5tZSRQdWImXRlgkhxaBGzeE5vb3TIa1Fcw02QfDPexex06iNOj4ULvPg7c
KqXhTRrWDCZrkxkGDr1zV8N6vm33BjD/aiWZdSM1JbVq2rbtePCX3cMQ303D0gg3
B4G8UYaoMv4wFxKHoRmxfieOcVLgB5ZEn9rpczQaeQ4QdBTyvH9Rv8fmtL8nLs9C
O1zaWt9TyTqTq+7p7eia31fyhsXrJu3lv4qhxpP3jBwzVAjVNPoHVTdRBzCpZEfr
7GRUsRxMkfU9EdOZCUurdHCL6hAKWiyojmWHKpBEyGw5I1fv9eMR+3m600MUJa9r
tfytsHp19C7jOY4Ef+pdMuoGAvozK/IA8wUet5E75l+pvI27Q4OGinTCWtJA4T9W
vdQ+3OhjUwPavFmDdvBKC39nYKPHZKq28W4fnEK7uRAWjz8tHqFdaNAlr9aHoYtW
jvmPrTqmxtSZeMxza4p1hoKC3VOl8PBrVb9wwOAut7mmTQOKA6JTnV37Mcv2oRq1
zOkgSiYyATLNz+TA5QVWZQArJZI88Ka7SZ/bjU32dN90p2iASxRKYuN1lGwUvdte
RTQ1Gabb7Krlua78+fdnlAwavUh2pVnwKZL8x0h/fi98MahtgFuEhRF3PezTSeRI
gwDCevIXQSUtQCehoyM6AGg+O2HOAq0jSF32XOduiP3/BmE17R2aipw8YyRZ86cm
YrkEeiXU6APuZSWPI62BAFkCsw8J80I95hikOF5SAIoePiXDR++hmrU5h52E/rNk
Rv3mX4WLji4qo+hrksD3A8QQu1Xcs/6abrfaPI3zs/6UYYE7m5lQWOXVMbXqQCDs
51Mt+gkNAtAb1mdCoPVLrqRqsoPFiFGOL76pBils8trFwLgistwHQ4nc99oSVWj0
pWXxZA2uJaCVm3L9Rw8ZObJnMwO2UI7LQriDzonqUz3SwCy4lzJ3WqT2S/O/tup9
HN/6NjVYadPJx30dshh6xwp6e4Q1Szu1HbObnPTRLS3x7M1n4lAbDwgl6zuaMGFX
0RXLx/52tuJWi3mghDbTJVX6S0fKRPLJIjugv07JJNWpIRyxCC6qC/yx4/17qhfC
HLVwSbsM1sry59gtoJQg9pfvGExzglymD6SYdOIx4u1H2tBwFeWxyz37OT/BYmR6
ijZVvZeboSWZcAcmwceu4Cj31javWQzdU7mjVI0Dsdcdm0f3BaJ7awZqQ56BfGWc
yIdbvGLu6SVzWKeCmtDPpkORgGpY7b6yMGPJYHu6oxqwTCiGcG6j1ulIQfiOv7m9
NjUgi7nWKgCYAxstG/f3HKR1wpkmTkM4GnK25p6xDnz0Dm4jG57EApCYx9TLyQZN
kmCCEkEaHEywoW0JYgS1TEKrUD1sBEO94CNMRYLcO4B1s/ecy42yl1X5hLHzROGa
FO4qCmTxZuli0Kjw91rmNOztywoOx+Goo2z3X0TgS394HBpcLGzdeutY3hU4GYVd
HYgltBQsiBGiNYGrKkuAY2wYzmf7yHi8tcajAMU2u4bcgcyJgGbTvAE5gydksK4q
4tR/etqQ0qw5QR/oCndN4lICLN1SGB4AvGtOmMebrmntnc/mZ4QA0eAlJ8dzqkmb
SFr3BKLSVpSy46jmESxH3TZZehFaq89dmq3GCHu4atl+pQXVDf+7Y4j2WciDNESs
4Bb+UjLiC9PPGo8+J88T4fgR9PPDR1IG0RscA5b6Re1PJlgVunxF5nCaxjGmAu1N
aEgNZ6bHEi3YUf/Ok89EP74R2CxO04AsVuMC7vqgb0d7orJPFzWqK4Vwp0Dn3rLR
CYEsvI05mTonoeJg2FfzfiQBP9GqyAB6Hry7MYOw2PBkvhNSsL6OQ4O7qQV/aVKU
71urKo///fe+nZbAAWT66qhv6XACAC8aT9aAxPgSOxUIcfb8TdRwbolm0H3g7VqA
rxlr6hKwDMesUzNDVjcGIs+M9fRTGrvJG33B4xwYZglzn08NhryyAkHqRntlkTvr
VdAZ95obg1hZibsA99IKmqzDTb2CfurIoCANQu8bYjuFPJ8DQDhzCUkXpfHZ9jb4
SbmZq1VlVA3ngqJXS859078FVl+/+kRBBQmPkpBqeYHUwjFT/K8h2peJOQud8ity
6FkHH9lkvzVfXgwHE52Trr0SopjRIpQcHnF0Y+kdytq8TA3Q8/F/YA8hU2lsJsBA
B9Js001abrx4pYMA+W/GS9uLsknUeRG6Sq77mRNa1kZOWff7l2ZXAyCZDhFNUvlh
dp9kcEUjebnXCixofdQeTunBt5VZcC16gnQ9L2uZOXBD7ZiU2B0WswobXCoopeeh
jlnvWwiq+q/Q0uBryF0zRgt2HeO4C8DbYGBp6M36aHkpFZysVg66+7qkIWHPDUK0
8XIWFQkgS121ebcMHzD3UEV7brNPJIy6W/cln95JWzRZzvZMaTWifkO2+6yGt1RQ
iIfiJkiOyw2qbD1LekLgJu9v4HqtgTVuMSf1Ob9dvAZ76oXG5FRFoBYha4skLBUY
nq2drSPlEYzkc5ctSr870hy8IcxPFD/m77ktgW2s0q9PdUIqcM5e54zmgeTLwq+G
fYuUJLv0Glqn74nYfwjubPZqdj549adupafiwuD7aonwMIH8/0H3kyua1j1A58g9
Wr3uLeNykrgVTIHiQ7S/Y3gMJIQFjTjQEO4OafsnYPiJgiwJ+bYknA0gqPtt9n+F
lIi2n3GJ0A60fY2hMksY8knXLL5m4Xnloqf02sRVTEZQ6n+C/LF2IRgwKMzZTlah
G8MeQzGZbJCQuS0pFi7p0Lemr7/raPBDgDUJduBVbWig3aQ/w03EjK0989BCrvy8
+Tsh9qjN3a8I0+9tLZf9sIRRi7OVWouXIWtmFEfVAoyQIR8wh79mInnNsuTbCrOS
4seFhMN1ITnuPsttxS5o4VdhAdgY6CwT3/9G6bKiC7Vo0ZagTUkjD3yQA9j4pgEO
CX0cOIZRVC079uqMwsMNZ0wbRmbO76HI/+QKhA7x5Kiko888qsToSW0UyxKzu4ZP
1R0eAMn1bPJpS9kPylnG8Osscq5D5pl5/V9kRVxQ1wajG+5lAjZf5e+mz9yLkGL+
YY4N817G/KvAUkPEljH/jIjmArRD0htXMm6KOengN/ZUFYa0BYikz+H1lzvjreDh
ueYfsMrWkMAROQrd4W3sz02r4QWleMh8g2e2pZ8GPPgdlQG8OTFdTrKkhKhL7pn6
2trydccHla65DP4nXBvhwC6LKl/qigTvJt42mblWebIc8Giz7mviOEzL6/nUnP5m
GFQp35F5MHa8dzWUJH6Lu6KMa9nJfUfFYDl2SOLN/OGt31MDXR3z3Y8ZNzxxZhm7
kPgTmAj3lzAhD/SGgmWsOqduQbp+0G2aMOTpxqcVX/UmO4iRuz5ic/pN9l1XpSQx
PLhGCigbpBfh76Cgi/gzUb8hHBvojM+pC3MYNaIoCBqG/4g/oRBrW7lfi/DOUxDw
M1i1kiJt53A5cuF6z5pytVNPv9YzuSA3w/NNwJ4x7yn0Ht7snoaYaTLkryLOu7dK
msCKvOjNRY1j+POAGbc3jz6vzo9z+XNXmVxQV3V22RF5S5tJ6HSxTkW7bMhnT5n8
Gjc4r9Zia5QenmzLnJefk9gjZb4Smdxu+sq/nR/BPJazCCIlNiM4arPsz1VugowX
1J2EQGJrbeY74kbdgpva36MFP0lHTwUyw3YR4xywd7S8C+t+nbGWTH9JCGfJQSwy
n3nLlgkUk3SX5zXSi6aC48IGncU7XtDz2o6bRW6t51DkZSHzZwQ+WKMr82tf/t5I
BcqPn/SFk1HY4KcOS5PvZ6lraKieZ3+KhW2FbTM/IR2ujbC+cwbpB/TEJ8588org
4VVPcOaSSMDof5IMkPKBNTMM7pbLRO+5c4Ja5P5BUrHUMTZy+7+DbSiR6Cd5ck/T
BL2SZwCYoWBc5BrkDKMwuk4cvXd/CImThjFbBuSC2R0EYjqPCT5TBpTrwOWydLJE
IQptFyeDZfi8PMfciJ4se3egbIihiiqBcgx7MAqLgm6Q/1uzEC9lQs90hW7AuY1v
Fp6GB7Tnm/vc11A1E81OhwnX3bnkymxwFlISlR9ezJ71+pNTDSjrhqhCv7G8JBLa
Lub2k+sTUbdkQBthXJvqGpDuuOAR7l/lQjQ83P9PymN+p85xWTSaVfUcvUaQKcvF
1qwgJWhPgB4Y7CvRnjzM5mWi7ksmVFdD+e+B43E0irwWm8U47szO8GrfMxLfJ6cz
XeDsSmVxYH++0l0D6LT4EPaJNemDTcgjchQAiVfOKrIjKOmJCD7ws5jplSoIVyxo
E9vBHtQItMshJde5l8YGufeZ7Ngl2nk3M8ngcMlPBtGcu0ciYjvuy4uX2RLlyanu
8XrhkgKOcBZF3U6/EHA3XYrOJeSQlisnb5e7E3hTkEWAK+w1NRLpQkjemWwWTzdy
fyf+0IGzd/a0FjTBcFKZnMzyMQFRemcT3JvAU57HzKtI+wLsM+czHMw3KFli2zQA
6BlfTK3bA5UQp32ByciNyHwAzia/CsXs2tmrRGinV38FFtoqDrobZg83m08VS5ZZ
lhtRQLutsc5I2WdQ+CVE2lxR2DVnoWPN4+Lj+tGQaUkJftE5E2FyC2i45kLopUhw
daxoXEOQ2srFT9J+UyQUnAlcpSxRXMXlqzoE07ei3wPksBAuJLPvbWu4DeXhA/S5
2zXwT343NaLjtQpIg8Wzr95epaGS/Z9J3pzKFXrse7MORXSr1yQ0ASgevp0mSQhX
ROtUdYbllHpvWVwof3medMzDxH2WM2sFtd6PJg2tiF4gnxjuer9gsWFJ2Yzbwfqc
k6UD/uZfjagPdRImgLwcneI84w2xmctGw03NHE79l+5ijZzYycCXwhkREYh6zRZz
lL4vtBc6/bCikR30tphN+sN5SIpZzrSBHTrfGnEveyTZWMR3PnYcvg/yhSSMtbZe
SUSlrc0ZrXs1gfx41IvkmJ+jsYeciJrzSvsL7oLJvk/7+arZphwVGgIFoL8/6cWI
kMP4rPjLO8tH84gq43EMbPvPgCk0HDZmzGnScgdpv4i0nNvaGbOGeoRjDYIsG2Qh
6vyr1p0+Rgq+2UkdNop2r9eyX+ndxuciD3nMQQsSaS0X0QFvmCxaSNWysINF+pdk
qY7rbJsbEGDIH1PvRiprN6+lqGjhAA9iz5zmNLHi/CP8CHsJUEeG770JaupoVdVA
xRFuXAVQdRi6+RAEWQWBTDSGeVrySelFErWu/JI+Kox9z96je+0y6EzfNRXxw3fK
DSQ4DFz7YxPSlz/4ed1kTz7yts8xnCVlfX0uXGWw8b1M28lwpZwGJKBdVW+bZDPp
vlB4kwr/vcsLF2085Q6SaT/3ChaA10eP2jZ/Z0wxGTUU9+gRCU9lqwB3xqUqXId6
9o+cm8X2WT4C7u/HUqaf4kkGoa/CQB56nvqC7j2lOvs9dKdAsg5wFL1wvVrMM97r
HVwA9bodj4s4SVgzr65ztO/6FE6mGWjN17yfB96eDfaz8qAEWcMZUduuQtff4Qij
kOvS+1zOn0r/9Gdiu5CNsSVvD8UV+5ziXbQz5F+TaVYm8jtf/XI/ONMyfExkAxIa
Cx1bU9I3j16LptWCI0yhnncuStf0RD0TKQOiYfbKWZUordDRaC5rT31whIAn0Nxh
eZB5Byof0b5MQ+whcNuuPdwTWIBKB2BLrPdmz8ODf8MOWdf7mKPjjJkL8epWvsVU
AHBOH7ouCtzUds2OkH1qU1l9kxrBk3BRPRaZqPbeHPy2outujSk2cmVS8rB8HAF7
mIHYYXyN2BTvkL+a/4zM2CQDOa423U9t7F5VwPLnEsqhU88OhEm80WJX3eDxWkP6
wgdXmz9KbjWdoq2gWQa33uYBQpNzmgg2BUsObpWoRlDr5Gkrqw2dlaufvI4Xl1Pj
54jAHc573IkG743KSVMES1HxlVXE+VPyjR7lfZHoPQtXRjHiDpufd3WPdR+IcUm8
AIp7z9cZ7vxeOCj5QLXk7AVowyzkhd4BPZqnNAvdDauynrv2hh0NIwMI5PJKEI1x
NMec0hr3PRiIhSGbGwywCO/g7/qwujTJ6kJYZasnb3MEIPo5k1uUCZN8gIkqvbTl
aPe6rY5lf/ClV86nH165igxzbep+zDpl6+Zd7jMNJKPUQ4iD4G06LkiLB10KzlRm
IOMEHgGWzHYqL2/tehmaTX9oKllL6QEbbr3EajMCSNVScqZdYe9ChYXID7AeDRaX
4MOHrpBWlbDaPutHL5Yad+ujhNRiMhswwE+VD2lK+vLvnWgC6ZAk5Ef3Mx7myPDA
/aJF8gZ+pNwHIyo5LbnqqQwAmEVuOTxTQdSdqK36H1kzEAcIy+jHG/yaFIc9gOke
NhTX2n9VtIgda39XU4Bz0UB9mvU9RI2KrSi4w+Qzu9KxoP4DTdGubzb+dMCsqnh9
wrfFkY64agj0/yevXf74hFBqTyvTp8vqSXRghLkR6e/jPX67GBUVm1fV9AVcT7No
HhBkwFaLWTLTrLVEVkQjSlQZL6LsQTpNGl+lhjHtkuSG1j+m4zaCRTjSsVKf/aQ/
BeNuAVA5qnKbBxv47DBsgdKbFuXi90EEwUGJLHn+9aCk/OHm0U6COxguxllOIYfF
VcVqKKayXEIBoFbBzq1QwwIxvWGUnBGwC8I5kNfU2TmmzuBSQNogbkr+wjSZ/WAI
XhrY6Rt+Ln6jJivgLwrieE0clkrVoOpkEe5DI1k1pNIZaRoPEY4UQJnRHrB9qC/p
wtXffTSRpgJkExLyRGFwb3YSMBVOfgh8llyy6KY0wvVU+tsC4c0apCvrLUWCOziA
bmXebHCNg61BJ9vA3u6to03mE9O5wxTwQNlOUDZiHikMx67qU1WdMm213tlsIMPp
UbX6JWG06iPuyOnfp/ecXtUmct/RvHs+U9hk4UAMG7PwcuBmXZ6eRwdqKUJPoiuW
+W4wHAg/TrYz5p66LpRJMzK7C8dR30E1H4DEUlbY2k5onIo0MD373zGGGta3Alft
7uJRpGXUqL25q7a4X4soeTStwwF6WYsLd1mQbK6lhhRqX9B771ecpGdWRxVewQRh
gk7dD8H2lESyb800U79AGAGazD0zfpvZQhAhSwwI+oZRXh1vbBJhgM9wslzvU3ss
hcuzP5T6KnoCTaA3vr4hQXNTeMA3YUXW6tcgz9dFFNfjM0rsYd0r8LXnBB73YuMl
AYhjznCLvdQ91MknYxZ6eM4ivSm9X9Ujsv7tSodRA54ukyXIzxj+qKDYKfAoWd2l
KAMRIKpxDg9Jv9cO5tcPIQhU4bk6cAgCfib2FNQKPoSjA3JEbCdIJUHikk6LzMhE
N5AtJ/kA/L9T4REk+Tfen2hreuzKfI0YskArUAqsKUJ9U4iI64f4p0P2L8+srSL9
HLT8oFP4D45VQ3vpwwaXoBhZJGb7tdarHqllgkmzBFQN0edJAgT1UGN4tEKP/ee9
OVT14W2UQR6xm+YLxc1bS08POHJ3TmHGOgCAHHT+xf2oWtbkHTsLW3NdiqFxDV9g
WJpGhP77iDjLIuLvHN23TaxFmEqkRjaYlnUJwb2CXlQh52vkhFDZMiso9HsUS4dc
E9WAyXgvCcp1zldJdyOqhbF5l9CD9yBEcvJBx6iT7pB4ZDcPRMoDKFPIY5IiDfUz
nWfRafRGRXppSid6zxXMr8H0mNvwoC96YAX7MWlPVCu/1F8aiEfn4VDCa5JWoQG6
pnbZ1BVtuFvc/0RZpWFiJh6GlMbRtB/jafD/hdip+OT2EH8wOA63qT2DQDFIxgk7
Gx/OBeWZSDWduHYmB9D4dEByeEYNC9buxvJxqjEBl1ccXjZ3cviN4W7JOg35h2ID
BkfWPD/7M82gkZ8o4kXjjw0bTLtWY6swFdxJe/IVrqzjH62PJD7WCRv6RYvCA2Q8
jfIcsaUrxuv5cmeG9QHqS+60FCEdM8J/vogI/U6vB+fRP9/HL8fuNv6S+3DAe0YY
SPSOCwJFBaWoxq8/sIFURKsFi9rS3FrUmWnCtV6re+wL1U9voC/xn/QUGHt5pyNP
1bypmm9o8AXjVk1xpUAQv9ADsxAuxowLnOU1HsTyNU/DR4mRVj38xur03uhA5Z7e
547Xx9L2ARh9JVjDysfa6+Xc7S/NB6qxqGAwIhULJ4AAXLym+d4NpASF3vyyMwhj
mJSBZXclQ1k9ywgmRjf+alsui2Zt//Nmpm6nhIklDqN8LNqeStPO7c0++Al6nETd
q2Vt8MI0Iryd7A65oxHNBbAJmrw8M+yY24pP5Tu8oK4c4YxIizPP2fC0riHLGjQs
cwfKUixwQK2V0ok844y3o/kKkoqC/WrbnRxPwnBCgdqrbP31oIB5LrweX12gotgL
YfZM0raM8YZzDYmdSXET5bl+4EHCpTo8SRBk+hUkgYZAcCBnaPEhOyYU0Otbv2d8
HwqWBseIPZoQURdeiiscM9Hcx2jYwTIf/BcpzQ/vxAbpUO9cQzOhabzci0pBVL+T
c0vdHsdVpHAiYqpRcwQ+kcvaoRljr+wqx0gyeZgWXXBmi9xJ2Qg+0QxlHUaZQGcE
MbQQf8QOvKzm8eAZPPbp2wQWSQ8b7p8A2awgw33CTCVtJvFJ4DSFHy2DBtXEmT3P
0MaK9CRaRa/pBTpbkUxwNLFY9YEV1n59CUi0IAw3ZfHg04FQHQoED83WJ1AFhKjV
7XlIOeFFIpFV/DBGdhy9pvFxgzSqyI1bjkI7OKdGHDvVzncWPyoKMsK814KRG00w
GZLpy2koDzUGNXNuUqY1+NT0Ff+vKxlasTzlGKqga5mn1MC32PGfCEUvhX/TiU5v
QCGcMyB2VUSHTLHDtCBOvULqbW4tbsMcz5eskqhVpSqmYr7Vx5F8mKkS2pbjT8zl
zhHWbRrsmduq8sR89lEzebDcMYm3xVgUR6zveRn5G3xzHNwkeWIyCkL/vLkRmVzM
MpFZTdn5cVapyzRONvW4i+gqxJgJOYipwmAyXlFBTQc8fEjGVgrZjhssbsAPXqOY
kcopr0zOfYlTKYhaA1RwlImLr8ovonYVAzcio9ON20VcURB4X6UvaD/TkpWZlWND
eBVxMkFT7Gx0N81fQzCGOPaZsDgB4h1GMBUsbVQW0P30ps3M1L5dvGL2iwmLg6/+
tBOcYgbi5fKzCwAsar/lAnMxHJgNl/NlYxuK5ntqJDeAScOvrlAeYE5Ekv3ywODF
M5YpxV06Kk1Y4wYo1H+yVEksn3ne7MPLGbBsfgV1/90ZQTL8GKUfqsDv9NIWn4GU
yMd7MbTE/6NB5cjPj05MiaOPK7+0Fcf5pJvyl62++HR0CjdV2NIicpCCwlAIKko6
8TPiQivphDX04ic9/OSh/4inDNWnzB0d6sboT28FuEDAiL0inswN/mVxqv8vZidW
I3WBCJdV5z6EWCh+Oc/8vlABYmtMFIgwn3EGNVM8wc3psg1ObCIiGbNqXgNvzmyB
gtc7my9bl5+DUaX9/w+7O0m4Zprm6FWnj67JxEcYYbxXY4lFRCZh6Cp65T0RCk4W
yVyWJK5x8BGsH35v591VaKzwb3GzQ/RHUUFYHdpE+0oubXoQjzYidaM7DQhdudi/
BY5CBf/lDtbZshstH7FDCgUXQ/QcvOkV17oeZVhChd8lfGuNlKlU1VYEb9IIxrXO
DyOdaVae8X2quBeO6Jq0uwyf6BoDL7iEEii8jPvW+2C+GQ/npqxKoyRnyM52hR5V
F3E8wPj1xaYOflE7Qns0mmCTSgjChWOc339BEzp87P4ltXxUWeI2V4eopyYqXZ6k
jKIFBXchjFsSMTthyEgWNKo1+0pRVbqLjPxuy25Wp2ghnt9jHaCEvk0l0QsRZYHG
ayV9onhrsHIVJsrQ9AOti8zXCXFYAVOaXMRw3WteYYRl+Xwle+ScqK+jJejlSMgM
9lsityzau3nI4jdJkjjznVoKsORObZJ70PNaQNgCS8GBmRKLJgHJPWhjZ2pkBzx2
N5rqKqvm7WurlayRleBk61vtOr98RDZp/kJ3OcTzFDk4YgO+8Trw+ESyjhFoY8Vp
tbG8PFsi/2Xco6VEA0LO/geN5puxUeZQyh0GD41VzUQiWWeQ7CF17BNOpLx2jnOI
R7BrZvV60TiCfePoewLcAEZP4hxyyOHIZRUl+yyRcejM5JdPIcMAHqViYZ6F2Llf
urqZXX7xeRqsOtz4xb8v/7px/ugUTcW8jRASnniQFBajbkeR7d7tWq6OLr1NPorN
ARm7TYh1BgxP6wf5JZ6FnkbTt3vhta4b/oCrUuOZGpieJ+QSSSAx2AS1FLRPYRIH
J9pYkh2jlNFn4FDbpuiZj3FUDt1ygyGJth2AC4Rqnyiz8iC2YU5QPzCSDbTmOXI9
MUHSSPTvjkSmK/LJY7w6cSP4dNbpwhE/+9vUBjhQcpBbJogUQYFasUba60WRq6W8
Zsxmg45yxYYhLy/v5ueE6JGw1FncIasaTGL/JCBPBONOJ/WZKLW3mI7ixf421tCT
dJZohSLYe956cdC3twCn9ADvlpSK6JzyX6DzkK24pl3hzOm9cflqNN1cc9EZBxsl
NuDmu3QxgS1Kv3R1jI8Rjis8smUCZ/YG3ci4kI6NGQRLj/oglMzVglWBv7zplI6K
tM4+bdVZeo5t3l/WAzq0G//Echtmw4xUrkqQS5OkTtjcDjYA/UjT8Sdjaz7D0wg7
1efZuORopqiF3nXPGRJx6EHHjOn4WkSNnUqR9+QQsgVhTiXPYKgUsQDWrZq/CTNp
VoIlMpLOzBWV1o1KuRmXIqUBQGO0J7spP1umRk5DlwBv4UPqycMDNwW+cEpnIOXE
hd16RdhMfMYubqyT1tt+yzunhfHqzd5jzYPBlNRP6Q1xRhxewF2jPL1dotw+DQKa
krCPyOh/KQbCcsVZtXFAcv1NxzI4l1qZLBs6NcnqVFAQVKsahLy28HVYdY5OBw0L
Pa1hTbf7Hr1WzHZ2QPm+srWahrfV5+hqQsAEsc9kd66Tgd8I9/qTSsTFKV4yqU1t
CeEE/sIOvukKDp5vGe25b0ITI6GE7zRVYiWGCUr2TXUqmRIzebj0Wmr4ZUDi5Xqj
QAOegGqNDs/SKmxQJuSinK1G19BblofMSxIs28uX6m/11ibcxReUGmLo4V3NwHoP
Pd5sXdpLea2cPvn3m61DeHdCsbWmOHTj4fZS/qsMsYTMQINCU9khZd9fLTDhbKsk
HBun4YcFPGywD9oRe1RJkCVZ/giSx8IXgKq7YQAGQRLT8SGLB4KPkEr+I9nVzUlD
HglE4dLg5OkRlWr2VaNUvxEd37baZU1Sex+DvwrpuffX5Iv095uKVUu1tfYieVxl
9K5pWn30yvVa70ekPIKtgDnblGcm6EBHanO2seWvM7HSJjEN9j9CNPvubyZlXtn7
WzsaUEfQVQ8F/PMbnqplqlKpjOiknxX8KdPoZFNTFUCdBpZYJQ4lbJVZXG3pk6ET
6Po6g8oxzGqIpVwSqXQ3ikTIbzglJ29XijdeqLO3bYZmjQN/9T6aOiiWHVQz38vj
6jTy7qcJ8GgMGvgPtpGq6Lu6j61LWUsPpqjZWqAZOA/RKnMQGv3RrNJgmIpqKA+t
eksaNS6mMGl2ci5NcZvkVe2d8AFGlhu5tnsJGqNXU0EZYQiXcOHfTzv233puZet+
7yHreOR6FfjCIuOuSxvTwujCF4Rn+UFrcbNWBk6SXV3Aog0WS/ediuRdCDtUpXM+
VHI3AWWjA7BEhCVVcIzNklHI0FYbLE/UrbQTfyvr9MXPYStAM5a/GKl6d0BEIgfJ
EP1Qu4fpYJaEj77LAECv3DQJrgTFgmj+7JUB1ZTIcmMlT7y9vj7hMEi5HRVtd8jl
p3pdq2fvzoNpNeqAeNsz8XJ/UOgbYAe2NqjLB9A85SrFVa14wsZsUiK7ZK4qJQ+z
ksHbkPWd3sE0yfgEqlo1VM/AYO173S5Gyxr6RiuC38Fn4uvD7JbzCF4l7PqUJHcz
8GF2GT6UWiHfV0lAcTB+F9dQpyAiLtvLnoTRFDjK+yJBhbEHU3Ll3n8YwQ2JlU2p
JUjNN4d21QyUYemWemhNteIhYFeekVkJ896jB3DIbLS0ePk5xJedEZeeEfMwrlil
QJuR1+EoJrYu9b1/YCMhMyPCc6jWwVqfh4om16nk4s4I5JvYA6Mcn6NrvMHkVgNg
2bClm3YwDUA4IV6p/QGnp1NDS4isHkoGbNckyDEy50x4GVoiSAIyW1QI1ZPJgrRr
5g0mslcLjuWnKMzld3HL/Kr9StuwtB836UwjDS+omlzwOIEwP6xTNwNkC30uY9iU
RAyDU34YbchcOsWCr/Pycv0IrA0AcLumXtIURF93Dy/A1MN3yjGJVZWIZUZcgz/m
Q7sf0m1UdKSPPMOfMxdSMJ3eediogtpqxy5WozJeOsRq3M1iwegFSfl7PF4CcBrN
UiabKIagNqCI3C11gt1zUXkwsOpQ57jOPzd64qehxcGF53yrQojFYRRyFFkh5kTH
VYdulS1vP7ktIzBhk27B5Fb8zkONFDGV5pyHlKPw7aU0Tco9hAn0+dN/RJdBVC5O
ZBHWxOGAMZQ3Dk1NRR+mSjWGNCV6OAUnZTgyaOaQDfBvXJRspXhl+oG4vfDLXFmm
wSzM5NoVsc2e0DGJ+yVSnBuLaytqYHRPekVN6M9N6UPDhPMUjNBrqN6mzn7uCOf7
MjuE+3FFqqK3lixUHD4qK3qFtlBAG7Bl/03Xu8yM4I+91FeYyfyJLkXNU6C3BVH2
/+/ng7e2Ci41XObdiHd3+FSV7OXUnDdvRqzjKyu6bqTXE+1SKHXvKI2CNwLOlBZa
Wxmf2ToePMfj8TMqOGfC+UQqk9hGVzjvFBaDuTKXXhKhCAK6IMixLu1zLq4xOg0V
tV1vCltHQeVOCfZVbvyTjUdOHNgsZcLiXRwi98dBkWK+hCXqCr2z7EqRAl7NHJtE
Kv/Tmo27Hbu9bTtBDjWOpYAZocHVFZVjmIF8i7UOJyGmSb2wbWAlC88rFSs5UaOh
LBH77ZPWZpVgnWlMIKQFSireXuJXNYyeOv3+ILCWu0m08ZJA9qUM+kNXg6QFm/pa
I7B7XnTf9pClSb0B8Fh3j32ZxR5rVXud6oKDFoSLT4FyCIA9AZaC44HijpkVfr0g
mwtWskbTcy1MTs1EG5MzATWSPyiY24oYUn4DA1JpAxEKloHwcAyFIvmY/TUm95rE
Uif5tXyHj7z7YtapgGIYwJXgmamenhFrUFkU981N+vROdPwB9yyfc80yFpdvhKUy
6blGdYMOKYf+RNIofrmJRP8MHR8M9DdgVJ64+Ra/nZsvsnVWnN2BsCroKZ96UPFB
gcr+Q3520vqqXVKMvR++QNH3VeTnkvUXQD0x6vc42NwtVBoD1jTvASQd/ES1HG6C
qYpvAoOd+WknqLW8/4Ej8F+rZR2366wG4zl9AzFEUxOiq4gKQcnPcSlAYCBSoSDm
ZyP7dW95ZFK5yzM14rqjb3bniXkqfiwp2S8NOh0j2h0ovk3P2kTPH22wOZE+dDGK
7U9LcOnfBPlE7POX0XhiE52I8R6PW6FQgnl5Sxb3nTvpBVoGowFMFxHI4L+edUus
wPa1hqCGVBSsg54L/K3B9DpW0w8Uvg1IXUyihYq+/poJKGJSGvyHGFhNM59YEC+I
jTE+pZWr5W26I2X9aGzxwVReWxQqiSMYz0vL3QaD/HDd7MCLqqZlfNBdXiFAPZAr
/a8wdKdrihtSzc5KXpi7AGGDcy9g0h0KMpV7HBXxuD+g09A4gZI7y5afN2XrPh9a
5t097lRUnmiKlBkfhn8f+SqNdw57a4W0xUh5nurT+ZeYkP879T8PmyKoWiRnyGgP
A6s85vpF+6qmHfm0XHQP+YbxT5Vc20yBEZmK0IPk9nyN2nzgSFEogc45c215dpTv
rk7bGrrJVT+v1IeHMJzDXtgrGwO12TUKiYARzlA3mE3HhPY49GRY1dou/Xwef6ZX
0qsjW5auxWfFgTRG0VwpIk97zx4/VKuqqofCZ39EWC+qSvWl4mc6+Qg/0E76ZYRo
+e4UKq6tLsjW9m6g9EwuCpByiUfluMbx5+mcRx7zszWmpSSS1TQjCuR2rwYfqEhJ
tdUc5GFEHQossZQDobd/uNB/BG60Sd6Uh509wb8gopx9IYeYu83V1fMMR5Ye/bw3
h8g/Brrc2XLPzu3v6kBA9tIX4+EzPUjg7VNHDqYLULXv5Udqoklsj8+qxLqnR7Nh
O9Wk0MgdWSHM6z3wK+34iB1lRaj8nXgtjT/CnmB7hu0RCUaZs1lTr4/DmseHoS+d
De4eA2htbpwUabeAJ7wJOHvDRAG/kyrNn989K0vRRhJvdMyEsohvIFdpKbGzX53Y
mDdDlN8tzvkRFjJF0PB5o212UhRAW94oIynMJh7DER/JWTxBGeKj0Ug8HWIvj6rR
AoqoN2P56tKH/i15Ddl+GaxjGBicU4tfBRFsq8nxZ7/yhEoOPoSjN7oI0Y2iP8VS
IqwjFCV2nX3Hyy5b1tp1qkuXvZifoDXL3uLPjnhG1WXrCFnLzVt+oEDpgl4o0KD/
AGaDkMBj0VX1z1/RyGIlpz3WPPh1150zKNyWygmRbr8DrkY0xi/Dmy4xVPnaL0QS
CrSoDCBgVaCUsdGY0rQ7P7Dn0LEYy3B3VWtkNwd7CEjIpvkUxHawdjE68K9Mmku5
EWLpEhIXyJcFJWvGQHVmr+MFvaswCgcwFgTikn+wWpoF+53Fu5TwY2vkTfJKwaMd
PkCX5GnueAIUGcA1T8MqLdZC+00b6OhCk9S985TXlRpShpSoI9Kg3sKE8C1a+CIG
stG3lmC1KOXNz1ZsuMW9Z8wOzrDCMc411wwttWZSnmGwZO+I5WLf3h5RL3TKemBC
CSZTcI9AYjdrBfgvZiWdJ0m0ZhmkI2nng7Je8rt5oFe00uMEe8VtRbgraGT2fA30
MHFv0t9PlM35NOO2zivvVbUE8yK4QmAVCpAeXxldG97/d/kF9Yjy64UzFSYF+fGl
TKUH8RgFV09KqSXqny7OQloIgeUBIAW6J4jINiQZXMoZBJaDrXx1flr4NFuC95WQ
ZzNsrJtF3Tt4192VEIh0EeHved8B//Gg9QWxbYckpi0X4ESHq5LBd6kCWIjlt4jP
Rm5DLnTyRuJ5mOTm67R0+qUqa4JV5Jhf2TWq1LsfKoReGyO7TbyXjNCQEnJ2IJOw
PLdFzAkB3/aPXJftYncUrr8gAxM0to2amMzuFxm6PQIenw9fSBE8WXkik21nxQw9
OY81Gp8uKAEI2rc1NWEo3LXexjOGJFhIBUdvF9hSb4iHXfbeoAFH/N+ca4WET70L
X6T+2vRKs7doYDp4UzznafF4d16OcNABNZSEjRUiDvX4zKdK1r1sPHsJey6e+BKr
mRtuA4pOLZOSrD9Kv2sa/XrCNmeLQrXzSIM30KOza4ipv9+HHzV0KcDyUHlgJUHt
Mws3C/7civCtJCTD97b0aDBy8+8/wpy70mY+g7141AMKPSHjj3Kk5Uf6hQrd90dQ
5Ul/2uwc7C0ovmf7pg8n/aZi+jhQ8A99gPyOFxv7YRWPFxXGT/50BgInZIAQ+lnt
1/BRwfrY3CpOK+IsOqAYVLjuS38ECtdqXbjfpKYxBvi1fXkpzVGijERbJBnc02aw
L6SYdc4TDSh7gWdSfDnJP/j7o6RIGv9bzZ7tWANuPgFQe82GKZBb1SuH26Ce4vr4
qTelbICJzTryzk0kMd1R2o1F2uE895383Z6EZFmwBOGHDP9a7gdbd9GUFpzCsiQ6
5HqjCsiSmkn0KWcEcrjV2UtEpZxwDQaII+uwRI0QKgXptxvvQijZB3I/MYgdyQWD
oVpNILkf4LcbT98S98Wmk76itsSqmLxdsMzYMbAD5Fhc7q3pJiP5fK+18+T78k3S
2pf8vErGWnhfXBSpd5eIaxbkju+m3/WCrU20mgKwFNQICmb4GFClJSUDrnKyn26b
9dkvKbColz5N5YUeSQRBr1+oTBaBHUSUZpBdkYwxnHGWwp6219b67wbJvybBBw8B
vkDbT+uaNS2WBwZb6LiiBphDyOX9h7D3175xP/oiuCgjFnWqWSVeBDPmidVspPk4
eHSaWX5toIcHdTH7n7oKkvfUPJLgNl4jTUwuCUX5T65/963Hp4HY9CpMCgzEnWYK
xugbTP3wI54fSemCTbcX71PBUJiw8dVzlo2f9I4nOt3sDhjnBaJcYL2hvqZIBMIJ
z784TNcGbRu4eEPx7ToVimBwHAzjQDDRUCWikQudhMoquHjTqElCEA+UE1AQRa8A
WIMhBIiL1/BA8jWD/L82YMqLBWH8xPPCwPGmrbIarZAvhOpTZN45A5/ORg0fpccR
SfGt4BrM/Odm1VhknDGRiqkXTZ1IsbB8wCZYJS4HFsqHAMY2vmFcEaI1u9bc/ZbN
6qQusCc7Og8FofOi9sDlRiITVhQqj+YYLnPmQnc+t/HrPn278LOxr9PZKCFJ/tDU
ePjUib+hkEhxahPAms3d25wv/mdrC/+A/qhulrCMOzSnJq8+qqWT5JE4wmf4o9P6
w9PN7vhLuv2C0B6GbwG2O+mFzmu1w9CON3jtFMUjO168YEBAUL/bnSPT+ToWvp5i
ze+Ff3IHh5WtD3CIlP09HXmY/sAaJk6aJpnqbn0xRvImG1y5r3a2ISVuQimE2eql
REu2EPDidNBvCWq5bGxJ6NQsbcD53F5yKNpgLxm5F3oId7b67Rjx4LE7sLtfjl0M
TzKnHf+jp30n8dhFcFFNvnTW+UzVUJnj/pps2myMdeXKyOezexn7Qx/tFhqpOvox
N3g2xPnvL4Vl70qPYgV3zQ0cCneXeSnQyi43GFgU5jSfe0w24hQO0DMoEIme6ZFs
H5bB8qDFghrVGTj2EQmeyAz9h+w9dOYaOyNVMZhPBdhLEF36cPorGNUA/rOGuB/t
ksWYYA0CQe8saMO/IspSibNLm8lDElKcAru564Z/Q+pi28jqzpptb/df+Huhl7f3
1j/xeX9R6tarYYqtx4gbB2PX0wSrNYdE8TAhJEfERapZdSbKF5YHWfqKWusp14nc
aBedj6knCIS1HbBBw6NGkr5eCGyWv7zKUpZw3jua0hjQefKZ7JZYQOdP3CRUnDF+
twKhKxxPBUt7d6zd+JUOK+imEjHzqgBakrwDMZH+qYk6p5ivjYXUS4G4Zf+veIEw
YZT4AhANvUNU//F47sHxC5nwszYmFCiEEUuN3P+egJL3JQwoeGwiwQugH/A7Bsaw
pOGhbL5VUBUaKukuKexgAVVRp4ISIGqAsD19506xmmQQ72I1ESmxD6EpSS76OruE
LtcxEFAebwHKWGz+nNptnyj7XLbJyaBJ52qrkGGSTSor9aCdr8ChG8Zb9Bc8vBB2
SORjibEqaWfRkwiSp2oPWZWorkyHbDVe0eoTEWExPfpqPKCp42fYP3O287v90sHK
CZYDlHLuvBD27VsQHIcjYhFy54zlYmoZZwpyDfFGqA0ZF1M/O27Z4W7WvoGQ8Y1+
4rM9OHxJZ0skVYcNvHVGzV6Uy7w9OEEbIIcDKkl/aTysvT9gjBT3qWeQasko5wvk
06i9DaSUWOOfYLimsRN1+bDvUfvncORK7mIwTdw2rilkpLdVcNqmdmSv5nCs/SJX
xBc9GaxAxxMFP6BKo2v7LXTEOHo2awTKaZTZMZAWuS1ekoBvjg8FSRNC2/lJS2oF
k0VGex6NZXFoL85SU1qtBDLlD+ZR6cmqy6KZtAMv0Y5yDDfJvcjkUKLtqO/c6pBv
21hmDsOUz6SoxcGh8ofEPrSy3szMmwJQWDt0/G4sbsFyMKVqIn2Xar1HqjO1SIOm
zkl+zEFiojyF/KZJ9JDUZ70aksQWGG0+lwJ++QgweJTR954EaBlz8Wa5fvu4zoIq
ySmu/WNHbPzDCq43NqVl2SjvSUW7aY2/KJiJTCrHzrs5NqDScb5NdnLN9LBIP1SO
J7Bwqk8KxCbjnHdRG5Wsnm24ut/ty7BqaS59WNdqF9MriLbBw9NZ/koqeOu5k7vl
f9lZl+n8SPIdpEgYkjphF4Q0IFpSDgJIOW2g9Jr1VyC9zj+l43tE5oe2nmhIsk+/
KR0tKC+1L15P5qrruaMXC4XdU0lwos5982PjruBrimPCHfRnBuCDia11PGImML7J
IRe7AJfryhZYqtBzRDLmcFPo14w/K1cBynnAT0KyTslCIGVzWDXxIteNwmVAaPYc
s3xXoAq9FcZUrm1wikssVsrDMCOnKyZdzr69ap4tFgsjx3YUdiyCTwHHSUQYgu6M
6vxSPC7iiihMLpZnUIfFdL+6/majkEqGVSyghDB+rI7jtqppMuhhhnAPt2msW7QJ
vPlNqm3li0EDEAajWhcDdIuJf2dxCMoEjmCKSv7AfgpLzFV4Li0Q0ALmuKYHvipx
bBmFJHxWtSixcqSpcEP05QPcQR6jIYpA7Ak8VFHszZcAWc0Cap6baunZs5KQhj6C
+g4bRuXxFQdu+q196Ls/pPKx0PS+6uXsQhLKttbAQ61atKO14/Bc1a6UTl37TUVl
4BGl5jkCx+zOhTwcZNw+ZArWvCeBk+MdTK/I1eP6R1n/TCmZYg3wF82ICZuQDZOS
AmwMf+JKXoOWlsEfAYNREIQzuu+lmbZQBoeqV+Lr1+zbCDC6VNnTccxg+JKiOb8Z
isxeWaz8EtDanNJbOlc8nfUoj/UjH9g5A3UFG/UMgFg0Np83X7n1SB1XgWVNlqh0
6AqIqU1dPgduM40DO6E4PG8yLiQr8jHwRaGqi81qTp4/Ek5wKCuSHKxj9Ddm+RBk
O6arOMTh/QHtgmzoG7pPmJ95y+TpUJGSuXGzZIS80dj1V+gHC9YSv69fI/7ZN442
vTUOsKLpKd2cmC8E+05bfWBSwaKL3EFunx6K36tX6ERBHy+5+kdLxOhaQIS/WGJz
6rabLraCCrJws3nFPqKi6vxbyRqyDktDkVpWUfF6E/faX0lwqmaQbGDxXL1q55N9
Kgmm+OtIzTUyARiytCrxfbiKsfXLJE8ATST4Z3NKXacYGxGz9EsDLhGcBOdJBoZ7
e/TRbMT0EtjAcKjQuG4QVj4Y1zWf5UDwnIl40ajKoaxf0yzvmEhXDHk+qWmeITzw
AP5yyislHkevMT1t9VsD3y57w0Fo/XJswtF1kClPMqDprUWAUywiKUzHZmDUX0cC
Ej8r6CIPRZEuZsJlFyUIGv6zAV8Oy6R0d61oS+MLFNb9Royo3+M2V+lmgX8+xPdv
xZH2PxuUpmHdDunxM9xj+izkZ3E6KRTFHssIhONuKoYkhVOrB7K/Mq94POYQNsPd
Ly3DmJpRBI0WPppyFNp+8FOaRnUF4WQkkOTdJnViioP0tFM4K5M30l/qAbRcIZ+b
zpOQLs1ewGIfpDU6hEhRZvyI2v7X4krtM6zoWmWezp4qFtiL9BWe2ioXtKUHj1pd
78nNxp50zlN4m28Pwz4j33H4skjtAosH9snzN848K8aZeEuUBfbupT6TmqAd9bD0
O5AJDdQXNH98HZRUD4KMl0F1uOe+Uw7sjTN/hdfCWPEzJMd+oSPr8T9GIUN/lvR8
m1s8KvfchYy3sL9GvCX0kPkXOmeLwTV6RzMgz7AIn6rHl+d6vv0IEC7ApFW9eiYw
pQnAry0X2YYgjLuQTB+f8Cyo2E3rIZULvFWa1mWwgpSS9THjqGwrs4a1sVT3+SsC
l6bxbhp4zK4QV3A5WWxpbriijsnP5cnR7kAd+7x2eC/Q2DFkjwkAYA3T4Q/HVRw1
KyGLhqpGDDowLZXWyrbdSKmSOpnXwEqnLesxAJin3zHvpN8xxrgQpF+lSkvU2wN6
15+z1UreQ1ixzHZCOXp7cjS7MieR/eYjxnqqLkVzhzWd8PGvevseFy1F6KYgnBKF
9ODnnYV1e2oZY1VbfwOsIYcDc3S+kuCktAsQoOevFhgnve8cXymQWieT/TtYT8x2
vnBIlhT5WkyGKYoyQaQT8HBVth9Mu92+v68yizKcQhD+yLPQ4i+T8798aNweXKql
YgxKxeaPEYUbk7ys1ck54BaCYKLfPG3jzJTR5EjVOOMYCdlApbCD7nnRDT8yvSXp
SqRKWcIdVnLhkmpsKpKDjfxN0HFYStgSDwUg03lNwCtj33KnOyUZ9s5+KvB/PC+s
9rpaDN+KvoegL2Q3yQjaJ/a4jPU9ktUh+dIf/xn929p7t1svmHJDurAULA6msbZd
PPMXJVapgM0kHM91kuoyzpt55Jb0KrI8JT21kyrwT58TMuugGAZgSIyLBwyy1Msc
Uhe+Rcap0LR4VZ1Ma9HaQSR/IMOldIm/Kcav7sxHSvavJ4HrcCbWJ9sRtXpcNiNO
PHtJKDiK6UPCkHrsEIuceWxhmSFeWR2qPkvhv1/itNG+gRsGUby6DfHYhR/lMMR4
+0tw1GpENNVmV9nxw3QksqdarO6onGI3zKRKtWx0nHP/xpSSIYzAwFXoUWoAGXCX
PvAZlzHHtqrGnaJInuUyhJAA5eS0uYRqQbBGAcRjcG82yLRPez7xM2w6oZl/2JYX
kmetIDhCxWSDAL1+AeBTR+Qq8nu2ZlSqXuaLrAP+Ls9CuTAA7T8xvCCLiNoFVnoh
Tzid9djPX8veCruF1AyYDrT8kuet3YGp34KGAgcF1V9gYpslPNzvcTJx8HKa0Vhk
PqMYpksC0Atj6TbmF0iodtpQAlU73eFRiEYa5CtTslsQlKsqN5gQ+u+EdqZUd8LS
6aeOc5m+gb3SD1uW6PnvPqVQf9yA7k2LZsH1pWiRU6TqdLYBXaDurw8rdeBsziiL
CSakR9d3Dh7GCj+O08YaTASENSvJKde4Dch1IJ2FT3Hl9gifTfL/tYNElWYM3Bdn
0eoTCUvDZJzW5svQLEMX4yLJ2L0RuuGJ6ZUXJFNxkceqiWxVMMDqnzxPsX6bkuCg
NDDupI7nNghVonmalcOP9H0uvfFpSI5PtqoA3/Fq00GF+mFJbkFNeyjtGdjMkzR3
RzSuG4zoY6dU61uKdnw+0gAfYFJOh1vxraDMuyFXgzboIGjqbb0WOB2eHZe9smbO
BEGN6AijUn92gGJrXKu8jFNm/eeZVCTuNiPpVfoGXl33thG4wIs6Jswg1cBn9OYd
VbSuOXRWaDtJGTu28mMmIRP7Bfkq8Zs3Vx+QsOkW+1zdaAhJAwQNyUiIcwZ7GeCv
kkrqzlrLpOgkIfdmH75hh2cHdiiUq7Yyz8wFMt4KlYqXdj9XfGGZ9ULcV++CpXs+
sPfszcF73fHDxBjIVlPdlK+n6nLjnOM6HVjQH56nZJl2RTD/oFTpb8JlLFRPN2K8
NILwuxPL5WFL1k0831woP5tFPV28X4h5T+CKc3QyT3EFhkP00F5ZujhGmeImmzZE
PJ7DlDS0v71l4vkdk+Sf0P4534wf1+tGmsXDBq67V+FS4Br3ukLPhGD5miwd/z0x
na4RwjF/XcXjAimDd2IPmdnsRhP4Bwd0bUNWIC1GIYtD/408U8MRamns9s6jy7fK
DISQaoGs/znhZ9Oz3mcOIazrcHcVAIZoLscn9q+pcwShw2fi6T7YS171MjN5hXpT
xunO4S9ZUO83ItZF1Ro3o7vcgpyRFRptILmlC+63pH3oEb/QNIlO8n/LRaXtJdE3
mueOyLwdKKHHtD0cbzxHmmoYhnXbXYz0kVgwnxKrjm+e4MjX165mowlzBCairTcl
Z00hOsHgSIyeCPvMVGzCANRvf2eez2Q9b1G796mekPKTM8RTLkGfkcCEonaGMteJ
F1byI1SdhyJwEQz7u59SKo8sX3AImgs0ndda7ZsdIiBh7oy9e6GCd9hCwydTu4Wp
Nzt6wZZRgGyE0RFIa6i4zANS9eOx5HsJ9OyR/sLHGZmHP8Gu7cNdPeIp2DPDG88E
YDgrAeS53PfiHI+4vqvUKrhKB80Ceo5NXy75vMx2Bdmisn7wSv48leTInstwQMjh
biLa/SiaxAtozjs4C/+v9CGv9k0VYfRQsX9e4u24h/bUCzd0LSoXe9AkccZTqy68
h+10gAcOT7FhW50is113LgTX2Apgs+Tq4XYigHG7k2ff0ZCB19HmCSdPGdEeSSen
cl6Oxs41mYQin/6IIKvzd0fp9ll9hkPN15hUgipptDS7o2vW3f3VaZY06zEqGNQl
seyF+XtgQVl9/J0uHknX0F8r9F+tmul2+6qez6ZbYaCq2Pp96auQRvyYQjGGzLS6
QF9HSg6qQfF9Sph2MeUmvkPnQZ/psMi/y6XC4ZYdvsgeJyZe9lK5H8iEN/qgZf5v
2C5/Pi13AuYbQEexFFlvHQRcaQkhxEvtmp71viwKrITRFkH+MweQ71YafG9WeklH
4vAHOdZ/Twi1K5Npe1hdOfClBto7GwRXCybz/dc1aV4ws3aklljBwdUnRQdTTpT8
+Ej5v8O65NeyCB12UjSdHHn2KuCFOg/vqzleJR2bQgu5sPGj+2SoVxvv7n2qUk8Q
MRZV25hCZLRchCFWADg7Obujmwe2ws9/J0pdIHuxwoFsscbMyI0Imr/FbsfwLtC5
f2IOeZfz+Cz6DWHNWaiKNEHdOBhx3veDeOQjM3ZKnJYQCsO8qUb6P9mvvpjKfEVs
rOpfbitskoW8yPIZQb0DmDPPgQWESc988pVifP4AKfIFG90kSU5045xadZGOVpGm
39CQnWgMx/02UP3mFeXyCytXjVvi3FH07nb02EY8X7BQqW4i2bwSOXlDTkjZhWk+
NVnq5k5HBFQEpL6BG0ibYhWKFLnIY8fU9SGYgUHq/2LMXBiiEnsP5ZDRXno3HJBJ
5fPQ/U/yQhl/dtWW1Lp2wXikJycnh3ignp3tsL1N1gxO0c/8fQ7+Od0aIc1X+plZ
NqduVU3WR2VYut90T9QehEk1z3i61vrBvZHDHT60gNs+iGY6STJtKUov1t8tOUoM
J/fAsjx57lpx/OnlWAj7G8RDur8xje4NK160D486tXy9vV7mgWUtpY+2wxoa3PTF
G5d8u/j5LM1r4xX5x/htYpmUyrmeH+4dY6CuC3sJnjRLMcurIHgEraXNJUSpQsDu
6fXoZ9sRxpFpFmzY9/szWuH9OhjJ+BCg/ZBF8RGletYPoa0/O0N2c0hTHNBDYBjK
cqB29IDkq3o2qlS3/dURSNgkgLcsDjb/gyXvdnpgv3I7g4wdMIfIEWxriz5si1S3
BEBTYgRjDH5v5dLuSagaSlKRf7SGR21Y+0cshcW6lOw4NVHUIc6XnzvAnH8ihmxr
4m98N+WyMDNrewVlKsreVwtyCdRQfJT0dP+d/s5zZJHGUwN1cFZt+UGb0mkXMqxP
fsQYHhcZgaL9gouHfFW/6WunHZ1r1YQGZsQ+tpjo0sGzSdREpgynQjM+76gcb95+
QAQv3cM2zhrrLofF0FShDSIkRGqBnZpzOJeOR/NOjRXIrTj/IwF/9Y1aq094aOBC
zirQSxyb8sLbINySReo0Ebrji9mVFx5EU3kNIRIdlXRS9PZLRU9ucka5KLVxelh2
MYstuhncUMec9aD4/W3ETSW03RGFr72UGQ5ETrv/cuYTv+F1u1ssOpSfx28bitmY
rch/YAzc63O27jx/VSItCKwm0weKhMxPV9KbGHr6Omra62x2d31tZiXxHaOVmKAZ
P5GxthGctvmz/PxDXAmMkcJf2zQJQeuXJuAB71BbhHSrD8swiL8XP7/hbYKBQaOV
qYQGJzBygjGUSh2HvbjSKa5PwuHy8ZPYK/3ldask2DGiFkvXKoFAWThAbZNJ21RH
hfsZ6ZN50KmDF3lpcwzvGZbZAIsBhIa3YlB8bQV7Je5UoE1l0banmboJISHyrfXY
RgM/byT83xtILu7yF2F9htV0UGDzrdmTmP2bKVH5zvy6mkBg4n3FSBpovPezfiE9
LaxspuTQbKIw7WP+dsVMjZZR9bRQwZtankzeCJFl26qCDvg81ju0vdkS/5KvlFzq
IOKtCIjMBja1Jft69aPz9/+cC4spnC54KV64fCLSsIsPNxUeVDl/NaZhVsHAVIQd
I7hH27DX5dCLY/IkOSK+gsJzfUbRVpL5WpvWLVtJ2CEtv3PjVgFP1yoWl37CTePf
PLcYJvrmSnrhnQqOH9KWw4KY6mJC8sxZ+mb7Pj6DBnvnyDJYKKEB/2tyyCcd9Wt3
WTbaDwqPDpFLeUzY64HdQZXn4dm6d8eZotndfyN83lNknO2sSraexqWnknwBMYVl
QU7LRvRgrB6mo4dDtZKS1ggUexIg31+6FHI7SEVXk5wiLBLfRSFkSOUl0p0BYzEl
RyxOVf3Crf85HfruhDVqkGpcUZST7JlL+kzA6S5mENyJOoCVKP24LMCYB2bPFfq0
LVfOiDsEJFYnvr7mdATFx735Sp8ZPV6DSywRGvJ7wbArVXGeXBrjIfZGdhGt/pPr
NZnthEq9SeKGRkPz3gXHHF4ncmpHVQoBBDdwIN+64xH3GHEjwuQwfVbfNsf9g7dd
cUq+11pzeItEY+UyH/LsZ92+epmgEntsM26kBjEK+xxV82lulXDcBFxbNi+nJaUG
N62253qoB7Yh2f3QcuO4LERiZ2VWCz4r9GgP5CIboxhEAP5MUUtkZ/uexfpANvFE
psnGEPuQCEuUPCyVSZWhX5vn3FNP0LDeOeEhjbJhym0Z/5/3CHf9fNawWIToTbTg
PT/NTRcDNZHHDPtXmTWGVpp2IDt97SBp6hzOpjUMXd0MSElXSi7KwdN30SQF/tJ5
YM2oKxoLIGwlihbq01YNv2R2DpUzk3mE8SJtbS9Cqen4wqM2KLlTu0mE8THJ+ptI
e7/NQggyDGor0g5WMOzreGf3yvKuYaueCvyjMiCuSuKN7t7qDywl7oeGwHVAqPhg
6yHwey/Hrz3+T5foHu2OSvxOy8ZsScEDKHH5cTfEgQkqgYEPqUdFBZAUVvVz5HIs
uvUbPbu4oAqP0d2N0ULdW5gNeRjnoWMKnREyhww8Yq6y6vk7pi30kauV1d76rT0f
chFxfhaEsBsvPQWABtj5JcicaFSNgsknRkPtCt1Jp0kyECDul+B5BGHZFvnRX6Uk
yff7OxBJSOvFOqDMW7sNQD4PgpyobVqCkwuu5YB/bUEkz2wNN9e+rutpMzXR4WGu
GEQ2Y6gV6TH0Tg9+HcNJafUXrsd82zJ+Zh9A6tuKWMs0nlPiWzF9EJXCYkeO+IfC
gZYkzneVt2j2FmZFIzm44TFEA4yJr4H0ZBhx2YAYyaojcupmzO3lj1i9yGFHsvI/
atEjPI/APNJ2jM9qO6bi1LmF6dJxQxQNLoufUwmFZZA1d8EYJ/uuCA4cPAohVv4/
i5TR88rW9PB06eAqHqVBXzNYbut7Pi/tLVzjizcj39FbrqwT+qYy3yoB9LVU5r3Q
ewQbTcdOlvz8R3pnan0nYh1SJdRw+njNK5JrtIO+rey/U6fGLZmqLAi5wDpq+LdJ
Hbdws4JPezuVfR/jI0TSdey4VJlP7DzPWqdVRfm4HGsK8Bb8QsKKxpZLxR0ub3jQ
i5qvFy7OaOQ3ypCm2UYwl4L/zCDPLS0G+UtQBCHDG0e63GH4QNkcbNElX3NHvpEK
crRBXPVEtc17PGS9hA20gtWxZeeOJcEl+SZmdpqXugd4kGIKGA39lp3o7vYc9a4a
fOpAwOJqeiWfMJg0j4V5kE2iRqdXtkBNFUeOMjATznePdNtgHSOaSm8Qju9XSU8O
ejSCe3iawlXjhaeIH8oGq89PAX4B7PtZJ74z3HPWoZ/QGFihUaMj/EUqEoZxZm3j
Yiu3brA3IEUrjeXwB8jRO7Dc1flIWL/CkCJNa1KAaY+0oaywJmwTn3aw0BDeKbEs
2Z4nEX+tzICikq+NEHKmKcfgbLLxSjhwLJlzuJjrqFa385HzpiYlHzU35YyWxRGH
ccyv+/qhXmvxaUKom63xwy9fZiJ/WR5lH7LKAsg5wilWZv/iUCQfNn31ws9qEgE5
eVvQ6ncaGksccvydVyAskLzZPdP67kjtftKTGjQaUVH2hGPDoHs69gwP3ceSX4HO
vGryMlrzE7MoqE9xrVWcOj7aiHSkYCc4SkSgo3xrUO+MQ9bgIpHzN6LNNfPYASzD
4iRm4mxNP0ldlAV9JkdQCS0V5ld7tf8x6HchuFG7gNIuOTr1hg/qRfJ5H3KpQv/i
TMt1fkIS0Yz5uAFkpVhaQTlmU6bszfwKYoaXHg/TeZ8uwrpv9+O/zwDhw7mv6lw0
f1peaTzkr6gjX71LsHBqbUcoCUpWDTCDm6LLeY29FzP8EeoHci5c6ajHT12Ce6MG
LjBwN8tbNf8VN7f2/QUyZTdcEEI4CrVTjxBH8RIW2uINVjo5gThc93oiU2WZexoG
i642AGLHRo1zjGbVXCiOW30YFyK+abfNQqNV+WZ3xSx52XXU++19PDH93P8aHgr4
MGC6UNfUJopr7eeyf6ckR34H2gMpHm9NSeQkeiPWmHCdxeofO18cFaWWpyUIgbbK
mUDw8PqE3QoNhf4YGAAbeieX2IsKKFO2W7LfPFALvrnbt8Ulm2u5rXUzRga81FVA
UdLidHVGiwpaysHNVZbeRs2g8wPmbWcE4WFX52iOy7G85uwXQkTNrzZsY85n4LpU
jLFK4whdFDcbeFBxEs4lEALLPSny/PojYO+coNr5+7ef1TyDmnTYXKhhkoyFpW9D
zShehVD3dT9PZ0ohcSpKWXdyLZILXkmqlsUV91zs2FW4R/O9a054rucg90tcqT2r
iJbshMrWyc8q8paVyBHY4MDHXGkxKUPk1RlD2u2lvvcB+joZxe8zHLt96szWbP3I
M/sbhU5aoHpfmkpuG8ktTt8ZEGte5z8Bv1jIobreulfZ28nUqfMGbjm4rpfkNO5B
tNYBXeetwbAPWI09WCU70XmyfWoKzeCmGfven7s226HgsExX9uggGmYOpyyStHkY
25yaUEpnEgRhN9ar9WIKGMWJbGpaGS0pnYJw21OZC3wT4/Q85h7/0TZqf3kOJBrr
qEBki0gdJBpxFuh+gT9hdY7OIiSMYfSb2wEMoY9T8Wh8g48kP83FaljvDlCag1xZ
Qeur2dF9Tz2hhDze/GUoYhclmrCsqTjAR+iKhpVF4IC4obU1ppx8JfB2FDjg1AKB
UcY4tTtKYvLRxcGvj3vHDfTfMdWczC7Kbv/mytoIIcUFja7alERG1pBUPqlCQrb2
y7Y14TshIXflFhTCqLlT4aftE3RvHBvUmyrSPZeNOtYxH+Yli31C1Q2sFTMw7HW+
lwcpI1KfLnCvfkqrLXCdkxrNQoSqDPutb0A6qo0T3SRmnICuWxeHVjVEftGZ23gm
4SfFKUSiZhn/zJNb+CzX4RPL5sIhbRHdLKlQiZkFdEQ17VjxSZxPkBFCWg11EBv4
jHbd8kJQsW2rujxra6ewT8nOGNVxWg2RZWOYaL7jvjuZ4pQBJqm8tZH1LWzzlyXb
jG8zzgHVXNHuQx4D+3WUJ6LCy4y/CQq0ObM4MM4JwxQPJE4RdZG2gfOJgaijrOHY
X7C1CXlQ+Jc3H++KwasFsEd4pliBBfcv+4lIL6dTsG4MFojuTbePdid9AHRmQ1TN
gy1GjUBMDtu27r7Bf8g3iP84Xj6pKgK+gHJarHPrwg8zF3XUcPYKXbz5reXUHItC
JiuENAg0A41Rw+y4lCOuPx2GlUspJ/CrgMOTQmqEujOnQK4SupgBeO/8LQpGO81a
5G0G5wAhf7cmk4QUK8S7AiWmeYDqhmWaUs89Bs00BlLiV5/4OA6X305lHweozEcW
wRKzcYhO/6nUMhKJ73nxCk6/hbXoekjEzFV4m+F9ltJaHKZgQPl4Y0RsIiWJns29
wzFv2mGVKRIU5HgZFEmnJU/VOLQBkYlM9ycNn6GEgPC7zsOE+25gw0ewXHabyE0Y
inW7AZkEg+lNQoZCGAcY0CLa8DgtAw94f/wHdoIBSd/Y0OMjUHKpDFW+wfIi+SzP
+SVZM5GSr7ODHHEd+M4z8ve5jbTo/NSTLCyuIEhF9/GRi5esys5B8g5+Uzvh7tt+
5+XyefWBgg8cgUTmcUlTfrZi9LCNtgjcAR+eLhKS5A9dbZvNP9i0imOobCAiDgE5
kTNRRBau1ml+LpilBpiPONEWnhRP1qIkB2+/4ztqegYcSi2osaJkKqRBTSeTdgIo
DSEb2Vxh+bU8sbwD2QJyE0UVdBxefcra9RiTCxjKgesgupb0A+ALPCcvWVY7wkBV
PPCh7bHzu+Oa6U1uzpisDsbZfJEuk5VWDpMDiZAU6bWWIHuVeVeOOJyd2oSG28HR
mrNNH5QbXfUTr4oc1tn2u8z+JFkeMkJSKh6cJ7TWZzwwJTpHweoKLmiV0gROKOIo
T7td4IKgG/INImduV/kwi26oVv5AWnVKh7PVaEuuHa/wo8EnRWlABsaYKhe+QP1E
ETVb1LXWGSPs1Pav/hilCByItvS5ZgHJQM94RgEfeTAbLk93dWFPcS74W4dRmLPy
0cQJzUz6Gk9F/Qy64PKWZoV5YazhCPe5jp629lYyCZu7OtpSwuoVsz0Jg9Z+ob6+
WU6J3qx+bsO4jMtgjxuPtndskwyPW2dPOeR0sCXRyw9kwKP29yuHz1v73Ls1yH4F
OG8fuAWPsWCF5yS+GlHUd003AqWjX8LQqw9/M7rR5e8Hyt+6i8NQq/X1/pnuNQP0
Dzt+mHrGOrCwEO3QlmmZUfmzG9AsWx3Q9JuiUtUQHcujBL4DnjBiZuNVvCs5qmxt
bq/m1dUfky1XNTrHU29O1yzYHFgVbFkv3dmoxk4mJpi+7jt2J1oVpJv5cw4sxrDg
REYYQqymUU+IGdLl32cyOklDKRDm5dE8mVO9Wh024Vkr94nRId0bhWthEUeIr8VH
k2oZ5Aow09Q2iegZdde6Xr/utShqKoUoJdnc31EL953nJc2xaT6EEL/iA0w+xNtw
C9wZ4jbNjNS3aB0pE8N5ZnIEanfw42Euxz47+qUAjAdlzsg+y0+7Wr85PgWQM01Q
zJuQ0VJTK1uyAEawA0pbKjV7R7CdItfIxRoa/odca8DxhnfCMGneJk/XZzGjZfC5
8nWTBElzTwdaT8LI4orXNt1XkpyhDyIqylj1IitFG3QCbD1Eeknl89oa1jnyUubH
uvS37t3qxgfaUv7jIoq8DTnk8E0Aiq1H/klLvshyS21nUABjVGF2VutwA6jT/l4l
kds4d9X1vwdpYkBaLkAdlLp2RyVL0gfuVTesfYZeM2OMgvq8S6TdrYlc38vp5yT4
HAMLyd1LZl9WH8nd8VNLq2WI/gsSrY/ey3hdHzCXh6jpAt3yi5ZXUSkQFQu8CL4L
S5db1NYpZFfi1dPVWk69VFG3uoeKBzOfH/PESdeazfr57ymXCZS7g1I/TVuizBVf
9LITGMr5PUBBKL+ZUehQnDHtBv2q/NdlirXSuxsDbxm3bkkF+xIFg2rmt4aohh64
LDMWpKnnhKQfjqqlEGXIcbMDoqnCsd0RDg5TEIghepgdrJ9WSCusawRqWW+ENm84
jr/AYJVp+HllAwhy3ieaSq7Er36fh589GZDEJIY9ViLJ08FAwj9GbydMl958DQy5
p4/axuTK5WBKKXOA0uWaeqGanM2vVvGWygGvvGDInc++tTPDwCWV6XaKlAQdFPvz
MekGUN/pAfj055PP3ZwW9bUG8wEIw6WbbGN0bu64ENBmx4jYQovYU+KYM3zvOlao
M4jBrmZmxLnRzmWaJ12npRYlWdVssq9LYL03AphAKiZ1KJ4wPzlxHyx6xa4zfOlY
Pagd9cMGWb8ChKEi9+M9L2gO/tdHqAe0a+rqa1bLrlw/+d6gloRJSPOhrmeFZE2E
yYhQtsw4QZx4k4TrteWoTTW+caD2Kb2JNW4E8SYManFrwt6H/bcJfDznlBJHxyDd
qLDdyKXli63DYhvIB2KXa+KamUpD+Jtd+n5kE5pt7fK214knoAfWyZ1x4QHlfsXv
DmOCklq7ESPe8WXQUoLcbyANeJSqXPfCtKlYCCn6YB0aJaztOtle6GoezZQQ590d
2uToV5uZxmRl814pq5SnXLteNNpjBrQn8gCKGKksz/RR2v77Zy44cEpZqffxsbc7
7z4h10Kd4wpUml5gBiOIgBzfKpwe5ZzBGflwbX5QHaWxzEVrQnVepwbJxsTFsD9l
ckQcRQ57kpbkSepKznQIThFD4WnREcMMh8e2e+boihvzIOYzj6tQeQO/RvcJVaRb
mALHhV3qwAXb+f2eH+nlQ9T41brQzt09Tkx49vt3StRZWxmNDUJUllpJbYIO8hA3
Vyt8IwxAzcMsdQNh4AgVKCKJLT5gWti0nzTekUq5XJr/O5gLaDhOjTX043Ng4+Sd
em3SJYQ4Xn+xtKFxFcw0da7ibptxk209p1/AT9oXbrWYWPq1dZNOLe6Y6Rlvu8rv
in9JfjWM8c60TBTqj5jKbYWymRTnTCXIAMOKjUR4eSMJF73f/Pz1+C/PnX9Z05NK
5Sq+Htv/t0hyzXngKYw+9Q3qh9L/IzMWtRFwOhY9e3kUrheqcw+2obNlZSr8SCXj
oRuvs+YUHXPQZ21eIPL+hJ0DJmNdvA1/Thz9XyXYa+tqSxS1pRso4gaO/9ya8SrZ
pA5qMrbUTBh72zWrLzYEb/nCfWj2nAz7tP063+FaNf5LOmTgSe3VXnhVIx2i7f0n
r1DUV6lsxF+K2NejQ05PiC4sAbY/kI5Ynw/7gxdmJ4r1vETv7yLAMzT9hLd12c37
cp5jk7e6VMs1iEa8oWECbWXMe+0O7iLETx/LvqlLsV2Uy/ZT4cD4enlfaId67Zqx
fxFodpM/WZ8HQz4Dj6DEee0icdlMXlnDhQmT7u+imPvWL/uxyF09AsgRd5zcer7S
hR5oCnaFrwBLIXvpHmeVxXxoQjoE/5yfaQTQmLuE26mlnC58ygdlbE3mSYlnn2yA
5Y4eB7jx6lBUGk9DolYGvRcpgGCN0njwONdlQm+vxtGkhhGzwTAuACQCeUhL6gTn
neAUcQLSMgYcxPDEsMR/lRtSnJwCrnHunZ9qtoRn2z/3AomQNSNOraP+i+tf7myG
dwNSRL8Bqhcrue+Xx1sRGcyEeyNGFI812kx3oeE7ugMejl4FBBb0youIswzaUiAD
kRKW9Vc5Iya74oR+LRQp6Gjzmv4R0d/j5WEOZsBSjZa8W2ZOt4bi8kGSavO1uM+0
xtnqnDb4bc2rveICJFgARykE8HKBGxBxMZx7TNA6DbrGugTalbBdU/G5NxlnvknQ
/qu/f0xV8/MD5hAmy+zWxukB6B1eQlV8TPap2e3TyTLleQXdNIGNeXKWNzIj69dN
ivKwf0MIJdCjXa6kg6G3WNigNP0PqfPB9Ll4m0ti7gEvNmtfi/w29oRZN6Ayp7mG
stZHDFZy4MONdETk4Qq9/3LLqoyueqWRPNHr85A9UKgux+sfms9jM9gADOGycjGF
DnD23RvIAWV9MpKz0hstYbuTi0idKnZnE+6uQO79E5qm/GIPTCJWu4S4r+cOKcM8
bRw0Su1gBggnKRh+afL79OWpPUESs6FtSVm5Pq6as/dkVqisREp5x/KX6O5Abg9O
xwOEfx0lfwrx7OhV52RyJPGvcAsZ9F3r18VGuI4D/BL/OH+wMaQPZOlybpQmPf2U
H1+s0NFmiEuONQ9IfWlIlCdN2De6qtdlmrlCo2kxsoKun9zQUc4hVMoFBIzMk1rl
8Ht9ZRMD66QNyLQS/WWYPuUzxy3pj5bGxcwC9o0pODtmGB7JFSXa8hHG/dfiEr2Z
AC/CKC18rnPToG7V0EyGLA9HWQYHU+I2n1rDZrHoHUql8bTOaBGjKKiKJyL2hmZW
AebrA2mnYO+UEBRnSknaIUzNeaOSljeZ8AR11PvIVrN69xKUj4JmDK6dzOvNJ3iN
7hBYchpTSLrKu9FE6t6/YiF6Sjle65Y0PRAgXrvxfDfFLjSpW4GJvPInPrhJp6nz
NCSjMtiVf/y9K+b6RyAAWlMXFEmTtOvPbC/Fd6xdITqWvHu39bXnPV0LlYbDP+xf
ADulCA4Ojj11DBd5HF3Y30ofTMlrNoK0epHiUFIyIzyJ7tzxQMOwCLRTUrDcRupf
HcWVpCRQJdbLEzyKZMD4RIaKMnMmdiDnB/FIAaVbuZ6BzYUYXIE4Oi8Dfj3ZEqed
VIf7ryQhh2p5CPBnHFJBMvMmD2pUiRjiHl12A8Rg+S5XA+GRVA1RIiarFPpd1yTn
GZTYgi1v9YZ95K372vKMu/jWOJvaihfgyn7lAUZwQWEo0Civdq+X/fjL0fS/mrS4
pG87tFfHpjrDHxRvLX80ltd3vyrIvvFD4hocQHYlGM83x6iksaJPVIMiyVGsUay2
cnBG/jALX0V4lnto6QqYYcvLyFivD9gaEXu9i7H2KGkZkOAVlOdB/oDiRCbSh6D0
Wm0IQyt9ib0c6rJInbfnuSexrCNnkL7BMdQavfptgcc/Ulw2xByhDNBwGisAoPWV
1gyjC9VXDLhA9czra6y+RjEy5QxswxLwUT40mYRduGmxSIHcFBHt5cpc0xkuNxop
vDrfwKmS+KwikJhQhXbQejetnDUQXmY4HEfKrm3mtQMHhaBjQ6A+SR7sYAgCXh1e
rH9da3mb7Jp/GABaAhpZuAFkphqGXE067i3jMdTIJJQckyNyOWvbNkC1JmfKJu0V
FwxciyjN5mDn/oVpmtXNaK9QHuDDs/z1EF4p/zv3Qm8G5AeVjLpDuFn+uAX9OS6e
kpVICt2zRzGudJiFWCXyvwLfnImJ7HT3FqT/Wx0IpKvEJUqwsJjXVxQBffSoek5s
UzippVNZBK/HjuBRR2Yl2B6LZYcRGX6sPU5Wh4m1PCgzbp+24eCF6KNgHowxE8es
7F/6xdPNZDeWNMMd0whMF44E5uQgFuj0ESvWVtNoFPamIfHM5Eq5vtPLApJiMO95
vNQ6k+WRFcy0rHRYQv53cayHqhJ+CO8OVAY4u2Q/yMw4fjPhPxf+h0GDGkoMR2vt
uvnl7P+d4XHEf6lpugUOo1bJ+qzkgqHP+Ki9tQ5TwH0+wKM5PCDj7Yp4VIoWaPIZ
zfMEM8XPdQAwMUXSdIZHHZUQBmvu0B6hlm64g0HAfknMbmqNsnn6qeW8pLRmZugj
35UM81gmOk+cFEJ3U33rPGFWTIOOOguGwwCH7eebchhC+aRlwtNiBE/DWzTZUTrR
gbBhGmom2y8SNo8utbE0aCxtKbl/IdiKhxri7M/u4lWav6JO8v4PLTNirUDRMxSp
wABzFExaPr1mq1GWMVZftEhBk5VWGk6aaptgWSvy1GdmxS8jPbcCxfrFij/pZl1x
6K1D16CXFA9auFDlBekFkURjSBHrDVKvcBk/IxGZzuzMJhoASnww4ZyRq1ctjs2H
pCuYpNXNMiqW7AlnTxKUP1WoZK+XdH1e/z4NxUzzdAopK5CHwMDDvWw0bbxUa7gk
v9qgd578OKHPMv84C6/oYzErBUngnopdcXdIylMpaiiSuIIJkNuTI0zpYi9sqLQp
hmuUT+DVjN9FgtV0JVHVLwrZ/GXM/jh7ZCEJEIyhqMR4zwiqKPIP6vNwhVh/apHt
AwpnHnq0Rw581l6PMkRhC+fRoB8QV/YfShfvpL8Uf+rywhIdMAih2Nt81z6kkgpf
i8WI1aP7aKd+Sb3qzaDqk7ynDqh+0BBx7y423iqiDJb6Jvp8o8vjwe+QKTFVmnOV
h5JjuC02zXtiGg1C05wARMwSI8ilE+0rer8FHNRvsc3il3sjo97W833/cQsvFv+L
KJRapH38sKTEEBOACOY4RlJeG4i1Had/ksxaqwGe8JVmplcWSG8ndGQQ4QsH/mPM
3+MHdPDfn+GVp9MGufQhgnw1N47ozrwXsU2YAUrFwD/DVtSq8sumKZsK811uheNS
f9ChTA3M5AKuzzffSZMl3uXZNQl/S0XqdINdGXEnTaUkzmeYvMUdAWkL1jCn6I47
6ODYAarNKiZDd4g3MDSK+1R/entPiQX36FaOIHq0GeJSNzq/eKNuky7/qk9wV5s+
J41wmJebIsDzPy4RP20of+d8QDa3X5CsvQvkhOBSj5nWfALDlht2MNeZnriQao/N
NkrEBzz/jbjcGlWU+yXG17gFCjnCLD7/E65qzr1812nm+lEsjuKR8y8Ux5vSkb/R
PQp8xID/ew5kudT344X4sLLcE9umgtCY9wnhztKppCVPuR2/sGnxlQkNxkkcpkE2
ug4FA5tFa6wi0Ww7cN/eHwIH0vTt3IZE6/sQISxmxE6vv4irp1fml5RHVku4D7Bu
yzLJUw2DsWI82eQnZSrBO9pFqpn57eHfaZj3UqFlN0eyso+gZlbccO6aAbFJD+Hy
UnyKevXoqWuxMVibylgDyHLAOW92SjB1bwk07FgdTnHWiULVO06hIh06eID3KGma
j68VGZVLCdPhDm186l7WYj0EOfVmRcWMtU7K1I0F0dSU4HE7X+KWICgbIUYBzGqY
E15QmQLxQ+U7wTvNTsvYeQvO8FcX/sD9nMEqKofSbvbmHkcZThjy4AVHn3bePwki
LLG57wfpq9JIxQSwkdmmGIj6HJDsNJD/93pSamL4GdIt2xvk9M/MpRTkMwVZa34v
UY0rwIenUcORTH7w7hO+W29uZnzLrHBEvBI9G35IZ/IltaOtKtkGi/vAH75IECDu
Knk2Dn7wrr74v/Z2+0MGk/97PUAz78qPufvIZEZsYsxP08T5U6TZoHB19FjvkiKb
84UIOUmVJZc05q63K1mdAk8DZkCPFnwYswmmyO2xpbxcXVBvrkHqENPm0ZMOd7j+
FtpR/YTSmqNrHErQbqzBlYtw/OvU91+c2xPDWlfnwqQZOYEo1mbfb52Bf/QQbvOA
HKmI+hFVz1AFtBgZOi8VPMwpo5GUWiDHFTpoqYqzWm2n1RTZrHG1LOEA936KrhEy
wgvhj/PzoP2xijU4TwvGgefPZWQzjF4TxWfuLUDRFOYuAiWRSiaBNlGxM6WGVxRG
7Uu35ezMVM2UTUupZR2BhOotKNz+TumkZRLaltF1aADwBzUp+okxUsAdNV0Lk5Ub
jhcwpXTreyu8aefaeqfEIfFLOstnCTzhDrWiJCZzeIUW41nO8H+n0Dg1wqca/BOn
zMaj1InutUof+m70Urb1qSABujKWqoosgvaLDGfC4f1T1ePsfcBJlW/RxL2Lkp87
QawZhtJMjUcZpRQBe8gKdEvQOjuRYHchyy54aDWCj21WanCzgJ6fHkdMa5VTje6v
Snc0sbFs67TM35Of7I2OvLLk05Wy0bQhW9hXgBXH1ZDK9qI0rtrWcZfN+aB8i+7i
0rL6a0MhbUoD5o3ESp2chGeoxaFwfWOdOdhMZ9aAso7wKUGr4sPN2kM8kuMcRwTG
xqkV1tSye85GVDz5p80CTAyClR70fJZygI0ouz0g98GT+1dl2NV+igChic34i/zj
QbTQI4Ly/OSj5KrpHKop2e94P2BTxrT/t2Y1BV7UcFlKXeZ1ZLSvxaJwtBNhMRll
MPq7jMupSGFXl7WhMgcJGNcGn8KzJg41k7GuR8r33ThtoYDD1WvG/2qQGX3ge82C
1XvmLL3FTFEzJJWo/3a8uSA2WFMkBuAoQDCtgu2rGLnj88cqY+MNgm/faI/elSyX
jB6VV0tLTkUOffwNI8ri9491G5NLcE/M2BpmRj/mNyk5IeVqE205b/5tpoG4C1cH
zWVCd6N4pvIpHeKlAKRzZkOUFyuSKHzUIs3oBYP/clDRQadltif8X+K6IoDJPET+
Phdh5HccuTf7w/5jDw1sHSXbwlx5YoZYDz8LAPWYADBNgS7o094IAX1msBrjqWzD
HkR8G2wAcW6KciCpXt76RY+pIydDZa2DMuSVR8H7mTjmle0PNo8ZU4lUEZ1J1Q29
+T9AlJoEykxBDN8u0oigWk3oPGZ96STLlYOGjkG/SkeNKjpEbVE0Fyzifmj5hQ1H
dbtJYeZAT7r10b2zLjmi9xWTGNrHH/Ri+Gt9tV2wU6HuJ5yWgvUHrG3ptls6besr
vboU0uIqgkikKKa+9d0WLQMo/Zj/AlzY3LhFoYzhshTuPnNJNTmhmck1CRXoeDbx
h3AJjsFFT67HgKWQ8yGgZiKBy/M1BAdkwPADvLrF/iU0gq8Jf+W7KiuOKS56jQxW
vre+bmHKgs8iMxTROLOh52vNv/sd3Rnhik/KN7keDj761Xpkv6bOESDsnvhA4JTq
nwuyXp3qUUN1wTWpRP8PMTrzbAjaBHMSJ/AhXN6bp5udk7GLn9Fa9FeqfzFIIlFn
Lg8Bgiq07+oNWyGOgC931yrlVz3tLgq5FLh9vvbJZ7sNp9GZJnVyVqVQoosgyIeD
47AEpjc+3AAM5Xd7aObqueKM0mjQ2hEudokk0Y1K9Axpd73pXNis17MYwyCtJdj0
3B1M+FnhmaNr+JJ8qqq5lGD3sIYAx5X+o3f0efs0ruQLmsuBxV1HBiJiDPkvGUaJ
eVnjKhLjdseyWuAnUELBA72505HYycdHPmhQTgeRJXH2Qv7S1+nVzaQVzXeYX53q
GlvbprXXarWdg3BC2HFhHxPBbONgG2eVf/3zRyIt11hsrTqU9HgMIvTO2oaOzuWA
kZkejGcQdmXL4Yg2e9CbFAFgwsMbEuHavr8ssbNLevXbMAmPQ0u0lXI1gUoe7cN6
aCod2+q3lM5BWXoLbDzV4MMbEWFOi6E0xk7iAlPN7I+q2yqss4Vjwn/MeqScvClY
EZBEHopF1LQG04mm1AA16ixmuFm47TENX9XwpJFjMpaC15VQXonYPrGm/cANJrFX
f3yGqhfCkuUevQiZJJu6Q46xPoM7ptkwBepSrW2Ugy+jmtqidB5TL+Rry4AxL07A
Z+7QdCia8g4Q3/OgyEwlt/kiwuyRZzewQ0RJeUXtLWF5xbzX0FxyGMePqpmqQ1Tr
hDRYDo7Jy8DLDIsfXIsCyyZIImDGst4Thozh/c4lxU8lHjAlwM9O1kRpbKm8mv8c
Af6V+y8rOy4UVtTmqx/YsAY8JO1ESfCuOclTQEyabsW5IxjMiCK+3uJFBQRM+bNZ
5FofBkPitJM8p8ehaasiKSRwlAox4oMjxzHMiPvPDFnSoT5sPVoVax74PpPIRGAd
VnkDbPkZzCr5IZO1RKje3khwljZu0FglQvcySYWNOUS7FoX6IXbZ8GeBBRjVgnYJ
iALUx+W3wEkVY2TcDr1LpnkSi+SLLY9K7wmqFlURIZ+DQCrm84P1CR3R8GM3uZg0
pzOwt7Ci9VgA+uqI3/sVKvh275QjDSTjI8/e7Zoh7+qxep2ey/OT49zs2Zuf7RjZ
3wovjZBog6cImOljzSy2daMfqUo87nv+GF3plQsNzPlSqaeRqylI6Xo+Q549wgnS
wH14r52I4zLHpGDteQDBgB9qqhMpYyfZ9T3OKvlWbnmMNlFRsJaBBbv4PUe8gier
2UBcs3vp0ZUShkxcFUqEh+nWZcQq/WE40IfOw5OnoTzvhrLhIaU5AZpJl44D46og
Fs97T/t9w0Ec/fiEh27C8gyVOj3cUaUXULNWx/r1MdBEbCeR3Mi8JY+fKhQLngh+
DH7psDZ4E6CHwbZb80PLqDkKR25xzaNgi6/Q5l/+6aiRe2w1XKajcnjhoKcjIRTj
4BuTXeg+AgvkIO6DTJfPt12WL8VSij+HQGIvnaXRIs4V1huLxqoxXwkzYYB3fUQs
PzxFGkYIfVhZY2ihk7TYmPl7QUirx1DrPnGJROyRfasKtO1kV/3F/KqfdHhQZ5B1
tlX5Iuy0xfN5oqKXw313lvPPnpawXtLSNGQmEj/tpNngxe1bc6Kz32du+kAGrAUN
Dq9/lUrDfB4yK/ldgYr4hos9BMKTbj87whf8FvgdnMET5zAB6W+CNI1D270RrSXu
rUsomBqNvfqk3ytoUouqvLkDAzjUDL1+lt42M7df6sZuFzpGlC+MMN9Yi+82cten
iwVdKprR6T0wEIKzxCKqLWHarKmsBdBYrjR1cLKojobJoI7HXtp/0qIGg0CSSklN
QcX2NXRFQbd8GDLmKRy+G4FpOd1kjEuWysMXzfE1uDrmQctS+Xd60LHjlZqeqflh
dEUlFLKhPBCKv9Uy0eUqQWwYGyYZOMVhcqgI8un9i4g5jZsQ86UExybzP1za4v0B
krC+4T70CbQ9+FuZBeGxuYEDaxsOD5jLzOkIxQv27Jm8LCoM3NoptlYtBGKr09Ew
EgSRs63b9Z42GrNsqTKFUDKe4jfyqRaNQOT+LCzDu7zZULnAx0EBF8s9RTPjIXd2
3DX+N6lL8oOcJQ8vbLvsGmZ7HqHMLQM5FIPhRIImM2moOVMnWpNeBaeXahsBDS4g
OoPTgtUqxjMkg+EsaEn+idFdX7dIIlQZG9UhfQb756AJFUMR91gYMlFDpPmhN+wL
wv3hsc/H7gINUXArUunQXNalTuWVA9Sos27KANbyitT4RDzk3wHDahAZklWJhYDh
mpIOzEIqaIazDG9lBBnIMu02KGALo0bNvPN/+a8qBHzHw0bT+IA3eapC5M0Vh3P7
RKJMt+euaMSA/O2zpphpKMcOWhUOxxzoLVGr3Z6TmUYt40bGE7jEx0UvZT9cDCkA
njevi8iSpNnVzaZroFLdFne9nj6UNh8lBV3sDGmcXbGEeywn6bE77DZlva9bRgwq
61IpB1AKwxdd++t+iO+RrpUWGU+X6TnU+hS8CJFV4COyDX5dO/HTfbPMISaw+pGQ
d1Yu8XfbpkwEIFGh0/wXBRo6m0A8xpQ2NU0/vrHJ6YsBT2wfYQhrcKP0rh+HFqsc
4Ya5xXtdU78u/8vq1WQPaIyEp3I2O5KbSQKyMmPpNcV1Pf1lruHqy+KbEKx3gvzn
AZy/FupaVwYua0M7WJoXFuaB2gE4bkIGXjjMVlvzJNNNRlUPg2UgG/mQR1zdlHwj
AWOAA44HewHSFio7v85fwXFTDsrpzqt20LjUEan//vkv9WULVYXbVvp01MC617yC
isBcdBnp2Mye2iAd8vlckn7qPxwLYjk3InQ0qQrDzdSxt0e3SzVV5hHvle5qCkxH
oauwy+EMDb+inGy3fB15lYCKknUx5KKTU4CKtAohnioElVteSKZRtMwqaFVdfW2g
ia8otH7KwEMKUWcSbRc9Nm7u10pbQfkX42+rIykplNe3Tpb9+8cpYjNjXhq9x5Qh
EYI7Hb0KFJo6pBs6r57uciAWEJrZdfJB5th7zt0yvKk9ju5obODwOhsp7qEPKV9W
BgvuB0SAIHUS9iW4FMdEJJMm/y8kuJGp8GmvUZlH+snOEkrP1Neb8c5M7AuzYgNU
XDM69eL+vtD7TgUlaWRPQRnEi8HGvJyXbaTEqoJ29eByWoLlxDtXQDuP+tkPrv0R
k8+URflGU7Ub7/HmYoUD0dblp4P2TxV6rfkMWGzbNf9gtJNzDMop2nsg/9jzIYH0
taDolfJ1hbyBHFDci7h606jp4MYJn5YRpX6mW85ma1aXXPss/hqDDosZs0DOb5Gu
n19ZQeiaz58H1PlFrXfOLz5Jx+G94Fo84s1iGwRF8E/j9+BgoCFVgCDTlvF0CSQp
L1ZJdGJ/bzoDq9zeH16CXLGeFRWa3cN/iOMvYhHB2NDgiIvZUBc983Hkozr1EzC3
jwo8RqSHTzmzIbMd4M85kJoRF7mu5PGjUTB/gtfUib/Slpn0yykazkLCugemkGY1
QiaUPBKxe0koAJSazIxjHenCaJR5KVuHmacoH32UePn1QScckpxzmXlzqFUxgWrc
dkJDGaa9B5TAGkBJ5ZouSl+rHF2r17xwDxOaD4ik+VFmWtvecCQ7GZ0TyRnYT0yE
f8ZQInj2S8WMmynfa17egMfpsFkyYkX/8ifrwQqFOUvjwEk86xVEA2D4YhaR21MH
KiKaV3BP+Jz3cNLE9IDWdYvoBbEErzlLGAl/zNwAyg16XoapLc5lo+3TCtuNzqQg
ZhVIA8NOiCPaI5pRwlbUtFgiZtN1AH2ls49B204hnfnKxiXwoUtT1ZAv/0/4JsZt
T8H3Uv4fFq3NwKZqEdXv0Ip4QMSBx3NCEHm8NLBf5j9Gt+xS95ldw9pWsT6j4mIn
nVQDbbzDJA4sKRdK1aOmt6SS+t+xoZy+kPWqVAdzyMh+Rfs3C4XeUEThlFdQyi54
ipzjjzSxrKEHdZxQQYPlIU0dc2SZrNjED/lWeAVoWPdFwHbgv2NCsYn94/Gs9aGz
FMP9cFPPif/mHbOyecpxeqJCXGAXDZHJ9j3A9njBCeWAbPb7EE52Vmzr0kXG9Jd0
0/ESAymXynNxQ6u7jbVBxrobkoq61EpSXrRCbfOaxGG/WPOonqUpTCNsMPHhPtsM
vv+vVVyPFXq4nfOhXFkTHoTFFDBI6YiJrLvUDSa4tg1bNF18OY6S1krDJvlyU/3b
cMZU73H9L2/BJ4eZRoC29Aa15TXLIZ9YQL5BPwnLmGHL5saXKCrfliqWIHafgwCF
ooHvapw9vp6EPRRMIxfQS9SACF+o8uZYMRdsf9NLnLELe5YRUzU82hpbdhycQzFr
5HLf92neaoSPONvguU9tQfryhu5tCW3r1cWQ0y0gRFjWpsGLXODGQWfaF5fvf9aW
Ndl4yM+cjUbee7sakphd+m6+uyhsFr+bnoMRq/yv7Z0e9tIp3mUJoohiX9oj0xLP
hysu6+1CdB4Gg95GC2KB0fF9INLRuuYcYPERVzDhl2fCReHhLoJM93rPZ4CmVVAf
HCtpLe9O2LMP/ba4J0I8a8kfdBNfl6nQZQFetP0724FTHWi3VX3R/sMe3eoivoXG
ao0pwDPatHA6yxpsy49RmTPVHuGa231w6iyorusU0GJ60UZ+VNSRNTCkJXx5W0Nj
Z/spfW+NYk1mI8GloDdbZ7efSCHoLwA+JVXXTPyrgrUbuIMe8JH0rDICRXWXdijK
XhSa8ljRFPmHPacW2fTGdvtQQf0KRWTOd/r+rE9DTDjD/6NwTKDyUWyXjgyLDbVV
gFpKoL24QKgC1OIUm22pyGaqK4ZVqZVVbn/CxKJzNpKmL2AtboXomfCYTtSRmYHL
4RwgPmVSSCQ3aiX6vjVh5zOrelXJxbILYrkmSvVaUXeWLuCBNFYsgn2lf6hroqCn
4pj1zI34xvqRClzpFW0EdF04NsnSOyUycevRVNOVUDG5er5+obkPw/RfyVG5JN3Q
LD3M5kiYAwfYqY4moaRtHJ4Hjzb50gBL5yfHT4ZIgQTrt+cvfQhNii96VsVRWy+s
4JRBviaoEQ2DTeqgSWssGwAXrXgkT6/IDDWBoUKdKdmFR3Y0dJRz80VsilxH898z
EsRjhgq6lj+j03CbeWB4G3TkGbdBOf/ID0yK3g4wj4Eg7oXNzmV6c22xM5sNCTOO
ktBAjgH8vctWH5AjP7yR5DeQGy7nvDrqjbAT1wzqqGSLIR57/hZQppVJJdnX/+le
xrioSxPGCsOIT9GwMU4h69l2WaZyX9MAEtSRDMUgVOI8wP/uvHzz7IDGyXCaTDCC
fkp+aKzhVs4gFdC36b7jxMhaDe4XBrcIJOyOhyZVESeIez3SLGrgdbYVeB7CfFES
7Ti8TpA1OMxhmaxqZF+/kRqRC/3PIeFkJMtAYxZfy6Rk9or+LexRmJnJVxwEiuM5
BWTeX7Ko/YJ2ocTiotWCqC/1uejro554owENaqSXxjT+cyr1BBXzfHGndve807QC
MFbti5F6NPHIYSOj2DsDcgFVGjrnnM34udZTgM33f3/YAeKcqj0HgSIsxI5qEfSg
NaFZ07WucQNTj32KZ9WQOS2pZoA3kK3CW+tX3dmc1L0BJFwCRRLGrQ2AQy0WXWaq
SmlKTfvxOtBNGw9HbVpdDggtOG9uNh2nXPxy9REaNTKOL/PBdc7tdt1HJHAAdW3Q
nTmcSEhaP3bTkLbJMfzup9goL1cGHHNqGjwVCYKKqlp+gT5iOiN1AI0e0WADUDb1
1lP5fuQAPOTPcAWKo5pRrd4YW3ySufjT4U4dZ0f+cOiPKYUcKEn4cStJVDaPmG87
E2IMAvyACT67eCj9wxt43TfJicmy/aOWDby1nHRDynb+4KE4m9Fzh52lPHHeQxUH
RYNO3UcQVwye0njv/hJa9DsclT9pts3E4A04gVdDJ32bZr/TytpPOmt5dNJ/jRzo
CZmxbqKL5bv1ZUQJIBhK+avngiAO3Uav30vB26UStlNdr1zWL/9oxMXn38cvpA47
nQRqawuRGTHa8L57yO7YScpf+8X7ExVB7g+SmqqMKq5Yq0HgxSV9nKEoBez6hV6r
9PmvSk/vM1X3bJvP6r3jeeOGLK624DX7HJ89x2SmvJwVhraPBSLPpEWLWvGqjUQY
FjN1A5uMzcygbKbwhB25EP6CCSKCz7Gr7yQ4shm8Nc0GH0u19UZqn85cl0vHx28u
dbDIY7EjKTlx4/1RykC6ssLs21yAtSI3L+cpIZWhLO8X3Q7CxI8mVkICDqvGjbVu
ave+LXOgofT5fqLLM1b50EeU5KRjR0HxzqtjKh8kJfxuDdG0bGy3ATu3oTe5xp7I
xburBnsPiFYTWIayKLt/GFyyGxyb5OtDya2Kj3VmeH4T1/259mIu/QzpE8kdVzW6
QXT1LEsAZWL0CFhpIIrw2oOmyITEgLDLv2xXgajeHevui90LmAf/65ke3dMUxssB
K6OxAOb/3C1WxXiP1+HvTV9Q/7GtaJXDFru3izWEMWMKyJT/bINmRiGwOwfqaIbX
19uKGT9RQzmzGEVSiwwWCYWuYHeJni7ZFYJGijnOhT/bnSB4OPZZA4VcU8GMomvc
U/G1yrEXl8bz9jG3+C4BuSkAfs0/ugCKz0CiWomTWoPy0b/+ItYub5C1n9w+Y7Or
Z43P3qKVMQnLcYnI4uP2q06xFxQX7Bb2Cl6opwvKCgISlHHcZjRkLLjRHVPRIR26
O6wmP+B7fiscxXCUDNgztnA1zY8dZIzDByABPd2TxxZD/Ed6aGBrwMc3bnmGD1BM
r36mSLihzWrf20nTanFUa9UtmpKhhppZR0vf5ScHMH8YcO6fsLpNQWOmjoYSpT64
g8p2VduNerUjxKw5VhXGdzL0CDNIeWbHtZD9mvBS+rjU1CE4KuVb736wHMsa9FHk
GbLn+lCP20Huy6Y4jqCNa0hrGctrbpg9Ez4hXWFo/IWujk85qZo1vftXunz/Wf5V
A2O6gnxbTeswTgL5J6KE9Hf3b9ZPZrCLW9p3Gnf0inbc7ekKA3E29hXY+yLqe8+e
G7UryGg2LPPcIAexFvzP5OTdO3SW9z7AcSkz0RYJzcTezceMM0MrU05q9O+AfLxm
t5Ze2cdmZROiJT8kzD4lK1WqDLqW6DgEHBS25lZmSj9ZXrWVXqK39XzzgqyEQmXL
b49zFZ0rITjzz9IDh2HjzJY6xsrDA8uHeDmdtrW8nqm/ZP3lMaVemDVO8eyopBtB
UwSlBpsHtjZLt6fXpg9Ord16jt/UTo1ch6XbGXK/8fIjcXAra4XWFsscN0Y7duVR
hZ8mkbxyv5rmz3eTv4gKTw11nvE9XdLHas1c/FIrTZVZcxpKrZhbRWbCFe+xjgxJ
VvFaM2KQrLKNZwaR/krAdvJNVVRohBBWPMIR9nD9CzTgpabPkRej5EQax3Pahk8m
4i1vfqdLAP8I+ctOq1BEkBbOD8BsLe7A6MGUiCCkDo3llp9/csS/q570KV3E8knL
iwUWYT1C4ZbcZWyOvXG9qXnLIBvAoCtM505WepRapGTCd451Dlz3bpCw+M89fInL
ZdFdmcnwohkKDdzS7vmuQwBv7OtwCq6uORLhKt8fTD+U+McEaxbIovhH/qJqzRZ4
vLVJYrXasdknbGkDE8BReJDOc88xUIIlNeQc5b/h3+ec6ni7DB3Z61Htad/VlNPD
55c62pmoHK1W1yZjF+Y21vO+tD95ZlmO2wQDWa+OV9ugVxDzp8YdKW8iBLlOsnOK
aqfBeg/NOaX9ZVd5HhBcbfzIJG5VcSBQpAIjZhoVdkIDvRYSsWb/gPXaUdlLx2C1
MYY15h+OLxDgd47URgB7ypsfyQ6xe60rfq1wZP7saPJmGPhVt2q+UB8raXrf8U14
/TJe9sBhFfCAI2MV/MfUC8FcOBFyiRl9SwdFv/GLyFLf5dPR5M7C+uW1qQyxz9Lg
khdAF6OerzIkShyRuie1OqaEDhhAIxIK3eDCFOthg2YrxP4PTaLqfCvqGPgZTBFQ
tN9rpigqpEl5SlG5ksggqeDpyluXzQVwLNutMWqTcek5bibnlLStPaUKyrfn9QAl
sP+j0Umryje7jKUOcxw0mUzkyFMcAiW4eeXyLzaOHfr1meXh0qB9W8NnY4zI7OMM
eBKiyusC2Gv3VLE7ueq+GYEyOicjck3sfOUhP4dT03jO/mlmUfdyZJC+fNjkDd96
Ko5zbYKBvhYigxLc1FN0Ld+QV7rU2JNUHUyU9xsCp9qsvuIn/hA6sZwFtQ67MUZ3
GseQJA1tdWbHYWh8eJjPIKu2O4gp/p6ByJ8mbdHyHnFN5OmFzHoB+gPmIoVAPTRQ
o1lsnyMCAnWq3HqEbZJagNj2SYNXILHtBH8OQTUVG1e7Wo3msaoXMR24rxX5nSLM
z/dI410oiHwz1sgSqeIm8Md8Y5yVYxm5nbiToweupeO3N8hzXn9+3xuiDfDgex38
1e9DOgnPzWgpTGIMKgmx5iIp25lvlWEnQoH0rUlQT+HXf/uPPq0fnaTvpbIhCpcT
XS72VZ4jsH2GUvbCut15/X6zjAg3GJuknCxWdILGYRY7tDLE4sMBGZqZQDvUgsGi
XPwb2+34rza9Ld3mBXgzAsUs6QdbxTILSR8zImGKkO4am8ULzPZ5H0qUoNclrgON
8NY9Y8RCIwbF9V+gIYwBGiVZ2r3mmunzxkR56hxUqfWIugbaP+xPTgovsAdxpAMI
kjhkVi5AjWSYltTJ0PdXtJqhnw89m4cYfoeb42e3ol1Y73x8V6U/0JwZ/kxES8bC
X0XadWF0bwxv/cRvTc9PtnV86k0uflyRc2FXqgr98zuT8yG0+3/pqViOsL/Ey0pf
uvZdKWJSxwmhOq8VTu+zAo784iHlxL+sjG8NZz0VFCZk75UnbYFKxe+Q5yez8PhZ
XutiMZFmZK90CPe7KVZzZExNj7c8MSd4lqju7wlFlGvrRHGwwr4FkbuWPOf9FBWQ
WGHjRpXk1gznBJYzAVWnaU77pS1SlSSe89Tz8Ub8TGAOz89gDZuhSOqX5jy13SvA
NDLSKRrEXktL41hpzWqNpOMvTtApSI0jUMq5fTSK/xky0ZkFFOQE+P3ERqk+rpYz
bXeq9hNIqeLL/uBwliYnG4T1tE/vJF4WjXxVVt3b7h/pI6ItGoeo58Pgs4X1LoS0
JLI/upO9OcDqXarM7lN606uB7IIRftl+iGbo/HB6hss6QSzMUSBFNPtiaGUAKhHX
DHGi+YeoMJnm1rWIIMUDsM8T7VTm7QD1TTxup8TLKIaOnnzFDp9+erHVMoT+c+72
QzJqs0igM7RfzTM3sJDS6x3v9Co0fJqXtL2loXl4mIejqLf0uU4cK2J38eNLDQ6u
qhkXkj4GP6QBjIIaDAsPDJzRYYd9ExSvyTUvvwv/YFiZNPGzbYFLMOB0L1R6burO
bqtHyYu2X9GnUrL1HdxCGR52p0fPM56n+BrbRnExxNySyxzJ1zuyFc5tQLpY2snw
g3cxjFO7+rxdE8YC/yMf4wRGH8dNgnq07Xk/b2pBIiBT+QbLFyrSny3+v6sYZHfA
9uy8kIITwIPtar3/pZ7s+VmEpTVJ+BHe66P+sQan5i/G2Chm342h3HOzhE6X1EmA
NErysqTCAnBB+V4ZvCY+J4X5MLlZM9iRGVQIlaSByOxQPuzR9KAaV/E8LGdiN/ts
9iEZ+X2au0wIopyvBXJ5D9uRbusOPvii9cS+N2djBPvaY2B/bS9kJk85AjQFVMoW
lEAFQtq1y1vU+UzJ31mxubEkthxBWdhoXo2BNvTMUVfg4N4g0Gc/PbX9UeCDpOfb
q3fL29n2cy3qbg0AjqpcJjwwX7TMcPbi9dlx0Rfej91u+eGiiLVWDknWUPtC1YFU
Wmz+1j++2Bnapd5mDHrtly5lVEqSpGaYmTwNz2VCdajCWiY5eOnjeRYjLLAPN3ys
Sg2rdlWH9me+WlVnJp4uQtG8iKibmYGM1BtlD8xJEPLWyAo1HXyKkFH/ye43PkQO
BHCzcaiHpfTOY2YkJyYTCHFIM8ONPqLJCq0VUpOyutZoKfvTQ1rtPoiRSmoWVDIE
MzPLTCiDqSRgd7mdhbXdb3ytv1BJ/nduu0uqeeA2c7vxUV09/AkXgzVN9RO40Agj
o4FbrfSV5Gtt756MEEBNfJb1aMmEujQi4CowW5s3cLOIvUkDPFff9rPAwds31JSA
/VefUItrft4qo0l/Y5O0qqaMrXD9yqsHa0j6moN7H870IgH1+JxhHQ3LyqrHMIR/
sXWp8oNEQW6vEd/3kTrLw87oaYEQk+nJOjdIK3TOYjDMsrKWLktSqqGL8rdaSO5+
8vky8UqesgNimPz0Pu2/tGavcWec43G4cbSoW5JRNq8mQn92EMlOzNIbex2/eaOE
6vcOXO3rOvwf4eAhFY/BnGFXcr1YdUXSvAoi11GVb9fW4BGrNcEIGQIRRLMrHH18
ZmQUjIzZzg3Tt8Xks2zevEyRpNSsXgjO44kl7y1PRRDGDdzgvPQaTdZLjdnNyU9v
UDU80AHfn9RlkR/5ZlRki+sJByFszIGY8UbRro5BJavYM+JhLnwvJ+sSqJWxb4Tl
/G9UCwLi3n+rc5X3UiAvFL7SAQ95JSHuj2t3CWMw39F7cCKukx8YV8NR4ZGv4gtQ
y2eBeOO4qlFuHHjyfsFF22eeSLJT6+M3T1GR0IZgbjw6VTWzAEqtvDrGSWOlmdXX
1C6qQ3VvrOabETRy57Uspe811R/BHdCs2NvNY1ammTiVVCctrku/yIcE3xMzMtzo
ypxCDQ+ThVrcdl+R20vZmC/NNKzuTqdX0BY8Vjx2MV/m8dKhtL6uHSqV6V7ZXGvj
XJB1y0RQk309FIHrVo3rYRulmKqrzVnke6D8qCHxK7s8e2B2LApiuHCvwP9Nnwly
4DfV4SmDanGIqqeg64IoALasgUDWJxw/80x6SszS3/ymnutVVUTcvOMdrxDW6/ze
emSFFUjv9yyDE20xaUkmN5SA0+DZf622GgQv0lTDCwnr6vnmWTw3PYwR+jETw2cK
hHJz+t7RPGElsD+BIGAuwDAO21I0SBEYcWLvUyBlQNlSG+mYI3Hi9X81QR7ICM43
6qzXXy811VyPlm315NRfltdlXSlWpa7skHGZszGt63YBew4EWtQoUNXJK7saptdA
95LhRDXFJ+UHnocEWTOt1tKvB6Kdx9/6gFCbfbR1hS8TDRPtpGU/oqMqSy7HvlR+
z21EDNEk/8kxJpIE99CUXm+pAjOYAI1gXeAnPJtOAOXHDnIsjpFGWuseCZ2ClrSH
Mky69cqVVXFJ8bSkD15iPi3L/CI6n7jx4WeqduPz7SY9cx49W6x8dnDi6ysvSDve
b+xdz0W2o2Rjxk94CbODaEwvFnPafGAX4kBtiQDM16DwZMzajpf65nlVVPltoURj
wOyn07CeY/HSh9SG0vUVjGBDN44+dgOqqgeQFZTFciJYU55939CiaePNCvhcZVx2
xPrTsThQJ0P1qG3hPjP+15AfVFOS3AUqpC8nXQH9kdYIhiGhwwSER7zdTcdePGOA
lzaIxUMCymmDf4BtmET2kIiT7K4+SYP9wjNSQRnAiTzxvggWQ8v9F21YQcF76W2W
zwRX1VAZgVYi3e483iK+VglzR1LbQE5SdVCkRGmgZWSth/FZRrQ/0b0pXXTym2Xv
gCC94eL/x3cZ4qAnepAF0ukzIKC4BK6Kp+FfGJF2kGT4/xyur0FmHpwKNAXLSLcs
OIuv/uSCbiJnk0/Bt8+BKVEQC30I5ELsAwiXp1DZeOplyB/1VP74Y1YnZPaYO1Ah
IdxtC5MOhqzDt1sNelCdt3rKBFISn+6nHdzE4e4UPSZPK83+KGvMG1lKuwmjGsEs
dyDakEwmtLKiDGalJKmpOTY4G1rkv6bnD40nO8+wTarY3Y4oNyLSevspDdWva9o1
4YDCYUAcjmKlwhZzpDlVZJGrHCFThwtgqz+tTHLk1DloRe80XjJl0EsOKm8iV5Az
uchqcXkMvti71Ui0q0N0S1U59IhPR6KeT2p992iCAM0CqttLhnw0HetdgUVwYL76
wo+DhZ3Gcwe7uzRWeYykNKCVn2OwjRskSvhL35/y1u+IymWstqjGvtA4LvI78IJR
IxfM5KPElyr5zDhvSuq9amrAPIFOfuKe4b2o0gkJoJ++aczzltsBW5923J4tzIB+
Vm2WPkNbwi4ZX9E3ATIswqfGibeF0xACU6C5x2ac+rDDReV3jl0AK8ozr8s+izBY
Quy537zxgugB/rP9NVoCpE9vm5YE1iXcCafnzkKjlFDaw2Cm2RfBHcis6+CQow5z
5c4vCa144fQLkA2OVNMCVSELl0BE+ODuCZ/CsKv5sHCCQBK+DWcV9VWmwYWWDKQj
eaPoFKH/ObHbVFpY/ORXFuXyMPeL4jUJSxEyMjsJwUTJAkXayDqi5ml9c/CPforq
ucA8ep0RfMQvx4uSk8bqwencBH+gOYPSoneokm4Tvw4yVhDsm5veHL9hWmVafl1H
BX//6nJz0bROZFuw4wN+I4dsON3xAZ2Qh8yK/Wi6f0LGLzSYABH9bbNySx5wffbF
2W2skCka4FPqIATmRjygFABsVRR1T139bRz4waaqDzw/e9i/doqeQ0cAXVymekBy
fszjnx3PV99RahdxvuZGQAaOF09HiaifUbc0zBi1WK/AQnht7TvYPPHOkWsaogeq
ZYf7B+BB3MgU/XR0t4ajYN3rZpAAwdcRRyzebTrL1FedUpgozdFcti5abcSC+hzh
71N7bDLPxP9nqdwDdUZI3lA2hVI9Ji5uzarbDekZ0Ch5aD1bH9RfozanzVpK/41M
DuOAFfhkB8WHw/vbSr/Vmc65TXElataQgMdlITZMva/+sI1HGNnsT4MNlQ5eQbvC
P/Yr7kp9sFHC+Cid0ukI/FRGhNhCKeu7tEeF8TKwGWfr+gy3HrWNLRhPlucILRuv
+fCCchuRCGxG6K5i09sXR4TfRiAkIWwfvjNSRl1tgJB/jwlC6uO+FYcBnSTDaFrD
I/R3L/u1v33DiRb4cqYGR7pxIDgGCc7JHISQoHXzP0NXymv3xLCpswITat0AIWrT
n8uTn+VDcZnrlu9hIUIoGtQsVULd7734N3kRzs4SwRjnK7JcfSmegLTe2u6HLrhN
EpP2+tcrWFnYD7TvYrcZq4Oz0uTb9mTu5aaogxztLvNq55TlwFdMIDkB7aBS9lvH
Tb5OBy1XDJ5rZKymZ7YBgT1mmyGUoGMOOOX+Y2h3VDXXRYQSZe4bl8gQis9krWMr
n+z7qef92xJXzAsuA7rRt86qjBnu/Qet3m2RrFIw4FZ0yiv1I1WuPRp4HYBR2z0j
pmu5wmPeuXLJ4P0ERmC9gDuGgNF9/qX5SRss22d60FHOFwIaPOG5DBdvsSIsVodc
H53hXRfZ7RKkF4zthuhIlfSxlp/VgxeYUPSaAwRKBoP/kPSOSc3dAcBjV5dj0Vu4
VJ17Wo9ELDu0UyW4oxkRXVDfxNxoyvpoJEseQYhVrjLuNti+fLplAB+uVi5qhB6h
BjFNR+avQr86VR9MKl/2sTvCO1+PWiL7ENmVl2pnn78Kj9NlQkUR+gFuOx0GD+2x
yk8fgBIO9ykgjz2946Hv0nqe2aKD2ap9XkeeKSbSI2vyelO0JVTmY5IMYuoMByP2
cBrg5WLkRJujvjgQ7qAv7jrkzWyEjVrYcTt10Q8+XxD6kYI66wKRwdQ4xI5qmUKp
mDCOH6rDz6gxZRuFiTqeiBL35okKIUS+bkKWz4FsBUmwNZWdp1JP6rYL6z+zWhNi
lP72Hc+7u7WIxgX0VvXyOGsyYTny1PdF3eUDJYG4mOo/upkrQVedPtEPuac6v5+N
D88yWrfr3uQkcaCo8aQNwGg4Pqq4xaCMiJKpvRKBTmwxaeC+u4I6Y0PmUfZ4CJRw
MUR1fi0MvBjk8NLF0caxhhOApmp0iqy0LKtAmL4AG4KpXJ7QWqznkOoknXBJwEv6
eJfVklVPYSnM7irQAj7D5QJelEGO8j4+c3WM9GFm3D9nHGIyLXFqEid1Z+HhSvI/
H/FFcgwavfL3362xAiMAUpJlG8JbLw63Mz40lPZSKLOqhvdU1d3OKrscs0i8nFxl
MvH3sZ/hYnFdtOKinncxXR1yATFL8aqJY8bb+kGEA0cw304tosVL99VXYF91Lnyg
MqAXX+ozBC2gO5w9qtsoIRr+l1+dssjPEoZsZz1jqUgaCU41+aeut0VHoZ3ZWQD4
t+9SAQtlCYyEMQH5y/m2Keq93HfZJdIv/gmAZPAP4KmP6IAuXmxE+yYMS6lzTiGn
+Is0p851Z4fJv00ikt9iRPa/mmR6yFMTPhxauhEYpvVHD+udHs4mJS6p7l/vMkIP
g2sC8iNTmaXE0YA3jdasUaRITsbIabTIIgqkLIoLtUp/vYHajwFTgtFPjOGXJypp
quEddXGQC+cZ9E5niwKhIIe2t6kITxHtyNmiQDia3IHxW984v7ltQYBtUOn/ND2L
fFRdWLjhtJ3v3ZRWFqECGRicoptj9ne8Jnc9AqhSH1hw06ulBMgGSZqKauypWIvN
hsugAr2TFxI0Fdl35po/aZxoH5b1E6j3EMdxqpmn6BWyCNTBAykmyesuWOVBRWKd
dnJ8aRWOTpE4xOp9Ch3NVh+al9ullxN7FnHMwfdVamNIxActj359/YQRIt4ShWic
aeQX46daljqLTra4vVoDD5mQ0ohQeIzoQWnVNtG4guh5pvMDq0Ccmo4Ojcyw+TA+
lTBNiCEenrHv7eL6y9JMGWOS3frrVHdbdtX4LNCAZd4Cnk1OJlXtCmYLurVjbmZR
xl3O3Hu4jRLY6kXIJrJkY+S9yUlpBF3/ByGdgiPK/r9zev4kjt/qNURh87THOwGk
mxl7VlVk/Ub9iySix8GhtsKCYBS/rNUKzdVINDY1J2XgvXeu92QF1UVpeDJaJFYR
ghABBAuamHUKh297oZuC/dBKBA8fvITRG5kSRlbsP6ttJv6GimLv3zQBaYCcsTvq
YvI/ThvvnDPlWkmGNbpUT/Oa3svEUEF0X4Mw2hQ5hjA2YOiNsxurDw9xnHDyJcea
psgamrP6eQHPBHHdsMDP+jE+WB7z/MRiFMIRsxtoQtsTg6YpxWA+osG0q/SSjYO2
eR7I5Q3R7kqziz9HvI90gwAB21lrWwPnZYDbJ/g9/svG4HtAY633vPuPTILkdyu4
bLQ4iCFvbmmPARBfHTNC1/HQTPj9ZCcj1FcEOd+jxwlwYFnmzi5LGTjQR4TFDNzv
grPPNhrax3qOI5rLOxmy/8fOzg+PQqSelPX3N0ZpB2BkiUGf6/X8Em3h4R9zuBix
WNDVGKfpsnEjDG+/k73qDxZZ79TpkDTTBKiTD5zzD8ei9h+dhS7wC0CftPxKMXD1
x1RJukx90p0s/2q2KJwKJrpHFRfidfnb+l0bEca17tngtZFpFZt6ee6JG5tJ121O
PQG3t8hF4PLPn6IpvVmrtXoNIoAhBYGyiAH1oAMaXycJd/co8DIdzTKp47bllPjS
V2xGc6ZssYTJYdUyrAz49bl6+i4dtCPgiA8oyqJoTNDmu76eqzerQPJDfa9EN9eH
0D5fumRoIfrYLGo6WnBvv3dPr53XNc+buhw+ZpDjCDD+F7c8Cz0VVakCgg3rd0dZ
GsGUOo26eA2qO5TILUtJF2AHv0jbJ3ByTa/cilqohPatoUhnAqAKZkkEVUxncJUt
NwQEVxXWURB/j+IGyI/GMAKwClbVYPjHnD27YqUzlecj+9f6U/ooKtzador7MrKx
36RhWn+QBP16x7Fc6jOjKfWh741S55b77iB964qpQ3dk++JtmFkXYCsHlUEy6h3v
+5ENcLyzPbti6m80JwVcx2EATeJTZhQ9+32GvfX2oJdU84xThElOA3vbaIERm5bv
MQG2PjeIROizR3jPZGTjuThRW2mIKMjqUfrHWJt/hHec1NdgVo7v8ivTfAMwNe4o
Dr9oDLjn/FTbP7z3HPCIDEk+bVdUI/PRfgtMZQqmXek3lJCy+yyigyWqla+cnYwR
RYJeU6mBK4xYwQykr5C00SfqFHlHqcrSXesM27wUbmibn5NzTfBclno+H+9HIaZR
RzUKQ327z13LCNuDUPovIpp7SznD25bwTeP1v0XQJKi+xA1qc3cSJw5olvvJsi8b
9j/QzHyTrbqM9v66NtMfY4wHt45xDjrZBmyBXcOKNuVzqvY8cDktRHRPr3v9+WLe
XYNf7Bn+a8LJ+aJDFXytvMfbnWDqw5RnW8u/pqkIwwqLVdwMhgEEyaFFKJYJraPu
5L14GWe56Hw1UPtv+stNaIqljQfpAgVh1P4fWa9anTThB+3GfRFVSTXCREpmcgBs
3OVyIII8EEEk7HmyeQMc3I//PQUga96n83dfikhHSLl2kTF/w1dxhc1x/A7vV87x
WIUMfy0/UaTNnwSMBcC5xls3lLGcuVapgcUL/OEIWfMnDGx5OuKJuwiI7Le3fqv2
VjL9MG8no82EtHlrwnFeUhJX6RGu19rQudcOSGfcuoUHMMgNHs+OO8zW8R4+63Ek
sAomuYZy7JFrl977HmjkZLh/SjHAJ4/ExOT2leS0hK5+E8ltKTNXngFX/o94q9yI
SIVJ14gGxGFNagZV09dFi7MrMQKOdS8rHqp9dYC8cbfNy+KRHvLTieleax+GFZmm
cPip72s6ITwjrrtSxnDlxpryhQYItPDCqiYPP3qpnKQm2HpZPaCeEjGNl2Ub5MTf
IfmnTV+wFAnXaV0JUVoNR8/tb8qvm1mOE0enzso47L9c9/It/tzMMH3eLjn1xu7R
qUJNUenPtxM02fzTuBWUbibp1hurNiqkVTZxxfP7LzR136G2cM5lxKKRb8YVeWmq
BJQuuhVcRGGzg3O6dD+gViQhaHT5e/5B1Yx0NVM413ebrtMpGkY4r8fqS23KaKkP
4XBgN/KZ5WJajo9AFzumnY7utu2M7gDCInN2I1Zhv6B+kMidkmJTaSC9m0zjbm0H
kJibZKw305nm/9aSi723FU99vbHJjmGi5+uzbSuF7sHhWUwx4kJlV/gxMcAcfd3J
NwV8m7nihIlZFck8aShk1ETnFbqFCZJPECvrmDhYHMZRL/nio2vCTvy2fcoadllt
veILJ3gCBvCaD7MHiCxAcH+8SoiZjGY1w/whhNKxfO5V3x6pifYqwaDuSBBxorWe
HJy4yPHqI5QmZ3hp26uqnLiVCVDAwSthrPpzgpICQzjyDwXST6sxYXl1bmXXQMky
lw8zzg9Q7QhONYJiERgfCyO883BRy7zS7NnA0ACz0Vte1O3+vh0xCBmBTgAvq11O
gWcaoqbJderHbLnb4OtD68WkvMW01mNy8FW4LzXwUTBwnI8Ewcx5koo0NRP9AOGX
DMOojkIyD98xpmbhOw9QFhgasC0JeyVq1iVwxTbFyFwanyYhlxn716CqbsYni7FP
ITuXK6NLeuJwpGnBm/lliXAGvKrlXBJsW5AE9n84CZ5ZoTnC8y0n0lp9iepWXiLX
mDHCkZAAYge4Y/SMJ7mVAbC90E/D+xgxKpxtn7rpKEpbnyPpsr2SLF9UAhSwecub
yriX9LExrGDWRKb0zKjEIzQ+pDz0hNbbiM5TmbIufgEZPbRGJI5nlb8L/cMI3/Bm
9ueoDaD6Ko3LpSRwu2rscrOPXHmafcAGUdBSSPCQOfYwsC+eKQRE5qjLLI65XxFQ
bbjpP/N2ELL+2SsDNShLBXpxJWdAfLH4Ka1cVUz/1yY+zcTusZLcqZG7z6AfaKVm
VPkkOGFAbRZVACTmeQG31ph92BQhaGvjKfVul8M9vMnP7ijkjthp0EfHp+ZCS/UI
expcGxLajT8fFN9PTXalpy5gv74wKuFGYers95EQFabRwyaeEQPdHkDxWf33Qi3M
YhCJeJ/miIQJq/YylzrksZchtM5vkPHDZU8xPO7fBrMuMlZyXZ27E3MRwSnICRX3
HXDq0XrMp2cPsdmFQ8WfYPapJm/HFF2HpVphAu9ewIr+HJW7h4cfMRuJ5NVRU4wm
qIHazfpb9n7J+4IaA+s9H/IoHN25H+lwXUPpaP5+mmz9u45JM4EmbfsuMg2e40ZV
o5DngxxrElpIh4wjKpwXW7u0PC41Igb7IkcRYVkmaSodBuijVIquMmYdp5E1ffkE
DWF776UT4RFf2yJ63BcInnjdElRV6j7DrpOiv333aeEOAtj0KJEByQ5Iu7fzmi+8
W7hT0k+JhOZbi7MjX0AlfmP67t1N5EB5L4m5fbTk8LOSsG/21LjGWmJT+/yPcHGR
jCEpUJ+Qm60eJ5bVtkQ43lWg2bv+q4iip5z93Qk/ySiUjAknrcnQi9bUzJT7hkyN
mLnosBjYQJLtD/PnrKDrSpLS4BFoUDjQU6uohN/ia4AXD+XVw07tFwehwpM7xzGZ
lRxTaXTU4isrqmW+MaiOKK+nFwu2+HyFsb/nnVm+EQVaXEcTAsyho8luYUEV800y
xzKlYe17caDUnJh6bsypFy6S0HgwNtKauh6A463z7gogqzT2fg7oFxacPBFdD60A
9Wpp5YH7xC65zkgWnDYXvgNEmTDEwi4mj1jfqvf82N2OYwqpryJE6ZBAScZto00K
wX2JQP4Ca9T7r7PvK1FG7RN6tvkMyWOGMel32vyO9qtpWvk9uZvdpB61w9/QuvyM
YpZMU9YbLE7RxH78CHwQfCCwt8mxiB1kO1IkHPcOC7UE5xdsg/oEeJuQDApmJj6F
LF+hl8BT5bRegphn/dc9b9cYasUdtKHDQtZUE7Np4fW0ouZmsLlUYHDgpEjebF1F
jNNO1qvRDOwcPlE9GlGngcboSGL0rMq+1CX+wMg+eZkYZCApxt5WFALEbQmlISWn
BG9zDzgC9KSmfJTpVQp59yTVCQRk8dxN4/K3b1yDD5YwVAo292T6KhTCk7rpLoMM
EpqrJT7GB5mIQ5tRyJ1W62OS2uvVrG+Oov5PLoWSWYiHcQvz8ddYS2fP6wJLIPLM
Qq9elTWA57ZOW9ont+qAbLrC/MdWHpu3iUyMWTUUBvaPoe3G/B5RC8rrSAVZ9Dvr
HtOl8ckODIub65nRvgh9ZmYyprVDjnKCpHYdlMyavEScb9uxdlPmL2IXZc3D513Z
guAQL5NsliFjxWszFAVjrcK2PE3No01qSs4SPvuoCz7eSOOiUTexFOL6eMhBVzJp
QbxRt7k0bseql3HP/PRne/IUm1x6cPGXLsGfK1Xw7P0ij2XLAQDQmKQDAJOeW4vb
8UlbRBKtFNtwe/s37qkRWExajIsXSZ97zABt0MwODtHn7IY20YRAJPiuo6hTiQY0
/aBAjOyqR8KbuUlHHGvdxt6eg4hu7q0teakvLf6gcUiI+2hiWhNAcvqIVyFJKxO7
lNqeOZ3BtcTyYlYQ1IaTJvuIMwKUuzCe+2s2uWPuHgdqk1+AlsiYMZUHVsz6SoWw
5e8Gevd12NgnXezTa05hXmt141TlTvHmJWm6juJ8C9+wN4bVfoIy50+4IZ1M+uxb
YWG7YXd1/kGGYrPB1zC9cwNIEGv3Q7OHdJ26EeTgLrphzmHcqaRBnSRPiwt6YnIk
EQLaedEo4J3KOkwt1OOyrjl0wHMAh4b6ibcR5k3WGBBoG+p/tvMmacQR3+2Qj1RB
6lYiaIpnqU5RsXJPsMWdL9m0EPUJ5aodW+usPWf3pMD76ZqPhaKVBraWPKfUUX8J
gZ/+9BQZTO05PevSO1mcN9G1+jaN0y0Qy6NLISuhDvPwF6UwvLzKKBuYgNZ2Dzby
agKRzwYVzVA8RXkrfNv77VSU3xAsrmH5tBvDvzBjdtYH7SMOzqGJ+o6DFJoMn3zi
RAf2VXlxIgiHIech2sV2RPt79pPIpTzGse9k8dDbiV1cxwDf53DWby5Emk90Ydr0
bKT2v4Up+L9nx6QLkYX+X/RPPYAJwMmWHOXNyNoYESIiM8KUPBtUIZRJg/FHxJgM
eUzkPenfcoSv2xUC6RtYReLx7zghPXraB0hZa+lAcCLEEntbNwrJgM3NXEl7qyLt
dWcMeL+Lf/ZOiMeTT9MWzD/8Hci4KNCnB03uIrHkn3O2g5qUw5gjMcw7EcghuzOn
UAM8zNYRCwwrMdt2aLjff8cdoivR+kbxjIiPAT65yWsOSlCQ1JxEMxOMDuwTUjBr
aLSphtG9WkvtpumAmYKNdiBbCOyfNBSsOSya+eYAH2TdYGye6JraEdwPbaBY82LM
IZZpu9fK+5Jb8jipXulV5rh3PFvCSKuman6ueC0JDicVYa4t6mcCHDPIVT3gO1rq
k8Pyhxzbc+LOf5TtbNC5lQPGrWTQvVgOmtN64BAwVwjoGv1IA4nPGwbQfAvlxrF0
TDYxUBd/QhNX/EDzoNNERHje6rNiJaOO3lAREATilz+jm9h3FxrwIQH7YAcrdITY
PlZnm60XRaxaED0ajrFDGJNckVB8pmDE9wttmzA1mCoQmpRJ/5T7UcRNfCQMZRV1
kpqgwVUuKedvWWAvihWBNwQtze0w944m1RVlYUvfSwRTZdlgoHgBeGjkymFwfbvK
v5u53JKPoxrObH06ihefSLjjkbMCAjIpzc9lCVHWsis2akOBycdW3F8OVRgmmouK
Z7txd/sO3ZZqEEMFH61G0kmrErwFwAZYNYI5GjL+xEZGm14LVAk/DiCL9WXvRm4H
B46wy1Y3L30S/gdg05N66gaBmCU5z1cuiw2GYEmsogDGnn/dT6Ht3hgUHeMWc4c5
gyeUNd2PrDReFuSAyK+ff31Q23MKPutVNTvLPmbtopXGDApqnFAOGqF/LyutIFqT
EP+i//a5bYOxED7tS+bs79IZRJCnG7H7iTOehziMhEh6wKyMrhrLY0fpbjgXPsB1
PSDL1+zTs5uuMy3NhAoSX3keRE6tv6EVw2youhMi+RDICr5lNtACEokPVsTtlVt+
LIopbbjm9Lcui0E4nTueGOEeQEYKH/dwN6vMYX/w1P6UFGEYDw0/n3Hfdfo1YxHR
qNoIDe3Tg3sjTzZFhGmHKgG/unXuxIVgRINV8KvZ0TLBMn+xEf27FA6Y74KPtko3
JJAEFuWiRNfh3Bp7gDu5j+lxZ0NIWTxL81TbT+zKoQrWQvlUu5xkuPOlkw9N40ia
wM03dChhefOgt2Zqa5zkvXRjkpeIgXIKM+d4tAqiDQKI/hOpDj44sYhdZEiaygI1
jrXNGCU8WxTVKTGpalRoby8CUupVqFMFyggjeVyyK1BmuilMyGDUA846WLWrInML
CW46PpYbpAKZzij+FULg9T2YLRGfNge17++15qcawwO9JQVpb5d7ptMrsOz8x+cA
KyDjI9SJ98GeCkIxU6fr4p3knvdA6jqY3XfH2PnSL8ty4pbkFW5xGPlNDh3r7pNj
4AYTJFDhKCY/+myWT5Y30KEsRmUQz4KXT8AZuBVOIQHecSl2cchxInF4wxEjw2o+
Ae3Qmxofvr9+GukdOsZvB9OdH/slZXLh6je75MR22bnhcpIip239ZvQES1+iN+jP
C6d8cwY+Utq8duN32daOeALP1aIZ7HsXqbhJzOif/NbW1CIwL7jTbPzRbhFoWC1P
Dmm9jdM0h8PPnLYRwwV3MPxxflGUUiRebZy7tGyhGC3CEO/JpVId+jsLMto6J7N+
5MSRs7akG1y8aLdWlRgBRbGSw/Bc8SpqOE+UG8//ZJjZ8FheU1SQ1ZEgt0O8CTlq
80FR3qUvxI8GDDfrnyV2VdCT11xB19z8/0Iz1u7FOUXUHF2VcBTQRvD+JwyEqyVb
HHlNNgnaZrHLAIeuoKXMQovYwLfdt+z3zX2c0yX9ENjsJXmYFvVvHsJRjTQRgQtg
4iqcE4t5GDr8LiwWF3lxHG6B8tEW6/UFD4YyXJ+/trNI5c/eVeFDJoeUL73vUGVI
j7JgGR7oc1nyuVjTw+Vlg92onDxe5wuVPDRjIkuomgPSDoWlM0WdH69KIKKBYYO2
BL1l0OaOhQ65Ar/TAVYxatlSNMOy9MhLQ1JgS6sHidxn02eFVKu8I6OJjXMS8ppB
63BaLaM+zKtobzxy7Jsqnq8mVUi93Wug53944uHUfo+prtlu8l7OW+SyMRtjE4kt
FMEbFNij0giJDfDg8OdwiOpQj5cF6pczZ1zhJF/G++UB7p0fuBsmHxM0r5mvjhNe
/V5VL+5MEvLd82ZOcg2+TZY5xqgIaoSn2Oz2hGkn+xaUwNXHd5uGA8G9o3N5Ea6T
rvghgsmM1D+6EOGRB5TJ4FolZYGD25LvYcnlZJJKhXTDZPf72d9bwI86HX8+Vzun
6rIyJ2qs86aZeT0m5xQffrHg7zpxX20ZuJBzehI9Xr6dlLnufXh933pZnHTpvEJG
qsIyfG/JZXIr3+mHT6NyCO3N54LzREaSeBqA4bFPuutMYmrAozEcT76T8AX1Xft/
h2rQn6nHKnoeeS38vSydTO9RcAR7iB6Q1I7a/tjATWIxZh63nKYl3sYF/dlneaRj
N9V6TJxNZ3ha0y7QXs0vtBrAyHR0PkJmwNG6Sv/K4mlp9sFw+jkL3RazJqda8IKb
kSeSf4vQ1bf1QHrAikZfZ7vzTOgixboGOROr27WhVk4mQ+GJXwelYPb1Ba/yRhgX
BYiRkShjMC4IOIGRQoOiRRx3dLwC1akW7LnupxsQPLwkkaCayi/oAkxMUGRsFxaS
ZnJGGPdA4DQlRdCcbdyEi94weMoKdTS4/2+xTMRMJ1CU+xXGm8FBi3BVayq5dlxR
FUEejjnQCiTabFUOXnKTsy/JxXU709FArSgHW0SGYhWYK2VVrQ9czOBvsPmzGEPM
aA9SnNR5+DETO16jJyrxQnhrfGeS2X92oVSzdlZoIYfvCsZg7rj5Z8pER81GODa1
FbTWebUPrEpxyfMxr0cEJ/wkeaPRmN3QpyleoqtcgDn2OqyhdIRgqDY6650QSjOx
6bw0eTWczut6R14UpmPpCHKk22ru5A43VfZPoN2pDpcuEj9gzzFdu8NIQ+6ZfBku
mDuYhA4GdZLASh6M4w0BGAPxXfvybaCTM+aAwRJv6qPm6XW4v4e/HYyi6MSjMn9D
hTb8Ueox60LoCGm1BqrPPipeCmnBJ4X4qI1mTp1gRoEWHFuhoJAea1Oo8b2BaaKW
s2qNWodk+jacIxpUza0eohO2bFqyX09oh20IuMkVScUgI3IchLCCLjlRIteA3CkE
SKO6G4y9HrTfrrU2uzI6QHrN1/6gdt0zmERZszjJ4rBm8eg0yWP+UQsHWY4ynEEm
qNMYIeKjOtcJ9ZioAo7PmE0lbSf4AxCm8Q0EBMxZb+WncnJd3d10zuWt64xOtBdb
7w95dfjPaKb+zKHEIrnWGlzmvwXzbIe4Tk5ZsvsUySuxINYkb0DAGsAGsMeSwzHB
JmnMTdLADg4fWTJP9WbRM/ueOMIn0uz0dN1Zn3gNdIu1sfVwEFKOeSPA4hTmm7Nx
a9dfUF/+9Z3bWT0/27c3foM0ps30bpqf7z1aSJwha1SDdGa2K+nLkEEkWujdYXR5
POKY+/EnMPdSj+rYeps0ie4Z6KREz5eFEkYO9NHPJ/C0wAvpVLOVugOlB95EBeIW
9JB5kiq8mrA2l2a+qiyxpbkK09U/LBese85aslTyHnTm082FKBja08t0QnFWImHs
fJQ9Wng2SOD6u/P/dpt/eqAcPgglyKHH2eXL3KGofIZkLzV+L9ONMY6XbeuyrYuk
sW5j4J6wgGxVHPz0zIBiBjGBbkZEYGG9qV2HFTVziwpr730VZCVSQkf8x/s2tbJI
H7YELccYEYo0o+l1KYvEXgV2yNnCRu7kAnJQ7xtZu6GkNZCAcIzpscsGFK6lA9Wj
ftFQKbWd/bXSiCrWIMN7Wrt/wBJkg+qLOk77hm1c0f6vFrQDFPdoVgJQ7ComNu7Y
aKrew1yh5LSKbmw8pam25CanjHgm7CVNJiyT2gXiKrmYh9r+44YO65PfIGj3Exss
Xq2kJTlQeI5IM+l2Cd5bsXV0zJPZIKLIHjgLUXj76xgziTwO4ExWFT4Of1bFuRB1
2u/Uv6NjMhNMFUSI+D95GnzH/HtKWFKMr4uIkyUoldp6IlfZO/+P0g8z+1Z08z9v
CdQxx18JjvalGF4JUl9wFoOhkYEiPasql15b543KyWHfbzebO+lSKAhvddmcl7XM
jh4EdXjeTJ7yW0aRbpm4L/Tbks9hawKFwJnid6ofey6RVwSEIyQ7EPrm4sbBIvpe
Cos2VQX5Eqf7uOazeMXalMFaOJTC/WWO6JP3JL/dKw2UsB7W1f2/qXhqrpuJXC6x
UtLKwEYT3JASXsW71m1RfTsLP6e7EzhaMAzzL4VsWAuvU0ksCShPaudEZAyHJzex
EYhwSCEbk7YQwGWXjz1ooCiM6xQAnNheFw5liVXOwxbe5JFA2Aj0LBfKasRdMg6O
lKxwlG093oT72zwW+Lss3r0kitK8nK3BuqGLQP1uormHe8z8NKbJnwJKd/HWSVng
ZAGginqjG1CV2Lf7mHGZsbFTCiA72EqQGQR6KUyOfTtrYroUmIu6Rh3mii2Pfdwk
jKY3vYsScbbBZkzrpfbfi1HAShHVciKP7QO1oP8UswPaFlkdlQovhtZgGGH17yFt
+i1/oJl2PGGdN9TCYw3hV5ctfAlw+9gPgHvwNuwxZeP1Qq33fH05QiXwLEW7k3MP
jva+bHxWntU/j2SM4dYdVjerPfe0g7L4vxwmMKqFy4LHPSumcfA5BOhMI8gg09tI
K+9h1aQaaDYE0tf/oMy0lTy3Q2MdMAqpl0JU6cmCt5DgvAjHrNfDgGv6s1kHxlED
gBbTDu1Jv2C9iTUEtdQvwKQM5S/HcMRlikYxriYVlxzAikn0i3Wu3kxtfg8k1bgf
wC2KJsS8x2ViThX+g3Y32+4UL1ulRwc9S3onpe0G/T2We5Y6v12dOsxYazuWHeXk
ENJ4mqR5/NMruNBJx7Y0LsbELwNazsZzfEC6sRuWk+pwfI0mBX9oMFMwpZXWNfNV
y22riPR2BCLMLaUkWZwsCoM3HYp0cT+amcvEDwauNQlCrU8R3IrLfC9zA/iYob33
Fvc1upWbny5h2ImoPMcG6ojrrSUyKJTdDFp+DJKrWqWyT3nhYpl2EJpxVDjFJ7nG
Pi5pWYRCRl2hXhIQM6AJS3z2JvXtlbx8qHQEgOCk6UWoNN7AXc5X5xvjmRBkPbsY
v8lSvD0PJMsm48lp8BC7HkEf1ZvbhFgSq/Gl9iu8W+PNktzw3DnvV4/cvCDbZoR6
+YVKpai/hNO2OghS40PVy9IB6DMBy0h8iniwckweDF0qBJMMO6K5vUbQwmerfdmm
WmEQaw0ARfJsPueMNUWjjEvOI7M+fDiviyHwQzbG7vWWt2Lfqso41Yj130oDAhPY
gAMjofDZsxNc3ffhKRCDUMddoXCx4IGVFUHdfd/1yxrqY5xX7vQ6nZuqd6jB2Xc0
/zPPERrR79vgzteB1UuwjQZzeNlqzRO31BKjnEOjRpDs4Efw2xHEG+V7eoA1R9rX
qkp/qOo0YaVIs5gtXGDGa7EvMDSG4Ut0OaNkpxWmd6++CO3eWWcTx6EnhtS9yXgv
xs100YGHFafUNSRlR1h18FnGH30rsmX+PZLGpmjzqcj59FYbQxl0SZTiUZ6WhQBA
q/DUeAQB2N6VmtTGx5vULrZkzJwr/Dp3ZbOqqviU/uf8HAvl6wP/qbNsl6Aa7mJt
zsyKLywgBI32rdJZ87p17+Da6/n94G54vj363DHwF9Tyu3iCQh2YXkHKCYfSsSTX
nHpWpiZGkBBg8fMfzfuhG5eM8zU68+Ff9KWtItRL6Mpz2HJjcDERehvDg9hb9j3E
8BbKZvCC2dnGLwTBxzvP9UaurSMXNzT8YVcwmI/we46mDdXZC+U6IdXri4VLI8Mh
BJN/ZQeUIS+OtlFoeGgyYTh/zCmQ+qeXX8VKzRX7I5NgUQdj4uKe7r0dMrweqAKp
Jxb5RP086xiJkGJEScNDdRlAYTFu7CSCyorISBJkxr4h+RJkBiwIwiTv8tIbZZmQ
jexuznCsYyGmtdWijzi2yBIyM6kCVxhZST9ENjOx/m/AHMgD4QHXAbscRurqfl3G
GGTvNsxBRsUhUuJhNqNqP7b5WIcywQUCuPzYxKfeugBmyX/KcIOX5DVUXTl8Cl5O
x0FfTPLyZr108AMRcdSGV507oj4E1QzLw3sdyl3Hfn30oGXfyEadN4T0pCi8/RIJ
8IpHlPHscnBD8WPvukCTya7MZWDLjTU/DvLHMGVVUxWiLRYjsRl/1EukLM5CxDBa
3DKrIJ7JkZcDKhScqMD7lvDrIvxsuG+gfQFY2Y3fuuBERliQ57W6J361Nf/Bw/14
oEreZeJUGECaLsI8+3dkt9x7txf3UTK0qZ74OFHXYDp4+p4lmC/XtbkzBdQ3kpYp
IVLFUQ2KmRsEE6KRJ1Z2Kl+WXhjXRAh7AiKJlEHOBGjJSduhOwlt2AjZt37fAc4y
HtEnguewQVDOGzur24Z4xSHSpj9kkhPDEOqN78HMTr9A0BC5EIWvkhuhfD6nwaJX
s2gud636f/kAVEHpSxdIZ/l0VJeGXEkDPDqd4D+7/48jC87OmU+TZ/2YDwVpIatL
mLMQZZU/MUIHPTzmslY083y9pImxw731VSw3MJTAO4ErU69ZMWS86Lru/deUjXuw
BRQQrymnntft+3ytlmUeaA41hzwX3/syexLRCG+I6/uv7N8PG2crelgHtzQ31bCa
+yGIQOBktKaNc8qoBo4aMRlHS5NKavKIVvubMG+/ZeLDWKM9s5yNPzEIQ8X9hspw
EhEfh8GBBCEn+tZliISjG2ahHAx92yBOZ02tuDI7XAZWh8zmQpzp3Yh5+l3bwsfV
rzhdRqpe1x7LhjWCOOLbqV5RvfwBhxzpQ1bDRg1STXNskA/z27OtKcBSgJkY5uWt
PRv5LtoGVznkezEMQkI4XMDNnqMhs/QlTnfjkRV9J9D5Hd4M64EaAvleD2ba+Sua
bz/mnWSGoEAG2pfcNWvPpAdtDSLCH9/QHJw07FopMZVtyJvk6W1PPIMl8/0MoTn8
4hYkeVakBeokbZYS/fuSBQa0NiZnH1gAovNsDWi0VwNz+Xv4d9G15+cICf/JKcAX
9kSMq6qOeBBpOzgFLM8AMUx61dpL3WG9eFtjnGahdaVmxqBRGZTAOBkY5X1cbYYr
Qs+wDzBlOLh91IZAFAgSbGp3dSOA7u8Bhv+l0PJ+6qtMz1ooQ2TNcAChjcO9QMnK
xcOEX9EJ30i1/tEtDFkyJKFCl+AXjQW83YjJblqBlgsiJPM/Gd65Q9WrmQTjXfM7
WpomBL+HoEyPda/TpX1pCPGWa2cdKHKIzN2dU8vzDn6kXGRouyXfR5Oc1a53gHOV
5nGK4qEuX9eujz9hguG2t6Sm5TO1ZTLwME+fT+vhtgI/LfpSAvObZi+gLS5XYkxa
nlXMFJVgBskGHTIB0PrGQM7vW4vlqVy7SfQNrES7x9i6+XiOUZ+FDf2mteWq6jK4
1fWM0VZqUF171AVZ51KSLQ0MgzeRB7W5eLBt04eb63NctdDzicCuwfgx6umVpxYq
OvuacsniU71Uk5o/w0MF47geAzI9uajV9lbPbez5vINYHjP8Ro5VUe/vuqwcQuyx
DNIr6y3kDvDxl2bPer+HerJFjGpowmSp7nv0yMz9EfATvIQnz+/M9F7duaX8JdLz
BbuVrx+YuD8W4lczZS9JulxmldvRbE4cBWUpRGcFaZLy4GF0SUeuZugsRw7j4FW2
b3927wJER3mywvrJiwSqjjtBf37billiZmsWj0iRHFnqTgSlDHTiY/HufU3RnRfr
hgKBfjRWN7koUumyN9A2flVeRz5PtjrwNw0qikiJ2FdlNalCM//p8nvDaT4+L56+
JYe4iJGuyK/oztM3OwvMnouEsXHlU0a/DDbThrvydiQDoHezZGOWznhl5R2HbzGb
xpy0DqJ8Rhuxq0FJQdRow00TSoZOyr1u7r7LIplIAk5mUxq9BqOYsTR9fjezbeuV
P95ZQWfjn3kb0fvwRAnjrwfSpZEXVmvy6gR9cLKW+ilWvm0Qu7M0W5c/c3yMj3sg
vxnmMy8gSLOvcvqvJADQahHWDgJCEyUf/ZmhSuoA04UDOgsAjhnJStp43Xq8RZ2p
VqIUB5TZb64/cltzqlVB8wQkF5uoN3aoTpU2/U9enfPmwWjjyqQfKsjR8jFtzael
3E3Y25vk3ccGSvkAU868+aTatOUWnvFw32wadOGqK+UGJBBTbbr4dG1qT70IeGtZ
i38PgtHN1Q8G7NiCxcXWjm4HvhtVkmHANoZG/PsgU0ZUzqIVAA5e8HpqTWsfoQR7
KIJ44hrVhOHZCW+ZTWr+/YVDAb12bPiQs0KxQGvAh0KxVSUw1bxigdK2nGMEFsVj
u84oXe60+LZ2C+OwMy6LBV33ibGufnW22t/eQ3bCKd/28OectEHQ26bsQYbyViB7
8bML+NywqI3jvJNHHa26RCuUDwcXVMUUwwI3jfuqbLDKEJxxopBV1+taIr23K/6N
rmRzoqTQyFqH7LbWoSfrlBnNlI4QuOUOqd2N4wcnBA9WYMq8nvTxRPgUH+Jrq0v0
TrQ+4jmYJUsscuiqJH8X91EKdHExpH/aXZhzTuxXhXIHFa0mmNXeFMpl/AsiLTjS
EXdMN6CB41qdwRr9+wb+FpfpjkAGsIDtKISS60sm3FhC34vcxafDfua5hL29dbJq
HhiIvbuC0tRIQVpzSH3incVjoFSWWT5jVHVxcdYoY9JMZpDJ/94ZwGA4gMZCZVck
0T7qpMIHFBtYb8kG3SM4M7KY6evluYX4bGgvGJPZVTENi5uUj75ndbp+vrbkzqt4
kinOrCQoW3WI+1pctgQK+TDFv8RkUHaiBHnkcxjAaTtCb/gW+cZlBGW26uHwkoZa
sy65wKVwegVs208f/ZH5FKv2q6mNAqPLjkVWVy1dRndMi5eJK4vIFcahbkuGBl1C
JCXSugfgNxJMri0+cT8JmDKU/Qr3yAKwJj2oI7YpqcCMSm+30WklXPKPzEqBRV6b
qXVK1mxFMCzd0u/6t2sVtjR2OlFdUXVRwEcQAXjM+RpWT8BjWCAgd1eJUsSEhYHU
F5erYByrjFdkNUgxCljZU5Cj05jJE3nF+ZR9tB6L6b/KU31+qDwzCupreqWFkJKn
CHTqKxuuMOqoJ0TMw4nV433fFsm6SAqCXylw02eXrZEuEoqHFiy16PbHHE8Ju4UE
kPtdeDgralo1LwtNaES1E36xusE34GKcKM4kUUx7VJJgOV8KgFgbCcQyTZWwBBve
l1D7m9BejwpIGnCV0JN+WeupdXJDXtunIsV/b6zpsmjFu89ojzaIAAyLw0IGicC6
NsHs3hN0ESKs0STw+FtKEmkIFuX+BFUMGveqdctTMJ2/WNVTe+o9mour45c+v4n8
6WGQ9ZJbZcH9Bm3yERoH4FwKnvJyaHeebttf0o9VCxWBpaTlQcrUp02D93m1RS+M
NuAnk8oXs1aoQf+nbhbTmX2h1pgtDJ37qk49k1SlfIZe3MZYSxhR1Ox8ZdR5ch0W
awjCEXLoRO/ItlKVTlgmg/ZzUHChdNMNlSYrSZ+Eh24IkXru//p2xrm3SlNrFoQe
TJQGhnzFaqAj6/fSzwUeAYgSxJvao8j9x0pWXgzMkCVrXWg1zNB8efp6Onh7820F
0uURTLI5J6DvW5XwtKFq2Crp9MLSSBGaDJt4NPMqX2hUTIRgpLbntFPZ/TH8564H
amv0FvI3vzKbs5tfwySH4/ZcDUrU/6QZBwjIXWXa6gtw7zCHjCf2g0OPqWT9wAFX
aqVDLYKGU1JPbD4eWPh/lhqiicw/uBXJuL6xeMP+isQaII0skpfNLPDEleqTPeeb
4LtxECEL0DhUG56OgGkrYHcfzX+B0IoC7/U1dWxiglsQRfsiCLD9/hz/1QT1UZ0I
xfW+Jo1GzhFV7r0MykZfhn/+tyryYveRU3Q/FRnTMkGdd8Vy3DoEfHwslp1rrEqH
tVR0RdjTM4s9jt/gJO1jbfG9QKkjMcfS6YqOP7HhnUD6w+jk/rnNsbQEaMVcFIKP
iZ58skeuGEZymzomh5iKfgGJm3x/Y1DIWJAoBIG84rmvTGXWvF0vjrBCMwYMM605
4jIvtccLWQM3y8N6eUm2ilS50LpALq0kG9emAADDkcg6P7hL7V/FHzjOnJzx6K1q
ab2t1BtbidIbvVd3TAyPixuVgF1ESlvBOQ/o25qFmLwrB+buulsL1Q+LLkuLrySy
9mg8nLFYPLxD9slIH0tY62LeNw2l1aLWPcD1Fs3Lq+0MGK4K3YtvftZF80tqPb6u
W/XCfaMOrROmnK60OwePZvWsDCE3S1XUgjszJ4nZZIlBKNRb4FRrlghLRcWrtdu9
0xhcFjRn5Awv2XRcnQtbV4OrMEbzjUmBAQjforKMc+NnIc0seY8QPrEz0bPdclcY
2bJTIRTMCCNmGUG0xP7bwNxXX/KwX5Y3RUzOXUjGNTDpbnsPsvK9vOwQ3X4JcAE1
vDwJrSyVSqzonfPLDcSLeiQN6y9BXhyliYIX815gnnOQgI/kuEGyHPVjZxoNTaP3
XE9F3LzmPvIh43DCEUEUfU2rY6WANTLNe81XuYvErXgAbf7adOTuN3c+c8SkNhAI
CKuFw3J//cdgwCCV1O/KyXIeXAChWwSxsyBXStTVJL4BYLhc0e18Cl6T22cT4ZFe
K9qMbyN60KXibbWqp3uKkh817ckj265Y84iZyJqVB9xZMJiFZLDM+U2YUejKmoBq
iKkfvWndtr+RBix6AojZ6SVOLLsFka8oNm9MiuHXBxMQ+0Xz6sJferf+qmJ0Wvf9
W+EA+/B5rO+HLzqyRW+Vv/sDZCQHP8/qwOh4+gU/P43EfC0CWiRXwoZmxVww3a7i
6i+bxBi7eKl8fLMmUoIEcMNh+WJZN6bVTgXd6nnVmyfsyWCJ8KxhhM/tX1XRF2Gy
bEGXua9ErC6JGypDAQAGP9xRSjHvlZ6NG46YT9T+CPSYZeZT2tohXPMWBbB9lhC6
doUQYhUzMcRPyqQN672GIe4q6bYYgkFcUC8DzVA+KzdBqR8+mIWOHV7BGsa+ZhBb
nztwfmQtk98HK6T1bUts6ez5ulsTvOhZIUfL0r2Cr2djW+Yhv5T+j6qEZpcJ2k0i
ChW4VxA6H+ucr5D66wleN3IHQTUz+NiAUKkpm0RjEI2CoPySEf76fuMFDVp+MOdn
WukJDKLVOxjRImbZ3RqDKCBBCSEJ3Puerd8V3hd/1JaNmZ6v/kQ/mv8BeamhKQvI
YkPcnBqDi64+HDAIoUytXYYPuL7WR5k8EMRo4D1RTtjGyZOWknVPq1NtgpXdLWbY
c5nlajxcpua/8Fap6d6L6hFtxZjNvlxFZcW+Ti67lhRhVUVWTr4yIj0DlTeV45Hg
XdIBgUFDpkYiIFThw0mZl63NculWV+EXmGZMTvnAF09U7vykkptUalUzF2g1U9Qn
IY7yWwrsMmKZcWdOW33GdD26f0w+/fneM0H3N8jqfeWZbEitxSCDxjR48v0cRJTJ
zSF4FaQ8xkHvOZZgd1ys2wyyKGsGJ1BxeaYzpuo5qAfmzFgS+DOrnhtIdPRcS/Kh
G/pOLWg4QQ/q4p/obiy9yXsR0RpkXWmTLwh+D+nTpt7iUzQYgGOyz+O5YcUEIVba
nNVbd1yl5n+dW1YWspfoPYubfmkvZ3wvamzpbtlNYLpMckG70x4wo0lc0+HSs7rc
ZeFaWorEI+etm9Ayx2MvBx3NvBZ52zuIjKCrOsFAr341+nRcJ3W1xl3kXngEwYMl
1TFB8PmXWbE6jhhriUc54I4SxPbzYoSEIhFKPk4qEYr8cl4W0wAuHTSky14SWh8X
+Ye1gPVwYTMWl7ZQVx+dj1tYB1j4Ur9igv0dOdmkvXTKffX3Fni0PQAnJsK2aAA4
mjBmjCSk3lq8C2jXJK/7/saHQx8FE3fQFatZFupymeS/Ll2UDf+yJ/y3R4XqTBad
YHGkmS4XqAQth9FXil0BBAqC9TqnKdrwLFTiCfXFjnl6ZOo22OQidGgidF+S/8/A
Gtc+HC1FKneN2LDXmMxPOA6dezQ/vevp/UV40LfYwv6MOMz7blfFw3kIBy0Eg4b9
Sb9l2rEQkGMvpuR823y/nA4q44gni/i+R9DKZwK9qxHMkMLrzx0yqkXebpAq7Yoa
lsSEcrGve8GQrcxKhiP7uAI4DcgFeiVrVoKdtTICiOosiIAWHbP0kI75pVx7TYRI
z5oUY43tvJ6vQtJHQBD/q2Fb+NMhR/GkX7/Qlx+752Qo4mh2fB3fB/hhIMFit8Mi
BYy/rdSNfzZkAO/iwXd3+h1I59R4kFI8ylbnYLKiTxjPrOo76nWq+BqwbfXSV0kI
Guzp/Gk6PayJnjox5YdqI+vEKUGzeBpBWKL5BxlKf0rVZE3fNXhDHI71/OiDjv8e
VxdbXXKUHMqEFHIzVEcO0c/WRRIN8hBy6sw7y4Paq+RnrKWzRmrAbIMrYak83k7n
UOPLe70jSKbPCeSduE1a4RWmQpfl5umlNPgY6V7qK9N4kwNL+3+oC7/aC/7dif9n
6kjEf/fH1ioKfNkZPQDdYFmAxKMofLZtvEeyr1FZAz/hac0VlrbaDtXPjyZZRQRs
XJ/EidrecwT/YJHafWi0/p38hBdgKphkVHUvlBq6DG+v3FvEYggN9VqcfV7Jslsx
9WbLlGI8KUPFkP1c/ql03U//iSnzFDPhJQ2o2A2tX7ESEMrd9HBgCWWFj2KzA9ic
SkacZte8O0n/kBl2abLLuDi6QFIuwZ/6lck73sDddFnA+NJHfa8GxzKY2SE1qeNd
3T0VtIgnQpgvGUTcsVO3BlZl4WzL2WttjD05Jcj6QI7cOzZZIXFgWFjE7wu8KpLK
FEp28iVJFBqt2tJF32xBFQ+C9b78D1kz9bzz5BcpuFhHiDE2vi66Wtp2Yjjq3cqH
b9qXLyu3MTomSFQYMpWVzSLja7Jsh6b5ZH7gTKucljsg7KCGkJJE+hNFsAS3m5Dm
HuGUWMJu7nJ2TyYsSN3eOJdVDqPxzEdbG/RClrwrNJ7FBoCM7ZXXZ7t0vXdDnQXm
6hUsuSD9lLKNcwPOo5dmcybfSOn4pumAjndSxSHp+4QwXJWOj5qsPOPz70XhXz6l
keSvG/pATqBlausqJQi477rS+M7Sy8557zGPj/W0lgI8s9jCxdrYHb8RlDSmZZsD
fmmk00OYjlsV3V+FIWQnMI1MerDa2Pc2ig4/fAK51hikzN/eea11ijapzkfn5ymi
6fP1YX/t80npgQ5iEM1p1+xfdiYAi6smXrTvT5wrF3k3O3KZFyKNQp5ivXBII6vH
Oe69+5LPfGavijHizrqMxFj925deKMF6dZLm8T6a6PNNzJM+U98jGTnnL8LBwgkr
QxsQkm9Yv5vIqcye5DeaA312D+D58RVg5i65p9Rt/hOEisuDx+BdqUEQVdhyTWWD
c1sHMk23p324dDQdUgrq0+MQ0s0Xipom08JiHM02ducR0dW8ftIms8UtT5hew0pc
n3A/tZClY51+BZMedFlWUbSjvDgo89qpE1MbNqnCFLcHPi5Xf28fr+JQmIh7+jSW
yJLXIxoDixoLsSuAZIpjXd/6W+IB9W8hPyStKpOdq3mwFZzvc2ULiu4phxHspU1T
Xo/5+e5l/im3lwh8H4aqCDS7/WTnWBWFeDp1yEGB85JOt5gco8HNUumYQ96GlMq1
InxDSHmZMO0k4Ef1Xc7L5m8EawpL07pqpZVqzBpucpQ8UkFeQHw6ZL3nO1MG7cFt
rOnPu6TRyjTzzlvyFFUpIkUKJZk61xRWiKUONO5xQlq0U6bN0seeTdLoNikM1NSF
yZA27BRKDLZLQFYL5Sc7lgtek6c6+zNa3M4nC088rC9gsqgfoVtI3q+KmdAGnd+y
ewArZdV4PZtyXmbNnRdf/GlejAGTANxOPueUMobOtIRbjrpcxSZqzWA/hDbt1I95
dmQff/w33KudT12Wo3qCdIJaoMjwgbsTwXOmxmzRx/lTeO+Oeygz7hKyyDDKvfu/
8ceXHlJhLpYwm/+MHOOAj+FR+iFhFv03nMs8wbgAEgu1u5vjxI/J7Z+nFtLVic6k
xYM5eiCSOYEtKQxQKoZgRmql0MHAxedfvnHObNKMbaT2dnoa4eT0X/CIGBSrl8il
r3r1HZyJ1i3kla9U9ES2vHyLfW8LS/RR3TfPQE75+a7i5pDMFFR1MBdseJEd7UVB
4Q/LoSiOSWJzD4DJTYDLYG0HIvZBU8JOmj2SbitXkPO+BDBgvZSXRFSXK16cDdrF
oFIxtEq74sJ1i9K16ge0mbwv8VASVt392zPa+gdIDoYLB7RBOkfmuz0y9umfuJFQ
eA/xdMtADfRvhc7NniChbrW/LRxux0PGNqJrXMMFzQPZMxFET4ML9bR4kxCUbrbE
icQnF7ZnnygJnd4ImWd0Vu/v8l+g/EMkr/5LEMY9V3ZxQ/TvbWKLWRaaVF0cy+Fh
6LZuXjPzfAlczE4SEsK1ewAzB3mek+R3zfI4gQGS+imthf9s3ZwtbFWBtKHw1PKY
tuizO4/5aIpTPE9cn3HX53Q3HhGlLep5tKm+XTV1MGQngxKXPMmfSCjwopnOpNJA
Olq2nesyJXr1ej8vk4JcB5ykWyqO2xr4M0YjxLgI6/uaziixGxblToifd12i2KD0
XchzHd7JraSSd8x2u8mWXOh1sCDXXaO8bMGUlAC2M5MnRXTSgMPwhheowPtyVm4U
pJkg31/8g7vqD657XYv2nhbzeA4chrNOuc9u6qqnJYzuDUp3Z8tlVYlHdsASL8uY
OQdXd9FjDTsAslV2IBltV51nZXuB5fZPhVucmd0DL5lQ04sKKL6UlRaN9N2XZDaY
23KDspIvtqNerpNsJLfdXozJTz5hbIzorBlDh++O9jwv79BzQrF65P1taiybgxlu
jnPfONW/M5aRHW6ahNb6R3f3uIAG/IIdm2PWDhPTs4o2bEI13BEI+tPz+gcGKXgq
6C3U3yNB/c10fZGBX3xKWDllCSc2p7FmJxDVIHzQ+OQbxwaAen9Sd5eyPSspMdQe
wF0R6CGLBjBFBffTWnfyl2mVzV0/1TY4CNS07uLoqeMHTdQLnUOjG/SABlxWA2FC
4b/oq6rlUJA0FzloRMHBi+5hhV6KpbJAf+HmO0t9RnJ2gQmV5p8k5kbCbEq/qkJS
M6MjSuyODUBFd9Zq8Ul5tWYDZ/bvoZmSb28SnZVN8U2N/RZoLS+3DrQM4/cKm3K1
S0iyersimTLLwR+sdnRH2P6cpEe7SIsyQvWcEm/fhjkFtb5cNs4BWKDTHvol1OwK
xmv3xfaANfYdHiy+BMKlzuPJedKNt+AGkUYYMNgl6S5BA36Ue4J0vXpDVFubgfO1
TeP8zz8Crn8IVKZSIHKGRnM4RvBI6U9w1+D3dwjE0h7h6fNrxrpHCjnDoE75pytt
Yzo+MTf3T5ExChO4PShorzChXzqqjGsSobbJH1MD6bDQcQdWvzwFRhG3rfltodmv
wgOwj7nZzrg+KkO9pMVG4kYEOAXSxV66vvuzbwTtLJviVWf6OWn1wQcngs5s12ev
GLyQnz2U290hHR6pUJV3TEmUdwIwszQJGNeQFMg/a4yKpFe/6YmBZyAKERB3rHib
z/4jpKVkmEOnCoLnwd8A1yWkX1EkHDY7oAbiaQ99e6Zsa+sdLUQWXbZ2/7JuFLjL
YcQRyD1W5ATm6gQb2Q+fQcsY4EGTqTFlHkUpunNrKlINOpBf54XbNx++gER8HUFl
VVX20l9CKC8va8+xyxliC/9L/0pcXcsLi9GQ1CYfiTwYZdwHF5hEvQyW0he2bZvb
gyZIVHHMR7wDQRMdJFhr9B7y0zwh1AOY1FId0hPr/u5qtDq5R/QjaWdwtXhVa8i1
i5yKw61Ypef7YSaZ8wZkAzZQksreQfJjvpvfOGLC8DOYbW+eaap5iqSe7uvHjlDm
likUTUnz3HKZzx3teTu+LQb9bgNOTkoHRJoyWdr+8hi2dT7wf2JduYIxCtBbR6aC
JynEy/56Xi9J1AE4Bu0N1k3FgquYOYhwU4WpPPHs2zP8KlxHvdiWURS7dQ/rIWZA
ixjxDBgjQ3JRzOCZclTce5EqyN272ENXywNiQMGxcAM+u1WX3a2ZC6HaQJWJ4hOx
9VRJDTpxaBKBbKWHDI8SCPrOpA4DVzjve09daHl05O0Fwi7DqKhvzZAqd5IT39vR
/cSETPuUJWBdrrm9hJw5yVaRd5cLfiZ99SaumkbtQk4rdS5sTW6mWsNqWoug9j6e
PaRV2pyKufVjtL8f1ac4ndhivZ1YT5u1NfOKPqVNEkdWMW4DLNteZR6ZWP4iuVKa
PIMbEaraCokcspF9EjtRKPWTGBrLR5BOCU/QC5/yLP8WWqva+4Vn+BsIyopMTXnU
fudpEpmXgr/aqBX5BC6o12is3NxtmaL4iKdIjh1P1W9Uu6qOPQvBbJHtJbZhi5Vu
ebRmqRW3+DPNYGpDeNgeGZ8WXbP85sm/Tp2xPQC53EJc68/Kdhl5m99g01Wq1onj
NsfQg8j1nSWvgDtXkZXCxLVSA588hzhaq50Sn0UJQL4f5kuS7KLCPiB5W9Vts8Q6
NhdFAHl9NGFNKRuwZm0bhkZwZiB7gcD4zruyCXQkFqUJff0ccjAEdb8AL4Wd3b9H
AJmHr6zNwQOrK0kk8lVhli5J57MFd9e+56Lp2LnhhVyvw/QT6nxcclRl5hzkuS/1
qTB6dnbla4ykqpMtqlFtXR9PIWQ8J3izv2swPOsry25nskiV1BH1gmj7oKFK5RA/
CQW0H/YLuuu2gARHdBhGcCfuafuEDUwXVE7AmXPF5JKa/13vz5tb/3VaRn+1W5k3
f2jOe6inuKG/9Br/k0uvUepYfCR+2t4vPxBLHiCWEbtGXpqmskKhahMKZHGEZB18
7jXxve/zZ6MfRzmnSfo7+wcvDjF7PW96l5hAqqj5CjiYKrWF8JysNpncTVFyqMWu
zDLOCK1HySGPlB998oaPuwDb7Ny+aSBkP3o+aSAILfBgxmxRv7EXru8kSPQszpFe
Fi/VjQC+r/7U0NhBbJ2p8J5uoqKfR5qp13DnVy7Urw6dYsuMa6yztBew4zzIL3Od
s/Bc7EhMJZ2evTAqWoyHxg+yCEmQaWH1MM9VySNbudfrkmMJjXoDDMpzcRfbMgmT
TeJeVFygRorl5ajQ0bUrxJeOr8vPbkmixKVFh9gzzcYji211GrtSpnjpx/XAy+iW
drz9lb0aiAhDn3lw0eYIz0xrB4U0HXjvgn+dq/S/ZiDbbfl8/3L0IUNVzlEHr8Cl
vVjyHHdWXEHxkV8fZqbUjXbm8PmPuAtoqgAN6ZanCHY8K+RrVvltOOjNCzleiWb9
BQXzd6K68pNYt7wxrtQsGyh7UDp0H/FvjpLhkyxQXu9bzsyT1SxTsTZRkhLfNY5i
ABsQIiRoWH+TIknRkYiJHppY1jWhINApHErB2UA9fqqgiTdT68gkMcrpChXLLXAq
Xz6C0fhrUDnUMxi0Q0VGxp2gs+daf19+58IExTaRnocqWPqQrYwNbyR9+BKLy6ZS
gP9HOXdbEMqnykttYxxD4G3IM1AWCyTc6ADyYUKZuFBN8VLmmoZKAp1ovvioFjnN
Xw9rV4k6ubyLcIk+JSXnNhyJkN9zpxi2RS92H5BiumQId8/dUaP5+P5Fc/W6EV36
o3vKZYRZhoec/WTa7myWih6P2eiA19EYc9RgDrgTfIgj+hzPlyHv41tnaYKJHVtV
YZjsGryA+MUtVrUIMvS89pNtEhcNXyC8HGg7OXWDuzRRCnYoHFkkG4Grj0NFvSop
lC1ERewmifEOj1MXNWWTGUVFb9D/rwVU44Eu2VBrtbbSt0E1eSmuOXBvacb6FidF
gDLmgEBH680ugMLQNhyPmWvATSo5PJJ1MY9igx+si+BRCNLp1UurDN+TOcVBP7Xl
3O7xCLEmnzFHV2KsCl6O5V+la6vG5dT21hb5jIDhMHvfraPvJlCYyIGruygDdb4u
ArOxPvX2C8MnbZFyINzlNx97lz+ngmp3jcrZ7Pltas467AmmHxO87O0gzi/Brtrs
Pufcwh3SKiQnpCriuaXsz7EH0LHS4tkb73B7hbL9VaxJYyxLgrqqqngqA3INANAD
rPCSBX6vVJLYPi4Lohat+yTTkInaRNkgfo7hSbpR/o5JfAd9DVQN2DjRs6pty9Bl
bArQ9s8KE/UhgWk9PWXbwhlpKT8czg8d/CUSqiAmVYJ26yRoWj8hzl+KWmvEAoa3
0qUtpehK0FT/eo/SBUtF5OAn0QZxCp135EHgrXdnyS9VGimolE93IOZBKE/fiV3K
i6E1BxrxmdH+rz4MB7kmiSD4NLLV5q+3MO7YX4kArgCnmKnZxWJADxhOhBwQL4SD
Xgo1BsEjz14mNDoy18MAILh/OSiUF67THwre/YcFnwmLiAkybScG8PgrvEplq6t9
x2Dnhqt8a2X4RvZKU/K+Ms9bhJgU1MG+wmOBZTrPJA6TmGu9K6to2ES7DQusrs0J
EHbibPXNaHLWNnntMv2y4myZO93hAbxema5EeER46wZ38xb7nNPcOIgYz2BcrUAL
xE63Gc6b+zYeMZNMJKw9wJLFqW3r/JUPRcIK7zSiuS7v3uDhIY1tORYdowlDkU4K
+oH3F/goQatBDQkV6S+n7G9fow9i+42/VQSz4oQbNPYZDc8I4pc81ok3SDR303Gr
2mWdGr8jiJbW7ootOecBJaLd+R/UMWIiO7r6q7+0vUvNqwdoNqbx5NhyKbJuuqe2
pNmlKCHFoLtOcfnQ4sjA9DT8BWisZou0OEFDyc8npxQHoSmN/qcFo1OscBekTod7
nJ1B169M9xdTvVIX9uaKXjAT4nc49YznapFQgHG4IiGGh4cxNgoup01Ih8nl1GoH
UsCAhKIi1DHMxbTi1livfk7FHs2LEAEUj/FMrGnmq9a+uXu791ph2bLCg/Cp5EGv
lFecR6zv4O4NkbVLumppl+jt2X5D/S4OiJ/5ExN/xYfaekcgpVIM7jejev3T0FJM
8wfhaBuz3UwhaWCLwWCotki/QLs3VABpI/pt+Vxq1jzmz6P1InV70dbDHfh/TubA
fKuLZwvWHicMZmR1RB/gJBepPn+1cMb4K/eR0xIFMuHGUcTBxuPXpC36XBwFJYqh
ljnaDm29F+JrcEOaSouFSg3jMruf5k2VqXfwXqb33FwULr4Mu983qFrSt8uK0kbE
YeYmMQK/2X53iHTWw/7ck3+DBzxKANZB1Rl3U4+zrWR90oWiyIeP0GtVUGesFzOF
ih55N3md+y/Ik8jfq0N3KfbgROavc8lI4Xd0+SBbLyqbUWPv9/P2YjDLMG/7lx3u
iiUiM4ebuLOFu8Wo3/gM20HENDz4hr8m+1DzLrGgL4i38JLQBnnrwattkaQ+ZS1H
MIPnN5b5dErX13k0Z7tdVSRBZl8Eh2meEnFZ+zo2/4O/gmahqSIDTEQmW4kJA1w5
Pvkbfojiax5MfAf5Uixj0vcQWdRQnUAnlFsaECETPIHIP8WVq3HAXazaFQH3JnRu
D1zs6M2ERAohT+75eM13dJvPPyKLnfhDLNZwgRGTTEQqyCr/ztIHC+nfJxfvlLm/
a4UpcPcJ+0ji84Hlrlfme6HOVvOMjd15bA6p5E7FgPdoSLei5VbQ44VIZNzpBwgy
fS5Q8Cv6ikJUkm72vfPu5/fNVG1u9wRSAb0WJPOFUWBlWkZkZQtdGsSfE1u5+L1i
RzEl7cFYQEG6A2X2L10EDxjROHcHo63ViYfnrZarypsxoZC9hDmf7Zqvbyjo0khW
ze+W9ok4wtZ5mJTQ/5SfLzjNp8H1CnrML52gBid6jBN2AldGdUU0jdUKr5gRSwkf
6Gr+EZKGbPh5qNQIwU+Phk3LiL+WpcRBIFk4CVSSFKc6AV8d+ua7DvjkIG6kyVAH
4V0xMpGAteD1ej+ydjlyu4VQ+LMFSV7yMW2To5SP0oEgGOQWbX+ztBlcwp3IatRJ
mAx+X3iu2EnrOqqRynMGo16+vHNLS3jd+I/2cUp8uh9hBIwjKSI3KC1yJtOCDOq1
n3S4S0CJzSUX7jAqfRUzpP4hoCeQ8OHfdfS5vlw/DiSRuUvRKBKdhKObxGXT5ryE
O94H5VbbAq3JWjrjQvXbJ0CeY71Zvc3p+mkcPxo973yksmOPg6qt97b+gR24lgeZ
jQuV90WUrVf3p97aXbwt6blWIKjgWUlk3L6xUcQXEZo5q3ECPdLKaiig89NFR+IH
954T0EsXlow0eaMwIWp867dxOSlb8xpdQ0vtj/iKHODGlwngyKVRC4pkXDfYrF0N
t2WShP5Nt7JR80GiydUdGcjxxul8zsbfYHtHwVJkJ3eeXNOQvKoEFJ1zBeoXmq4S
XJqYHj2E/IN3uoykoZd93/qETtrd5OIuXmT4JHkohcOVHYoKqq7fVTMJjv5ZH0CN
fbUqdQjPW9RkaA0MLCy8dXOVTMLUZryx53Gmbh3lYzAULH8pQF3qqmTGpkZbxhh8
MZSx9tSeWnjOBHY2Hw9su4SnYc1O3D3rw06vPo4+tJFQtbpQpMc9PSuy0PFcxj3v
01+pQPQajG/7XCO1o0xZUAQyusPg5ng4EsTlgVWCff2J3FxfKQwRhjjdoXniYSyb
JwFG167Z0OFyFyo4eYehM5cZpYfwzlNebdTMrRX5bq3FkwF83t5a9RemqR1V7XzU
BGODH7ViATlgvo34p32gbxyh5Ugx5wMTqRH6cF69hzs91vzwHcEJY8LnRwUgKRTy
LLSBqdA/Dj7dTb+XkpbP2v6oTyArh3e1USmT/Ro5DHOiSsRFZGSWsFrqBcG0Czb4
W3EwbcUREujrr23GZrKrvY+QlEGSxmLqdQa7uvLzblZ7WZwIAqNmBzV6eaKYDWc2
YLagGsvXOg5v7x6ODISzaHmXKbSEUw7oPsMAM8cnkf09hsez1Vb+c0LI9mawKdQP
m+z2gCUbU8H3u718goiilYa75yuNgemxpPdUfwrnGhhJfDfOlZwWy/N03bGgDwah
cbIa1JR+sv85g4JSUd2VLijM9c5GH0u2pRTCgTBJ8nbmQpC6MD16VBt739Gynoo2
4b3+PoGc1WwMKfmJS+9YL1Wq4SowcCwaQ2eisJhH8V6C7kHdRyFMm6c9BH1GO1/5
xgzryfPhiNBXUaBI1MDd9DGjX6/JTWFbaDhz7K+nibC4iXY7slB1sJuseojw/Dpb
kX02OT057/7xbPyCfZ1utqHfFDOJCWQy7b/APopf0nBGgdlBnyMCLskMO673APHZ
o1jeBNGdJ07VLtubB/fLD7bU+p9KHqHP793vpdEvjWgDCdCdwad6F89gUuVr7YRX
zqnEvnWP7mWFJaE9tGp9c+q4c+xujsrALYmpduWbuPbAbPGTPBALVfnQ8T60YWLG
rwj7I72XBLvpDEQPE4oEnUygOwGbE35wCmCOORDOGAdL3RlRuvz+U7w9iOf5yI82
dOnCxG0IH2R6IAltUtPPjKieVZjODoXkEP6LNJ8ZY1yFU/6mTmWYt158oWi+hnPc
rxEqfqP8B5PUItGRYrfc5Umq+uvF5k9xYex8wI6G5vQ6/TVvjHXVXg4zTjTB03DN
K94hfQ+XdItta/qu8WoOSA5icywdopxi+kY4UvexIyzhHmwc94W73ed+vUT7f1LC
YL+3SpD9L/sk/8CFTWo5rR1amVqRWDhFR5oBD+bnIW5tQQoYI++hmsHUPggeqCqF
C47oU2XnJ9/gCFI5Dk7EkSE6pYWVm8PnhBd1COyxpJrrv1yPKC1IgrNKuD49c4U4
IruY0+lJsxImK02Yf9aQ5Tf/F1M7mDBYN6EzCZWZV8zbqxR+3Fp46gm3DAQEgIdl
wgnYGxPa9FHB8Kj63O4GYct3dEkTNHpE9zgpiZE0QEm86mi1cjek03v+j1n4Snr9
v9k/+IYxRTSBKHZPRf328K/ekgox9QHEpRzQjh+HYCHUTY/lDoj+olt989pjFIYe
CbfCeUeq0QD+RDG7OFt5i89daQAbenHhHHzNR4pOA2TNfHW+r1pQnuS2ajip3MKg
s5kr0STeKs9GFA16Uu2vWz5y7RzIrPfgFmDk52Bo/Hl2UBt/gGolAIlecErS2seK
MUDQohDdPO6d4m0ULjQlBWi/2nSYSXC+dphq/XchGXs2F8Hq5VFC86A9Xo5209KN
R3H2ZnSjUxtAxr5fOXg9wSPZJgDM4c8SAvz2I3LyVen5G7tKcNBQqaxJb8HRgM2M
nlvwFgZfvbi6uhRJlkKRLMbPEznX87dAo+mBAAwju58cDOM89fZL6XrXSeBBjQXv
atE//uct8HxKdU1sEmpexP3W1nEwo3AJffUIwn+OdNpbEamteY3jpmyHKYF4abka
+miJ98e9FC+5se5QixOO6y5uBQiGkRzQEmSxRI1gcjAyRVMMtO+EKKRC3fBosJFK
+mnMZJeIODtu7Xkqv1wz1OHVU4h0qhspOQ3UzXoOqf0uIgqEjTrboT/xSy3G6r/m
aMThD0JQyPJddUe2A3q0JnPIihVYKZriNq4HozlWTD+rjbpx7C9+y69aryxF5s7u
igZQp+YP92UzcEf9Z6qYALPgMbCMSpG9vKP4qKOMblOi4LEHnN0BJEnLTgc62HyV
ccEXvWcJHRrQxptV055dSHXo7Imz+zewgKcSrFhqxtf8g9Q8+69hWFs30lYvLojj
lVEEmJHcfeYciYAJtEwMYiZOW0/NUmSrP2RbwOsYoo5WP3GNA3wEMMKUim4iHBZs
ljDAdTRMgYRDsalH8CBgJivc1mZpcs+Jrho37v+uIJJXlWlWNMT/jqymxoNOPu+P
e4zAfT52KZqQJRzSo+5tFGxbUYqfdCMKemUQIGtfubp7JT18A87z3sUv+3MYVMeq
yDU81gaxPmukmrFkDUaxcVTJM00+SxTKlUJiKEHvXkqLh0N8xfzZ6yXjX1wZlqnJ
d9WIhHt2bPwWNviz7wSlcmjkau0Pgrpk+g2QdQmxFAlUzDCbsG3kmVB6PU+3j8/7
nFPtkMVQ+re0hOPksjfJqC56TvPv8Fa7fsD3ipoB9/Pl/+9hKtVHh56hFcpBPP4/
DCImhwejSyQupmtCm6OdfXyRdoAqvu5YncKWqZztEa2K7SyqsopO576/DO2iH2Ql
sfIw9GG17El3zbFpVMalmkxLN6eIyHFrm9/LPWuph0L4BaqNWNzj8gd4XA7foQn9
Oad7OKqHq5ieAjxc90K22kDdUeaZ62OgVgwtsTejzx1lAoZ/fvRMSgjQeVs9f5ah
Arl57YsfmBZUuyO8xwQMD97GfRZxtkI8dfVquLm9j9aJEfrDOMpAQBdtDJV1gYhH
awqeFDICtAOZqXK+Z5qoePnaNd4JKTE1s7/FibFKNDE2A1BFVIMOOkDOTg3qiH9/
s1nJSWdYGb4S4sMRZQCPtucHzOXA03ysyubLw7kcAWxNGF8Vu0wGYR5tXfV1rGog
Xt7K+wW04Icj1mL87olOF6/jFfPb2X6QqA6Emu5sK1RnKnuyWF6Ae9yT1pBu21i4
2F4XtQxS6M0eWJ0Jno8sTKb8/nF51vmYVLQIKDD2NMOwA3EJqAZGXmjSa8mtcZt9
rGVI4/BeIruCpZu5LAe1fZgYSeq70QENMe6eQBqwRaireqV5qXUqJu1zCtsV/k0Q
kWjP4yk/0bMKFLgG7GHBUXoXVubuG/EHMVWrPCgg+5NFoBRmUSWnW/fyON2hDt7d
KzJTrK59XpixFnh6pT7de6vcVtydy3LS6VyGH4xWoEva5TmWtb6kDr5K3RsDmaXk
1xKsuSI8b4HnhVAXUnW/oaZC/N1eu15yIl8J5Kh8iEwj3HI+Tg/w0dPkojfif2m/
9eGDBzQ3TBihG/Df1dVeIaKcuCG5SpblYYcLZp8QVa/t9MkKThqhugadJLRTMzkH
8SUiMEdIFpl4LjCD6Xbx9UjrwhptFbav155oqagLN6AZVA7cv/cdR2EEiBAuIAI/
5KNXrDBog8R91z4Zq5qS90Rl2i2nlDITHj4XLb/QfJIr8FvW48aw7/LMAj5yLVpR
FNXLvCoPKMBwSdu47fw4COxzm6/yat7Xuvvu+gzpQE00TRy6FXIA5B32t/XeVY3h
tEj8DGgGkql2zCs1nboL7yOM3NFSxiOuzThhUXwdNN+fCg7TYIjIIeDyld5w4f/U
vVhJk2GF9wDDknFAvNnxBtQU2H7OFaqA9mWWqTibTnvpqMQcUXFl2HwX0yMjQ5Hv
MqC6RawKdY2U3nyGqcTGx2k9xX3PcTGE7pzuuY6jOnNA+JV7r/S9KoD3BkwAF5xW
9EuggYk96eGVOtsce2q0bZ/NU1APAyyh4UrhwwVaH3fZsTdqht9jpW4IsV8pxK4m
TObd3wS3YmzdqgRAooyh3PpXLKtMrda2Sff/SjNmV23axELH+qXw58dZEhlAE2u0
+GKMJVMqQrQrGbzPRklYk2yGYVweOF55pNn68q67QvUWaox6ajg/k+7BKGI0GhT3
0o2aQeu6Hn9dk2ZUePmHZlWXa3FQXaFPLUQ6QnIBGDgReqngsnzQ9K+qBrnxdGVH
eZH9rYg/crv2VhZzN7pCowQLQyjP70FBQF1WKqVJ44NR73vlBLyRoiAQ+bMOJ5Jz
5hOBeNDjjaQPM4wlBAABEYxi/RJ3cO15AFF9L+OmrmaP2+uq7qJR18MJsn5SB/AW
XTGNXDz2WwCJqDlARekR0ZDQZwd9yDibEdIwEbCFGJ0fNkY4g+C2P5HqmGoxejVk
HT6mvp0RiuuF1zLbsf4PH6BMHEWYvin9e1AfcOGgJZxaf1xcjrAR0bVkZh7G2VY3
rOWHdFRBhGmunhlPYbkJBZIsIgveYPnkmI7tQv/SFnfFQtfjaT1gBKutPWKeAKvK
eZJ8eXpeH2BrscesySn8w0ozYcssvgwAInXpGIlaZBwUIDpUZTpooo7krBb5Lgn2
V6iJgpw/oApBHTcHiODFFJeXNP5EJ5fwIP6ZW3hr41B2LtwYaWVpvkc6A+U8PJXZ
RY+P2DjCJNBbL6MvqjtA1GDRQe1rRAAqjFDVlk3IcdcMMDgB3SlyMNDuG3m8YdDm
wfIR1UrEg6B/juI9aU82ZdYd87cW0IQtVZBR0ysqmzjSDeYzpP488g+kwuYMRY0z
MZ1ab7+Wq8p5l/dvr9B2L5YYIl6Hhk0qhSnNrNf/tqPgs5DIyY558iBgAFE38X3P
gPi29QnLkIW3+8iyETmXcSlRkVpmz+1W7r334zlhNFsYC+1Gt7ZVpijfSL0Eyida
acNePJlb4yGs1u8ZdZdkqLMWo/3jFiCK+a51oNvzOBkgBskrm+Z2CWiLEbxjobO4
aSZWx9MML7S4JOsfTx7/AGOH+oy5tFe2QAmO1l1sTxkc/TE7+rbE/lQmuVw9obIt
FIg8mw0GfXFVMa8iUwSRIdSV8iraunlVHxD8Hryl1JVIdow8myMUE+C0c4lLonCu
pw5PDeklephQ4QgRTgHARJOHJyhhyrquFxxeDlX2bZX9QLO3fl2mh4p/7AYw+wfo
Om2WN35hfuuLsjFOOxD5wQ6LpP+FrsUPoLWsG0iY2SIpEi/lN2NKSpIxGr/xmlzR
NtcuZ5rya7NUEbo8mH04EjRSRW/V/XmC4mitj7qOzreipZXNOVV2+ma4mIU+nAi0
gIHqaiq7kziWq5qU+T4XyMAb9p8MCt5am/5rE4GnrFYKucAkItSbFSYxB4Rt7qhq
eo6/+5+Js9kHav2lfJ7J41OkOfP68ouFL613gLVz4hwgv9C1ixZxbNpTurk4O/3J
TJRI5TTGcuASGPAerYm611Ss9mWGm0cyBVVOi/jfDD1y69Qk8JNFVSV+2pdIdKAx
4/765gJqmUa4Wu1jzp+4hQaevm9Rb8NUwe1ovLiXsEDEKiZxJNek5c+VVwTiIvX1
7HHbWxraq3BUvsJh/kYgYukqMgDFgc5f23Pq0WgTE4lE2qzSVL7SxBR5p7FuHUzi
X8f4nzgtv5FAk7slpQT6V7UM1I8Qs6VEh0ujPJCDTDMisvkKs/Lp2gI+oo09ksDq
b+LRJoL9XQq5Piy/iiKOxGPRiLqdtw9eWGkv/hkkeEkPaneRy+oO3AOZcqL4v7En
kxQRzibs6Zjr18SGDM5TQFJBnPH0paD5m92Iu20wz4UICJ4A/e+VW4ALTynZkXsz
1QpDfCl+3LlWtSnMw5Y6w9gUk5pM3JbXigx+Qkj/t+BeBML7CjO9d1NbsYjFdQAn
vVVbWFloMOi6s2bpPlByHUaATNkS5dF+hVfddkl/rEY0acbXo2oEL4646cRoQcAx
cMQFt6bVTDtMHH7vydfOdiJxuv76MnsSlUzAmV0H/8cpOMeTipZfGsUtY80xkOi2
h0Emg4KoACHtdvd8cI/5tEOPESu5BS98lVRaS3hPx6odNOJUzdtdlzEJpTgaqmD6
wSjUdOVgKfD6BjjmEjs/JC5WgzKK67IPxJfVp2AOfu0Ea+hG9DPLoyXWzBkN7PAV
p5C8KpGqEY6NcRiUeqmjL0D/wJhoDWrKYX0OT/HcpCa7UyTeOlLjP7IE6Y4vRQqZ
4+5Ha/YIbI/8Jqio6ckx6o5AA/NdnyFdDvEkZJ8RqMdtbwtL1oISAvZh2JLjeONm
a3XhGhF6RzAV6VisjQRmPKW03DZmdbwT+dfMfV32UBnZC6GHl5iPplhp6T753nf4
tivIS5BlMBxuHwCHKeb/KLr6hEEwUtSGzU4oxMduxgwqVJFeY4RPBoNdtY3UgzvQ
KFb+VEpcbN8nzlnbVaePady3WAG65OEhw4BdiqPWt3FOqcBCmA8dyZIUUW32nyUs
xqot3if6zpD57Su7/j6/joEYIUC7ZwTXOjp3xLq8YLcFXPegu5Ql9xGdWwgv8weY
lUcTUjZt/n4CRhTXHk95IgSWbFNgiqrKe90AceWeaZO8ap/Hp5nF1lTu3cJvObdy
74Eq9ski9SKvaZzHEAdTFqh9z6Fuu2rzlc8rxlP/6J0+Cb1+i++x3+wQIm/rENS1
ftOOytvT+Z7Q/0DYJTuAI8QxAZJhmPX/zoG2HQIoCkjeHdsEENbEij7VgaluAXOq
mwkNLyQ3QuoJLq+K2B9NA/CG4R+TVynEC5LQPwpixdb0jtRi69mvez4/LTsLxb9J
4ohxAELUA5rjqccJGGjB2rB2JfH1vWBSmjLOiAvCVD1f4QpkMcrmTqMeixgBW751
V7uuDZX71TIkK8EITjE2oPx2ORy9ZN1NyQc803GQDo1AbDc/oWK1UtIiU2vJkXDa
zPacOszQlZ4ah4bBDxscPk2uK/L4dUl3IYqYGJWUBgxzDR2bCYCsqqXojCCUOBZ2
O8L/AUdh5EmM4SuvJ23X2l6f9dZ3n15D8RRyj156OmiOawuu0TuI2iCKMNLBpm0F
yuD+jQ7T9fP55RlvyjvgBTbCR8bLUAi8L6Crt5Ao0tXN99G5z0N1pzZnzy5y8VQd
XikmXR4YqZJNXxLdgr9YZER3+E/z79K+GOaS0NYiCeAaytNDhY5FNOWWhW3Q9KQG
yT4vdIFqM10V5gWuZov4sti7wSdD1I4l7VjHqUxbbXSbqHjNsQ5meVactZU8uMc7
ipFuTwzL2uh6+aZHFJFFE/ZT8fTjJ5E8R+/PhBhqMUSn8fjNdKpZOrkdCUbc+ZLW
0Q5p61ooQ3VbIY0tmQ3BCKwFamOVhaMOXw2/qXICmSvx7dlUMKvOfb7/BZWFP8V1
ZcycI7HsF4PjdfpT7E2egXNW4E0kBvGMIKp6IfHPGMs9Ks9ZcF8raNj9gl0h0pv8
PRY/vxvgp1WLJnGu7BWUq+kVHzDhSz1129Na9mGVDOMqZZZgjq+AncUwJkrPauXR
q0vJk/jUiircBr0noLCP6kuO3pdSe0wztbVCFLm1Hi8s0fFIVDrFXDpHZTijWvnr
SxtebKVwxlAafsr8NFQgxrCFfb5nu5OVA3D2Cs9A+9FS7e11Gnh5IlzkjLyOGxLz
eK9uhzuYIZv5v6PFiszXLtmvQpe+si0XG9qYov6ieCJfdGnRtmj6tCXWyCSWAsMm
F9+mAD/Y/fobjRxipLHc7HGlFLZro1RYsNwBGU/aydmcVqDnzPeUsO+0XE+Yy97G
jHut8xerUK+rO5ArAcT1ABIOFnZ+ryVkmhbK/odFkmAp+gVxV8FJjhjV49QokXCG
NvxWBbedL30ZgpIho0rVq77emBtdVx2qizERWQLFuFjNXSTGC9va/mHeqcGB2ty1
vsNaJwednlKZnoBKXTJWoGbnQASCgD97ExZPqP1AUD7GKi2dW49wY3AvUrcxfcCj
0EerTfXUAGqwdeIPQ1+OSgSWusnGTPyazX46Z871C8N/MnaiScuV66lWmNRK6JW0
lHQdKBBzAJBm6V394qIBfFFXcBz2d6Y1ChlNQrYjZUftcl6P/0kdJP6Lgpi0QA/6
mwzCgu8kZ/XXkE0BO/2PAIqvdxNJaUlBoPOUytSnk0u8SgMyUSrYhDiTDTQ1pL7a
rOq0PyUqa12Xy9rBQ70QsyNQ/qxuECr6PggCtUhGYQQBE1fMf/IA/JsfQrOnBAmx
IxN0lABZoQhF9L/40vk9pn0wX87czqnslg/XxCkTEkNNJwAj/qYVMJ7IWmT86hJr
/HuHzXmKt/Z8FN+c5/YMyhH+6I+Ut+Oi1rPRLUOOBUhfVnB8mGUHzyuBdo6sRJ8n
6qxlAxNabjGVb4zJpz7CyAQDzsU7Yo9zSznLWWg5c/SP/J+K162bnhvOLQxgfATx
bGi+rJ3EvUQoUCKhpdwJqmozRu5D5BdmZ39XWDHfD59cQgNCr4lzZwB48ePmkWD9
EpK0khSrUUbsLRU0V9TRN6MYuPMxHSlMssdbnJsaS5N+GGbQzBszGwXV2nT6UBHy
rrfTvyAxpIA2hCckRs/xftYzGGcLcmzl/r+e+AhGgK/d1lrSIC8bpBQuQyS4NAMr
Z2Zy1Er+7YFTcgQkKIQ6B6k9J0kQRbwIkDcNvsJZbFAakcIOtAGM6l6aLMGyEWWl
oK6zIU0tZ8yfXlVDO9XE4SL4xEuN3KJibh4JM+BgYoYYEVdvJGQZvbGT55nv6pIl
PDsT+7ggAnaXyesRQoOqmuEjjc9gCqpHEJ7OZrWT1Bj/dVqSEfKGoDaQbvYSe28Y
PAyZSkDb/+A8wYbdOLLWj1F1+XbJnB0V4idChtKcrX7m8bve74xfO3PwY9m5vJ2E
nHhOcG6k9pCJ+yhPsMqaXy2jYZBTdVx4RXmIr1ucJVlIbTvWKt8s1Hj0kpSviQgo
ojVS33tCfHH1m0WD0lJmQrPa/xuTHilHEFmBX2Ccy5eEOhcuEVjYF5h6fq/KeeaT
fS2K8bCQKLhGLEqv64QR4W3zlFALLh3rC01kwBB88dEL8EGv1uwdQAa4YOCldmrF
566akf+Ee7zYpsfPfaKF+51z+87zMKdORVuvXfHWr8EW06vAxvNGj/bE2PnFv4dz
ccFn8bH9dQ/6rUnVJMG4U2AvD70lMXwysTOa2gd4BfLPJ0bDBLHvTHA/X8MexidV
MnYqqr2xffZpLYjcRKihkn9EW9wLLNlDpxPEtMNoJ3ZFw+yEnXuoCCyPUL/m9FYv
HAi0umaunRcP5dK3WvU10ee/FikCkRi+9OaOCYDFlFJvxO9O3tlEPkhMMRQPTDDy
6mmOtSZcpCOTJcHMUhGLjzeh8VThRjP7mb00tk/MOhvT4aG0yI3o8M6APvxICRGA
N/11+ngjVgmywyCYPxC+rhrxlON8GYpWVQsCtvO6Bh3vC56J/SA0W7By6KA7x5wo
PbcsGPaU1WZBNrnxydYC8SBsUiRLJLe/RpLt27rWCawj21ymd8jSZfayIiEOsJjk
TgtbYxXXO9o5+azPbCbctPLh+YGJnFq2W7XZMpqOBcwX0spg7qYGiKnfrrbYI2Sb
t4xUzIGH2ARq/omx90dgTuxS2qrGeqeh7a0dWUVJdKgtWuwMXGhrcC03UtwPA1vC
TgRI09LLalAufTgeyOxoHVKm4TwFuNt57CDzsHHEnJhotT2u0lvu8aGOWk6InHob
OB4B48GBIyJhrnJVtlYPnEGhH7fW264ry46AZhHwnAxelro2s4mrk4EqbFessF8x
/eswFapVnCZ1DHroIMs04RFLNlzRQ2brYyO5/d5pzmYDjHhy7cV685rH3Z75D7gf
Vq6YM8kNAPDurnZl0myaJ454seabwAx6Nf9o9WkBf30GaFscBRZ0xHGpIRE/Twus
UOdgkiMUa8Xb6GhzOgAwHHDRdLuDCeO44R7aQDtO6MeUbKqTHjMn47I8N8e2tzQZ
JgKUrJnn/jH7P6AgNcU+aiYkPKRyf9NqUiBXCLtJl7M2rrfihgqTP21dKRz/0n8K
97RiCz6AVa7d3qswGcvj7PUYKQDHFlQ2yGBKCQ/xUmL19obVx5bMFEZNLv2PA7/e
+jIiN/GMxL2rT9fRHXcjYqFyHBOvCs3R1LPhoRAQiRWfc5N3vjfPbeKK2HnUIhtE
kuT1kMJxNEgtDI0DNrpqO55j7O9sGWERUXUgRYgRDdoipLgE5YuBfsJdbjtnSa+N
7FtpLQNYppn+wCkMIotXk+UotB5nYRyBtNYr3IGkuT4LssetkNeYqI3F5HKGKThM
jZ04okzBpNOr4C1WeXTMGmbSBSsL/SsL7vsBTGFj0KouMYj2J+yoG+Mib6J7vJCd
I0JebyYTd0d/pfOQQtLqB/jhVDPqRSf621EPDJgwNLOse2xjM814ZiNgQMJEjrbA
IGIjpDJW5s/bHtWJU5pubQls7C4sgPnErj4WL7rEoAR+obtxJWsTunGDfVGZ8gxm
Hzr/Xc9akGDfOWPMcWdejt5okCJ+3F9k2zTFQXvUlGel+Yt67sC2nfD7slxmdX+S
feCqTodoFJt19mtgkofKfAiOh1PrgB6QujIwVZ/lZ1HwP9A/FGQy7FbM4ZGAaKGb
olrZCmJPkV97jGx0tmXvYZnEjEfpK1c12xxqjdzBpJfCZjoWYZDbM9IoQzxCE8rS
LBuomJxKuiai7aUhJ+Uxs9Oea05mJ8CzF2BlLLxhDIPoIst64jpMXZkRltmYorz5
VeillwjI5esYuTG8jUGDAd1+ftE/qg8cd6DNP9gOoWRX/tZKpYBDHg3Rgznv8Fdh
5j3h+CG0xgqliL9supXEt4vAd+/w9NzB8vdDuWngu7ZPGLOumODCjaLKGQbYfpGf
9m0uksDhCrDOsmWyJ6yyURR325H0CqXBMIOaJVJ/Yoz+nt9SfquD9y2PFGWr8gD7
6IkubQp2EMJ45zgAOEvPgIb6sLGLOvU+vclZ9nkTSQx5I4hdZmEqGq2fNIQGd0Gq
X4RYJUkiGScpdbTEjJuUDQEBG0dI6MVsl+FDFU1A6zJLPU4hgxRrRHGUf9GX4D/X
Ur2OgSxzUN4oh8yfnBe6NpUybNPJzP+70Xm0dmARAVpxb8PUZpBbzGAfCnnAbN2e
GzDau/ibdHaeu8Gor0yKMzLHALyBLsuYmThMbMHqVN+bAftQuNRjfkoviQQ3LEyh
wq/qdEdpkejWGtQvakAJltCFVxqEGxsykXR0ZzRmxk3EQdIwKQJuG4s+7Ek+nUm5
hZgm4TZZoFVSv6REumqrEJGGiDQWjuvhCz4+Ha/RR/KSa9a97G9rJTQCFaaYupqR
5MsBg2Vwl9zgWSUKaDJb8qNxaRh4RF1S38o48bDmkuCF94ytiozdPv7uNeYvGsbT
9N6FzsCIurffTm+O3GACRtaUh8grprfolv9u8IxpcMXZTeM0boxZOhAGK4bn2R/H
HSy86DZVJV3C8cmKUAwEjEBFavy8N8TB7j2TN06EyrTBtkCWkCInaePKdBawnPn7
wxfI70DhME9gB2kGTXy9zyMUfI8RtBg4Ap1x3n0NIWKi+ATLfKT/Srduic/ufkpC
wxOP4jdHVxKKgy0oZV67bNq0b1lna3yVAjYkbb+BC6omJkPVLAlDQS6GGc9i0gdS
uW0rJDvbOIT1cEv+xzm8E9rJi461Q1Ekl91Qp0/SF4/eDGPdDOjTvgQ+IGjse1Ux
FMp6uOh3BW+kFFquQsPXQdpJ1glPxJb9tW8KN1J7uYp7z7niO/LjOHxVzZ7ePhSR
iNE5lMzGcx9+8Rbx1eW5k2+KLWsgIYMC2edkTET2uhBH4qnQ/XzIg0d20dlYRICF
m0dtXi+l5FCrpis6+mRf7g95TrOaoXr8dIKRuRH7W0hUGAv5arrkLMpTWk64ZBSl
fsdzGJsg88uSJRsm5uEM9tJHGwEwuaYK+tJi3T6F1k824BYRUYqlyNxkR58CJ8kH
aEn8Fv1cKDkds4xOn36pVnocPgzpRDTwfp1p1upmNYvBCIlA2JXX2v1cFu5W6iDM
Wd9GKOjmxcHMnX019kHm1MzQu/W7KEe98nog3JgUKTBKZ/4OBWXZMXOja7k+ONSj
EI32zqpN9XyCss/pCow4xsbDjUJ2tEpRLQochn2xmCo/TNp+9MItaU1deFWMlf66
DMYogjYsMy9knLa2yKg3mQUIM+JK05j12pnohz7j97dQWDg5EwSOXHJP0Xv7cXFZ
So306QvlWPuh7pJt/mOnWGfLtGbE7nQTf/hs/ekFZliGJLvBC5PqxtvQXKIxmbkk
vSiE6xWuhgRCKCGFpxihk3GdkoSeKyT25PEIViFDNEWiNdWRQB3HM+l0XGzoXZSn
VVeK4TL1D/bl04G8NEfFGNsg6/3oefN0y24qIID0RslI8DMEeBaAc5AmkMLBaTsn
Nx1h39654ArWuOGecsbrg7olr3hd1//p+kfmj0ThgA26Gh+F6qbaIm+3ooHYGG3W
zuJXBWXSwoQ6DhJaMsjcrTSS8Ouyl8m9oQVO15+paqioe39ewy7JX5Em5Sm0WQD/
UU6YK0bZ4JrdOyRQVJTKDC3f/Dry7VUjgFZrmAinxeNH2nzRsryUcDVbpcB6qWrk
oPB42nq1/fXmGqecwbLkeUkPt8+HW4TqMjkVnAbKEu2mak14RS3zILqf/DqS3MdF
iWWhwz5I4xY+CwoiRy6tYTzY1+c3nOLOFQbXEqQ67MuzcBFgIzkdnnma65xlaG1B
ML97j3CBYFVq/mpIQPaR6eQ/M3SZ8aedtf1KAqDfrxAgNIJnQ2A4j0ED4uGZ0i35
eFSwXUIoIM+syWuQebVL2vNi9fDRqsBLD9Zh+npyPivLv0JeMQksegyT3OaMvj/b
tS0mu389prE36u3R1BIuadDhReqQsOcbggl9s1V/ueBsOpSMNH4pXnLprDCzYaoK
wNOwoZ1edd7jK8+klet011shBaHS1MUIWgdMHs22qQwMhWVnVkv/iQIAmbcLx9tE
I+jU78zAZhIkJML26r7sPEj8K+Fcsh6aHnF/dhTzyMU3/oI/PphwKDwYdTZr97kP
DCuM02y9I556C2R1LNDlWp6mjnQUFKsZRhQxMihi/0k0EDlm5VHIdNMxrHSaX6v6
aiYfXPD1tHT5JMkKhRLvBzyVfg2hqQ4sReXLCbR/OG3Ln05ExhbkNRLRbmTXxwMf
9cp6nQ7+wUDxrmEutn3ni3kd+fVLpNOk6EImdRUVial9ygB5+bW0PYWN4BvMVSb2
JM+YDgwH5fDB30ZLhb1OgQ/Vpm8D/jDV0G59K33vwY43VMSxQ8Eiha7pMva6lty2
s7gLvTaiXkApLvfO8/6a8pD0TatNad7iiyV8GUpJV1RCBMYCHXlGfE3xuzH49idz
evKFfuttZwtAAryvzyQFpREGsnFWxxJHPanKPtY3DdVPUG3nxYrfZmeh4/Sj6yxG
rx+EO2omy+8FDP62feUxaQ9mqxRJjOtiLMZYM+5DTipVXUDi3455/mV2fqjhUwPR
hCRkPmLWJhegLa411bT8CVdKmjbidOAO3+NVWzzCKn5SBkjM75Wvhg2Sc4AYEzSq
dzI6pLi14e7az6i7vRNka3bl1xb7Cp0cJTqwG2YOGYNhXv2RqdDaYGvLmjG19vBn
OxFSHr6BvC1irVx5a1QAculM2fQ27fGXJEW5yNmuTRuwpW6Vi4H0ZIiwFeeJjl0y
/4RQ19b4xKwwdmyTe/BNjYWO/i8B4vJfIfXvTdZTiNgVVKtrHiYrIXTkLJzj44eR
VvH0ZTafqfp2jm05cmOzdEu/wNMEbk0IVtsrixpTVFjVTcWbd8BBNgmfzGkmwkpw
I1pSIUc1R8hvNRBk7HvEr2p9IC2vOELK+GJYHQ1YfkuZr8eU0bZnwWXrUDrZlcGy
cX+YE7h2+iBDHrLTPxyMveOOOV+GlyPWRkTSOAxrC95LQEI/H9lwHe9sHa7m06QQ
d7UBZgoWGyvaG7vBfw3qKniKLtxWviq4a4XFx8VTODay/sHRcgY0xOJLNHIwHwt7
dSaDTc3lCLLgLASs8qKJSMbsMz/qKDNub3JsmCVN2kJ/WDyNnivaJQ54u/oh+bf2
btG90+RxrX4E6BJvrgIQu+NWTJQG3ZOS8fLzwc5mKBsUc3+GFemC5EsDaepsndV9
DP1NkrYWln6toZsXCLMoNEaKUWfh/an65j+6Hjvo28HotUx1Qk3xwVQgRKMhSQs1
RSEMbXH3bP7V1SUDlND9caAG2MLA2ZESP/4ivnoGxwkmIENdRshOefylwQhNH9qX
tmgQ9R3HK6SJics8zYrqM8qKG29+FHUgTQ92S/f8ArYcRO/hs8xyhKMHKVfa2m6a
0O/0jrGhrmpJtGiRRS7TeUhZMeRcCDAIBs9umvch5BwD6mcWZooAWgJxVCBGnArC
pJufVIYd0IWZO8XAIoWhDESRfDVfcB0Dd7IB9Jcm4mNf6OIKp/8gvqOWbiTGToB9
K5PMVWvBl1expIq4bDuyxCxqDfVG47cv+M0ELMYBQO4tFZZpgrOTyjy8R65nsQGK
QwPtsNv223hE0b0UzC/GbkuTIIteQZIE6XKBD4tZHqIFgJU0D8y1jady3BRw1lie
zFjlXep4G2cUXnago+vuLVmcxR3iwVhMavFVp8DFM5fdcWcIweB2SSRpby5f9HuV
um/bVu/fAU7nvV0k6Cc3T+Z8NwSU4GCZWSusSeuQi84i/LL2U2dGCj24DIM3Ocxi
MKXI5N8Kg+BKDsI+Xdegiq/9/L7AJ/s37CynJaT74DPFXnBCreY+Pitq3+3tzg3A
Vs7J/bcA6jDv+jNNsM4pjidWL4B7PQyKH/IMy2ACBSDEZoLnpaCNJxByfy8G4dop
4WZsCjsGrOhiCiVYpf5jZWHQPN8TkwwuSw5nXb9SHWMbTdHNhTaZLaQdGQygBUYm
aMQPBNq4p3gpRDkpVTvSwTze7bF63WJpJ6nwugL91dUAqfTsrpLrvh4rewwPJm9n
95PPrDIRpHI/z6w03DdKnV+pxSOFIWmDZEWP3O7ty2hIfFSdv3kkHrVRdmzrElYC
m/2aOspBhNAiKWyapq5oiVNwCJ2ejUNmU8IVu5ZZDJob34kfn5hsh54I3hybGIMB
QHXabfz7jWiv6Qrm2tL97rOUmrjU/BLDq9t12126PVDA7akYlvNr0gl/TwRnnG2a
scw+Ji0MFWY5oe5wyDqfQeaKqPB6DtzsRWEYpAONqDXsJ6feie+XQg+z1dfM1quL
5HfN8WMvgq7SJjDK4geAFBbWODc8t16479YCCM9QUeIGiEC/32pCIPcxb0vkaDdW
4oC4y2HnbHT6A4tpMzSJTt+bZfF2kLvOY8TrKcGUhIR7sDfpBb7ipjO6oRQQWrkV
79X3etJpa+iDNnpzZY1avbdNLHkbKYyvQ4ecRqEAy9BX/NbJOzClw4OBKYBDSsHa
yTfeLyBBfmLcOQ70jvYiqMJHtFGPBbL/+EpWkwu8iwc6FwiZpqdU0u0cAw4zW4sX
j0ZjRSsU9xa6X7Qlz/EzAQXxbfHX59gQPhCzVy9dKtkyg6FOrZf3mSHJ5H4UM64A
l1MUsl9An2eh6Lz+wyjMt4FtA6+OEKeI/jsIwFe5ujCf7uRTRRhEimediIOxU35j
CosyAbmkHTrebSoe0uOqWqzcp1dZ7FUvwSvWKU2eUNV5Wa1MYi6QNvzgz5MnHW9j
S/dcetJJTZpBZY/HiGE2aeyanqiidtHFi3Unw8IH0ZC8+xSng9w9kHK0lio0c5q2
N3m6AHhlnF0rsohHKw3+Osz4ut9yDqO3IPoQJFZgZN7b7Z6FdqniPdJ3vPYbmoTi
EOHrFXFfFKpSb9B5g9nkyCYJwNcM9/nc7bnef0WK9IKs79pQSX6c3xJhmojxYxL5
Fo2vVNDjQizgFufiJfq/bHC9t3b+oFyvyyp4H6CP+YNiYN4C8X8q8oqeOgFAayPF
tES0qMVP5mDglxuF1EDk4uPMjR+dJEZd5Srp45Bu65y5Z4Wzdguk7ehzWkMJG9OG
Rv8FZPUkTl8IXQWB406Keon+7Rtu059rpYqL1w2llHA2UYbsVw4isdf+O4h+Kvu9
QMUHkKML0Jt1HpmhO4/7x7srZxMWDEOdQl/SyA5bSIwA0vEKtae8Mvm0V7VxClS6
9bu2xtcjbY+MiZzN1K6mnOuJ7IvoTCjE8JficDfebyyYAyduSEMlfVxJx7mYqBG7
Hw3Kk7hE1zvmaS0BnuyPmH4WnVJx63MQLGAap8G34KUfRRA9pCgc2l4sjH7Qsz4M
lys3n8Ez9uY2QjZrWNKN7WyIeJt2ey1c58ikye6zug10lUl9whn9Ig+VjamXRbJ2
QSVYwW9p9GOKIJ7cn9tt3Dwzs0cF4YnEUU3zSEDKFzpBIxqNCsJvyZzm48M5cezb
5fRNvq6vttKzlvc9qF7aiMhOgcSUMGavOMCYk4vVj7Nt9SGw0Ar+wDu8t8KecwUW
gJn2rWdWlEGxKQytBxFLy4ERfEtsIMCIwYn7N9mArEYFCwXI0rFu3blmZnMgkTAE
ls9ylgzD6dfHW0sPr8QCp/eewE9fsglK/WkiFQZwwn4ICMRu9Hpra8+XgKTy9S83
fwrx0l3b+DC1S8b47PyZTZbjAQg+3aYyjltfHOIXAcoAsVPRbhHjrRgNpAVvBMMc
38rL8i2Vn9z/1QT31mEcIIxh0aVvHbNOH/EEAruf7xZRr1tmgwSG2I3Mwht8bgfs
uxWwBZUxbndZFKGVoIfwwy5gcnBn/dn+77lSAril4oVOSsHKebNcQ1wIbdMMJCoZ
d/UxBiG0IJZMQzw1pHNqv82wrS5tPDO48VuelMRp5xGQt//AN9aTgEZupFoqE40Q
beQda2HfeTa35+k01HoPjGP4E+5AGzZykvZyvGUf5T0TDyKDDUdxwIF5dKKfgONt
FBUnLi+UsrgNP0pE7WU0x+89iufmaIHg6uqKaF9WMrV3yFzZxQG+sCdVixhKK/v6
7C9yRS8FgR4RgAvjxAYcwOBfn1A5/p3A7BR+vc0w2qzFJ4FGcmomy9+6fe3rTfdB
Cjw+M+hHYm4xLivj72C7RgjUamXz33v+ui4BEc3sIA2oe1p8cqWYQEtZc3JU8lVu
IygTwzbw6MOvPJVQp2ZUActx2f5VaNo1NxxDgDI1KV2hcmoQToYT8EVV5i98UWwC
Drm7GaLhXLKjGzjYSjPrDS4LPW1qn+fkA5CnlbLy9w9OPNaPXVKM5tsdshw11zNV
F9qy+03m1r+ViSOHNe6x0pKcn35g6ADAwJ5oe5Id85p8swKW1zYUQZSQus2j6g4T
tDpVMCtD4MTEa9HtkhJYFTarsVNx2oXFBdG0SbdnulNxxX4Ea/94Obd2meBlULlG
H40SUUKoIGg1YRMj/jHwikFuIbMxt3QbSGpI0dB531TiTK5rbgWO2JDSA+JRdVfN
iLQEM+TrZUV/5DNUvV7K9ahYMW9d+rxFJELtsGv5cgZPjNNmiLa/IdWmUduQqwgb
7UpuTzAIQ2k1A2uliWMfGY+bXkhA/g1E/slJxBLFDnHC2ivMFM/+aax6y3zkSrO7
Os5WA8EsI6ZcAFOUmAGKpPbVPpoWUMHokPmkl2N1ax3GxCX0tpI1Z3hZAtfQlKqD
2BO8k3vXSuosWnhmHW8s2eTOvBl5EiKSfGS86ygkJUU1J9Xckxjcrq02vE0a+Uo/
J3ZabhWxJcFdWnAbCkbiVNDqf7IR04aMdJLZTj1fm1Q54PR3GhwIiOt30lTeO3IT
qRXeUP2J0KlCF+A4Y8XLehUKHGtnDNkaGP/omehrb7rCEHkCZr87USA0xvkVE1qM
38kkF41u260B7pAIvEc5pbWyHRnAnDDEG96i430Cj5ARWM2MmmwGDn+JGpHespHH
EMzzta1nugXk2c0qRE395dF8FnC3VHt7dHeO0ohUdJWpdhNt5ZRhxbCdahnRdq1f
mq3thG/5GXx9i/jFQYLcScuRXxtVnS8CDIYe8HBm26+EoEuosTdj+OVEnfH9HXDv
GecvP3RE3QmcXa5NqfPul6EwOLC23tZaHF9PBa2sPCRBgMlF5N8IpAFiX+yF8QuL
aWJMBv6wXQ3d7heVaZ4hMUunsDOMyqi1uv5WBUEH9AeZFOfG73BXxDV4EJTN0S0n
6w5q9J/UPtE5XH+oA0tb2IwOGfpOBIsyGXwNhE3yEcA1ckBqY3+ZgLrRU2MtQGUQ
y9kFRF1ffISPed2TKfglvpXBgKVYWPOnnnY+pOxuk0sjQiKoTXQEQ3oZ8yj8fQU2
1AiDU+uJcnN3mjqw/UEi7L343Cdq0kbpDX4+0y5WGXOSh8xpnonjnRiFK6X9a5Q2
u8wgd08zYp5/rOaWnyoqXnJ8cAqLSotqPPiQJJIn9u9wL/UpERxSA2U4ZL6SKuJw
l8BiV7jjUelEiLtwufKWslYx6mRImbmVV8a6kRPmggZK/C3k0bLNBw+6plWQUPus
Uqtph2Zua/phwjN2SfBrWooWV80KRcjRXPnwgoUEDu0IjJKUKOl3WyuAAAgxelTz
pDqF/2h+LAVSdB2jGGZjG2Sb2xN8PDkY5BWTj37n57N3yegcvFoUH7U8JZxegZuS
Fo/fuPS7h+5FHwGUGkLKFGZdKF4iBpcLglP+GsKUzEWa1SGozNBg30ClgNFqPCPL
ZwxbCbYALeipvIDmXqxGTsFXKD49brYBJwFmufuilwCsUsEXeCnQRL0x845x+Zt7
fRoT/k1nQR8J8Zw8UYAnOEnS9mM1yG5v0Bs/N+46Hzmxg6qRv5ZVqZfmIg8EnUvr
6G7hC/VC07Wrwi64zv2jNeldHCmSXAXhJpE9ICvMTmWu4WeZAOyayY6nC7K1qlSy
7+H8TpQM58TUtyIE2C3jYlxP7yFWMnp0DYsLVINLCurdfrl9Pl23u1ODyKe/aJF1
AXd79o4xwSqHI2HaomEgoXWqaBrL+WLkVau8B6Logep0CkOsjolz7my+mhFkmgP8
nhLQrYedN7iivU07OAqvbXrIDWe7hJ/JZK/ZllnwRVOApesjV3ZxsPCbDsO2PHAF
Ty4+wfe1DWGk8eiEoHWGTryjHVasvZT1r2cuuUTp+6NBCRcQ7oV27ZpoZ+h8vvay
NodS6uMmWWGu9v82iSaoNnaDyqAVEmZc7iMwuuj3sqHMS4L+ytDkFxqzBI6zz26y
FrALwhHfFuE2pD1caDD/lv7CcGhm3N0hQqE9qhC+zmKtEhWYcJ7mj6l5T8tez4uO
HJ6kiqREGFVvVPU5LXMpe9kOvHMQZjReFVxjt6cIpa4fSWHq6SMiez7esXiJLQh3
twpb3vjI1nNFcHJLb2RpFQ01JokPi5/u2v6X5R5TjlWp0d5SR7Q5fF2tq6OvJzho
HlCbEd5P7LUhlC67BNwM7OremQ1eQvB7ps+J/7/csYLhHToeAlarV/W5N5bkwzxR
Z/9OoPkmzVVOZlM5vMgbIk2yxZ0SjtNUEJ9nQRgtVpE7RGBwVAwvGOzf3VDBrJdP
9uvE9cincAEOCR2XEhzieCe8d0perSx03c2Ec99c91ZXgl9k9kM4o8LAb8eGQMnn
GJ7MguKX/k2PCAi9+/mD4EceB1QdMlcceyWFjSxr60D2EdZ3K/yVUsibqQd1+3ZO
GCotnFsSgMsi2B5fTVrHQqYgdqqzCwTBo4VJt2UGvM7Ad9A8P1yvzroyLJJePgsB
flbvYzOmwin05I4nplK7eoDCB/AHGVarT3DQvnkOE21Wh7tzDluJUYpt9ReO5yV0
azaabwggNiDkFZM3OM5IK92cI29n3Ju8BqUiyPxfY13XBgkNJcj70s4EKS4Xe6A2
VCsl7dWO2qaNnlpI/TeHyIro45mdhiGnjytgZZIM9aBuobdge8eKAr4jMRIYXV+d
LCNzkE/I8SKn4TxMocZUcmGTVFnxz5deMcJIIlAtJ5hRDz+Jwk4pTBjwfeyf4DOM
Vr07yaIsqVf55IXq7LLCx8zCvXwls94x7Zdh6deWYPffWlDEC5A8gpiLYShGKNqv
sUNVkbbrUl7EGhHjMmGIX2gkEZiGHY4tGtQTdcxXf6jjLlwJWRJ9Bd3U3J8sk+t/
F6yMa80MsiU9B71HhdEtPF5+5zW2ycO3AuVqEqmhXu2DrcUA9NYpyBYGRv/F0nnJ
31+24hUey9EMUN6KAh/ZL7I8frlUxgcK7lmPFJ4J1eswrTLUI3oO24Px/5vYc+9g
NKH8IjJ17kXqs60rMJ0PO/1+wKflWIAU+V09fOqb8Jomd0fcmObSjrVTzCmYNNDH
/9L7NLubNLNcBNVm6U0hJylo6aJWPWoM5IBAKoi53SQZFIf1wHJ0uVp7CHcq55b7
IctMwIoUG1gWOAq8GRobAHFEiiXPqOmM/gub0efED/DtAxhLnFq2JVJ8499tYvpL
jhUalwjVBfUes1UihCTycJYLaSPQXhF+9C4MH/hiOREN2PjqdRC1FAgMQxS0xw4Z
r5wQDR1XGdl2sTXsjOIOjExgb+ZSN62KtGCOcT2O+uT9pludu2d4i0VyGohNiPag
4EUmP2APJ8iYxRvqBXx82rfoIDu3p9joDdUAeSfWiTFwwDrym2O2Am3o5qUu8qIj
P9Qo/hwWbA0L0Y0Ov6DEcMLgez936RoufKieK0vnD0nm0E+3VvJaJa6JwWRK4K6G
3yugAGD4BsrBJZ3nZGj3+V3OK6iZMVNweQAjR/jEloyrrxNiDJzj10tWh25mDIml
1GSy/XnaGciXKLlvD3WDBAgmfSaHxieTxcRp4amWmqENO2po4VN1QY5Fjba1M1VE
WBU9+hBzzbd2hvNeiUGngPhEqOmRrG6MTOf1t5vAc0k0yL2Fy5IfGMNNBlZkvt5G
BCzE2YGeTgUf66Cm0udpiC8tuA8sbCFIOMnJi7YjCWzQCwb1P/E080DnMs+2rLc+
nDPempmV9fMgQaSW0Aa0gyxnkkY8sLwsn46HJ6oTAF2BcTRHdtrqnYuOi0G5guM7
qKWHaT9puneDa4+iKbfbsDq+AodmvpPzdu/0Lgmpisi5aHXVo3fsVBMxfEExlpws
5+DUcqXcTNY5QRzVUoSGFa2qyR/LOc2wOwf+Y7UF6M/3sbAiWTewdsuh9p4MrCAw
0aBcGvhGRn66khn1eqiK1oWHYCwp3//ItToaxgnEKG/zrv+erOSzUKGaNRzE8y6Z
RLMwKezVOqPwg1YOLCip3VYj+Hk0RZMLORcmSN1emAKqXtF55hrr9G+WAtJQWHhB
+r5f7YZYNIRr57NSEw10ny9ODIhUDk5Hse0VJ8MLiK4RY4BEdmWVprYFeh8mDZAa
EhA6DmhKGFHbMQb8acw+ZlJ7K7dw8NHG98jx+6cTuYmXDi6hQdgy/OZ6hYHzhBqp
7sD6VVAFR0x1CrNHMsmq7vEbJp4sU4JvgjNKbe33UY75DOMqgUJ3xBT2QgKnPGPX
8V0A3FsBSpIbkU8eysA3f7UKPErD59j9tPC5G49lV7pk0xGC1wf/tVNc6haGwoen
AtHaKVNhZNeRTUqg9IhOuzCv4PNvDQImkYp3It8MOIwTiuH777/BkCLtdNQ6niv/
DrRob1tK1AhNtmEA2k39plQNJ3s8JX8WWKQQSww5kkiWfCWgGC4Aa2tvEqCKnD+t
qT+BYMb6hr8VxegIFvuKjSNO6u3ObiouBhXQi0nkkFiIsExbO6tu0GhDEa7Qesz2
klTrBc4JzRD9bzlzmdyhW/LiwXrtjvn/l7eANFlr21yhhU8HtlyVcapblYH9dA/P
zfZTCbrI2FRcJzvUHO1yyOiE6rF5UGZYkKvlsAxUZpG48Txt7olA+BrpMMPBhgec
6ptnGvrvBsBsDeW3Nze3lyUuIAhlBEElqwi1TofZ1BqAxU1QHr6Xe/eioVSuDvB7
6Q5qGovMMFw4hKildAic5Rhi3h0TqNVgwmqo/Wqt0NvRBehUj2NFzOaa2b6b+BvZ
DvxeJKcXCCuqBI3soLMY3nPs1ZvnMH/BVFOK50G0gLg1RbCdHFt5QzR8X/cy6RHH
KjSxHnBgjCd0Isn010Unklscob2jY+3qWxJF+DiUebU6zKskDLffHMx/RESFgpte
yT3XCOOa7o4z0Vy6SFZPbPg5TCaRajkNjFFp4SzbO7ovWq2t0OTeLErifm7zWhnY
4faZZW/x6lbwGaA9wsqClhyD2e1KedyTPu6KkQrxKftMyrtd7xf5ifC29ixiLTrq
roteLg1BIJlftk9iKSqlMFDMFE3DVsqksuvSkKe9nmAQVqCRLBoQKTvcW7JgOtyv
AfnpoderB25KXMN1ueBUwW7tp+F7WfzsDWh4LYYj6mQ0eG845DjmMdJVr7wKE2O8
m7YDY4I1qYfK+OKWwoLOziqBgPm540Sf1l40bkB2XbV0JKNZd8jz8v/foJ3S8XDG
CWYX/3w7Gm67ZIvqVJL5Lp12iIUbgx9X3Ig0GHvrtEQBIp2Fg/osaixiQlIL1jeZ
rjJFh5X+r8aNAcTXzyH+66MLrtvnFVDizeNstOej2mlWFpcRLCac6v+lPE6NOz8A
LiGX1OArRJXKe1IjVs4fMySBgMD5Qnt4fxMU/cxp3L1DsHNl9a9AdPMGBMltWWmL
ybQ2RZEy6jMMuZZEI/cL/+8Tz6Ia4dX0kimYuXIakbGe6ucEN91U0j5x9uOvkG85
XWhT1w39//t1kZz6hGL2pTR2UAjzuF5AVzkaibPFU6vS45UR+SqeqNd/Lf6YxFhC
8AUlRpaqN9powJLukylRmjYROPNN1oezu2DxKbwQfWBbjf1fuD/UXxsBsa6PrAk7
GigyesJWoAH/8Jb5b2h2Jl3X6DFjcacshLYt3/EQpbn71A6rM/h8Knro2eiHP9Ku
y4Cn+ITB5E8l98uGr2iQ3e5rRzWcwAQhvBd8FMM0TsBKCKW5/T4xpv7b3wcJefyv
2yedGYzQCh9vJ8aJHJFYRaUw4M+R8BbEaNNqeLwr++sPLdih9iTt+w09qSh+wF6C
fcelzMjYCQThpaICvdJFGrABfjjy1aQmfDvgkVMx1RP6rEEEb6N0pVJa6ISlf0+H
qZ7jtoJYjpXRB+opzLq0M3AN13yxygN/ToSd+8E4gW6vSza8BZMOkiU7ynIGwz7c
tpAQusqKEwKsvVCAWNGsJnm/a99MDHCGXmSvbgkI/yOJVv+NoN/aBtULy4lMEmI0
GCh7Q+y39AMe1GouZrDFHRVeDBvMFssZNLi5X87uBOBgfvkTSU83vEE3NVQv9RGE
/hetrGN7ygh+B05xVyW+/4R9pz8kDk1ptOv3jdLE/+GNYy/UVSCwKvMhkBULRsLN
tjV2uQVLaBDpmqvyXBQB3btmI0bwIkJmJlO1RkTzOjPjeMN8Zsp0iGZEhUrj8Pwc
i52N56kKjn4eb7vCCf6oSuU8Er4ss831NuxOmR/m9q027aOZMssyjOAfVgA859LZ
2rXjPytSAxHBgDlTDYAhA+ikmPiLZazkxJHKpMeKWiqchHe6q/+o39ZoqYOf31X6
4spVmhzjPlqJSwKy8O4nnSrKfcu97Zj6pR/Ng3+nqOqhSfVPrJ15lfbEXkxDEKry
HgMs4vuaz93UpRVbxHBt0tL5f7E83UE236leQNJrsjIbUD9S7cbfxHKrYaGIWqGk
5anaSJFr21+dUY+zeoIWyDw62v1IdWLKie+32/R/MJ3cR2qoU3BuKt2wUdjpn6Ws
gvDK8POfb11NFEWSBNamCVNaMXxUHMMiG1etM841qUBPc3jEdflzbLOcsNhfYsFY
sxxxOPrdiYgG/sNAXOZ18PQkhsAQAhcSxfUvCD+lwKe26k6ixVmL7iHT8FRRIVwK
jpULo3r0Dql4If5OA5tSHYxB0ss2T81OqHC4EROBO2qamzm1FnZs9KtZYinIIofA
McPDDnhb7xc9PMpcx1lEe52CfBpvmrQRJiLs0Tw729281brpsZagWpRDp9S9xKOW
EYRVN8o09NpglV6sFSKPlSmEubh6VEKiRDOURqHYria5Z8N+GymYqjRXskRvIOQv
sYsZclVJnLmogWigVw8SD70FlFfBkg4bKybW4WR/4uvmc4YxJ4Qh4w9mPbCDzVmM
PrYG3YY4lbBuSX/RrbohQoLUb45ULOccIY4WzfgTjtUJDXADyJ3JZLGJzpcbq+g4
7RjTBVTSs+j6hJ2TZAPuDwDfpnAxULgsOCiiyGoRYWFo4WAVX/G3CfMtXawpKSjl
pv+NwwPnw7Uw1Q6Tn19AMwTk4ql+NMGWuXl85i24+Aw4P+QNgRRLkc6MAKHbgm2e
mOuI9vTvOg8Qgd7pKC6EFypq3TAuRcnj9US4X7Fo173/zaRL6U3d76WZJKY66aFo
cbxEfI2Np02ghpJJ1XrFQ8XSBxqJgXjUR1jFJWgNgu859Aun6LZu/bxagSmeEcL8
CgfotH4sI0eBqD77IGGqjTKoRF8I9ZFpb4SksmMdEjAJaidK5hSIS0febbGCDDaH
g50hM5ABaRjxoRb8da1fn30Gpr2iTInJCyda9247S7Qm8M3hLZdePYW1kkrZCkJ0
q7bxQ2/oNM6FnetcDoKNgaKiBMkMkvvz7Ab5Y7CJVUjW4ECCxLQb40cxv8Tu3Vlx
lyqCEoDLrlMch5Ij55P/oFQ9w9ht9WjYhWaRESHMhWbk1lpoRHZ6VkHwL7LV2lOI
VdI+iwJjJSVFFdSLicWkmZqqArbvmtby8N3mkZclKhqNVLEppkWXOMR1Znv8yAyy
vRtnYZaqh/DhmfjJ1UGhGB2mwdCjRje49gOPLte2CMFyxAaiDYcqaU+KeifvwUjW
yyg5SWVhWbf9t/6SswK0FgxHT3a6yBy5ioYiWIaHSV5ZK8wWxm/daoGpnbTTfQsI
fiM4uEwJUj9MlJD+RcEqQcSMwdZ4MkNC9QYjG0gRsEx6L0wpNeNfCW3gcWA9iRfS
8U8ikpe0KC2+hWy4fiZl/oaAkSrKGUqGZiscKQAZ7rkUbr8wxjeuqLZtf9G1GDBN
DDrPBtfxlW1W/WBCrfEBwNS0x34ruNvA5ELYKaVZyeGaEhhHGBc4FOLFiaAM1D8D
nBeJYDR1+XTlp8RHLTN1Un7HIln3oLtrtONA4rDbMRhQdW+D5/465P+XLlxeEiDl
mjWsQOCqdZ4MX2Vc4mXH2r1aCoIBkD770zBvDK/9cHHAauJJYB2U8/p3bNQQHhIs
wJBS0wuUhj7R3kyMK+Rz72DTqtK0nXi2GxRGZFRDqw6dkKseyH1YiCvZV4VWJkX3
QwwPmU291hbt2afy0F3rz/U/z63blTCHnx3gsWvQw9gKF2EuqkZ7VWbtt7Tk3/Kb
ZEmEzJ++GuxdLgtBzNwC6U9//K03c9M9lOEKqsKpNESk/YLot2lUNKKjRA2L6sRJ
8nwHnMGvVvC3D17hFoGSS8bbHLvKAHkKahkI7NfQ9NZIiac5CMqflnBTsIRjejsS
fVYctXGt9a5k2DTRHOUamltTf7oNYs0PfPzQdxZYDrsP1iB/xXyMf1rQOQ9pZGhK
MjqqVu23fcmveV36PQYqGXcPvKhO0iV7g706RkG2yLP/p9RwwiF4HIuIXhn3bELb
Ug6esC7YUNMtnFjtR9CPyYhS41klgrDtJFdlyIvXZbVvcn46f+cWc6xw/TiVtdbL
xNTygpCenUWvQx+Gol29Mg1SFBgwfp4HZXHpfNirYqX/u9PO2ZDtTTWlgS6J/tZo
NuyB+4g+JDX/o5uM3LQuRKDRPCD1YO2YfGYBS5Znz9wcQZ6Os6o9W6v/pUchAnT+
JeJCB5fq8zYKMSbrsCGm61Tk46+6ZbMDkuofsm12D9/IJJytzVSgEmPBsfxQJBWJ
qbiv3Pz0bX0gQSUWQUKOj/SVGzXaz9ownHBdBo0popf6nUggkZNBUCL/NMDFwO1Y
Mp+fAoQ/FLlPH4btyQCD5pRwpFIDMOYQ0x6UMQAa7hQOCFf3wBADN+t0+IgegDDJ
I8M+9Nh81tVgGff6gsM77YW5VHjq5nBe+I9wAIHEFB7NJHc1Vl8+D9sSfiGv8XOg
pHoxPpj7Uxaxd+LtpZ+tVu1alhYMnesMeUsrk+/uiSZ2WkAihr4laLCUYEP7vo7p
pT//ZU8JQpIwCMaCbyxTcllb+aBRCcyJ3pnro+ERGb/SCATAdaITXH6nLtkqVvyM
oJoJN7Fr4wstdEMKSzgh2wgFeu03IEFhS3/X3/XAWMyTX6OS6L69MZBIwWUDpYdp
FrFr4SOZ61OWP/zAb8ixCb1ft5F7nQVuGU23Ogb1BVl1BDIrhMFlNrdQiMNjrz9f
1uA82QffuDYe53cIHvz9Du9pszf9S7ILt4IKoluPtgvRj5UoAGuCp2mUywTvDA6z
FtiKJ/2SPz5UBEmw8GHklX/HmsxWAS9JVnGIN2zQxAHY2rjnEZ/NkiYqaNYYLIgQ
k9FPiTC4p4bWGf4m2GSlsOltcX4T7MC7jA0GXP3Km3TrprQ7S5v49Yy8xybEHOF3
i7rg+sAfQNUkK22QhpBzIuHbvCQStQuR8thaUm4/yWK3VH7cJ4vU7iGzeHRfxSbW
ANgBfc8k/Y3TaCJw0j2eOKB19a0Q7wY3bc7qWpZ433vg3dqaz9b7zNRzwX1IHe3i
JMQlfftY/yIfLcIY+DBWVj4zZdHw0JdiOKk2ywUJTM2Wwen9GcPFV5tfX65iOVc/
POgu61++RCwZ99wGoW5zX9S15cJAtdFADEplHQEzciPELbOoWmhpxqhUulJTZro+
n3hLjqob7psnUeiI8PPRS0DTbgNcdxloeXE1/sg/yNouivimDrFM6wkelqprE7wv
CY7hUYcxIOci8L615zHm7cSXUx2rBccQJdVmlbm5jKCsBNnDcyfKILkICwWrkpXn
U3H6x9cczlHLsp1rK7WfDDTOc+4+mVGAspBj+nc/CB9MNqMBYB0ha7mqNhAu/jrT
E3sITC3a0J+NfA5KWIo3TtX567BY5jJoFsD2v3e8nCqLogByMbS3M55tm3EaNFrs
dxs/7vG1lhGIGPswALX9C969DjzMMAUij4FNyJ5LaoqGrgNGS7Ddtxq09fzkRSeL
/rDmrr1M3p64/Rkw5UMHBEaEuWuVqm+ve56mnusQw2RAY+Z8gcgRhMBkoQLlxuTR
Z3FdZe2OT/FPyz3UrDTovL7ZpsUcBRn8sXZBLQG3S2EpGefjQ9GjQ+qD4gVUKd/F
QKc3vIsY+RkDbg8QBy2PvOLnDKbz+v4HUnPSuH0SJR3FCrrJzOM0Trzcctpq4NaZ
1OHcAWYGIW/G6dljuducTbxyNWXaie+gGyRFY6y+hyTazR4uwI8gA/od1ptKzAeN
xeABYnXgunG0xN9efIoDJ0INBs5F1mw38zJwk1ZHl+nzBAbhiYfK9AD4/Xc2RFAM
WeNdnBZDgYcDVntCFG0v85C6sna04TsOtwGEVs1xMGrvOUJsNfp/4lNdmPsh6/iI
A8GQhX1HH4jSyE1ETnigQQtq5dSHlF3McBGFup7Vcap4cQgg0t+/36Vhou8Wljnj
pypIr/+Q56tqR/mpkk0VfIdEXZ1WjbuGpPIQWoOZC8JciJcLzxuZ9CbUcFRMsAiS
LY4kq55Khdq5vm6VhiymFqTFVduHswg6qEHwdRnlrsQhwUKK2KBbDA4sXgDNfXKN
De+VjKKLNpT7lUjFpXts5cY+GOxGiuY1Jj6Xc04WTbGWDwG1XEG8NXyskHTXCimP
xqDQWFk7qY6dyAAl7zMMrc68iX3r/jviG1doA99+kh5omT/ZmR4Rz2lYvZ+/QFzK
swBTCtztgDwWQRuIkkg9Bob6U0GN2B0J0G7xeD6cNgiD9WKWlvbrtEtyUmb8DAO/
pf6xX6zNL3yEB5vIus6DiSM0c3542zVzc9DFKhRC6KzsaEOgPa0yBymfdHLY/1Ed
puDVRjN5RhZuZq7TAlfcotbzemRwaom+ithSjIvcV3w85/NACupC4tA95ZAIujiI
ReWVnzyP6b0WluhakPpWikYS6UTzUZvyNPy53bR14PTlqaJ9js1btU35L4LDXuzs
omxItQ2k9/w0QvPyFUn2jqp/HST/Cjd2y8CqYoSOUhxaaFZmQbbdpzN+W9M0QYi2
q+LxhnX0vtlTPzfHUdjhirDRI14bNrHxZJ1bXuOKoNuKkUjVax/VW+3SIhwLg3Nt
c9ltFWWOBChtEHdvzj8AMVumJJZ4i+TOxCSAiUBge6EnpY6p5NCH3jeXd4QBzg2x
JkkTlfQZh5oEOYlR4DUyIVLgFQQmS+gLeZxHplq64wCOak5BJLCDzsAoGnXIqJUc
9SbaVO8r218NHo29DDhhD5EyZk5dhECNpv7idEmRIEa0oinzC+Isaiz481Ee1e3j
VCfC0IkIWBIzj8Z+dH4wyQlTNQuPof+Vd31cZHARkHfc2n4FXmCtyWe+366ITdAl
Ig3AwlyYhi0uhAre9XVt3lhFPCpLkc5EjcezECH/Zl17AVOluWwORujytSBkzuAl
77Rcq/sjROv9p1o2GedHktbjL72wqsQOO+1+B7brWN8StBCezvIGUoLoIwMyjMSR
M1hXJCCZeB+QkKzrS5gGX6SsnH10abVOhIXc5/JpaawhIEFkfHSPmA8+a5J6fuxX
iJRyiCoID5cok/XbHPm9FSjyjJiCINXTgixsuValejI9qY7KuXzn/qSSBEMgHWYn
mpCnD1X9aExrkse9XA5mpiKemu2JD2HZ581d6msQTm0W5tGG24WJZGRu9XO5YIkF
AfdFs9X8MWQF6woX0tGUvnhwViY6XwIBMD4x7ybyCzQbVuBHHc4djMzqPbfG4j6j
v/f7LH99yQMc9C3xciwEBxOkLSoU8Rviq3FZtp9YqhFVvWwZRrTrcn9Z9yIAZW1s
CvbKkk0Cj81vu8VQYS+7hshn0EjhzIVH4KyimVaODUccirtUkQBeXWH3KlCcd6JM
3Q1BTeStzlNdcpo1pi5rUH3bl94+msk68ATAsGHDNupxUQjv5+lACybYP6cYU66S
u87qyBfi8r6gOXThkxupzWe2dbJ4wy2YkL+CMGATi4aU99IpSQWEZQlANUbWSVdE
/MejOcT1B6NlyKXsqJGSeodCyNLVX7npg7tPpnj6Av89nvEitjKOqDPFMULQn2fX
BaAxR3cuuDz9RfT7xs9kyJOcn91eJmCo4tcgUwbtiLroNHYahpEaZPNiBRkXO7pd
2X/vbZlUf7HzTCkNw6WVPdpBJ6KFPMUYgBeoVqQ68TnlPK6QP+4+WOuh3LPb70DH
SicDdr3Ntq6t2udg9YlVL4CujJbL3nurjlRuNfvxPKs77LNpJQVNfFzD5YPs7+Vk
K1Whwp0CNEOd87uHjiFngxM9eXlvSK/skdUS5NqRs8GBzmgPBZ3mfmju60CNJEUo
bWY8/B+r1rROZsQuTXoyUCStGmUyz9Yu1T1zczoDpFEZi3drpSGFgINOentN11lj
Grtbzk4R8dFxaKzZLTqPin271KtdRzDQdye9lcgiX9rCyICcOBB/tcYNF3Yap+Vc
gG/Z4JPk1oWUHSoATaNabGK9Z46zqPlXYQPsKAw303goP+GLcWDTkdi98ax7lMKI
Au1nb4p71c2DJqZXorJhJkEGWrxIu07X1QsxugCwHeRpI5onPSMFf2gPlcr5U5dB
NO9yxCpQdLIlSzQPUKNEviVGfs6gZYvInzFGzvPDNmbWHxPmWbWoJxDCKJIgOpoe
CoTuL4KulJd5e6QE/nYNTiYuaInclJFuBlRCpLOIjGU7mjcqzUI4yPyiLPSAnv5q
Er6UkXQnDKlLQ8mp3/nIssBijdl3otw77h1RV05Sgy7M0F9QRGFQR1JP7zPkgYwf
7FQmGaq2QPZD37rByHyIVClkpq2zgZoBqZArxamWtrgcGu5S8fOUagcNbDnuVzwp
1YacIZdOT3vgbPqHOTxOKcsnFueOpVZdSIbtm919e9EcIZLcKVB6Z5DXmaQQva/t
1z0VWkGr77ebWHdsb+WNGlayNxVQuL4pEBBu4jzjUSGVy0tDPS2VqFuCqf8RaSIJ
bQorbWaG305ur+rSUns4ws41zGflnbhVvki6f8QFHncEACFGYTiK7hfP/IhSL2mt
ohRSEHPmCDPN6jxUOw4voO0AcO9S+/97OqqcfCUMlbJSuGTRyMSUmoOUBXOV4QHh
c/TnH1TEKYTT80g+vcpl/AtEbarQdoLuKMEPpOQFzLpG5af9O/rHGELuiC4+Yy0W
xCbeoG38VYn+14/CLDJnpPYV7WtoEzkh9pzfModAhjfpeL2ycnUDBOmBl1j6wvEo
4bR+4GM4n1JJLlTajt5VU9x+8L+h+sBCjaq0VbyWJh457MKOkdEt0RTr9OpmSJEL
DaAOYAUn5nv3Uz8vsGwC8eg5pYTnoXKpCVEfiRt7+9Y0X9VHTGdxCuXC8PozH2Sa
gsIHBuVB94z2RZwe4TU4NiA9MDgjzec4NNU68n6q2REI66Zd7UI9K2h68mn1BVgt
VAZ/i6KzCh3EN12mgXsWQZvnVwgC2/xEtQbACJQkmr265zDrxJDUAPXpY5sGOb8k
CMu/1iXQzAwSLWhOYGm3S8wjiK1Ew4Txh3nD52rszLBQVi++C2fsK/9/B/TlfWEL
TFfYzQ+wLIQ3qo0UmMWWO3MoC44BL1jp25YwAERBEEBkuZqi8hEOYTnERyI8AeOm
LUyFadNoV+06zehvGNW7ppaRsZBMjz5sz56eQJTZT/klJGxQRDiEoKKiGU32HUUQ
eQZIn0hC0BcepjXCN923YuN7yDOYYFaCEZMItBLwRnqviukatA7oB5oTWscYo3Y0
qzZBAGVeisyCS5LT7ZNERw8+EYcw+SYxgj5E+kcg3gY1wZJ4CS81qyGJe9LzIvHV
IXZAqJgch4+Iv8pY/3qUqI/PlvqEoEXJTvb8msCcCzNc2wQpgbzpThiEryCT5l1X
hKb/GUl7cO6h0+lwK6ERas400bddSWaqDoEC8yev9rskN3Uy/zEyRLuD2gh4O2/8
92Rb/BTjv1EI8LiXodonBbhG0SI/N2yje2Y+4QLBIfQYGBkFH8YUMEsqwTInzVD8
nqAQ6nCt3lHnU0ZgzS+6gcfneqb1TRq0Y+POX7UtXob5L7VJImr3x8oqWzd+7IsD
5tu2SrVnSDj2MwQowAmaQAXLv+jU28uQpDcnX1/wZ5wPcFyT0obRjGz5qAmr4OBh
dn1IEPe//n4Z7NVrlWL6ShLQinDKwLU6wNfXUA6XAHfHy8XdV+3oQS8HKhiaKqap
QAKJ3GQ7kOMehBEFFrf86Dsh1MRBeEbHHK4N1T+XicfvvzZTCz/8xgxqEIedpmmb
eQrsA9WWq955eNbpCp4ZmrSwR/y8BGa2IOlWqFkzK9dzP/38FK9TVfczY4i6Er1k
HRu4fD+d4LDdiH3Ory3nZj3ZOBTWfT2FAV+t4+W9XLeNz7gXah+YquRQlmLGJ4J9
knXruP+Gn2GM2q334Cg1U9Cf/bBXljNG2ibJpeYdVT3EDOsHYX/bZ3KfWcVmP1ZJ
/JZ42X1NbkUbYUmmYker4yP0dlEMcsIZT1j7a1YWt0By99CC40yQ9vqELjDKul/6
ARZ9EwR32JeDcpfAabXNgE8+znHAtiWBZTk11AsvsVR8Ca6fuZ5yWJm30/EKaFjm
PO5reMUqSohk2XEHivfLS9TTeqbUMuYbbebcZ/RLjdIAtWG7d7taLt5BhMxIC5kO
6IDDFI67b3UYh1gsZ8BJRXD97xrV8WK7IwTGv9edyNybQQy+258yDpV5fO2fw7Os
guo3VYGg+6yDngZHzkA9bGIGHyEEauBky3oxv6eLLPO1nrSK0k5prHKfTphs9A9c
YYQHXoTsW4ghL3usEIVJPj5vrdcS52DZjGF2BkYwQclzBpgeDnG+IrwEniqhlKh5
M87lyXIEFhUoIh+xJeXiR960oFueuLBknTKbuS7cCe4JGFh8o8JDD8GfSzdb33C1
DBFaQyjpL/NB9F8l8UIZZknWQraJI0VZnnokiWpt2rYuBYndVjtZnEZ0PE+k78o2
emqxKgaz+yhd3NDCLCWXWZsa7RBXsSQJwmVZdXBI2BLCAeMDoC+5eJM61eQd4CIl
R0HxRxU8hPj9SKwEHG+kl+UydmQKcSDcTnAISQnEz+ZKg6GVdomQIrNBpNQmd4zF
0piujUygFBDwX0XGfQ0D3HK4YPB0qnf5NpTEJfckUZXrEMb6AdU/oDCi4NK0sbBE
WX/6dDl/TO4XsbuDHlWrVSSC5I73W1SpTGX2OE2Pve6Cq99vsfBAYiyX+4Kck4JV
rvLafn/MBoGWKMFkgfMaNQ1xIl8/3zo4u0ctZwSDBIaFf9Ry/eiZ5HRQRs6Q36vd
ic/OJyiQkXDStsr+JKF226iYY5K6sDW6WYEZG2Jq9EHUuSB24EhDa7ClI83k7quJ
ATtOZD6f15JdEVwDfrpVlGjYa/CO37Q3bm9CCIOWgkqnYwx918Da3NdZurTiv9rM
s5s4kakPsMyiVSvfBJoyCZ+EK5V0WCD/qaoTmc0yYGv0UReIxnmxeAtW+SxPCahm
SdKk+7QtSThmFsWsD7pZccumj3nGRhs5QvkzRZDGFex6nWLEIrUqCX2Xum2nVxRw
oqCoaviXyyXxAzv4AaqyRTFRzBtLEfoSoWVmP66QhjlVlO5JO138uXw9sNDQ09e2
ClQIfg/43mhA/43hSvkb5gzaBIXjP5/5kL4SC+Dg6ywnrYkiLWCMDz4Mp1lbHjxl
kDoM4RPSsnO+5EN0e9TqFVbSxJxXqqEEDEYDr0LOOdkCklux1K8DB7/qFEek/7c9
McAs4BQYuIhhpD8xZPqGvkRnWQ4GaYM+2imrzftdrUv4N3kCsfiULgJs8yWsH/3C
zSxiAigDIerb569EgBQjuwK5du+aKU8jaA18nuRKp/ZL8k4a6lYC8WUJ6OeyEptD
xk7hZPZPQu1zk2FUPgNam4pLMy74gGT1vv5HDxEBma4PEYUHcDqQQ9RnWwW6xwu5
F3ynDZbGgWw/5J17M930buypaFNSfh8h2C9vILRYjOjfymeqi1ugYjZN/ikqsdpG
wD2w5T7L8L7vn33rojsQoND5NlQE4bY5MoEeTeQLOiI/ZQMUpd9JmmZL24wSVA9a
W8xwnUXTJ/+rinBlqo4tfQX52LAr0Bt9rPiqqGDtdks1LAdEisizjWTmJH4Ht8IS
YQ0McLUIrU93y0zJ0rvVzt7WzxKBpghi/ymHXGXUWwaLKFtncAESgVKgLgal1EHr
6jNkR6acOEV9LQOxMS5rWZRU4+in81XtooED2mV4DLR+7WS83hDZnGi4drjklDTk
ylqUcp9BdpYL50u9k+7jNAWbymRV/U6vcBQmKgtG5YS+eNUDmNwshNKBm9CYULmC
hL1Z2rgJUywAqNSagLtAnfj1AkMcg9EzpLy0qBjLCYDSRT9pm4hD/ltr3ibvK9Ha
2jEyFuD6ndlF8JzsvS+Zr0vs7byRIGd5iFnSRhxJRlZYFzoaeuye/8w9w8ScGT6u
MjMQxvxojOHLAW+fSYmnKJuu21bXbpWaTEvRoM2iP5+6+9AEbLEvXhEkgQU2w1tp
NrgGljVw4Z6Ct1+8oQJ9SW6qKaiAYdDh2m/6I+VgXPIWibOX5Csn5NENKpXTokZq
66eSHyzlLKGBY1C82I5E4MCZU2c90kPyUKHmUY4GSEYqX/Lu9C3vmuFzy35TUrLa
jgC3pUM2CaRZoy+CVaCRV4hF/CpTPReftW4xmC6T/V/PmFjybdW+FUYifSpAPRl4
UPvCCVIEY3b0Zn5B6VgZOvWroV/3Sch0A5Nre7EBvDpdQIJH8D23MbQbXDSOZw3K
pjzuqjZaV58JviSqqgUZqEPb2Dt5PBPawRIi/7tQbxIG0KTwGy5p12vTsEku4tgs
BOhdQljrK6sUPd9685a5RgzHgQpzHO3hVhptB6dqK+eDgvfTt9KkbmQALuKCovME
CpAklw9JtsT4xuKK/AmJC90hpuAKaL64YbAZfih2I73WZlnIv/MCdlMquLsV5MOg
00EhrYFDI9q1Jn3qJZfgd9aXE9uCA9S7hoXOUj2eootZ3DCPY4XoGz6ocTyge9FX
3yh3/LFvWVOPjAhWTpwti5griPbpWdeExILgPmmZoWF++YfLZ9DtQcy5J8sjU1as
UIHmK6YnwZVo0uZ+J/N7jSVzHY7fn/buloKpV26CiJD88FG7+Q9FYOnsUN1/XQuD
CkjRtJcln+cKhTZ0B3/92DwLQlvY/zF0fSOAjEuut5Wnw+i4Fgwv0iPFxaPJmV7K
tbWq/c/nbXMpM8Zkip0WiDq6n+Sw7NVYB+a1gSnbAL/YmrnyrYe+2T/mDoYQgm5o
jjD/ywVw12Kknh2eaxKuTw1s2RnUHq4JGYxphP+a6J9BxBZu7ojTgxKA5zxysxJY
vmmstNo/RDrQ66TCfOcDuv9lj7KfepwAC7isV6mjDu8OFi4IpCJfqdgnVBz/fUkH
Uk8Gf+ebRPw0vOwpivLiV0AaWxCQPn3uzFWu9+REZj3yoHli/LhfBtxL9eIAqmzi
U1vhmrKRYqzMilHwo135Br5e9WktR+jSQX1d9ee2Y/yLTho/X45dK0o9hiz7CVO7
++iy+cV8XigpIGNqZWTX2hk61gZIQlt2Mio+TH391s5JbKDBWJ1rYFFk1Qj7Ba3P
c6ni4W7cKMjDyu/Hn229ji8FPX76VFeVMzowUkS1BJeKncGlwd5BGZ24IAx3cTon
I2FwQ1VvYF2wC0/6ddX2RDmrA1j9YtffZQpZa+MjxVYhSb1N/+8COAH65SFIvXY6
WWyJeO6g4wC06XsclxHeGh40h8AjSWkp3+c7XsNI8htYmW9WhLTSOza6jH1jorUe
PPiWMiwCDPJPM1uytOblsCTR1t/76XFv/+OfxF+A/Hw7TBP0KIfZi45Cl17Dx/wn
T7nJnTeFn/40JZuSOMiRv7qWs2mnHM0HF/HP90AycEdZHalvGIJtqBcVyUfI9Gvr
ANYXTPjbfsRwtalLo1tOf9dmWOu0h4gbSCbXuNnNnWenVMYybghWUQBGPcclPpwm
tKEBbo6rJWdKVSFQuj12dVX4BlF4CFbwrR53+sRbVTay5vjC2vteIBJ4Le6ORt5X
UYW6DCiYEwRsFFYexdc9eYeurF2i8VDaBG3pA5jr4oW0GxuCkBtzwhGZj8E64272
giUrLodex8vIu59fG5rxL+Du9MBXBD6zh4vAjtfvv6D17Nlk8Fi8Cb8sYJYLPy92
LAYJHi8Vlz0ypjtPu4w1bT8WEbBR4Ee5RKz1xfNZZjyPaq3gL8uP+jA/UojumhPJ
WYzd7dPUOZuSvDFmKgmkPLUyOXqtxmW3teiMSuRcgOpMsYeUxmA4OiAWwpAlaONV
MMuhdgCwv9v0Q3OvvapGlWRVLTlQXqDjSpDm9DFYm4vuCG955n243NYs0SilHw6c
o1/q5FNrHrIwnvLKXJSZWUTKjvagdUjd4Wwzs4PTCizqcOcnM8LNXBU1Lc/qRHJp
Kezv0f/+7omyPeoIb6Ap5+RBHnla1/Zuz8uHuJsHXIS4zCm0DjESta4ydDeH5Yzy
4cQMIidZCdZ3oc0y5cgNIY0yaaCrVBGfCgG6PmpmUeEigcb2H//+Uj7cRyMIMnvi
zCaVxMoVQ+5NWzRRIls0iAlaSwPeWYSyw2/XtCmnO5LHJS4OWCTCoUCyTgo+yQZj
jtnFwzcrydL5RnW2VhX6VMwd5E0pQGlcX4siyg+YFOzMRKmkFPUYNXLt6Xsc6UJT
GXOaAFKWNHDS4/bvr1J3mrS9Ms/JK4egOgwGjzL/rrJ4p/nOk/ctz61bqfxmlNTj
aWfKOOKF078y6tr1ryEwCxjlh3inwzwNHOd8evQinLybhMAcA+0RGkj09s6MaSoD
otI9M0fu46H6dfVxWbDoyXcbOeRT7f5MCnVrqYsoTt+Wp8mOPz6CXUH3FphQ0epg
9UmXY5YpaWr+ijgbT1A6iB1wwOJKpsfdHmoN9e53LXA+/gAJL3rpS0o9CPj0ONcb
frvsjvu94DUUZzm8+5I/514NJQ2DTiYP39jJgO3oYY9WMuIaN4NuklBeDpzjmpMc
sOp06ouuo6zNcOXpyspAJNANfbDUafV/rPJPgpoFE/QwbeOSDordYbp+avEMrhL2
HRHkIVRFuidIICdmKRZZ0BEA9srJXTjfRXAd0NUbhJ+p3/5HbWT6IF/q0edasGP7
NirUDWYc9xP7nU9kzaK7KlJNelu5E8GG1az4a7Hzm2dywCeI4MDkFC0Jzpid80yy
ubjWjj73Sq1LGSdUVPMs5C/4wFLmn1DpEconD45ULyg494ilPtM32HFoyT80lu8x
O2mZIcadBg796cST5fqbMslTv4JBNP+n3sfbWxGcCsAhJdiwotObRO/YjTnNLEKR
of1pqm8msJUC6zWo+EBL2+QgcqCHj/R7seRnmhDqwFNqm6tl0Vw/KjUOirhIwaS9
mfN/c5SfL3J0PwF0o8RmDGu4/pVt3da0/RqRzAjeB2A1eSFGHQtYbyI5dv98a2z7
vDrWPtb1Ihfed8z8Q0sz5hocH7V5f9W7LWyF1xvoMF81DvUIHlajNnBCjliaDaoH
eQdQBPpvKO/xiDjdT9tltNr1TRwwaagPghYIqxzuude/lDXVZzTmIzVqPU3QUpki
SHiz3LxsgdnQMp0rhV9y3T2IrKhgIHWn0Z7zoYuxBzhBq3s2GalwnMksUL5w9twt
jIcumAV/uoX6+9il6Z9H495ndxIvDurLtKtHXau/FuA7JBXCo30Yd4Ruli5omOAx
KNqN1SKtlECNZbtVzFp9NRCQk4wQjTF00TumUt2H+fets3xAXUsRZZcBdM241/fw
1JwZlAlIV/gPAiQsUbEBTV3QDPqWyVf2R1Z6TUiTnbeoak1nBRcz4ylIWNJI9iIP
n7PEAujULegp2sGMw+cn4IaVnZE3WBD3/ByE4VQd/IBA7YI9hxmkPQNPZvZ8kA4c
hIhh0R9Kbpulb0NVk3wqaHI/HMXcOIcvdeYreDR39P/3y1c3paK2+HQY6a6ytW3w
FkK2RhqYs3Urd8pS2gXQBt9Vijrs5xwHHBunaFSLxt8BLDkn9gWfbpjT5Rgkzr6D
M71MjSre8CMOyzgtLCtTLtHMKl08208MN70C6C97kHAaCAa8UO1UoVEGaOhgtkyK
nAGDaLriJR65K0oVEtZvN8Ini1bRiNRru9YFqyq1uV/2t/DVIMsEuZKTj2u71U3n
naJw4N0RuHp/2cISmobQF07aH8fwbUgtxLXgJlClHFUkNwbVE5AUibHkixOrDKUU
8Eg0/s75wOD9i2keV29tLd6PsfRNj8YxnrBqNDNIclyP8FQJuQxS4gO3iCU+jV9B
6v5QMEpU8IGD+Ho3WEco8Ow1WagdFdgV503WPtqChIhcjro1PyYOhyuDKQMZAdsx
oBlCaaGBhUVbaEpJIlTJoM8Ipf5fMHJbLp46Rg0yhoRsgBLZVyR2wwE0lg3dwYiZ
JTi48Ecaxa75ZlSHdAULMPG2Jksj+2YSEi73ixymiFNqEBufp/+t54Be5QbnPdIw
NifbpEW9y+wJRoW0+0zfuMU7fWzf/JnFcUvcv7q3zQRyQCqBqJcjNILAEsuZyic9
d/8QFtI5zUZmT/PLGsDwliy1T2tSqdTvA5/GBVOS1nYPInUSgXQBLDyBcyHCm7kF
PkYByoexQFZf0TfXIrzVg9yG/UdSdqJjEwmlsX9iIcX5A7Upl/ferjucDl8hwzS5
/BeEo317UZtCmVgFwvuIc7ZI1DUoM8wMZKbK42hbr9V+tC7Ot/Ff2d0IMLfIgEf6
ZbtL5cTV6trO/QRIw9NKRQ+KyciFrCRT4c6B7f+/+7eywrpHd9Opti+y9Aeg4Fc1
8e1Mk3V/u7vwczpqM84D71I3LKdt6hqnQwaSZ2TQHKd7CN5pjEZAK3aOklSBo+yk
62uJ02cOrPPzlsNYwrxM/OKzhXVcZUxhvSrL0sxkoTUPGV/lWEtSb5M6aD/R84gQ
SFVKLgq5InATr6qpljVV41OLikkmFSb5AtYbK764a7+KwE51yn9tSBZoiV14xmAe
0ofktoXwDsN8srFFaT7wgLijJB392cX/T5q+3bDf7rrvu5/rk/yl+s/lZD6aOsLj
cy+dWwBTTZjcjzv+SDe7w+fdxkU/fe1TQIV2rn1WcmxZ6Hzkvi00vpsLKVmg31Rk
pqOEeLiFW0aNQNH7qxHoC0NB8zfhmn7PPkvZ9Fm7Tb1jOdIG3dyGtgVjksrMlprH
3hCtJK7OisaM2m32pDJlwPxlYb4vEgvHWWUXAv+0H9rC7N/WhfeRDMzTI62bK9Pq
4X8eNpGipsPUkVpI24FuwnyO+BxUP5SP/o8NZAoT1/TiJJpwUFS5JGiCTb+o73sP
Ji9jftMj3DudaQmEl+Hv8sYhFfL5DL0NS1FZCkqIviv0PANuCNLb00RF7TxEHjKi
sUxJLJIXk2HhtQD8ACDcSplEj3XcX66CozcBsuWbsKbdKZrp73PTNdVVhz4Uz3Yx
kW8v93LydOJ8Wjpl2/zXFLHO7zofi5K+XJbb1SRGGJty1jhVnzqm76owGVICjE2K
UeglogO3WkU6+5X4Tf6IgVswrLqe+/Io9ZjkVJi5FsetCM6gj93TpJkXwXc103AV
Gjew2IC5ExVUDoQ7EknIqRkBXT2XNMsIIpTFORJUCJBSebmxbrQ+v4KOKJOZOwzU
8kOBHTiU/5dFG9TUGpHeZzN+1WTtStnJJHeAKV87VR5RKn4jvmHWoEtg/hgNwX3O
ojpSpvTolqdKA/mp6gYnlZGTdtKsLH3zahd4VhHo8JC4qwLdI/Sib4qatfjMtvi9
a+RT5qWkTPqM1PyEHCugRnWETgtFlMhCTiz/DP2UI37dOD2x5GFvqOi4vIy7XkTw
TQIi8JfhkSV/pmjHjDwqrp8VRLNT5bmGpwSCxzh/1Vjg+6o0PkiYFAxKkdfafB0m
gK/NAAvqZuYm3DCiVTNi4VawgqasIE5somvhhc/JC/daq2AvCInZX1suGK/3tj2U
Gw0wuxDNKkRq5lcVrBIbdUn8ionFyT0dWaSKJpcMnHNVPeS3qGt6vDa5m2hovyIR
LK9aPsQdgSrCAsjIpFZDXmnFXz2qdPowAacl84f32lqexf9FepFUYfXSDfNjsISh
+T/gtZTEgj69eIDuG2kfXCFkpl28wbYgCAMCwCkLZ8FkSs19dGhclPO0yqpDHgS/
DYtKhQ94xMTCPIZvQS06bfE5uNoRjQ0Oi5csA12bD2XqxbyqNvRRgSmFMQSSD1Qi
Tpg445MhjzCuxRMnt/ez45/nLFlf0dfYZK1DcMM3D4TfnnPYsCxLf523oyIX4kIt
Cb9mVqLLbLcj3NAXxl7+zcKW3lgPK9PQZ58ltv3LwJLIKHvhDs4UtEsXhHLS1m0V
Z2zLDcTUDHXBrFk0ePv7vZChEyY54sR8mWk3GRvHF//ec8dRKf31KE+oSmsD0Sax
geBCdUjM1pgWDpEX1Ty49c0EWk0RdaOY8boKp3vTisffAe/0vR9ymouPt3u2yhmF
0M1xgak9Bb7Kynuk4WAWE1Al5uiM3A+dv49ASrxrsoRrhO5hSZziP0dxQZi0QIpJ
A5VPqQW/0Ntv/2PAnmRhyV5O0iyhNwbNX+LUalKm/x+l/NRSb4PJLIszIAYtWpfF
Jn4rjwjYuzcwTt/2RezIjMgEOOoFBhsvxNwOTsm5gpzg4n0UPrC+4lxM2wd30k19
YI7sK/o2h7sNpKK8XLeTm9O+cLvYP3mIc+cvmhErxnleVUtKXQKTdog0N1zbqRsy
MLdWMYWQpj8gCtHiFRPzm/61yax9PQvhNbHwqur8dsaGA1GOeEzVef4QuHMr4UHJ
nYp4vkEbORUtJNZQYChG9w2n8yj+98Ga5cXOYuO7iE1TZXwu8aNZCuTwxC+W0TYX
ihOnCvH61DecbiS86qk7gebdIbB9gVNZ3h2hcDnp2v+kuHQH+CggtHUITBGkaI42
nwm0SCDAJIO8BgbLj5WIb6DVpsuglUE6yE0jKXTuSc53HQXYPjKTU27NayHQEoyz
l4oNy+9YEFt0Nsqs1KBZhTYWMVeXuhsM8smcXfYU0VyhPjOPQ/09ORZSD7o5oxKh
O3+Kf35tBxK1U+VT9a1nRG/8q9kkgXSID6ydyej/1eYtfL7pb4aPdSP83QrySs2K
IFj0Vp/uxy6RhXX7TbaXfaJmHBciQyV6+2b4ILelLBqXEc3SNgqh/0D6plxfHQbe
0ryyzEnYBeNuP1D/IQw/aJKsXMr3eHtZKDBke6Ma0hl1rIyall/UbuLokDTP7jx4
LUbb54+oFJRfr4Nm/DaTPVdNiWZz1rue2j9T6/5bx15a0nyVpNXd31+1Yy211OF3
guPSGKVvnf7AQjXCatnRST3sCIeXPimwy62bhi33fHbMMpja/J0DMX2A0/vAKPIz
97Fg/mD5rhArf3J4bIgpiFlK8/Ejj3rCl4vEhwCT3FWzgvDcujXoJMtpXaFcq/uV
EJgb8wdkX2NFF21w4PZzNr3ioJCduGFIx+tppmYNyghnAUzgG1RXw9spWkEW984H
MmrJQjJP4qOblptXZj9/ksxHn5KXtsUmhpFpe4Pwy54tg1gARSOF0e+AC0zykReV
c0IbaFtkfY8h+Gpw3iSLlN3yF98EWDp9+rt3PjTlGb8oOWahUvJO+BkTXjTrWl/r
V15SXo/inhtd62XreiKbAK0igUTw/wjOVoThO4V/Ybz9nYpxPgfkPcKyDHI2MHZX
Grrru7BUjOH1lOSySWikwM8HbW6LsnzAjyB8Ns+VpLardJz8JwwqeoJOuQPrrTfq
xVbwpmFrtQSwDAQb2hPQDh0i7xBr2LkObs6K5BretegUp0ewm5lV8yUD99SPzxuO
hr0o67droGGG0pfP8fnAQFlVJNkJPXwjA63NB+PksVnLHu2AaaNO/18SYCLur7nG
GrF6GJh2U/J1YzrnuJml0FedYv1MNDFkDBQzhyFuTAT2fYmjBZ7z/r6LkfB5lSDQ
zWJstHh3Qe4y6cHAkmEjLxln/M12C0Vl2hRqJgBcrRZ81hVb9S8F71Hq9Sak4GKu
M66mINqDMCLh/90lkpd4/yGYDIOGZ14flG6HtikuLm/VOFTfJXvmuLU9PKjwDu2z
f5FiL3TwMYicEorq3jZKGTl1UcXStXTqFlZ6x65Xlbw7DdRMmnVVRW1Ye5c8PpcT
v/JYAvxg2GCqWrr+LnT7+dJ21TKt7kgFWOaPI6T0JgQLNYO7vYIPfCOle1d0yO31
uTCxYbLs3FJMU21vRoIAFxy9Svp1h7kHYX+UfkqKwb0mvO3MJeT+8UXhqSysChhZ
cXbCLmxAMDUeOQzRH8dysoEkEy7+y7dqmHp7FB74muieAD4bcdp8a9HdI6ie7wAz
tP/CqGpnQsTITvlnXHYKG8BK80slBRP+ahNgNIJ83svUfS135o5l5J0jbzuSo5XJ
5IehlnedCntUH7W8GY+HjNed8o8lKKYmWLfqDewT0PdKKFPqMjVUGa4CpI4e+Lf5
jjOoonQ9uV9eFlAYShNWK8Fkei1W5jUj+zVmB43LuGXBe+TYNi2oz28+TfCDXCpl
VrYfMT8jNrQm48aWkw85dS03ywbMn94xlc1K6GD5FzgQ7rfeXVFviySq1I6DvZEY
v9kX9/AZT1P+ifj/7cTIVX9HPF88Srj/dLzroktdkrP8zgY2dY5re6b9pIazrh6O
FfRnrakZId/Cqa8NfrHmkbnnP3h2g3vfhn0kFmeN78B6qlFaK6AFiQ5cqfJaivp8
ze/RHlBIplo23LEjHbxu8pCZGtlarS9DjaWqrEh9j5klXJ7kfIcm2Pou8vecytmS
XhIRv5EbYdT/CpLV6c0dPoxScFgg1cuwRzYoV97YW1uqZMSZvD+vxt9fCOKnQ4w9
eh+TkRyqZOJoJ7+MKkg9ijilavp+WjxRd6FGSM6jMa2QXoHmlRCBEQEbrlOVtxnt
8zQ8nQLfzQLqsdpMPHsbNZ8fgv3IDa5hP7fW2CN2UFcUAnMLAJpYZoHTo53dlxHU
RGf9ac5gqPeRoj+U3pAVv+8ctqYJAfuLYrZbbO08hB8yDcDScdInj34+j5oZjdmj
KpzRgSXilGUy4QJjtQPxMnq+9LtMZst1N4IOzQupgM07aodgjHww3RtNyloxBP1d
ys38Shhyifm+vde1IQRqkvtK12dSvGqXOHyi6Jg1ybIxmNHYeiL3UQU+5HCyq+qG
NUo6sqMWafBDvXDEy5XHEDwvla8VrVkL34cNk84xjR0mNTfIVgKy6cV1n+qdNtRS
oZ4YrswZjuOg/xSK5H8JnthdKvEjZ8H/oTQAd5OJNvG47/cxiV0hNBwqhUJrF64z
Q6Kf6ZcakfJSeIJcT/3hVDtZ34pZ49yr3IcryU28HV4m8FA+2d+FOVgarj4eFv2o
5PZd/G9xT5dzqLJ82YlruYWZSJL7ktF9JjNqT/BH3FQG3B8mzixSctKk7xHXEWoB
GtVJZMjFPeSdKW7hvYCAF/CBkPq1y+4BhI7Dg4nNENIGDP5tGK8XlL5ZKnuHIdT6
WCuUSRhYRspmpcioGI5p1uGp0yGvNPAvd2nQWdr3r/lGTCuhhI3QrXvcUS5d72ya
NGNxi1ejBBlF1VuGXynqkQ4Awt0QK5ZGUWiEOyu3n7jJdmVo3//R38mJGzMjSoyh
Qj7roNolv/e/gZAHnr/QmEBKWBToPP1WPTSzLlhx/ijbv2cFlTt989a5EpuRgpBD
jnUeb7ZHaC9GNDf0+Ixwqpi/cwZIThG/ppgaPzMUvOdyITup+Wrp21uaWZE/ytmn
PwTQl66ZR/ZhhnwbODFO6gmqevM8sEHKoL3pgCvtS59/sbWP9teN97tJPkZQvjPG
7JgqS7siooAAHf/hRBaQeSX1PJbgDNKkFpFfTQFJkexT7c2fK69gql924BULE/5I
LvkCODGRHxFFhH8ln5a4+OTVoVmL5KRj5AA62lufZfgFKCAYNC0LrgQa7DZ0feJL
idVrXA0GhQSB5cLRHQIsPDQpT68S99g7/3FzxvB/ItivAsdyxvRudh6DM/sL0Zex
RapVRJww/fowanyXwcHsybiw31D/CFup40pYD3+LUqaSoxGQdrhrGXealKyVUmI5
892jaWGI6287oGaqGpQES9fVyvNHENgQwCXRvyshkRA9Psvj+/i5uvu5kyDmTPkV
AcIkSEWOFY8lK/+zUcNWSYxwYqILFEo0PfzChZ7QbMmQW1++l780woEyFkoBQ0iu
NZiHbIKTd8PNtO5e/YqXXlvK0gq08W85KYJb1uAslUqiDn1/hL/IBPymTz44vWrA
YTMPPsAdgDGlvhz008wbn6YUmRo2upP7BDzlcVZFqWJqupZUzubRyk1n/XSgsZaN
q6S4zxOjLrjZ+8bDsfVrnkdBNwbRyFG8A7yyIQIRpTQLBX9ZJcX/n2hHUcUwq2Cq
tj4hMBllCKyql0TKcqIbTF8ej1cAkKSDqP1PWWkk0sXLqFQjrfgePf0zA3PyzDb0
iOPPCOsAdFupi5EFSSzq/5cOvqOXZ0ka4kb5XWJCSkZcBcDV2rPiMCVB3UX00LsZ
ojWZ/RyG9kmhxxK4Cc9oywEkgo6b55aN4wzSyCKMV0oxfreCgUoenwOr1TMDR/gZ
4ojfhWrcBzZmJSLctc7NQ/6BDca6DSFEH11uN3Q7L9GlAMUd9+36s0QE3UzOHcLB
Br6T1jXc+PbLHfJhUkFoatkVL7XVRta21o5AQZtdcc1S8wcT1gkerZF7ff/lvqWr
1rAsbS5ipIp0cWboZfD6ldX2B2D5PidZy8IO4wuELVcD0hML196vVNFrTS40e7Ck
Uccb8bdhEo6YQ4xFLAtG6cHWN0eGsScKK/L7wtFKVyb+kBS0MklKFkJL5tymDq71
L7yy0wAL7ifr+oGl25+By35lQFbpHrRYcx+Qxvm5NwlGFaN4MzFeNCYTPgYSMrxL
mUqp5U1McuMshg+WyR1l/v3xx/hzvz0hpwqHrcdoqWbu1bDe4y16U3kccNV5Q3Dh
g+lmh4FxMFP5QsclNJjvETR2GTGMRAklNMxflXK/gniT7WILhBoQAKbK9vkDAlch
sB2vXwT4NknSZwhzcDLn0BSvi8ltErLinjWJoSOM8efeMYARucURVKVFiy0iOTCB
GMFBJaY77M5V1Y2iGZv1gm/O8CbcgCf2SI/IQofKVZkLifvFaidfw0ECrVHw6Q+n
DqYufLedSvuQBf3Gm5pIkf/ov1KCwJ7McoSiNoG/wGpUF8Go1AXjJ+v+4WOJvgfp
WI8YOWK5wpzsaNcNPAbGpgYbXxYEMPDG4q4l/4+Xm0L4goBXEd3gNbmEI+AfgbVf
D9Qt7rBYoAHAIyojpN6o2K0p1MCIt1d/mHPtB3gvhz9h5bNYFpt/PZSAkkHeNk7l
rhVVT0+lwF0eJ1LT4Qge5R9jd4Ei5+IjzmnEj7/V8IP/SR302u4HFKVqpPD8XaAZ
JX54bA10WijaSuZUOE3N+oCSwPWfxN/HznOoZomP9ZSFurL750hWJ4KH2RvwJ31i
cedWv/XOifLKkLbV8/Ds5fPcM3V8K+ympOUuJvLln/Eq1cTxssYPlJFWlfkHtoHB
P/xIhNvgSkL9eaNNP38f/o1LoPISF0lFbuOM9bXUUT9n8q5wRBr0seAqCprGngn5
ih8zcdyhzRdDs+uJEeKyWOQap90n0f09fSzjkIgq/B+Ia9VIMUM+19QED0EtgJw+
O6/Av8Yr+xWfsh62bxVxQzTl9KnIsGKK49QfxTF9mlPT437iJKn+s54XmhcyVB8s
BYqfHPZzt4wgNU79ATLtkz/uSzstI5f5pN80hzKzF5urrD+fiwb9bT00TxEsI9+B
srr1FFvoLyMumZrR++fSPcxiVtlHGWlAgkiiDgamjHIHM3f1GLeMehHN4qMcJ1fr
JK6NQXbCljUuXJgIYA8DhDJPgvQ5Onm91bCpxAQAAhJfqCIG38lFvgd8nzSePmHS
Wqe9EX3mbVT7UD0CjNtMVZCl6PL9vSCWKijIIXlWT0S6aiQJ9ggbem8Pc1EPZXKX
DCKWCvHkjkC6v3F3Mtx8kY7s4+JzXXjoeGTBXyKlnCXojK1zvAxUTklkHBnzhQln
b58bCRexY3REp1Digb021Ld5usfLyMhhuCHSaBpjW7tzsJY56xo0UiCyy5Z9N8r8
8ZehWlAtT2qh9AX2yK9Cjj6DpVxwSecT/U5bVFDeKADyrtCFzX7pgiq6KErHAfWc
T8fPrjxe+KpufBE0WR9yjX7qknuu3HvZPpQ4Qtw9sRWCzdFhOHIPC+YeCfrnUmDo
wohDSnUbKbLZyd/Sm7LHmaXh/V3ilhSpjRauJpNI5KEIqFAl4jLotsUUTWFLQngU
WjRza998gELPDNzJ64tyGz8VHseU7N6i3+RnmL481WZ50svFxd484SCmRob1+3lY
5Yvk/OjkL+Qatf1Xy/ujrk7oDYjq9U7DLwR/tW7JfxYH1IVeGUFTKdea/ADVZmcX
Wdx8/Akwn2Mwy46s1HuB6gTe0o9R9kLYZHS1K9ad8hEiFL1/JYaxrRwmnl6egoxV
Gb8f5oEUxCiOlNM1IMfcl7Huds2UFPRtKRK+7knO1dkQtoSP96fdoKtbp92iqQpM
GzowVJhfbDPP5nHqzLdRbN0YP8mVjGcw94vugb9asbBpShyiBrjLlIk6QOmxZHVb
3vvYxd+QSM+KbNPHiP5K7m14rR8zUcB8++eXK/0EyMjbFjI7pF+nRqAksOqfkf7r
n5JvLkyb5Oya4xs9Y3IFmF267cTwowRKrLw03duI+/OtziAxk7T+TTNuGRlE0k25
lX/sSgRUlkX7gykAxptiMiGzlnw4FQVRuFf02bCdg0VaKfchsMFBqmBFCLvA27XI
Z4ZR+9bumNoUNzilKO0OSb6Wpyu218WRBqOwvj17R/iJdP0TlRwAIabZgDg/EtJF
sE6EFqOSwwUjcBvR2esf6UDBWbrW9Q3W2D+GhwT5LH145rVeom6qRlSsvNSTotCf
oW29DAjezSZ4ZMTJgp2cdciKU0BsafpYNhI47NQicJGa0I2mrlX289+8280O6xNR
wPWmYHsCbheD5SOrTaYHXMws+LPoz5mTqpalDo3ucGXAoVzEMr0BkTiFut0TMPwi
vvNTnAi6d4Ukw79jWCP8s2MnoFvL5UJi5f+BV9idzVQHBaj3az5Xp2CwmN4kHLAU
5Izwq3yiK+ENSLyB7Rg8omXtTZldvRGkhdSksFVUgPvf8I82XgerzREd36T7lih8
3F0XWr7xTO4cOs/gdrPnNvSjheYUP973zB9wGcHryUcin8xp2Ae4bfIIOstZPwQX
2RTYDOShoPzZlF4bVgRIIc+Tel+W9Hr25V87giBaBexxGPO7J7pABVwlpu/c2Oam
DJJ9TsYgso2SX3XujH0YfIss/OkFeYc4DW1OIZIJgEdmc01wUk9O62VTB1k4gane
sOs4RpCNjg35Qu0EVHlSebk/Xtgm1NVewg46IKWK17KIkhqu/zV5n0joKHTBxtg9
siTnE2vEe6ceXQGasK3t/DSvLQXGS3C7T+aF5rwUSIn7b2XuNIpkV0mYksi6k9uw
OueQx9EQFLGzb0LM4ttPLLht2LNn6aA9ygLtwiZkOW29Aiyb0ZPQWJ8aJcVsLLS2
4lSTaEWB1ac2MXssbpCEjTZap+Lb4gZ3JXBqt9wGTmgaFuHCEH6cLKwpi2gJ7tVj
+hjokEfJY9XI0OS26bg30hXNnk2UqmhlisScfal2o3ZqMws+Dll1lSPSEZzI4TzA
QcntPhBJczBLzD8GcCmN+JcypTVbbv/OUKPjQPiUNxU1jsYlc0eLdmUqE/xpR0IZ
TYeE7etqcpAiLTD+DpWrV6FhlyGa/Z4AYrKk5HLW+rVqp71HeK7B/VWS18ofCbrp
EWLlhj7vMuyHE8wpzWV7P6lNk3gKthnDUzclb4FzFbqIKTWGToGyqbfEv/M5OdOr
I51JudcLKFiwbc4Jju2zum797m9BbqVw7hcIEhqe7Ge7wA2RVrK4lla29StL6fET
Rs056k4rkl54/J97BQcatntJVzWrkhfp9Y9MZWWdnECLTBR+i0S1BIW0ImacpP7B
VdB57KO7AYuSgyiin9f2xB00whZSliVRfniB/EsjOhCe+GTedgz/9tEtb0i+TUqE
VUlZNlVrcj0KbEmll02g2BDyQmUNvw/PibUzy5iXkEZLK3R+rFrbaA/RIQt1bQSg
r7cjN0tW7uWkty2kBsCyypYkxiNxWNxTj5sLsjww0XSCdjdIbZOW76DFG+DipUgl
uCOqwDSTG2q74Z7hBLbwTlD4LB1zCgbR1obkQJ7azR0lsToD7WLTWz0C7Zs6gDk1
2fuFZHkgu3kuRJ+YbgtxX0utdqOJH4vJrhgyJLGDA6xLd51WNnWS/bGjGKIot3JR
NKSz3FPE20NZVtjvW/ok7uE17kXkyriB41xChFzKrLQFGmqZVhgvUmeHIw3XenLo
uH7PXRsGEu42tS9C6Q6/Xo+q14Ukn1xQi/DA5clAYSPx3P3b7FgpJsO0fd68Xm8P
5CAzkTjW7NA19ZKAR8d+gKA2MEwEdPbuDqaqe0EXbKq6N/teTb4OhnbkdOZxiQ/o
OXVcNohHDQC0NImSUZdTwAVfv7Ve6O3A/DBb3Q4mjKTp7gMnsIBJC0QtmYRSPkcx
UVWVKL45KHYCbk6Sr+YGT6JQVjja6r+61hq2tJuEWNYBG0X5kS6bB2wXUJpQ0gmW
4+wJODyX/DzEIXHlbfaWlc6HCc/3/QikdAFTGdWRKCWH41SduwoaOo4dSLcG0qR8
N0qAWyW91OS7paNPWu7aNd750L+b/odEKDCCEQY/Avb9YTYYarumCy5AFMAvUb5a
9qF2ZzpBMFKdnUSQek/9cHcQmD3nSCa1qlpnyKxBOSZ/pZOZT7cez3RSt0yu6GDz
YEQxdErd7lYhq8h8q0x6+hTZxhVNMUAmDcy8LLDIz4sgqOjor8CJ3/8g/Ft+8Kn6
v63FcfQ1trDCi3LJIn/aQp0IMIw79w5UrU7RyVMso0fzdqDYjRYxtzTWvVb+Z7lT
POgGDF7QKWIQyKsSoIb1TvSqLr7w/q/KOJY53fkvrNRTX5iNzzR8tWuGO3RK0a21
Gy6BnTO2U/wfhsyp3OMjzlEyLkNwEeczxVBuPwcBSstKV35oWcnRCyfRiax8sPMs
Um1EaVTErB+5K6ki319vDQprFtASbBie/f18+shpqlT/VRNEEHlbfrHOgHzilZfF
qtvgcr7bXIifUfVdkOl4hIdroqXPjHOjYptCWe+s6YRMglcEeOL2F+PzZlBjpO44
sE0SZYQmEyUIYVsNVJcARb1GJLssXqLccgd1Gn8dDC7oSav6eFD32nBN8jdFSLuu
9Jc9st8yCrBPY/FiZ9q6LE+96IGhRiMddOk72rFXIeP3qgKJZljaaarBStgzy6kK
lPe9ROvr31ViFYsUQZfH7RNhgnSur6Bz+mO3Qmc6Is29B9KXKsGdGSFJxDxtuwrZ
06I4TL3VKASZy+69YUb/qI25cv+ISWph5rvKEwyzVOZgjkkRZM0+/0G6pPg8ZtCu
HEKjRo1kNUd0vl74LZI2a/gmqlDYBbqwekLomQkGYcYXlaE08WZl0ulmrJ9iVv+q
eVZ/0710RcxgXycDHEct+EN0Rnn+b8jLJeBFrz9w2BZ0Xhcu8Z95s9wug3lbI2S4
4unUmhEnAUQmEEg8q5rxf0ze1ZfbzLDyIR2OQxy+AhqqjAmPpyNJnX/acaSCRKT/
05H3/iQmhxJhXkP1R6nihmbmAdVfrN7er2LvPO6qTPs7PENzZ2/upZZCLVf0upyN
Iq9I0QYoev8K18BoCU1oiwBsNhHiRb+W8mNiU+x87RgiFFTaZCrK3KhdJuatION+
wEek1MxNfPp0vUhsvphUmHmUYT1LDjACpcCqSbKE42etn77ESI56xilOS4oT8Ghi
l6dOMRdWdgLAkpaAgXO8bmNFagGgVW+HUFWbHHbw5dXalTQpD3E9xuB6K+vt72NB
HeZ0cbH/rkNN+dIVc9BpSvqqGJzHRH1v6ANqQ3PBuVNZ6DHTiUHFJ2U7tphzEwnp
o3VY5srnF8Mnwmz06t+t4YYb7QZjeb1KFnrgsXZNoXXdLjOvcJschO0p9tTRGEAT
Ct9wnKAg+fVgNoa+3W3nkX26zfie7oUsxO15tPxOHhL4L3I8ZAUvNfu1VNhN22AN
BXGSBMLgbX45Nhfk6+e/JZxuBRK/j4MeyFXHDdBTJ7fAw/KtS7pUTJvDBxlNYtpe
TfYcVOQQwvYGbkzeOyEnDKYHrFD5zfsMOwezXI/6uIkved/zMG6Jc12YR2mriyZG
WV7kMmbywCZgQA32w9oXcE/O19z4RDOTZ4BpM4nx4cRxaSK7r5yEUgQkkyzje6EY
Ru7ygC5tzPSL+cflGedvAz4oZJetO1b/lnSdti7T97i/vhrVqWiPIVLowCCuujQC
bNZn+l5tCrjMrQSHVF45boBipAnva0uMw5hbvx8fEQE87THCZ+nLFDE0tkxx76We
Ib5Oq/VTa4WFkvG8WD4YPxQNlVM0d2xegDKPragcOIxc2JnfSf1hbau2mV1T61f7
+a48m1+wvsOnTCL1J9JjXQeZtx/SPE2PIePGSgaOHO/9TGsNS6Vtm0v+Z+xmtD5O
DA/6r3XKrJP+OIAERcYHQR9IBhzXRenIpMqs/L2c0OWPE+6tvEnQfxSPFFIigzsz
nEP2q11cKopd1T6oEzckT6N8kgckFS6fmmbCLDICTdA15yG4Ty0jaDsCw/ejFkmj
l8vWIiMcz8mQeMsc8dC/Zvo7EtF4L8JzJRIbLmgoHbLIyFV5bzEcd6hBGLUjpkZK
e5fVrRxHuCXnnEnDT/HtzO4V3I3yFviv/btvwxWeQgfuTlQhy0qgP4jAHkqD9kwV
gkF+mXpxf9Hk3fCg3SqJ/0mDNQEzrCGDZpEwZe+gGS30ge90J5mXcU903yRSZDFg
WZh2jXSnom7EeQTeS8YODJwryJ9Rpb93OMRv/SzETSHbOUxnKz0NDJgRHv+w/5qd
UZsqqamHdabkWgjtQTLWWhtjlAALGeBwpzOj0fApJ84ePjlAgkD4L1Rpr6aQ6TOH
V65ZSjOpQjYaGHJ3WgdmNI/bzcRS6X2utta4jpN6R5QWx6tjmYxNztRxorUsT5XS
knmBO84YEe7e8tJDj1Tnh7ceqa5ZYjwLJednxEWQq5F0sH5toyU1jdI5uqJHePxI
BZr+01WjoivlLYnuBd5VpcW/dRxRoBDbk9TeVO9clykvEwu8xLbOycOdFGf09z8M
5bk9s4e6AKOK3WpZ7WHJH258qKGGnVE2G3XyEimv6MMTj9Ltw2iMZf7u6Lq+8Wok
ZuPsWNDJW8MlsdviCJ/XRQJNPI54J53a1fkFzyWAUz3kKq02zi3BUhP82dp/D/Nw
2e8xgq5T3ryA4N52DcvkeGFbv2z76sfMeiHzGmxhPoGpeBORrwAjXflUTmoDPtK1
LfGNrCmx8dp2G1X6rjz59LwYPdDEHKaR5Y3QNuvh0HJI3XdhE5MYbPLdZT9kxtxD
WK6Qhsfq2hkGOCmVPcFnB/g3OLnAmgOJS8Aj+ibRMgKb/ziaP+ITif5YEdxu0Q5p
WeplzN+CeU0F1o35mwOBK+bQq6Q8IWZFNOTQGDLVVafN+4Pp6SB4omLHaE0FGk0A
T2MTJP/1PacExALrBcKgJ8uxkh7cplltc/lSoFsgP/x+ceX209c3cLSAk2Yy7A4s
jtEsPe1EolAdSmXXSnokoRNrzYt7LMexUflpR3LbOhCH8gDkVly5bhauHlLsJwQO
tyJ0IwCzEG+bKepoOKhGRBgVPEZx0SfGeB157mKG8PNXDflDNL3ByBjlLaBrRy38
NB/+7QGgtWoGoroRx4hp5tl2RBgnrY6TPRCIVHpROcuIt3itM+XOpEYrCTTaU1aL
je9HEaAbIv3jj/ONeC65Kp2XDRQH+e401jP4CkITfui0MheTo1Blk4bTcaMPGMc0
zRYO6RYPRUoELPntsP16B36XUtSuwMtXBurngMuMML3EWNnEFZ03zh1GssjvwWQW
XWB/2pLNGAIwbQ0TIDXKoTOr/GgZe1K22X/VB+EUPw5Q8Vxcqj5+9JiZXmwkCuom
N1VfawX4kFwc9EoOhNo5IMFO1DSOrh2LyEdR+62O1s9Ezo2FeDV0u3iCi2zhiB57
N+Y61yBtSvLYG0soUveItxZzDRxzv169GKH5fbiZL5+j6JBMd81FbKXwspX97+db
CMKywDSHoRWae6KaGRHStuIRPwB412Cr6nNQLkV0bItqzHVje7tezeavHEH+QWBy
cxP38PCIJuqOSCXpGtRs1OsngKwlQAJEhcbrTrNFYzo=
`protect end_protected
