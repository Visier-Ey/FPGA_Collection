-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
aFuzQtfW3W9B1xz4GQXp37sNyEcAVDCcJXdsf+QUcxVkzAtjRdknbGA6YnZQmJbZ
sX2/C0ukGt6a7QcvCZqKKVxEQMQiCVAtyIJ8LSc7bO24oKJrIHzoca2z5Ji9/Vno
IvN2X+JYZDUoSHMhVeuIBwh4qzE/4NiRxtkmIPUJ4ck=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 13035)

`protect DATA_BLOCK
qb9+Tgg5I7igQtS7VK0MlRZ3qp5WzwRt00On7S0kjeGHKGgDSFTKuvLeOLn9hNAh
tt4746NEpCKWvg571JTrL2uRea5+dF03Xy121l3f1zq0Hx38hwFOts2Dhmx+TocU
JkgPo1th8gbVq8ayvX6a8tpb2yJuLm0+k1nsbxT2kOCxJdiMI7ALqJ8+EhwtJknd
Nw/JpD8LCJ2EBrozjheJdsVC4z54lrdeBfCzOVTOBFTUSnUqe8qGroHk+uAddbFV
GjmRV2nXuf0O7y+M5ww54Us984MbXVxXZzxm0+zdG3fu2IoSNpuyD7ltxRmcDmlE
z481YQ7BgRtflctrtZNfH1+EPVw0KguQ5+JQoScXKmeK3IlhCTLs0bKO2sCCCBRF
JYZ8GdmJslCBrOD2r7OqrhTmAA/YZdhAkNUaeCz/rMt6xrKzNDp7AnJdNubHpHAp
diC/UzAIAxR/HpORm4CjsZ5eHZIizkfvC4tIKZ+pstWP76Yfp4JIu1nScJlSlrCo
kx87Zj2kiVeO4hbFHVL937G55eX6S0U6puBDxVFRR6OS7Pjrje5fuaklP9X8unih
Qxt5cIxh4QJADu6B6428h7ahfoC2vfZppSxiJQdNa8hqXVx+BK+z2upw6w5ByEV8
1+Wif+eWg4VCLO2MHp1l6VXLYTKg4U+dL51DJ2X6g+0onstlZHW3iy5FCiGYx3qB
I/3U5rEGt9Dqg/3NOi95wTwUKuyridDWEL+j2woZOTdnMX1QB6TbUXT+99LhYqKE
wQkX6lm61LaZ//mRbjjl7T2uhjbnSQR1r6QYxtS6mH1Z6hoCDE/cwN8ezuwUx/SW
s6hQrkXuDZyhpSYuhf8exRo2BvDmteiKmTnJMIZKTsaRhvBYUHYn+PUwK1mMcz0y
GjxpVlpx1FRi4O2gySFpOVgZKz1uCPGlz0gXAoAwhRF5IAXHKS4j6Z8B6YaGWnJ4
5pxSDBlVoaXmQ4thv96uW2fquskiBCDwGMw9v0v0NbX1EW8dMTTxUsYL9RF8Iz2V
MWzFpRq9S1iB83m0s13heFGyFRxKpQH1cqeK+UnPlshInVKFVm6bb6YUu873D+Hs
Anr5Xi7zY2CQ0J/XidIMIJlngH41wb5Xp7vh5YKegjuICYqJyrbCzVhqm2gDbGaC
RrcTcP2vvLTNnf13BEcBr7vIr4S2OkyLqLTVNgnKc7TkYJg7fiM3i1U+X9nvdnEy
Xfb8Q31muckR/g5ED9SFiZj8I8k8Pfzx4eprOUHspcqC0PY/po4nYU6vFvYilUCc
3lcssTQDng0bYR4osgVH+yTY+EBU2b0qQOYxXxe1KQxvKL3lcu9XQYXs+zvlfYGl
X0b0r3IoBiDeN3FQLeOMURP72KR7HsEDixjzQ2pUPtZu+/dzUJQ5wC5c44RfcMT8
en8dCbYWd8paooX+zfmToj4bSp/xBd8uumwnzU6OTXL8bBic+PkJsuQgD7VbuZ0t
mS3O0jEfdRgwYKZDPaod96F9MlrCuEvYV6iI9xZk7nrdLuwI5eOE2+EB7GPAl34J
FJufEVbKteZ9KwMeeQpuIR5aC0Ji6zyMvp0O5p+spIAiL9CKFm7kIIEodKjUknKc
jBS0u+2U3VHNNOPjp5IitaXtoSgp91Y2Dzkshq5A6Qy42zB/cdZ1Zfdl1RlXnYvC
kGfd+MfZLUCJsGqAs3vAo5NEdAGqSzmn06lMFn9G+Cxdl75A2/+VXM1zg6oVaxdz
zvnZMDqxZ8PxEXr1P0BPGLLJsF27ztK36unbC1WvKMNwQihaR26JfgP950sbdU64
NkOqZoHMGwniA1QtNzITSWfiFfsPsWjbThe5/OkEfM1KDq2emU4AiaWfkh9XqF4Q
AldSCQp3V81BmC6WPCBV2KEADYuox4A1+xkx1e48fJLbUzVNGz/copCUMxIpFFi3
0w25ZdQNBZTNGimxRoixX8D9MoKsnFD8Yqqz/QtgtPCoMnwanmBllYn0SNH5kbQH
7p4tmse1KE50kUOjfO4oIIProDUuNINO6nJgFbLIzsrUdmb9XGlE2tTHoYqwg/Ni
Ih8Wt83fhg2//HW2dyVMCUAT3Zk8/H2Z6T91Kec0EW7/39V0MabS1WYvysnR8R92
IkTz0FL0/0hepVPT5mGIUcwnw1uls31mcSBCDTHH9yd6zrrO0B2woyZiOjGvTXrU
GVkCwXRuxa/abO6x3lLx5hHE5FRFmd6ImmOQnJZtuBhkspdh6TaA9Qv8CTu4n6Hr
7OH2QW9Np2P7eyuIsPCvIwj1sU5/V0byk1wVDcdCFZoJxMUG5IBt9LHlTdub39Uc
ycLtxvimkMR/zKKaH/aFGZX+ABeErLKL0XvNpGjuSRCRTj8OoTm90GLfDDIrzHnX
IwgsVtZsBIQfac/xunh4u2xN4iLLjhPo2oeQnCnrHK9+6zeKjjFuwtxROvL+IWVc
7lm4SzZYAl8fnR9XavjxywKu2SQYFuOfBldKnI+Y/uoEOYOiivwJMHj2iLL0bbh0
JVfX9Eg2JSyslIplowwHPub1Yec3bOGqyeKJyjcGwFWNqaopua20/Ss06CgCIz/p
Tgf8CJLLlUs9wFyOlZl4NON8s5Fq2dCFUDKSWkKI3yhD7phIdqKR/ImvczV4IPUT
ERbuVok/ZtgMo6kjmYx7Dq06LGxEgf40MyWVilIUe1zi5gvHluvlU1xoBFx/9h+j
5RYSCx/D4Lm1owS3DufOJo2TVzgq+qQySaZz06MoRzrMPKj15jPbGcPOlro4iz7R
urXKMN48ET+YP6BRSqT8mlB6B08/G1aos34Vr2qJ0b/F3GG0CMXH1nvZudLBM0v5
ig87EvDJ+NnIEx/GDYPk/kVk8MmWyTq8Qun9RiTQ0/bK991nvuubOV5fxCdnR6SI
fLFSwPjQVdsX6nEA1GhVOjgZvDbtw7MBMsY5SCg5WdqQJcCom1fOYCSHPgjPkngJ
UDtidXnIB1ndfNL9T4A5Z1VVkuKchBJF6cHMIxHnrCKd3jkifPD0IWyaxPiOkCbP
vq02yqd2toHdHww0czr5/TEZdFzYFSw2ix0nLA96h/rRCRyYtJuXfl32zV7/8cRI
Cj9MXPe9Eb58QSQCer8UVdK3mbX37XFVlBcarQV5D4kv97VWBRbqVmxS4TEZRAxF
h1Lg4jAh5iQ80FJR9dsy1qFdm+KGIPCzGAA6khF2KctlyXi8nuM/8fJtizcWHu8t
zP7yrtxYivBl01kfhv7GnmImKVLedPFWvb/ujpT2l+bnMekse1/WiXIMGGl8a9di
xYPNx9rZd74v+Zp13ag768H5pZ4L5hYLYbYl/XxUqw3pbqV0O68KwsIdolqFpLPC
UX69yfMkgylV20/d7IbD2CudQxbcGyZNOrLRuHpaSHvrX8IuSt+G6BPVoekSUfpY
buXomwglvB3c3fUo+vRs72o68TkpktTvkgzrJ9BvUykF/SwC2lx8RiCg3BRpbXNQ
/GSXxumbDXtPbkIdLbb2iCRV1LNkcrHUtLZucNXknmkNfIg4b9h0CVHuc4oZ1SWW
D4zq4rhBhPPUCWB385Vr4RJFaIlSCjyBkzym+nrjuNKNz60+WCR5R+Qg/NqEWlTy
OeBxGovVJTr/BExW+ojmGVKy8BefBO4aUImoMEnQfOHkWYR2k3ue5LJKSIn5MhKb
VYsPHRDkg63KbeUHPvIDiq8Bz+xk8gEoVwBUR3otq/XUC87n8EBpIr9BxN8slrDw
C1dpTxNb1CnTcMmZ4az/32l/l6muRb/B8McjNdJ7GVpSd6tnaqa5IsdsT21tMMrT
Ie0PgNHI0yydu4ZZxW8bPiTs//JAjaQhUwClWQIWFv5AHx2w6VDLVdWHqYDQMy/v
bzs74cvTNXn+b7qDhKfHFG6FLyFgi1rKuzgkmiZkGpHyXdK1xo+nfcG04+DA24OE
VJ0DxoYECbh5ANOyeJdmzgz+3PXi64ik562VmZStCVmdtzdM2+gGiW81wdPaBk3/
PxRzHDoRV/G9ULq3bM00w2YSp4elLDmFsk+MrvAuZ2NFHW1sAdZzLUv+DM0HCrlV
mS8a439BSiUJlQCbuSkPjSOxdGTVHojsg3T1LmOI3FDEP5EIUfYN91FBZ0KT/Jcd
g4j3HOrKQE4Rl6qtKNvP9+6U5kNEKv4jxv9KlBj1YTkOGUSOvuPGNEZiH4wl9vo6
11MJlFwrm1ZUIJFDA4IHPMydCF1d02VNH77qHTFd/TZcvJHmchgXm/JuUCAPerOQ
HCj5VNBvNPrkP+vBC1jCXXklQ4jZGiRv8guNuvgmORuIqluB/TZh5VQgqKWIxED1
/jqA4dnYTU5YLEn7DADyff7npKRGQp5LazNmcN8cBmzx4XZYzSNhZ2EWhIl5p/HJ
NxQGj3ATjY/iHFlOxiTdFMwaIHWIQqs/fBvp5lZ1upc96mDKLIF81dllJNIIKfcH
ht5LS65YbbLDypXIcUSqdJ1Gd9x8yvrKqq2lTYejmGG1+AA2ldc9KDeOQdqiTOhF
uNYqH531G+VEDHZOrPT2WGZQ6uz8VWUQVhtGoBO0Z0aYesELL/e97hMMiyhDNTzA
b9EVZUAq4ZjYpa1Vj+HStAOPDMokAjIkBlrv9SqZc1p6F7UdCqH0KDYGrWnqVHLE
M4RppPEPDH/0TXxpBYlJV1lBwIbf4ijg6ooTAWk36ZIpvlFqDDXiGRIW1ubE2s8v
GNZ/S79n8JMBFQTy98cyB08nHMafmt9vk5Qn7DPxF91MdqS5Me4xRsnVdISbv+Fr
b60GTMCm9m1dUy7u/xHcDMJsFhPEQFG1kbtqpEUxA2WJuLHJxZjvF6OPe//UJJzs
kECnWNm+gb7lP9rUb6nCgs72qCUsaTLy/k8ZqPeEEJxRx7lV8g0gOAcE7os/rt7h
Itx80H1qrjUw5ng4YXNKR6vmgqHO8ZnfIfk4jxM2PSQvP5eK+sehPzaX8+857Kp5
zt1NuRrpyoOmG10UXCcaACwdLgVFXQoPgS4nC+0mai2x3KyTFzKBlsFmbsFIw5cs
JlUTrP7XLmXu1446WkiKqrbl4Nk0mh7cqzgrdIKCfvEemcvbVJqHhy/egM1ZXrfy
6CqR/wALUym74fymleECS3SHRmPN1QQh7Azz7r9MSZJUZ7SqlymL2uO8Ij6AIizJ
QO4/yU3tytCbGFOIzXCgmPDQo6RRXq2yOwZ1BEweXW5V/sjYvafYMud82FXXA3ym
asq7aFQFJ3RRKQlIlkFmgu27h5LmlOM3fJnlgA0gM4owzjL8uRcXwOb7NpKJJfaW
6MVyC5b3mple5jHc3K+xz4nwbTTKkHBNGy0c8XSlriRYtC6GfU8O09XjwtA5/h04
mp+aA+FUSco9Ch/dbHKhmWUvqQfgC3QuJ2sTVfz2aOX2kPjSe+UK53FTpJEV4Kmz
P2YtCX0hcw2fl5AvuA+leb1s5QiXIVfmfN8yiWUulGXa5VDLxBSt/hSqly+9xExo
SVMBShv6Uf7D3zEJvCiRAo0YD6hFLtGwfYZu0QotZbxpoZkYqnBUyUkF4lx1XekX
LfQ4rQ5l88f+BvYbWNy/68W/B7E+lqoWRD6oipcEDWZfXFVPadZSnDjQhp53owFp
+d4en7Xl3qV/OfTZCl87sj+GNIjQtUqxdqnX/pKgpVkr1s8rNp/WlUuyjWMjsFYo
CC9zWl1rChhiTYoYiP9618CeF2m3Ex9KwQAvOB3jyOCwMFl3NSHlnmpunU6oj9mo
IK+w3NcPqa4LM7qzf/3ZEpTFdwvwHI0b231WO9ipAHF/tSLx147CnM3oUOaqPzMI
7Qdz0w0fdDkX8zXDOS4HLxjgEYd5joN2xF5FN0IPkaVzd2yMcvAAlKcEX2GcR0nO
AFjD5Unk2dQDYBZ57L4pFe5GzJZUTqifCpDNEiWy6PiEdOiyvRdiWIUEPDAu0OZO
f37kVhv2SE5iM7JYG6CMu2VWhHFsf3IGY6mR3e4P3YDix8BmTyXrI4e/cgXgE3Mk
h/D5E+36wmCb9RL9Dap3g+wEbFPA/7elo9Y8yIoCxTc9C8/yQdd5lKfa47bMrV9M
w2z0f+xcMyzZ6+cyZG3OAb3gfqlZ4dNRlIO0fj0FONpAHitIozS5tYb4iTboJ4qL
JoJLEBkOtql5VAE2euwRsyliXLAQ3iHQcgJNtAKLzxoepWOmQeBJw9AY+udLg5Ja
ctfyWHQtu3NQmnuZMPVXpwG6/wsH4FU6bS5kPn9FAW4z2cU6zdMxRKXVxMZs14HE
N1xmIuxBJkKxD/BMoCW7rgy8RgE57aq1kdjyIoyVWnTaWenyD0dfWj42NooOn0kV
xEfD4txBDE6LMsxnpR0QoTKEpUwa39xSl801SKfQe7rP09+tO3TYaRKXijFyKHzP
AteozbQNPNROxLtaTtThXM4OQ2ggga5Wv55ylKV0YNsOU0f7A2OxLWv8rjatgId7
9JH2YlQrmWZz3nwYllfOKRHJ/icY+DE6k1+wyauWfpvtr5pt3lOyqiz0P4pecqfR
7z70+rtbxdQkqnQ1GLKktiDMT1qtDzZHGmQFB8hhf8GNWO09qCfULygilawweE00
POc9hWHtRBm+9rBCGCxYXwxl3CaN/1I5jsDRRcyocCNl/7cgGRFhWoyERnZj08RX
wVrs6upzyEHTrJelY5dZMWvQ7v6yhKKN3NvjKWYhnNyz01Izyc/eIe7ubjj7U8uD
EcGvlGjwHMJlL2jfbKB48qfqgCuNnLF/OQAjVfbKfBAUKJcIW/KHpVgupEJC+3C+
K4OvhveB02sRuIMca1gL+/c1j7oWoxto+/u2gUAaDvFTU+mSPB3cB40Zc1jV67s4
geHcE0gPQ+FwC8TtZvpl7m5vx+6aKURuyRQvgfr5FlxsxJmhVw4rEqZTTI+4m7qr
du8SAJG1ePwMBnA4nOWarZIvA1Zyz/SX9Punp+o4CBuD54+FaFClVEBYV48q7uFD
tMiii69NToKD0KGxpMp81UCX8sW0f2fhF1Z35CLjSbdTHlb1R7dMJzXkDexdz+b4
TX8JYa79VDslWfS8I7mEYhXAoCBSyZjO43KnFZBvD5k9eCozHt4rxFd1dhCET6Dp
NpPCiYs+16bqxfRJoey8davk3BAVigyvAUDWRbtIpW1u1WwUIKZbB2KpyBmbKPaV
0Vo1gg4MZlGKpbI1zdo4g628PhoTAz2VIa5slW8UpTpYXy6N7K9i+GvuZGo/m88D
C1H6mv5YhJXPgHwCyl3mRgw17h8Xtnp7TUDQ4XJSn18WSN6oqvBGeAn8keSUKkRX
q3TKdj5G+8WN2D7P+GmKzSHwU27SDPxj9L0qKJ+L5YqxhXlI4/ZUT8mcIhqr/7vl
pJQCK9oXrMtYFPb/m4Nddbkn3yhpAZ9KioyN7A4igVtHUDLFYFn3aYixf12+PcO2
QwGaA5N3b5uL31wXe0dYUeDiJmwNuNoLL46IrQ/dycSNfdw0kXO4QdbB6W5A6yBB
pvO7yQypCmKAWOexdeNsl3CFcnMXaW7Qci2Ia5u4OViao9D3jUPhfn6GEZ3OZc75
38ZeZpMEkC7Sj2NXjsMxs6wko4HoEgRfIo5E4UaQPCqFYzPrJCbY7bgL7EBTxjxH
TSpAz3TgyzVvcvcY3CqgQDT15HFLJPC1vnBzBINfYGNrrNQcZP1dcF0QNqtVXreI
GHWu3/k2QDU56YZpCdYtHLXZ2lcYi5Em0Z34eEnFBZiPfd/2sLp5AMbrLoic0gEb
PJsBKf+Gsf57OZT6JQwigdkaBj52s0PFWtyRWE1SH5ATB1yzDoX1wmMb3XSp8knr
qsjhxGqM8YbwKOSR9YZMOs2GBh5+2Uy7YUBBBNbP6YkZU7oZDT4Da4rmb3oyAlxE
Q+sZXy367AKoxoc7tGHwfqXeEanXtr//BjLmwQNISmp8/a+UB7SUzUkUmAD3IZiU
iAR/0OtacfXDmrqWJbCadNSK+kj9oQSp3xv4oUtR0qrQ7dpcOKkrW25/ueH0vmd/
VbH3y8bJoQH5ED6sSuWvWEuWfmDUXwCc8JMtqS0driH+FHoOR31JB5xMR5DAQ2/Y
lb/erymTmDwdxTphuz7hxW0vVSNgKYq9+qt6LBRU4wW3RJWDGA5Vp238mL+6iX6t
CPt+nunYVxntfcQxBLVjoOWNblTvmEDxRO2+mvrxGXumHW8STMxOO4SWRGHcaexp
CNLSa7ZvEh9vpmtVHhozsfAEhREHNc77FPzjS5uzPRuDA80l3PmofRzphNuduncs
pRkOX+Of1e5PfrmI8BUI4gqUKA4pMpkL0MuhMl+YSgnjU3NTLgInNDBz+BWe2lM2
kAzjUMq45CpnG/AJbmO63g25us00iFW+cf42enVZlFqxzFh5lu6czvwIz/QFrqGv
byLMS1h4l9JwQhHzxslbm48VDIoWuUlp2RhwNKUbHc/2j0geJjzudz9dziWSO+Li
9PCeIM16cZy3pJl+GABpEsbrjWxTTD9/RTXl2GFyzsq0iFl34ZiXVOMhvQFzxhoM
r5QTR4kauUDs5kDWK0B8OselufC1dmuDBwYzR7gVgPjtP1vW8wBRx356EN9qqWr7
/RoGASjNauFFVEWsjScVLkxe3hVHw6Ok95BCE8QQK1reE8ksCR5bdLDabd1532Tw
QfZG6C0Dl1JW8zoSEY0ER/7PIkPWpJCcipx4oOOBWmJLRVLYpx6FL5O5COu51pm2
t3oNHzpbm4htUyiJSMZOoeAfVH6mk4aW7CNGzDjnMomlWM0XFEYivqkR68exPCRb
W0TlCGOOOw8S0bhbOFV8ebhvei/Wg6MHUeD9NkWTpQqLLbrMDsWbCcGiA4Knq7Ob
k/Y/Svmj0bFIDSGZqNqMtyynY+fCdN3Cj/yLdwEUsvlb98GUcgeytPToDb1HpiHf
4W2myKjLPdglozCBXjC8AfBPFYMBtMyK1471NsV7ZcUcRxZ+nXMKE3W/pL/f5Dz5
Y3Q+CNVbs1S9kTTxmqzko5OIHTw4OJByr4hoU07xiF7UhHtAcEzzW2gzpWzveBJK
CwSfbTnWAU9c0K8voCIgoMwoL5aqr+lQghltNPepYT2NnjqzRxBA98RBTDIXY/H3
3jlq2kBZNnrB+7ESYOpZq69gkcNYou0MwV1gWzla5rBhXYiFgQwaJfh8Jl0bt7CH
uz4zyRjLYZOcj/hH5hTqsfZq6JOyFWHNpGN30QG40pzN9Go/6d5Hgzxrnj9fnn4F
qMXRlv1UdNR5dd+dnkbhgVQAmVkHHR2FOc23zVnJrOqwtYC0EaDBXi19MJWlS53V
PqwbZfYsAsLOP0zjVI0TJQrDidHTj7OoxkMxZPLFhdD0Jril6iXqc/H5UFlQRrgS
TkT5Oxc63GAsqmRmQMAljKPXjQlWjZQzEPPHXF2Y8qoiGWUGJ9J+JLDj9+52WwB/
nydgiIDMY536IvSpl3jvFLtOLtXP7HgB/qNWenhiT/2pZw3KYcCo4S6OIWw4DSZ3
/EPf12TAjtH2+P4rHktBRQLlGXhddoO8G5crSgCJXo+rG3IzrHIbJx8BA4kofsF3
8ZyBTzKPaZxpTYAXRlhXG0kqeC5jXpIuAmBGsOdycqkf9wvVTWU61u4wXNpobm8Q
jpbWiI/DDzZ1huACTLHd3KF7j7VLSKFDY71NJgazNwulj7Ey/ZuGBaq3/fP7Pzl0
jW70mmhYZSZhGP3hd2/qBU5WtGsSUV+bQ/AaoJ/Q/4Xx/rL+SMVtaTzmqAQKLbQ2
dTgbBiun5gg/Zs2SuUf5aGSRVoT5vuo+2D1ykSRFukoypDhAXicpfTdUSy3xYM61
ltTX0fdCXKKeat+CARw6EN6ozk6YdKYYvoQHWCDCduwh0+uFSn8y4CB0h8aYnaCl
vGZdPTTEuUNUXXeodzDXumOohZtK5q92WbKpGEVb8vnWih4aTAQfiRRfV0VDEJYH
Ew1sNoaDztHrOCUE5Jf6tVfrr1N7zHdM2HR4XnssXW85+ELfMrez9niLYD6BIAr5
OjjJRcj3dLyR6moY+KZs86hbeZhzCX77KcBLxaTicdikThYiJ427yclcE0IaDVj3
4QcCuKWMr6fftIBzX2CEx0AHlo0nGiTAnTj8gh2znMLawlEywJf1Yk9eBUrPLbum
Z1jBq6aNyr8EQSLr+Nu7rAhHxsJvk5Ty07jn3y3uEu7KwevhbE0Q3NHkk8KigjNC
PA3ghkPfAFl2kxt3HV4OhqIFWXxbuVN5bRp6xDDM95dkjYblVnhCPK1c0is0n01e
ziACc8WIZMeQ6igNdxhk8Z26MEaRtBiMs3EjvKNge3D63C5inhdlLRM5zwXEk6fA
VBbayIeSjCs+q60bAMsusmg63RuSkpWMuQ23oqolWFVcWq5LwcT18uZAVkmDd3FG
1qLITZ6rDfrtj+wGcAaItahkTRx/mLE5TTdghq0fUJfdNkS1d023MsCudEFQj4Hy
kqxiDK2m6sDyAULlvTXVR10HDHpRGDBjKBWY5Twjpl2792F5fp+L7LzDH8Oam1Ie
drYJmAxxpcvDhCbB6a8QZfuLAnXXX8GrGgSiLuVHAABnRCTVhOqgm0fMp0qJa/dr
eN7BWlgArp8kEkkJiaYZWbZJ2LiaqxkSrArRx0Jx2bAqyLmTMZzBuHkbv43C7nOn
nEMS8kZBvaA1Flv6YpCPc6oplvh/m8GE9mS7PzLvPgDmAkPSx1/jLoc/ZYAhm7ju
KzRVahxxi0KBe5Kip3tx9aBQizKEE0TX5CYMlWCfmVv1EQ1ER6CPUj2+IHvEb+6E
bhI1xi8YVkFjqD5dJ6Vzx9Y0a7EdpO4V3e5Sra2eu6jhtPQ6bWa77G5MQ6PyFZ34
eliPSpdBNF3OdGuMEYPCKzWslNcLyY0EzTCB5nM5/zjNZb7MUblEli3TPBx6QVSR
qcwzu9unEUPudG++YnVHSlHf0CasWmssTwG5Ne2oRjNLV1c30FOUln/+B2FW7tzo
uRawEdHygeFkGujNEucNP3GLDKE+isO0IDAuTexPGoBuy3DWTo4Gy7noGBtSOjPP
vKRr4FfxyhuAdshsFtJxBXsxx0ZWdo+lBZ9p8VJnbIIQqtwHLa04JHIDR9ZZDx+5
WZWu8HmECM6zUnv5CmS6N3B2Dm9lbsyiYxkQMHSzYtFdg+2QWo4JwXeGveLfzcW7
Uq3GYjcLURpHaEjf3PD8z0gCenvpQHVom4QSoYF03TDA3S6pQ+KcgkH409HpQhB6
xy6+nxWVPoo+4XyKd9bQh+JgwOTKE6sog9+MrpievMqzsVUYnMCKeDW5EvXeLG2f
HYx18KEJItU+CRgMAo3zHHYxT2PdL4lYL4i9ReJyP2BUzRG/YmMQh74YBT+e6vbZ
+DtsKtRVgq6aVPMG/nNqNwwtQsoiCFmXb5w3dMXx2LdOKtE4gen1XuBjkGYCdzwC
mnjB3qt7frJkEYogd207ObmVU0ay4O58lLE2XzGKOsCfXWjPYyjK6/Hjt8SkThPL
ERr2AGh0ooYghYDPkOyy6oL6DXfZU2AD9W/e3IJ18RjR9/fD3lX3h0vNQiHX33IK
hydeXIpDcp+/kFFCz68iNV8g0ey2C0NrnHbRTiMhXs4pIuD7PI3Vg7MSzOhF5WO/
0NoobBUYVGplQl5l8QxZ0AZGIJVuaoYmV5vy2+WgcaXe/jHcQFJh1D3NMgA9yKbh
itL/G79QqUd4hjDmYTclKlLAC3up8Dy/0YWQHH9yEuKp8OFXS+yXnrd0my+8txZI
OtD/4SnE9cNw4T6wkb7hQaPt6HX7yOR5c0jrOmWaWwGdQ3RXKfRDgHUG4mRK6PB4
1umT5GSN9CSkj9Ts6SmqANzmNKtTIPSsvTlwTDKcA9mW5V3aS0h17fLzbtIfDfrJ
6dMrZiavR+rnv4D+uhKcYJ0/fEIkGuOPnh0rp9LLdGgXAZ0goO5eD0gOxdgBibPt
rv459TNBnLjW6sLDZzUApVa5AHg2nGfNT4pl8U+je4UzmoDmLuL5JC6hjSfKazdw
c+FemXC+dccO7Yw2kC6YulQa6OCZdUjdNYus2tpfueWrJtpVwXb0Bn6E/nrZM6sn
HJHUlwHmMP2Z/W+HXj1XwXeHZA3kepsWE/l+5XEONT5jObYMtGYfyFidIzQNS6qj
17a8caO/Nq1NGj5jRzX0xDbEIDAZhO4SKK85F8u7yM4IXT0XLIwBud1kZX+H0Tb2
OD1gpNsZF7+UJmAKrQMfQJZHz6sVp5ytqcasEZ4L/CR8jhDfe+YzfQcDsqCoOfpD
qbEdSsG1T2NH/efY09NuOHAQhIFCiVjAgZqb+OcQWoQz9iYlM+MOSQrKHICIhWGi
BshnlEqQq/2gMq/x0Y81hXONt4451H2npeBWOCX8zFzXLW6ldfscOe8LnzgNDzET
45+BxcVYtWD0lZYVqI/nMSsLidfAZ5TwLkxOVgCB2jMoMeiE/1k07rECmkLhObM1
uf4kJg8S32IncAQoMpx6v7pD2/CVv8GN1uGHeOLGDYem1gAr0q0VWDmJHDAWqbZN
4zmDKvPgX8HuwABrlxBK9BvQDoFJI2TDqgviJkvMocQNcUN6z/tHW+4JC1VLLyPn
DqSXdDp+LEOwUgem56JWpHmBANej/CiYQTzw2eLs3KOW4A4mrIEBQG9Sk1fP96AM
WieDzXgBpGvf+PoC5JQIY0q2NJpBVJJ+p0kJqm26aXeH9zwSDntDY6N64D7IBamD
nje2mk42oe9d1RuHn2zEk1Kq/zUOqWT0CwTFjbE/znQPyOjsM88jiXUf52mQ20wo
814Xac/MfAVed+Fc/wHcMjT9I03GJGgTByzBBTly5VtLYCNd4KtFVbaLII7Jl4di
3NwNyCgjxAH293XZgiV+ilby06S4lZLGWr0ul6Wl+NtrHpggg7hB5nXf2EakhHAS
1beyyjfpziRlTvrK31Js/jESkkEpT01UueY5y1Stups/ngz34dxnkh9bnTl5jfDL
OfbDoLaERwYKRczJ4c9/mQQodBCuvW32LtsA4yu08YaG1ZYTTLCIWS0gkXgi9imm
c7JwP6DHAj14GEMk4XoqJzydKRiWI46krxeAb9ynYC3AsmkpVBc8neZaRgbXpZb2
WJS1cT7c/1kL0ox5C/t3EupExHxUkNC0Ij9WGsO4tMC4EzNryRCjnyEEOcF4Oq4I
7rkAEZ3dCqS/AXmPdxdq6qv9DtjeAw8F/hW6RHcRBhE5D+w/Knw1ccW45Sf7Uf4P
MsE5Cj7Bhk+OJQcdyCT+VO5hLfVxWcPXMnuInDsrd+kD466tLJ1ZLPMuyQunA/C2
122eCLyNcNy2t17f6z9UaVsd4yj8WLAfECO/f7S25DH2psEtWV7WauCuULOdeMBL
FRuJwQr/ivjL+F/rkSYO8k670KDHfN4DrgiLV39dJfgjRslpTKr5pBT+Yh7Cwu64
5GROB3Tue0zbc+YGD/6Nm1JKUIUv8fR8UuiC0rwr7VWQ0XNQxmLCJ2qA6KEkF3uE
iGZUaPGlEGfkt+3L+CYdRj0nfAKYmsa7oqVWEUsGWHFJ/kScPretrl7AuLQgMoCd
+lWavzkypPa8lh3LqkOYj5Saopu7zh1itIIi172Z0dRcO21TzmOFPVGOOcYlEMaa
m3jM4tStlJxtN3GCbwFJqk0XyMf+q7yMiDNvUbvbJpWEBSEbQXK58mh6NJbXOcW+
tHRGH/TNkR2rnHyA4MAnGY7MRe0SSgwciSEVdL5W0N6zR9aImFuYHl/Ewjvxp/0H
QZmv+HGXQzUFZbp0O9ckN8hAsRvudrps1wvsMGkRs9TLk8n5JqTJjAghHc1XxLZu
KBJx4kUAuGMQGhLOHG8+0EDXim8Nrq5KU3XO7r0gHWwCuKQ/wcR2JE2qK8AwB3wK
cVZ3FzJft3qTJWg+/P+Nhgw4r59b25VPXEHRQ8N8q2u3uBPUku2kgw3Nxz14ZQCM
lzZLomYOIlPFg/dE8Fai4qV7AM/98EQUlnLTxpI4nbj1ldhh4kWdjub1qyZBonL4
mYwMKeD9F3lNkVMom4XsxosgF3GVb6x5xUvGHwBDUNt3BPu3HrzlGgvW10qYQuMN
py3b7pzjcPKexDg8AbiWiHl7xbBiyb4pxc1762ycNvXIXCcOnzdCMfP7+bhI5pYI
1Z5+hzAX1fJJsSVUp9m0CziJBDiVF3UlgzGQ99r2YcUm8a97HdWqKtIudujMXO5c
7b0OV8PRjkGMtc92uvAZznI2TCw+k6S6+qllBhtHVG5GTpDgH+cepV1DO0cOnB43
qsIbpjQzd+fdfUwQ84RCFcgOXkJM3ulgjCW+XQ4Oatn9NfXnYilFf+srKBYa/M21
lPbk1bu57FMmHmluiMiQOZcfqmjulX7vqe/imrscYUE3WTHBkYcavqPSULGR5fnd
kF7YzC/6ie54RqD0HLnitjsbMbPDLPq6FG52ZrefEg0+3wobkK4Awkd0uuaYmVI7
i6+F2fhbdJcb4D1pRiZ1ghpnYronsI5ibaKg6BvHZqN0qmvGetwBwQnd39c3Y2sl
/5P8gZ2OegBJBsnzPw+OLslvMVq7AujYUOV/VQMcdtSDXnw9XMIln+EZcvNmEN8h
GrhGjQ4H1h6rbdgvg3pHLnIfAYijVrDvpoHdPDInGfFRykVATccfEegspf/H5+5j
KhonqjD6PQwYnt6ixqh5SuQjksKl0hEWSDkWqvfjdFoTEqBVEe33Zo5g/VgBqd4y
MOemQ8QqY3y7uQ+Ww/EGLlclrpL+ISUuixiJerPb780zH1hDOMZZUu+zqc7TUGn1
qgVdD9APFnqZ02H7Um1xf5Uus1IsmW/GqaUr5RQBwQV6DfcJs2L1sik6e7JNhPE5
lusfLhSuNnHVtziBtgxqp8l2jhjDGsiznyqT7KC4hvYGHmZszry+88J7j/iHzm/v
RnVKmJx2PmPhrHfjqHRKzwLYXwu3qSzFZnSW/y4BY8fCaKEihrJuBDnoXrpszFwH
PIL97ATvDpKuCK4fi6rfk/4rZdFClq6nGlJRDeVULcnZGKmqHL+I6UyxC/Lpz37n
ZOWAop4DkL/0st4Sk4382MA3QosNLeVNcvReeZrS51QvWNeYuTytkhuYZrURFD3M
DKQtY/vGs8oJSzekPiWeCc2r+TzeRMk87dyKe/0A8QGW+HT6j2VgDylICBwFjJlV
ZWy6/letPi2QDHK+hdCkoqhAnx815sQCzM2Jj2hYm19lRJGE0NwzoGFvVrvzkkGL
qz2jPdQ9kKgvi6WtjVCuA8zeDchpEG4XCXjy/LUpaJFK0JnHEmFzXExwxCzU5/vw
fVCbOaLLx3EvOZUPATlrokfgAcoDh244iqTOxA7SOGcxCqN0U+7WTAX9VHNa8HAp
tao8nYQPctfdJDAPKPtFYcLUFJRKQBG/vIqbklhEY+wRSm/P0edhZKH5T0dmymZi
Jefv65V2dUSCcUolScpZ4+ubYfVfiO2gOWbLJrbwLIG8veV8aXvQzC3ijeuBs+WB
BwaoHmj9TVtAoQ2afNklIXEEb2NZmHL54DsXYl9pQrbLIdDvDyKsArgzKnII2GON
jWtkKbImUO7UvkaU+4eBdBKfeC4lTTnLy1UgBnMiZpXE6KAW8vsA7rDhhY81F6RE
jy4YMRkJa11NRdpVReIqUE46Uq0VJTDgiF/fw50LitZNrtc3/5oABigkp/U0DY7T
rggeOJDhvgH46+ss64tsPwZ1+RK+2cFq6Z3JOOEbw/2NG8wGCBsfDMbpnPda32sr
y8aXzSIAmw4u59YaFO5Qh1mViUMRv+g6FfNJsSezWsI1Dnv1JZW+p0RFgSu1xEKW
eVeYgeKHHNT4Ae7WImPA3AbUsT5aVLSGlCmFMzO698i2qdZBKKlG18Q8UuhW91mq
KrJnlEzmgAqc7MHoBUVii8hq8ekEJaZ1MYK1o6sgtGKSJxdISfqYaDwloDDZHtdz
XTgjqa1sKV2AWbVTIIq1RbXP2cYRcAEpHrFiplhXs4F5K1iYYNh7mTcVScSDsZsI
v73DB7wDKD2UnhULCB0Nh0BltLBRIP5ABt8A+nbJR79BFAeQ3yLh6SK8HO66Gtby
YlvdUhOQ5/UzuIAjjvUOWnJyQE2hGH5SJmekT736T+s7hXdPnMMamMHn3wL18vPQ
vhzG/WT9UPokA95+lWT9lj7i1U4qH0zrxJ0eonX84CLdciLh4xdYZfs3sQu2j3zH
kvXWqJ7sl1z8x06SYGxzdbYLCt1r4lZBKVkPT0j4lvViEkAwajnKCbKukRYSyMcd
Bkm/d2kdTyUjjOIuebaUWfcCwBx6+eFtrOcw8YcjNvdmUpG7aUaPp5kRSpujHYiF
f8FVp+oPyQD7O9NXhq0/fqjDQwSLPWYUd1UdJ/4wzD8ifdgxGifC53aShzoNGw5s
Ad0hRRfp9seX8kKIxaINrpWlvMffNJRArcexAZ/litvkyTTsmgH/3K0RMT1gj6e0
Ik5Dueyfm0hfE6vO+4SZYqDhuVWKdfPd4qtY/6tzr8tPmeukMXUxky6AuCJWoV6K
NfaXNpQPKawMP3RkthMfTgdUyMLxi1RcRrLmWyWZIH5M/yetM/CxnoQ3iCEwx4wM
+M2iSkX3fGIU+qRx1G3U32zryKaRBwegQnwzhKG2lcWH3WTi7LiHCwZXNq2vhUUN
LvU+wa4Wy9+Bwyp3o6CsWu2am5EKOyHYH9ZwX2DlEElqBX5fONz4UbKQIkR5H5lF
DQsqi91W9MGnhqImpqny0mDsYe+lbRz589meifSd+hIeYBSbbHzZ+NnOfdzx4cI1
K1IhhXUWEhaModzzlNAoMPI53hkty6U0E+Ey1oYapmAHiZ6bAQFht5Eq9FBJesQn
vzBSvGrWmTJbL2Q+irF0Oi9AqHHxHD/MWVPX97XQ9J3u6D6trKONauzD6yeL6O4i
pRvQQ93qIldUAAn3mxMvNoKNKoGof/BgUOKJbPHUDX/8g73LrvIxF/eIn67H3Bgf
4UnZUzQE0KA+GlbqsLFO0Z/CuQvvXYTaAjB8uyDQMjRXEp9I2baX2l+ZgL/0To9r
UoDULUQ1PGPYFsZyBCYoZY/luzrgIT90lejODEh0CoLmF0TrwuO6Tdx9U+7qHH1A
YMAFfjvQ9YesxBaIqwDMSYfPxHCCN7MefWhpecoFfbOY4zCgrZgsg7R8O7uEo2ng
k8hEzKg3T50fer8JjPbfk+kQRA0EyFeaBbP/vrDrz3rm2ye5sq0FKnFxU5189IRP
F0qgfIS3I1mxgPF3K09qNBb497Z7F7YvJK4qDbnIfCd5DCYlieHkAO8+NtKfM716
wv8YR9gvTig1u08Zd9NPhz8/jjUQ0+88VOSowwKEezCPSuwUIv9V+1tFzoWe4hgU
xyaCTOZoPvQL0DcxacBEMGYL7C/n5Y1uf0ZcQJzii67aTVTmP8LOF4+GhcL5q2Xv
5D6pvOW86IWzqe7RVX1+sXt7RMYYCqG07v7nPI4Iqhgqm60pybdAglvsJjuY9HuN
2vf2YeBhpHwaC0j0bB6DmbHzwj/MKzh5thm5a+KcYUOeHtu9OnFNsRUTgpsEykSu
`protect END_PROTECTED