-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "N-2017.12-SP2-4 -- Oct 23, 2018"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
x7Js9Gig+lmyYjWH1CeANSF2pXcD01ScsBNWYyz+UseQzfxqvx2hDftibjIKAExA
uSxBSlDX5XgA6Hei0N44gSFskJ7JV5aBiNX0EmCV9rrbExP7X48yvszrF+Pkcfon
SE+eVLaMDfyiLTbX6YMeGL+QSqi1TklX9K+mVUQrZn4=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 11552)
`protect data_block
BaZR0hGM+pmYtUQqFNBPh3QZigJbSWdB7Y3CO2A3FuyDQRw+/fQLrCbullsRAe5b
5AzSN7Iwk0wNTEvmYSY3bG4/WWNCrbW8eXigFCXvYuFLwJ71dS6LNausWbBNI9yi
53+dxCd+vkPlPMhEBRVSUMHXRrd+c93scacR4wRM+qkCldHbZVGxcnqqytXm+60W
HS37upUfdcBABQl0PZQK/Ple8XLzHOefF+nAKsj7AiMHn6QwgCYeLI7nOFmev8gt
ew3WRQDl1WJvOZ5MPt1Ll2aZt4m1SqwHOixSAvoG/Nd/XYScQrLnQr6AbSZbjblK
qPeZuiDMIoOC3VOXTRqLGaXVwZGo/8k8qGG30sjzSlVfkZ3nNwLoZfyyXBsTMxS1
akY/J/GfM7fUJTS5zRlgjZR+1eIoawaKHh5NlBSfr/TSVRplRbEHLFyBBd9ZVkoC
vfhTjnVozpUup8PQMv6hqlpaa8ckcqYd91/XB7XN5N+ZmFIrTsLuWDUk7fCI64pe
turZfiDRQgyQedRgC8gjvVRlVZigu7BK3rZbKHJe3hjyDVT6u20TcHaO1MfPrODD
Z6JNCZLe5rr3+3V54vEIgmKoam0/yOoo8YsslH85kJUM/og2iWra1pmvqVXKqPV/
Shv5g+r0U46VMyYiVUXkd6yjn+tenSMlkPbjtnh+Wsh8Tmzsmr+kQpSItEQYs9oo
DdZ7jJWMrcr+K/TVgSTBiGPUf9ALzWktyRyG9rw8urqFXWFpAWwVwZyooYFzc9x/
27iQEwqLVPdkyJiSywtxdLICXikHR7sQWuJtPmJ02ciXnQBLRHjhm6qGUBf9ZcQa
PcaD6Ti7TvjSZzG2NAkNbvEYFrB+snE5i7am1qel5NW7WY6P3uxFD8/aCdsRHLvB
m6YayFvnnWk+1Z31ItU5C5luQqQwLxIpeqq3H5vpIbPZkh67XJD29OThHdss8O5R
crfG/nd5G521HPCG0VKBf5JRZ2Dk8gqNRVIDZtTMhELrbl59bjdWbqh213oTDPlF
D596kM9VhYmIQcUsjzeKdc79jLnAEvfd1VzFX/y8Gcx9qo5UcsRHbuU/JkUta1UZ
RtU4CqrdvSs7MmzjpqaYr1dnXQGPAp7ZIsiHjfkHtQ4ky8AlXHui2qmMfGLLmNOB
3XLckzHL1JMpEHss5evTmz3w9m05fLQEcqyWGESwMvLluwfdAdjfzyMbKtuKZhz5
5ucDQs3OOLH3kxBvAhMU+4Jk2FUdgNvj3x0l3vlG97SFp1hH/GM19EHW/X8NY2ME
ppqKUiu5u8f9rIJMNdrF7/hFBniRqWSyjq7r+ZD4IvcByoBvAj3Iu0r2ExMOg3Tv
036yW/TVbNqVmOi6PqLQDeau0Pt3w2cgPF5JZUzUcqOGHtIC4l7qsGvRfVjsT7uG
ZsNITg0RMi7NHUvJokSO/L+WnW3efqk3Uy6jkuoYbb16VMX7u+v+UmhdYV4Q68UE
24UcV5NaN/W6Kwn3s2tTIZ6MdEFo0Gb/rntDG+C0UEapdsIpUPk4lmrsve6Q9t+M
Je6nMUoNHffcymouBQxnFbf55A+DCMC/b/lAKkhypaL/RDv+FZETlEYwjvWVRdid
QvA90EyQ+PB59M1D7WR/wiOOhhAP0P0PVsq3DxdW3G+ufigxTnbXxyb7D1bKkKJv
SntBNJx2a8Su03Hb9Try6JcElOllK0YXamiWruuglYcAItqIxnXOlCslddXtWw2U
lTDuFkIntmtFDuqwsztznbMcAiRC/FBo7RCVU8pt5F02SPtLanUJJhkbLtlx5tmf
TrLlXXN6p0JGT0eP7uLa6f1Y8MGRpoh7XYou50t9cMMHKVm8oVyTGndbEI5J7gKN
ue2Qzme3wh0DKtUiamIvRLcxJ+TA5XtMP6Cd44So9EoiOJuKJrkwaS6O2qRQRz7Q
OYV784cbrCMzBmOnXCpbNhVqge42yiomk+J/RLKuxxcRCfkA1XHZX02bkTZ+v7yY
QamKhHSVpfjrQRyRnEwmXd9ErVo5ydoMKbelV9Yw2G8YRVBkWu7OOBtnOHej4Wuq
iKETrQBYABBsZgfHkcSHpOGWfM2p+0oqsXPkqD6d5rtUxcdEPgLpmjmdgj6NYlT4
GFZzL+bbFDgQlI4ORX7+HiM4FL3490D19ZOpIb1ScgE4p12Jc6gPbwBdzNrr12n5
l01I0xqgG+j4DKbQf+z4nb1KdCiyqwkqAuFnLsgVbhVDriyjs+VU69P7CoVuur7P
g/55cVRpKjGkAFYvaMAyPzTKeq3o/V/wpozKBwCOqsEL2x0uAak1UiYutUSgneeg
CJjtKYtphOBhEsJVH0T9+hDhFY+yT9yIsK5F9a9uEZr67Vz6m4amoeuG5EqdVupA
mt1O/2wDQZ25Uv0eadyl1QVXgBSsEJeMsjQrmRvSyn0JAZY+Qv4Dxz7asCfnNETn
5s7xBIuGeMmsF5yeugMoRUhC006KmSub5Afs6NhZnATvFzTQEM+sup2Fo7tEO/mP
+u6JcHTcFH5x634e1wKi6Ndq9qM/Kjn22CX+jklQr77uau8bqk0CjE+nvge2PzAv
2bH7y8fGS/cMeCSoaGhRchKfVBQ6MryhvWkn/O2WHuRTzaZRzF4f1dvlHBy6d+Eb
yL8eXc/63W+uyvx1prvAPzSu44lwAh4vhiSK9kHHjE5mU2s3DwoGIIwGsI9FIWHb
k4cxRh+61b26gNM2qtVDtmdWeH+EpcxO3j4l/ss08wGdBt/QlBRHsdULdd64k2Id
TgVGL1z56Njg7V4doud7TOjNqotB/2+ey3sPDrzknN3IrqzGw9bPVxvZvlBcimxS
RAFNyTfZE6siWoS9SltcicKqOGUraLMG02R7HuEEkXaiw6CFXGlRRMtoR0Xe4YdD
r24NZoUlhjuuHS9u31H7nTpmLB7dVDpIUyNTqulJpiFLXg/EZVJizvw0l+NW0F3K
VSjVqamDw4Hq8j+QneVrdd3BgLLHY4wOv0Q4Ln57M5tFEPeW7ZndbT1Jcgy1jH58
hmvilQXZHjOXNqGkNnBGZahTdIgLRDnLHa1BIUCQ5pc6GTqaRWcU5B/6RUWHm0vJ
vg/qqNJieQ3fAS1aACH3aFN3B9s49aEb0MCZ0nJH3ajuffvPzfTljXhJ4fBcZheP
RX0rs9DSh7DANLm+5Kb4iXsLt3w2DKZl5xDPTKksK7WI/4FfIBXxUMvmoV4aHKbY
rE7nx9qyxA7mOI9Hw62V5C4ZXgjeEqYdUwWQQd5sTkI+KeSNZogxMtItVNKciLGH
cwuFeuO2XGItGjsnKEC8s5p+TnsAtEvaI+74fVZPSCfXAodBhXfjwxSYGP2kNHdz
j81dWS7jQMcTj2qMQsDxOa9MBhhMmtkkvakFpfcNzeKjt2WpTZjDxUKh8WoSTBBH
RxhjpigiVyWoZiyybUIQGwMLb+yAxhy3YkFBs7jKl49r4B3I3x4hljI96ouygP0a
KbYb5XgVL6rGeZJ+0nAJ2vNe5GeIlcl51iF24faWp8PMH8NYCG6mU178Z5/KwI4n
dZJ5pngpthsq6Rit6+dHqs29lDS03IqlpXcPv6eYfAsWUDQBV+B/rZedTqDvSd+M
T6pQD2I8C9ETMZ/JLoMo6BncRijIfqmxnuD5iPfSSAI5elvyrkxmiNE18SifhhqD
e/WsUYLDijZ1V98l7o+XyfsaAjEjjUKsTrrPLfK7Yi4nN1y6bZyksfgoCID9a1Vs
5nm6PdluvlUfTNtQq10VdeKR6BrW0mrV/Br6W6eack/HhJxS1xcPiCqAw/pOoMPz
93GkAwVzaLSOguC6OXK7yUJ5RZEKNRJuX4LygyjFNszhoWDb+pNwJPgUz6uV8pJv
Eu71KTZxljpUrK43uNClCBmO+PmM9ACaoVO3poSaBknN4+r6V1E/dimVfLc/33lw
X6Zc32a/IKVH4HlTplf5Q1c3RZYBFWMJiSJEB6wyuQG9WDcToOtKRzSdgi36nOJs
wMliG2PhRTGOcb3TphhYS3AO/95fW7tq+GiSR8KuH4NpX3Grjy4mLRGnEuiOuAyw
AW+/NR+2U30NiZYR/5sqyaEzcM/5CVy7GVTBmmv1rEWoOie9Glao4GVUTwLIwHup
aSap6eSlIb/WCMcJe99YrLXScgdP8jXVQI/L4zGNIDi7LGqE87iobg/Jt9RBA+pP
zeZVUsJE3K4HnCxjdvIYfxzFDhWFHcXTdealsbRn1pqusQeHYHAp8yal5OmHVoWU
Bt6bEHL5hj2HgOErzPq3CD04G9TcEUo5b3hdr/q5dC16+TLQZDWFrP4duSPgfvDS
cPkfDqbFoUTIq0pVUf/MY3aUetkZf3Y42MSh1QEeO7qLf7ZpwdNbIzWX5ee5f7hV
lT2Ukl0h1yzHit9WnHcfF5uhop2CeKauQwjJt70gQs89JfpUqAgfV89H0Gci0rnK
7Mc18m/UHgd+ECcIAvWsOlKrokxebITEG+0kaqdujq9nhIt2hxqzi7R6L7poQ2I9
BIjn4HfCNwyZxtJf9M1CtI4vDNyU7+7k5QAkPBHF8zmvqJfWJhnXOjb3x6Dcmj68
OQMQ5ZgwEikFPej77mTIfUmwhSohdS91+q8LwmqQxYJAleSuYUXdKE7QNUZIcBeE
s6aceZaD5jAETJMhQ9Iiel1O5D9iRMvZen2hEIIQ3Eu6y8JhKGs2gLcEFJ2ps61S
/uK1ijayd4+NsOYTSGZQAG+W8RPRFSmz0P9ZtY9rWayCRC3Aobem8OKjTNPcMI9X
w11V6ScG6u5WABlzYUzPYbC9+As8hdDnRJ7yt8dcToEq/82SYB8uGpDn/V5qeGpg
n7OQ/DOt5rf7mugDC8G16jKqSnwhqAksZ9jiu6AHnWieQc2qOnc8g9jC/34gDM3h
2QmSyjvLR3suBhf8ck51GoiP+h64KVhf5ghfr89dbE90B+FJHEV3WfKYgWFBQ7kQ
wa5UNQzD2MnGYETNK/+naLfxUr601Ygmalxifccw5m/oXP3Za0SDa8aRMPZmUW7n
aa1RAFT2X8riD+Zdknr7LISLwIbzSqWP0HiKaPKTZ3GDD/iiVm04tV2wjregvats
E6nr4+DZvYPGZexHiszeh/oMqbzH+BxCBh54OGUyvxAkjwfq+9NfIq91DfP8fdJ6
rG/ilnB42POd5joRmt8sCJh7U/dwr5wfmGYjmqYlUMmEphq9l8414ScIJ+zT98Qa
KMmPJjCX+90dU5CzM2GyPP6pgSK/pKmH2HZmvTpevdsvsTD7OgSGShl1vc9QmcsW
QWUq8iifGOMRtIceD/bZwXiQXNgHkUQQmDUsJoNIEFys7iW+WViWLjecxSUH+guH
jev5pa5+ho3CFpgyHxiMTetU2PazBEste8g6mbEfsYX+C/0PRzAR/tSq8ncbRAJ2
5H7pAhiYfDnd97q7xCBiSpQhRZBVXs0yyVTh1BdElAFijUqgmZkney56lGHO+wtP
o2PleNVtBU62AB/6nijz72L6ZnZiSWjpfCsBJ5FZot0xTnnsriJXmpTvpg3QfPnP
i+X6cFyvkb/9plbpgxqLwk1PLYC51Im/DeAG02a9ir+EcT9bf4ByzCSuPVACDvkG
iJxAGVrQLQa472HmYDn57Au/kdijmcNkRed8QcnCEts4ZAWTwiKjbkz+k/9vrjT7
NgjeHpk1m2xcEeyWd7QDybOHDqyx7/1kmR2rlumYHJa6Gw0G9I0TFoO8cPOF5N/v
nap6lvcNAz41ntgCdB1A+F9vn/nEa+ahSJMxEl40Ecwdyn5/qi9/pi68UdhpooUk
yczS/bIrKDpun9gUBRcFRF1+6j1mZSQVh+e1XoeLT8jdvPQoaE9ArAW4qLBmMwRf
/Qv7utPrd34dirdFMxZ6Hd2Y1yFfeGGT3+E4O7K6HqTu9XDC+LGrerZ7JyNDHEY0
kcXuTPKHfcrQiuGyWBFCnjbi44CbNZuo5ZV/ogLn/6hBd/VK7GmNhNiHEeUWCRcr
5RmQ+EAzyOgGwFTE+3XxRPrzVVhmQKcXhXaBuXr4A8g0WxcVgJsRmisQ5ssjYrSv
+WAajkSBIFYNV9mQCVKFOeGUBv27y8dwxCy72PiTYKN5B0fz1EvtaTFCLNE/tA/1
D2OjCz2Lio5pckaNglHzVj1qCFnR2mHSmoHES2HCKaIstu5XjWGHt6edhBH4ziOX
2z2UYKnQ8KPU3gVCxEIZONwH8EMXWjQLJh1EwF1RFUB9mU43HzC35KNoEElWXJGq
1m1D0XwLUDKoQQGLrOhvCWkc5YUhQvT+Y9th0pxJxfaZqUPugtvz5QH+8jZzz1VS
yMLTfZ/MsuBJKhazZtTCPv0UxdBZtTSSFZve1wNU0LMc52hYH0wowoEPqwBD7184
ty2O3CNR9dYZWFiRyttN1zTs+eZZvPwNXK7wGBPEz3ItQVM0EUPD6ZUIi94jOqQk
TTzVboNOfRwdfLSFN977vbY8bYXARYZGHxQXygnIUmaPlfAlecIzPNHKc+iLmmHV
768QEecke4vlK6C8eIAsQO1nIei6uPCyLROXsfMEuJ+AQ48t/7cAtDHYcfABdgt0
1TG44fa45VDzUKzdWg33pp7UDHqYN9/uZdI3Z+5eq7z/XkFbgj7yJhCRlAi7DroB
HmxhEz04376iRuWP6z3klLE/5nTY+PjZwC8K+sYmrT/IBEosW3IZ6RHQbQugdr1A
23j1DAMFtujAPybUy6olLLaoyBJdCqOcGNpdR0fEYty0+ztKF/OCRg9uSAG0ACoc
rRHK5XPvnFnJjolkIu2XMUwfMTb/0I951sWu+o0XKPgkbLiyz7PjYJ4jt2PJ3eEO
gyGlSxS16+rjwwgWWQ3LGkrEUPdUrnHmDAYnxzZF9fmTO6lTPSSO9MrQXDUhZSoe
Q8f9vVBDM2HrJoWE9o1U+HRSYspUE+l06TPVXR4liyENGOgyXzYdbuB4dvnKRgSy
LIxl1Nnu5s8VfgqJ19r6ggtTUWWbfK9aSxdlJ6UzXHD7duGNqayQ4cYbhCJD6zzf
OJg2GGUT53Nowcbl+/gg7giZLbfYeI50htMhuxYs5pnPOAwNLhxUF0iAWxj/xJDJ
Go+tWgsu4bs8zeiDn7kvcdFcE2Sh1ygDQtf4xl2frAXEPFkjbt3MwuyM5Y7FjXfq
XGprX/EH/cRKtyMMN9S79UDgGa47vA7tt9w0yH1K82x1LB9Zq+U31C5xEiGaJuJD
5ixdc5/KLyJACIiIk9ceCCBmzN8BN6yey6r7xqHlC6e7a0VnvUHUEmv5rb6Wg2cL
N0FSftJYWBG13BOXBKFcGD8VLGjYPuqAmgqRDFobmzqydgoztHhIQWUqIjl2LsLt
pI7BZ7YxQ6fETExXm0C3thWvDzTGzWr5Am6U2eyj8bInXDHwprKWA+3PdVTIiVST
HyPlgqVSF2FGkA4mdWMPJ10Ork9XqGM//JoYo0rfZTa4cupkH+/dvLHamipX/vEA
ZfkaZZ5PXkQeOnfZfT4aiKy90k51yWflyZRHMkaGw+MMvvDgbTfqYtouKkpviRrH
AWvoi4xlwXO3kFI54D4NLhbxhBW6Z34+vRBBJSHhhJH9FXxfXPCQkurRNlBThN8j
/6vu9F9GtolU46V/AM270/iCQ8rpsmM6KQWu7OK6x2Ls4SQ4N3/42uYCgNCLgHyt
qlu5cUzqIl/YBZR9HMr/f9haXIJ6/Cu1AY66R3zZq2dO09XLN5NznYjw2yi0hvK8
BXLSoz8jgh24rqlvG2Js3KLysvTzLVVa0pdMhQJsPzKcGJJHzTkFJOv+Vu46wyBI
boKPu9/TUPcPqRaZIoUPnA2NCXZJ6zxdGhRkXS604mbSiWHP4OtoDIjnmOc0xWvZ
+FpvAS7tXXKBSxqlTDjIeCfkzZwD00YU3WpXHKhhPbBl1y+IME9SG/Z25+wdTTiL
xKuTIwy69rdH835oBlFJaHTzXGlD1gTKev04le4hg8WsIUjeV0unyR5/dP1W4wD9
ooTwyE9qgKXdJ9fXrXAGIgg+R0FWOYGVKDzVMB2LqjlCHDdoLJ6lWgW6PL3V3rQ9
TbrtjSJF4crR0ihhnKXAhnLsmIN793SylRpZ87i7qLh8slxIf5gasQ9bgoBmYjnr
NmP9gdU/0isUseFl0+4rlJftF267hIKyHuEqwnvnNORGnDppXajCSoMpZcAYDLVO
oXMOysvjUlGoQZn4DUj9NzwpBeDFoCdlIkHtZwzOhs0hoB18+l79pGEGwomkgaGV
/VqOUkpZ8woFgjXBltEo3i8x0o3z+IqAY4csx7J/PYgI5fhxTZaeX85Pu5XBH78s
POzvZJzZ71EEeWwC57e4SVyQR/UDrmGM4EasBF/HWOj5sOynSFAS80NFzdrYZ4H7
Ylb+ECMqdkUujwj3i72RAqsgqxa1J4x90fOuR5xlw2689p9v2i1p4lBFogqZ1HG1
f66ZIFqxvkSdgqvgzevBH0B3I6kHLdS/6ko1TPic8CP9cHN6v32dAVPi6NC9IDyv
xQXfzFCzkfHmcSjWf5quBg2WKCqgIsZzCZZgs0UvbaAtTxE+AvlBuwp24TwR6i17
Wj1eXsDaQiPwY8ooyQpCIOTzBdNLIrSY6vGQfds7Yhi7WXUn0x2YFtWr3eOKaNSN
DZI8Er3nw2RLyAtupxLMhWrvFh4Laog8xTsApFFW9rkU0DDBBF5vFeggwhR4xbWm
hfUzKJUP7jpG35xZYBHjEJ1f5UHFPQ7+abgXHrtWg8LKPxwQChy7pHfJpA0bcbAr
//i2KMKDsMyRXL9eqRuQ2Za0E43VazDPFRJww9fI399DE1KbcYRLpMqDA8Cq0qVB
fB/6t2+RZ8grtk7ei+9yK9BHyLMdIOBF/7tv46jxmGhDqNvWbz2L2Ptl4I8heChh
WUpENaP/AKCCTNhiyb2WIgrJ/vyzAiRN4Inbz+//DYQGltnvyKU78JtSO/SZPdva
ftVsjZZpMo9fGQLwzXaqtPkMUlvZpimrILHhovuoOhfnrU1dptX0ORdi0HO2/soc
4igUUPp/G8e6Uns7nuvJxljBXYHRgQsVTKHqk4nE9xElKsc2p9GncvXSyBSzAFJc
7+SUQCBWi8GwMGftpigovryOt2uH/TKldoKSCe7k8Z8cA1jKWHAs6zmrZebPQJHT
dN3HPwx+R09iH82C3Tcndjt9PjXg329Z7VX3n8E0959Lx7g15RpAWYP5uc3vYcVp
mviZMNgP+Z0G6WCbEKrMOkkYFFy8eH/YY+KiKyzMg2wdA/TUUhPYpVBSAwDp6zW+
ypgVL4fjo5giwfvgHiHtO79fjtMuJ+YtJzU7C9iOetu6JHF8XwPEt6VSmBHwc//B
eev2I0331HMZ7CDqdN91LF/hFLtyGlbFffYUlDdfA7zfHYzll2MtSbMkZufLKWtp
kokQ+0YbFpiZZPHlug3ZPOcuM3qv881qNyqTb8Sf16b/HguVZ81j/pTj4EuLCg8d
YoDvv2Nc9f/crt2JEoNI9mRBPZ9rtpstWYaYrd25ZGyZ6ZruTV7ZTmcIhs4Y9m8Q
bWoyfRKisOYEk8fBtGpYCz0ptpYEzRfnU7WKyGNNLTgfJvYfrdJRTGBYbF4YLDT8
oyf5h9mzcZrKDtZ7+WRV5osYmBoJGBqZ2uMP1RRUtaHxmLAyP+UjoNdZdzV9O3if
envrhwcX25E1VeycbnDXOUT1AmqFCqilEXNsqVr6asBmvjd9kvelHKk5GjGLwelW
zvcsZsja3O3nheELawhQh4r4Oyp+XhSUM59FAufDR9HVuOz5kR4HIJm2+DtP5cYd
Vdw06fRmHEEUF/kcleX3T3SOrzg+YMt/+RSfI7N23puwC/+Oq1Ujl6e7teTGmkpP
gYk0mkKAvVdOM7ggBIOtjTYKmhwnIJ79Ox9YYfQNvOSgCmi6CGzGLXibe9iU508G
EPqv3+XV7FHZh0VrrKcbOr5Ra8DwkbHRdca8oNOqfjA7DnnwfJt0fZB2gbxXLqoZ
/xyWniIAYSNzAZJ4m8XTo0xFGayciLUEJ9paVh/w13Px4mT9KKQtLeXI6Rgf+IP4
oqP4a92StjSqADhfRQ3q8nMqWPb6ZsX7uJWOI6n8tudXWc5S/Q75N6/KmSNxnf4q
8MCk1gfd9blgsmY6WtFQiay0h/X6IXUw9HP+12B/VdUigUI2xseQxdEPJpPsFlNq
wII8RBAa7Vi4aXes8Kvt9AUHjwMc2FVPYKX3N55GPEh9pEw9DEDWoO0cN/cXJ1vd
Dh4C2X7rnggB9O2iM1BVFR2rS66oo6cutfITqMwwzyHau+lm/AJ2YxMYMSwisrCT
rcpEguOeeTogUegWc5pzV+hLl6nfxyICYuYBWjOq6/P2W+C9ssSI5aaGIcYlXeKn
3MzShKkCDTWl6+uEnqpaPqktnGn/2aKTPMbb2R6DbvWhnNlt0tVVLn7E1CI6A/dP
My1rqbsYJIHuVJ5yQekkBe4iCiK0fWWb1+/4co5TIVmCv3CHNOlR6qe1xfF0C/qG
xChbGJdCXEC7dhaEUlBue3jTE2JsMKktWXctPH1roTLwYqWO6iViWN+HVaLyWtGR
riOgoFA4IFkjJGA6cW8mVORRVjj0kYMhTwRny7dgb50CDwsQYzIXhHJzeURZ4xm5
grqCe+1Mhnccx1wft33LK60tFMnVainn06OW3Ms1yUM/glpqIH6QxzfSK6kEq/wl
+0LeGZ7+UFIjPVcwp1rL5+6/5Yq+3xI4JOXX5mwVB4dpjkQ9BVn2mohCB4GHNNHZ
dWroFtP/riU9ZHr47ul3w5HRi6BrQO9L0Y12N++psZ0baVfwE/EiM/ggwD3I2UhK
RmkX1i2YbqWWlxguK1kblmPFLyFR6kD4coxRrIfjiw1ESUjhBbVsDJ17us5UNeoA
0zGjRSYyQd3U0k8TH4Xn0/imUXJEefluieepajKtAD7dF6M5RHo4sf3WMNGf/XYy
mM4ycaqaC42AvsmF4PukybdizBY6H+TtLX0F/Qs/zUR3U/SU+2OclNqF7VhPIEmN
ayhlMVaFKR5p3BKCJJmfABcFCCE3KuAaQCEzHSRS6cgNxMsdvXWwMMGntZmZFkNL
N+o5q15g7k+wrhSehGsZx3rIh++43jjS95kIVmeF/bNuFqtDwbTdpf6OMZMnL7B3
cG7dqxVnOUH+zQ6//qPSvUxb6Ldkv63/JQ+pNG8QVRohgzrGCBG4d51rIBcY3XPS
HYXPK2smQYwgJ+5IRcLfi5XSSbypw1mns7Vx6jy0W2m7Mad0wbg2zKXh9HcJ437g
oWtPEU2iPA9DK4CegCHTDk+w3wHwX4z1HSq8Nx2R1YrqV/k5Kqd0nHJL258+wk1o
nmUxvAQJ+IKlFFPwYKl4RqOpifRg6yik39nv8YvGd4TL+aHtKuu5CtLZo17pWpQw
DUi7t0WQSZG6/J/VxBMvsx8JWF022OBz4W+RRksC9AXQ8GkNQcV87w8si01yTkR8
4P7gwA6VmU4WUn9ca5DjrWytfZds+njNxtDG5yV6HcvciNqqyqz+w4E5AvSYejtK
Fc7djHABnTyF3Or89bZorGouPIYXYIX0rhWATD9weNOVKgBjb4qTwyF98VRIgOBO
WPjjhoq6rBQgt1J+kt4OsXbxvKFW0l8/EoFcyyDhBcjFloFEc1LuaqFUVBRlINWY
tVpqWj1lUhZeTFdOatAG9RT/62ZrnAVsV81COMiaJpRoLVNCGO68fqv3KZ0TC+C8
w2xIwQT/O6P4CRJl3LO24LjrIazYkrLncy07o+5lAqGmUqAYLeYHvu3173OrSTd/
0ns3qD4JE6Jzdqyr2nBgaVTs+o60oukfuyYoRcO9G5IX0VLGrw6uFTqPG7KjiAYn
3Owc6xuocj6uTFjbuzr53NS/VguQFKDeaeDu/lyQ6Og0uYQgt0/HN2x57jEemf/j
0zIzzXytVwVfaLzY7YXmhuadoXZQMWMz1niq+Vgtmuvl45Y62VTsR1b28OhurBSn
ncCn4x7+PaSvyuZhZjx3CEpVfm+rJ4woLx0iCc9q3xcJolBVnqAJcT7pFi4fLBjr
ERR6rWJNpLr+DXpuUzZg1dhDd5+CaNx5EVcd45slv5pCJhZblxinuPL+oY9Ho9XM
doPC6AxJa6KSNOjwnAEuPBeS1vVP/IQ1EhHmlh8gfLsVLt23lPz1SSC0EUtkK586
kNWjjv25snhUvEQLZuu2N+I0ZkUl0mkTWCTc0DhKxOHEaOR5lCd0+n7WSiDwHiM4
Nm9YQEDmSec519A3FOXXiQNERdhC6BtPS9+6Lywe3zacBH+HA6/2QD2PCvffV//J
Je4GQ1/qp6x/2f4weOvsi642dzq1vA54gHyDDNWBThgtOi1QKlhmf+nvAqALzDFT
0+OmKwvHjHlk3AlRCdeRId+lX7+smFz3td2V7jwtvISk6cH7/yF0zgnFyW6p3RSz
LlN1DAYqSmOxIsLOZXKTIxAjp3fSmvQnMdckTQNicOoB+FSKibiQQOqs5Ml3QvMT
Gs6kCA9TINZLkWRzEpCrTFOasVwXCyg2pu0tLR6i/cx2ctQl8a4iEYLaSYYqV71O
oMupJwG/gTX77n6dOSZLF2TatNTvCrs1B6dk90OqINGubelPzwc2YUTHRsO01qf+
Y6OAjf+JU9xBdTRtBGSg0EPDkn3YWs/54KtFVxk7ulakBMYGK5TKUABTb7qxyaxJ
W2S+BGp6CFZnXC0Bz4ZHjKx9DDMga8kgbqoCQt98vXQN+pzRPoIgIkPkfw1a9a0x
Qv/wwpqwlom86IJhn2mXy1ysOf14b3ss2lq0Jy8lJ25F/gh0g124Can6d9HLZ3el
1XbxQ5C/88RpGJmm9VC45eZFew4v5XHg32IcfZipyDIXGl4BBRPIT0ti+IMGiS8D
gLiPc1Nu+eFDfmnYGmYmiIPd+CpO8wh+5a/POpIkqQAncTJLt0JZ9sKwVsLRFKaJ
9UrS9h4gznhU/2n4ZL2sPWy6Q9B/BxwqJFNZPH2QJjIlX/z+j5b/IBHhkuAzQrFE
64TsoJZF48Uh6fU0pxcUxNH7dqJR85BgkeskyGhOkmEif90NiAvHzOvATBf8do7o
JU1DyJiX07GgKsW+xl5+c1rHc/wSdj9AUViLvpYgeGhd5l0fWdkc1X5QGSOqoJ68
SwkV6hQ+djX26MuIuaquPGwwjPQrb36SOutBtamj1OBlA8KC5SMUQKQiKXUn0/5X
mp8mVNVsebyrMfJFnhKDeBnnqsAXuQfd4Nx+c1f5lskBVvSzjXRrQPzlcYbw7fpa
0+IaVht0l+2xXUwEmqTDWSsdUWaVa+lPFvaR8xJVMbeMIoo79Ahk6ZGe8Sv4h5qU
uUn8EfT5PNR/MhXmVBCvv0pf1FFU7qnFmww0qWQI1ptSHr9Y42ltHrlTqXKyzMBm
deQIGaIk2x59x4WZiRq8BcouPmhZIfeq9sdwrtwfux/5O3Y3XR5c+HngMqqyWYIj
lgUkgkrTFFk4xT+u8Kzkh9STVEFxJTMYGmJcm+1ZegGdVoyAF0p3wbQvxViykNAV
wTwHaebT3s/rOLtqj5+yBeqmiKibmFSTpp69IHjqnD88GFKiS8wNkpYk3npykNjZ
YlbUED7EslAs0hcMawiRjvqqqdDofyLFj3jpX2frBJsjIBORPgD8bmkxX99VP1vZ
3sO4muxGfOIdjNGmt3WVxI5nHY3qSZIf0ZV8ihE9yTudsiKHeXXA+S+1ocR83Vvs
ncmQ23nrmzlDFQXXVDPLwMJ9t8hOEEt0A1rGgDeZntNR/54ItVPXZM/JtHaXJ35G
Tvts7fwTIADkSSvdKmTYsjSfo2ZwzaQ4HX2zYBejFYllqyQdRgHTyOtWLXufFezK
nrKV3txJN8soRoLUJkr5LuNBlzFvcSUzVo8E+NgFuVwUNDR6UkGrTBF5d2P1/3Do
aafdR6d9YizwwS3mydKRZH1l/sMvcB0wl5PhlTRE2DVf+DoKQBv0+gJ4NjU0NDXs
birqq6fNQe4fqRjlb7MZYB4yhkRekKb3XiYAAbpFY3dZtNizSsBSXBEKtt7RktR2
SA3dd/0qT7DoDh4wzGRmJjz0tt1u6TbU+FW31vlXYcUmhRtHms0mBNUHbBb69+lS
eaSCMJA2/hWB1N/4aQICHkAQmnW7bS3ZdgNGgckU5rN30/lTvaRuaBqSTmEmH6y+
WYHKhFiqa8ALmOtI69CUjdRvvFo0a+AXMSX0O9D3GYmcTKqjNN7aQRKYqTeVQ3j+
T3H8V2ZA+GeNi33C6mQ+F2u85LAefYlPmLud93LZCMugP2/ja9xqPka27nI0rjiK
NUaogtBVWRCrHunzAo4+ciF5k2F0qMDwIl/YKqiN+fuyANF3jDRrlhO8Rhja7ys4
F8hOnkq4s1vwLq5d1Lit1227EixJYmdktVB6KlSoNrMkgKIK0RYU0x5qzka03usI
dc3QtFbwlRwgNWZYW1qq3WtHH0ghe5QH3nBZWLqWVUCkZY7xm/qRfTOoqB6YrQLE
WuubtFzkoAZpW9O3swdN+QUy8CpA0FwhwQ0lTSiyLg06uoXWhn5l2Bqax1HsDgt6
0/YvRkwVX/37uTFrOBBGqcSiRN7igHCBQQk+bl+rGnk2RdnlWD0RH1Gk9MNcx6ST
dEFuzbepSgpoIqn+zgvdwDE9nyuH2ZCKc+nf5DFuPgZEmGvcpTj0INa7Olwip4fu
G8W99NB3wVtoXenUSz6kGAViOJqCAHGATXvWbD6UQi9JjxAJoS0APpq2i6BEhlW8
/Xd/stA8PeUseMg1a9SEGvC1DTabvwtR0NKMsR1XI+2TQPsECJMHSRQ0flqGPia6
jpRYvJj3nnMGa2x0nG85nraCJJ6PJE4w3BU6maXwANHaqaTBxb3FScS4eeHRzeuZ
xLD0+LdWQ6ZeCLMMH+NKs8S/cmitayimTNHv2oYiJmhF4Yu1DHRgvCXlVndfmux8
N6OJfnxpOgCaEi/0C8EFEjYEhIa9P6k0pF+d8ZIXMNuu+jaNphrGaaYqeFsy+MCv
Ygug5k1So+eLy9XKaPq8TIFEto6qXNnItJqeF3IbHIZ3ZpLJLKuKO5g92pCRFkqJ
mmF8FQUTeCRlZRsPNYjyhKF2B1+2CQFtXzOEhxUMd+VYOlEoE4rqJda3dsUos8Vs
UykFMkAHaBq+AxwYL8mZD73QelXkRyh6ew49W0UJdvd5KsS2li7SOnE7dmbQ8kV9
zsY2v2rg405eRc3i11oVtCVxdVYbvS8X7QYq/8YTa2m/u37hG8ftdn3pcdZnjk+v
7CFyHF5bXL1MNBsC0Iq/G+TNpaSDtrEP33nY2h9s/GEgRGxhji+8fjH7UTit75Yo
dqVkr80xCQLXap+5zNROh1zLt0SNJnDJdvFKyTYh5wVT6vC0jI7+t4sl2tGs3QYy
2tRQnBy+sDlQSDkEBtWCMj08TCgH5FVWdw5ITFU25OMwF3v0oMR2NJtoIysMx3Zz
/pZRoUYLYrjutHAsVOYOS0SG7TIp9u5UTeZLFVNx2Mw=
`protect end_protected
