-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
kxDq2x+b3dl185sUuBVglsJiYjx0ZP19fQeWe6f61E7WFgrKfpY8WoDR75/Wh3sLrrucN75Ogztm
Vnzp/PnUJRxVE06WW1vNHD1solPa6WFXLDzgr/+/SRUMjel0UonVqqGpKsPHhFzpJd5YR4osr0L0
1QAidd4D367Zadu48YO4EW31JwQa+dI08VmmW7wYx2m8plx83DFUwJ0KOQ2guVEcyNfdGbeJLvr7
+67JoiwZX2d87faeGhmYj0JipOpKc+C42x4RnbEnc3nvLIN5NcNmn+vziQ/XEC12DGwjBVRuYZ+c
/8SwNyT1Vmw2/0ADkO1TGUhHoAUzLtlwUdzsbQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4672)
`protect data_block
vL9GefzSMjx0qlm2tYQ2V7RoIGluW5SFCJbp7OgT6vpjsMwN8jVR0Wv1pIZlaFWOiMSYVL9gezdy
GUxVc5kD7jTfqjFcUi887nJoiZbn6wwlsMiY/QyvSsUBaBmPwyLNrWtW3H55i7d3sxB2cU7EEt2I
m6FndT2MykP0JjaALq69N2d4Tm4AJD5KoJO98faJNwomhY26WfdfvyqtJzcR5pXGfxd8HFHtanXn
ebJCBknN9tlA48md+pLoio5fWg1bSudhQndGrwyRucbw4JiuZhZ4wzA6HMLtvlk6+jMrV2A4K4FB
if1RJSYwqWFyCsmsQskJxsf1UvdcnQbRbQALPsJy0hwnoZug92SLfxQ3n9qj/LIGUcmY131umPmi
aQ4Bd5mlobEI2WrvY9JMIpWgUnxEsZluwAyemCmEosdBK27yicko2G8/LEPRBpi8ZbZPmL+dEGh1
qjCpI5PEHUoiHMCK6/q96+o+Oh20kS+Ix4UVoUtDJ3KEJHrlpCC60iyt04+eTQP8f/Byr/SaNhsj
X9iFTC3UtY6lppLTjMvCoI+e8q73B3z9vaksBeAYSihfL0YihBRPJGbXDumcdAoAGnNv9QVa2mM6
2BHhmNi/Yf9DES5XR986lpuiEkFhMiRZOeM37oBgg/uBAeYE0s4AAQ3oh68BmAmzk2Yc4e69AiYs
tmzQ/iHY95u3LiaWHJnYYbdtt1l9TKIavDwfoqxsoHM7AbWmdtlUGYfPYf9/YTm76csK3B0BtW4/
VIaBsrOtilM9kr/ENVpZyc5DOOk5s77THrwacgUA5+vJrsrqPFH9ho2FSch1i5iHVfuXz3X2Id1Y
Z9hvoDM5gINvhPwybhp6KslSZLW00tgNxhyiv+itZzYUrSHJQottFAV+4FhhYFvj0TqihixaejLl
2+ax6a+qsPMiayGFUZhKQ/rgpK2NIQL/C742JaM7fh9fVpWA1Dhgkq2JfYDQUAjMIYM4O8Pi3yB1
D25gtjmY/xhUTst526Gba0LhP165TqEEbHNUbH2003/1i7xQeJsQTJLFDI87XDFN1ju91ELF6/pC
yCeRdZZKnd1uWnTALpHAqItGWd0mkuS4KfRgkaRBjXe7Nw0EOrWqbL6Gs0+lb3GoDAf90mQoNDXP
RS1OQgZI0l1+2LJBTVn6aNPSCq+OmP7xDe5lFOG/UDMlybGoF8gf8F//O5Ypox/l5EmBJgYTA5c/
qdEKo6UN5SKpIp1m8SJUrDCp3wq2GZJNTa45od01sPLPA8USkP236kkfTGcBtTxCiz2t3O9qOUmS
GleuG9gZbs5YMCzS1ZNeJNGssRMAIjsZANQGq20xQnRDF7d8A7O8eAZ6xVR8Ug5ORysAojvVGdRE
karFBQe/N3wwwS4f8hCwnxBD/YBY3Kx7ygQ2Kn+TSlYf7XFJ+qFeeqz33xOZAYf6pt6qzZXMBPzY
bXQoLZ8GR8iZY/VIa5Uj9dXYE6PmFajKIXr2awEjbHu8HNTao6CcD8tfE74UchuyuNMOdcB1LShQ
2qRfr80pX2/e0ynubcofBUBUvrgE7inF4zPEBSHMxMFKQqFVXb6oJeSqo3vOv6Y0aVQT7G61WSjd
jIeI6Z5bBZ0+2WqFMBYqMM+QjpK0bF8EfrnxcgxWy2MxOO/S+nbmPGUCfvpC+m+QGz+HLo5QnH75
PGG70M2nloHDUoeOcrFHyEF/nC3QuKsU32hQVAeDxYRLZWr++vO4WmfRFC0we6fUcjXGjmuyDbZZ
sEjqN1ZDdduPjqAGcVC3z92W+7KL9GQhAQ1EqjAvewEPk0TlnfCyL2VoTRtj3nzbORN4ZgIGUgLz
oq5DC52iDxTdm6cB+w4mO9wbtgSH/W8G/wAHnh0tP3oX4jj37u+8JoPy1dAHT/m/FbSt/ccrfLTT
DRQdmkfk3PCsV5aDhreR3tbm9OcR1+RYtn1sHUUmLw/MMuzLI9L2yEc0l4q+808Jw/+kzAC5nzXM
Tz/b9RkTdADh1hzmlgN5YPwbheNxN6kFFigYtMix/fOaKzhGTQcd8DDTCgPC75RaOoF42J6spmZP
ig64V16wuGkcBC4W53HDv6DhA5EBiewVhtrZIOMy3dhkffOqN42/sGoLSEQrR+lpiCzViBIVMKLb
4sATyvsSaX3KsjsZB2z/dNhkwVQF1mvtWqqZmFK7oMaw5RWZta/CaSh9MFOs1Ocn5b/H2EHqmk0r
R2sIkfKKWr4a1ZebaU40zR20uhdE8WLTL8i1ipjUtMrRFaawbOet0krSCRHCN4ggPM+SotbrCOyT
Mzsudqve3O5qVJlf6OEqRdVKVZS2YgX1jpd4iBRgvir4OHZaxMntZi2Y1/hjv3KYtZU+MOy+0ymM
BNmjMqhxBGNBn8sFCZoiJQJBVbBaQnpGaFHUplbv0NbEXXdB1BxBLqVLQR3Z1Le2cFjGoAdioBY+
DdHP+lPSGdOfnwVX8+oZly+I1YkncxOAWvi8IccSnekVT+cUSTMNy5bNuBbXsmyR8OCnDWUjqw0L
UizupLA1vTAyqoSGLX60NXM2hNGdBU9IEICi0/6U1iam2zZ9HuIcVHVoA9gRkJ0YUfvT5dQCTK33
CDfpsCdXGvXLYCKFUEogU1s9DaqKXYbo9wUufD6ri8ekGtyfPTn1zktfWvIi+x040bHlB66xt+yR
jusDKMCScE7KfjBCk94SSdwchvk2LbBsfnAzUzxAGzGq0t74OzjRVZdWD3Q7lnisKMcyoyEXKYQU
/wOip0x9HeVxxktM/c5YPb9OvX7Qrix8ILmwHVy06zuwFm8kHj14r0Ot8Sq/XO/vB0q+Ta43Gktl
CXlqQn0FLjWZ3z75WE8kuOpAUPoM93bsRG2Ljxcm3oS8z8phD6/qlmySycZXjQsl1gC25zBWCBA0
7t6uTr7BXiN3/NGoGFed0Sj1Qw3dw1WNssjojVCmzCiHcxFRJP9+zIe4ZhRILytlxvJegOcypbAO
FDhIrthevFbj8wib4IpwfofXHwgVK1LhwUXPpQC+HhEJX1L3MEi7Rkg+pjq5/F2BPULbRoyNYbdT
otJKnOd9pnffciki5BZfWn2uqfId6kBem4Fd8nXKFOc1qvzPUfyMDWGcVC3XOy/eXWpCVvq04b9d
7RVy9PFdIJOBL3+2uMufCm2Oali3jT/w3wPOeMaB2Q6pQ1myABUr5reQ8OeLY4BzIumrlHpqqM8F
ez1J+ooWz+O/83huKZhaBwqUciiSxgJ5do6S0C+89enEF3u9OtOBK+SMyJ335dzbDFZ7n64Ol8mZ
+MvmEWo8cSBKLJho4qjFBbdoVLbCSmoYmTnj17oZMwz+pvJLKi2kal8RvC0OHQt5GFYznrLkhLF7
cTSAzO8t4dmI1NNkUTNVVrCl2VJXXrw4BUSLthc0iZJ5A7BiweQXuJKuieuLxLj0GNIaW/zxCtD+
S4E7z6298k0R2ptDA/CJe9lYKtKA2pwJYXcdZnJbDcweTKCB7Z/DufrYYDn+elUIRGgzYbP2V7ff
qxp2mvEgO7q41Dg1fxxciAqp7EXLB2mEIEydw8oGwQg8yPTbs9pKfAoq/RieGa/8L4AOr0DJ0OIq
pJ2D8IEtuXdN3VHY50mCqfS0AqHjyX7EospUYixC8fbgn1KQlU9mxFtKR7mqQ6upXyErE0jxXVVa
XfvEvya8u4zOXiwq5wq2b4iuoLXOgvOpP9i9GXCFVwwIcsbkG8k5uTOZhmAquyjJrDOE2K3Cn09i
Zf5rZiM+PfTfWt+MRZ03Kfae+pbWc6MrinjnOmtXlRftFUCTXaRLlUzW8yFiTAcHDpz7uE5Hkhix
0fvZKZxUR9LpIyW27krrTTzSpy37qhtQ/NSAfiUHBVsiQFmWZjBOOsjVZKVsSy7dyloZNskZOrrP
emdGFoOxgfLoq1Vr9TLXjsweRxso78AMWgaCpINOt7S0M5mG9SO5UfwHcGWeMV7XZom2NFVOq9pa
q8T5AZIrkcElvGDJttmkWP2symAqZG92OQVKRiwWyLSn3mj5lBRAanLRI066a9jGSZlBkfEZx9SL
nRb71TsV3LdOOEOXCEgOxCV2ocrloELYxM8TDmnjqPE4pABnDqoPKJJYODSbjI1X1rO/WdPJLDox
X2NSOztTmXkalSed/1h6+jY1WDMCVPckMg0DcQnHCoWrYeV/YGYsR1b44tzLZEdPKzvrY8v8q4kw
PQ0Bgqz8Hd8dA/gBl8jqiDQZSRRUyNu5Xm8UdYAahfpx2pTl8qDaaKVv1hfqT51qNDPEydthyWta
ODUmVCJvYDHQqpukC3s11r3WNDAw6BiWdRhAWcJDD+ZeUtYmCdYd0A9uuLuTJadZ9e+p6mfVhAg2
nBp8IrxIRfmRmMsuBlXQ4GpLKp0JyOlnzqiAEtUlyLmRbb4cgY3pY289fg71H03iq9nUOln9p05A
N9jyQhDkh6R5bwr9bXEOy4avTAm8g4m5ZyzX0r5tOiBRarYTEAhL5pn8JG3GQgYoASqOgK8AbNmD
lKaUpcu0riPog6GTDjGzZG8YQkxkb2xWtci3EBalchnoMGC1YRpt8Pb2MSZ0fQq8t9JTeimMesAM
cLyUWlylW6X0NgHkZ2g2MuqPB4eqHmBQ+z81us4DiowAKAhkxefaKs0nZlOm0CLssnI0VoaUyrCz
QME9K+3wUpEfDh95lrhCJZIW7mudm6/SRSbs1j4bgYbRDhFWL3LjpRyKCu6++XqDBIXI9uLwoxrR
Nq9zXH90B6S0DbmuKFfb6MiiTEFeuoI0g1DawSD1mEu2Z1aUEU8HybFX70fyouuiLYvPWATVenjM
vzPs4BZ80r2/9qYsp0LmrYNsimSS4trn1cVoIltTelBavSNZWft4bgXjmni0kpNGAU6D01ZBaOkq
bzgIcqqbta12bqAahoiIIOqhByStcnJpF8OX0GqU33Gd3WmZutF09RqYyoHLT6ZRZ75vJC4ClHSe
977h6uDpFbkuBLyDjRZGTzT0101mN89iMfBjcNmLxFIxjIFyPW1OizIP2TGsaNdIyNtbxcbLv7MR
Hw7Lx1mo3Z3NNhQbbBgmUTdJFZ+DntZvXqOoRoWwWbE21b0s2MBGzmK4xDKnh5fv/itV0q7Die39
KtWgvPRNv3eL2KRpFEhKjydmFKObjr2VEzCiBk6KxE6U0lcbSsQln6/Yi26WeupHcQbL5EzQee3o
XnH36e+yVtDR2zFrc/GoLrUudEuAbxIuahb2rq8XXlzW8a8SXR8Q8vZqdvfvSkJTwII6XYUj4Eke
6FQla5+C2rd7EJKiNBgn8/o7YnffboyBkwCJ+Efs+lOgxmbULN+fwKvA9TnfaCDZlcz7g7PrVMs9
NFaTfiZ414FmVIB7n+DFwuzxBRuXuUbjVTjnggwDOj6ifVkbsA3o+qLb9B9khTA5Bdyj2LBCieGE
dvlyu8bn2PYhjK6ldVEgZ0bGNdnN3gzRDemuS2MWuPb1PPkuxCgJIW/7cWipeqlcNYmfE108IlBw
4sF9lk8IVcJMa5gHtS9m6i29YxwovonF416WK+DkQGmVtBUjODcyYhzduDLfD1eqzfhu7dDpbDrm
91jkdCWyAGiaMmFbMowjVQv2hTEiWghHUL6FxTXfxz2FPeDGjYPj4qIDsw1jOTk86x1dDFBAxryo
vDRcy9edHvgvqWMjuorN8AU6x5rxOklcojTB5DI0gBoouvId2n5EYsNJHRgJ2mj0Ge6PWBjhf16W
qgFLUVM5eptOhUDmlDo2xs8bBGj6H2qo1QMIG6DuyuBSMdbZQB748GnQRoIc/ZrUOMJTm9AgHaaH
dcgY4jWqjce0Uepu61GXv+/VfAWK4Um/jdEK/6iPfNjQxXrp2Yv644JUsZYWZ1WVE/RRXpMAjFoC
VI/qnD9paiXNCMBopPacCb2Cs5E5DLmTn6lux0QqsTWu3jKwF+ElfECfKY6JgRpPMmH3IvXzCmtP
Px5VJt3QRWI+HUnOZVphLyvUlh7AYjX+W5nN9GnAhHh3C3FuyqJqjq40WY2olGEI2dNFd/tb/ByI
bmCqgtfg7JEpc69hsRyWqZCbSfCYSGhIhhnXmfJWTWtauXZvEb2GT8Armho9jpgRAgbut1ufBOi/
SXhUjUfs721UpJ66gp+mYxTPm1REAJ31CjNmjGJ5PZtBjF5b849bUpc4RGAGJLdlIs5HqIXaL81i
yE20ub67bCorx0TCY8Wcchr0gbZcfnStaGxC5msagnjYIdtbu7wSMVCRTXWdLOo+AB1yHOm0+w==
`protect end_protected
