-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "N-2017.12-SP2-4 -- Oct 23, 2018"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
VCxkLBqHWxEheFfcDkx5EJyDBHEuZ8LuR92NLRHyZiqaZyccZuLv+IAc+ql3Gyb5
hB2Lc2t+SPmhQwzenoTHbkshRsQv2Xmqex/Yoip5zJ4L2LPyD83mje7nI1aHt9nI
0FO7ThjA5NjSQsQaXZc2D5GNUEg1GLGbic863k0Sad8=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 16528)
`protect data_block
Bqm0v3p6dSCff6cvHstHXpyFlCvBsgZs8vD1LBkg1T8Vd0OXq+jLJ3ETorAJZXZm
NICMofM0QM0rI+dMMyebJYqs2KDVvgIEFWFp+E8eYM5eBm9AGXOw1wp9jzYccHFj
jPEmCPxb2naYoUR0uO6f26frTnO5TWgcWYy+ZvVpAUyCNpeedoE3ohGXFHJCyYbH
wypR7dI8ptihx+zMMaKPKXx562LWm7+xlhnBs7bdOUFd4UhIWwAO1E7Mr9bSx5hz
eOTblJPJIp6uU+suERB8mzudS2Xp2FM4jOuIwc0EC3h32VtGQm0bi33GH65ck4cq
gOQYh59lQS6S1HdL1wNkO/kRtVGsGk1iARup0yxWzQ+zAIzo/UCvnrLdUae8VdSP
Lwv/KB5UZQUKUDO5lCTadDKgQGzQhkkhbBjgqtFYs2SVha5JrZPwihJ4b4hIahdx
LYuMd2/K/+ud937fcEXnRKZ3in4gzblnWYtWzwllzflvU8GIs1sIz0Aht9qYjfr7
v7WVPN2zhtTQJKt3frG7zy61Elxj3aYsAPUZ6+hOa+tBHQqoc4LnrAis/CA85vav
wQkiVkzkKeh86eBg+IAIjib/wYkLSXn7FwpMCC0tqXOPGiBUFLjBFYOqORWWuEnS
wLDlimwbYZzf01koQlCzXD4lW7IvmY7rvhih6+K1I8rUZfl97KJh7osbafNabLNr
hLj/uEDwXT7G2KdGKgCGCk1ZEtT7YDS61EM6Ek7Khyn3W3CS5vmZ9oTX/uD+zOuL
vEPtGIAD3C+DMNJWY12SoXdJn7OTVzm4lY/TfY2Lz+QyP+6PsEjFcrpyt89Uz12U
s5yUJYilokYF3Z++fe6lJS7uch3DWn4T2XswsI+oq5Is+27K+d6FxOTlKZSmn+Hh
Tmo1JoFlcCPxlWuKqL7A6VUD0M8Pe7BKGo16bmvIkZ+qpjNAy8mgFfvyGrCpNA1+
5CLdPFFg1ZQkjSQbgjteCOR0cC0lJibKs9NNxkj/BxCZpQ8PVPChfQOAEERcVdsx
LJYNX8dorXV47pDtkuOdi0gTKlZKIHI9pXeqF6u/5B8OP9Ao3GrCRt2U0ed6gsg4
4XtiClKNojPmfcmhoFjZ28CgydCtQkLOI3Oy8BR8dK6yq6yQH9oVQ82VNwrStcai
LJ9Hvr8SNY0PfE71n6tzO6mg3Mp8vj4FYIF3Osn1BuKWxpclQVcno0IjlvNs66KZ
HtPQ6XICDN7kEuI4Ogxefuhd55Bk080pFNtsx05QRWSSHha2lDArO971CAzUaRqQ
ysRX6z7EiI7UCnod438e4FI4pDkakp9Ivg6KUwYOmuLP0JdcLFI3iMn6Esqh03wc
YRykH17/8G7WHb/Hzm7cK4woloTOc8/U2Epwmm8HVrqHGkOMX9W6KcLu5KgR/wyW
999edXd7Am6rM2g239mnfisgWxkZM1XHgS7lA0g2smFEJ/RK7N5B0vSM9XlIrABy
gYaFICGumkrqe4sqfowCHiHpu/4V1/gOKTlny/gebE3v0HZTnoPnbiqldkjimZI0
FU4OgPNiNmgADr/FpgOc/SPYa/3dOSvVdcFwwWkQZV9jqF8fPLleyl8R4oisqRPY
tbZWmFpNg+n9MHY5tqSTpymLxdYqSNaUmNQexarFCRy4oUItv9MPWovqgrkwli7f
N3nvxjkPJgVtJTBmj5nrBKt8ky59ML4nMRDOk1UFi5S5EWeGvuWlGKzaMGR00Kan
MGENPLXk0hMKSGvkp2ldI+O/es5v7VepeNiVMh5IaBLVDNSBi4NQVl8jatJcOzyz
jzzZ5RHnWCq2UHUF8ulwVUPb+3BrtSN8MSC9q8oMrQDtQCSSdKu09MuwiGsqXA5G
hKxWPuh3EjDQ9fuskTdKuPwg/Gt2+yRrsGvDTDM3DNLg4Q8WD+oEYHa91olr+udF
qP/GpPiIHSsevfJl+JiYfvEGjzE2cMxjDG8FI3c0l6dt3n1WBTAd9eoGOF3hTS5x
XhA8I/Ewpf7Yj325mXa4f5+UoEpn1BzS/doEUnOVHZroLjs2wa+qdzREdIa59ocO
TxrkuyxwdolJiSDThzjhBgIR+TGbVOUTOi2YYemFiN2ogCq53d6EdLqzM83LkQaj
wfYrpvahR8rAkvj7EN8sNRwAdthG+fgOfwcOi7P0bbQrhTofWVu8t20MCSpRZsCO
r9ZiGf/bVnK5nOmLzYqPsOeMOVV6BHjLPfT6HD0iMeib3+BBYwz5jqb4y2C+F7d0
2HLKoVIdirybiChsk4ywxejUhszE58eoeomMH+VGT6XywzkGWVfGN9o2XiyNpVOc
Eel2cRJGOF9HgNavH75L3IrwuG0brCWx7sByn4qVpMpAblnNDOIyjqqRIkQ+NimU
aWaeDxkboB90TpxWPGfJ+ZUyc5tDr/DaS1rTjxznygCTQ+UXXwNblrfHPs2YC0vh
2M142XV39dqXe1n0fhPo/kqXBHlDF/klqzsevRqRVswcAbQJbFkT9D0aPeQK08PS
0vVfYFQcfWRBM40lS4iq7XwSagoqWqph5yNyQw4hayttIx5TN5MK3glYQC4QJcIA
QZ6TPlLxv4glPFUBgjnUFj8H3bvLy/vjbDW21jGMNOr/VLFkaxwiAj7fiBmxN62M
BuZJmFb5K7suzy/fbm5xL0VL9DUySyQvXYWyGhIdLE+raKVdjbneHt97ScZAXmZb
dvIQyvHbxI4xFFXDX1lc5rviaoyKWb81iDmxLINRZxaiLb3xF9FDH5mgO4bcEi3+
JH011EHwQaFbSG3CufX/bowdlp7FWpE1DX9wJ0i/oumQ+eDUCupqR9FmiendOS66
AxeLJX4io9GyDYCOsXk5wRA9iX1rpSV/HUOOm4NdkszhY9RP/7eT2FGKGxayBvRW
pN69CR2CSi5GDGhp0Zs3GDAenHOFg3G4WvALW7F/rJLcqb6jgze6y/MqPGSu9wPt
W7QuJLIXAwPGYxtW+LZcdkfLG1Twq8tsVqxuaaqm+T+dMtg8GcfKzRErC8pEKima
Rx3MXbM+2uK7ci0hFfsCH5IgljwXlOjHO2KlzV7EL19cWg30Jzj6dwpaGC+CTADv
guGQkIz1j6vuqsxfTNJEnSWBQ91A0PnquR55SMgZfbRYUVsXcrmCnRhU61eKV0I3
OmprprEJ7K4YUtua+pRbxB8XbXkyRDNWpPxNhRn9CGmMBpAx9Udswqn+M1MicaUa
amLsAO8wntbshxPq1Q199z+r+ilGzJGBq1J2B3LZYutZPTWIFLvOHimws/QYKAj9
ThtoEgiFYCl5ky+P2h4higr2b4xMbSJJ+deDrDE1KFiaZ7T9glAHBNaXYWpm3924
jYniS5DAfOHFD/gpsxWWib2WzR9Tpu3NW7vTMwxfscm7tNzMIoBraIwOqPuUPjXx
9k5ybstahZnrdu0UbEVD6rErpEwBKeEFlrH8w08ze06BpIpvIHbjlfbV6q50Jhy/
M4esoMZ0NBvjzFziyMlDL0Ccuau7lHL/f5LrF8BLad6U0m0J8AbLUnX4+ZliuWSh
bN0Bo0K4tvXJvYPqjMqLlY6HF1tXjXP6bTe+m2scPJvCREKb6daaZylpdA3lcpJC
lwScgYwaU1SREEJwMfPI1+uBMgFP3ChU615ULTMuhOXujCNNYS/AA2i6cS+7ceFn
0yDlk46Z0QVJtFSPeHIYzCOoWuEq9vhj93MBNUudZjH/kBiJFTQ4YJZP0PnPE35z
9m3+S13BcWfWpklBzthZu1jnZ5BI8qnmwW03DKbbAenw8DrGpLOGg2J+97KbX4XY
dnZkD3ohAJ7BLk85TwuX3SeIiFE1YZER75p4gzyw6iDK2dK014UWUMtNe2Z1xliC
ea0eZXys1NyHHciOaSowP3v7Gbzt6Ua/1eSRnphnbq5fJpHa6BLYwIWzudV3OZlk
nLyOHQPqxGgLPwRbWGeTAQUif52AOBLsgAzU3lI2M61muyUJU1bJvecCZrUXOYI+
l+dvc6D1F+9qdV3oeF5cv1sPJN3aPT8nQjaj15qjLfqkNyBv+ySI3C1e6FzOBAIE
x/kAiyoxAG/abzxDH2PbSA3IEtZz9KP1jnM1Bg3P5MH8zonBla2wp/YoUwJCdJ9e
KbSKgsk6p+wdH7ArLPhAY9tYOmtkG88woGsnR5EGfj4Bgke8HJfds8zGxnxij4uw
x+X0GJEnog1tM3ivR+3nCFqwgc+GZepT5Kyj9zpbSQ1k7NYM1p/mGLR4HRRFzzN2
xh+3z3qmTkZjfp1jlCg7sArr5DiqfcHMScYSlQqGnwbB9nUmUjULxTuSDV+33O39
I/o0HUfGic9Vy0ACKfsYatea0TRy8/78YkFwpslc/nizPbcxoN9lB3E+tbaBKQh4
5M8t001VPBJ7ttymaR4LodNjdSoWm9e8ufeFK7mvzNxr4yhi+7ZI3GeQnPiCHkoB
i/3yg0kU8uOia8a0NVcIXCnISptWUDsQxw+KERnLqATGLP7trXYq/nUsgr3aeFO2
b2GWeuKt8K7Amv2JFeqXxEhhzB6ct1aZyo90RXM7y2VL00PZH4utJsIPR7qFoI5M
Ktg2VZOQrkWefKrVUOrpp8MZUdEXG/+t1/GZHu4OIs/wsIY68sG6FOArI2rpQP//
ZZ79SkPg2tt5d9yhDGKdPI73Ke917roSVmaG7xiDtGgHHJ4CpUjaMd+PaOXoKqxB
7hXi/KLN2mSTh1HVvREnU6jiRaF1RRB5AR4JVe1VcIf63uh35HSBCJ5dRKXJV3F8
MBKOHbCoFfd328RM+Okcm/B83rQCwZNnufu7eXRlnjWbnkA0DnmKJJb7jOKYQbt2
NuTK7QCLvXsg9AQf9iZ9GFeAHJxXnJO9TNQoH2ySouyI7ajKJxOQtTrZD/6pVrer
83uJr+wSV0rComr62SNpkHrnkacDuw6RBOD2FzOE9ThOg235sVXnQKGSUsbP43Yy
IdWGo7j0RPDTMyOeGx0TyE42hRctU2DFH+Ug6DdfazcZdssqJJq1IP+Xki64lXDT
C3ttSct6MsJYOOQKiz8uHuqa6zKfVjXvx3ZAfUaPh6Jc5E5VKX8hr+MCq/fPHX1E
zfORb0aJeQeL7ntiaqerN0KqhPYxodAQM4E4MY+JfpU1qtScSaApRIeAvlbnKfBv
mQS6Ubjs7d0oL93cczqy30fGgXamMNWR2O+WXvHyWldj5d56Xud/1bwOS0WGFQ82
04uWVVt0UTfzO1LgtWf2BR6WJ1k1PmsKnQz484a8oLmJujY/yT2AKPQU3MjNJ26b
yKpbUjXzne+P9oV7Ovo2jzqYb/bYMbRI76/KYo9IOepwkfYWaMUAj+xRvzdeMSkl
diEmu+GXNchzwbRefCYR7i7d0ZXNL8YfrJl4nutLApT9ECBdrKtSstNHKrQ+42Xw
nQTme0vMARMKrcL2kSeRI0xZRHnnrOeIOXGLYyBnJdYK/IRzcqOzW/mc5zZpPwIp
zPchqtvnY/1AktoP9GPsManFQswEn6KkpUFYqEgbaU7hZ/pznW68mnYJqCDdWsFd
iWKRRZez5qVdNf1mDQrH2mjyS4N1HBBJOXBJ5TfEw8EqGkmnBbGtVwrACyN7FkXs
6kSiZwQZG0bYYRK7GQVNeVVJwoSRAu+PeEkm5dG3bcz7HnkeVUuzi+SgDkwhsUzn
/NLx9KSyVZYNIWiwoQGw9kt4CDsX9AhGl18lHD5KRYdtdtS/zctwrBtPI0mhixvl
hdRoBqXJH7MHzRYGRiFa2S7EEsNE7V0dpywZo/oU5QOn+up8isWi/ocDHVRbHIo4
cF+QU3RLFlBRkrLapZSo7V/FTazoGDbC/L5eK5Hp6YfGj3iGOdwWrP2f9rgdlpMo
t3OIQ0K5fxh7ktwSjrWh904cLIHJlQDvuNsu7DhMcd13TTYZfZhb9OEMEQ/cFhvS
+lJM2N7EYldKZ0E21i5zJsYE1E9TE6gWMAbm3GuSw5Wi0xLLFiBQC07qg+MoWxVr
QIYKhu7ry22UtjkMJwAHlNWV77Az+3vnK7R/zSlx2g1fk0d3Bl8tivDx+rJwCyqe
jDaNMrd1fQEKiHmFs43LcElVwzoFeVIZi05BnN+TtHfNbRnaXqoZeGcQubtRvR9a
E0qPKtldkxnWDySvARyFU7hZnBg5t6LNwSykLLCkXARNDHq7Fu3OTtszWJ60Z3nI
uCt35XE5BxUESVEvto7aqP/Y+bjVz5h7OXQFfXH39HkWeZfdplhSgRop/2xtYIqG
24AR+fAqmbxYYt932BzF9ueQiH0B9dUE8YyldA0BUNXMwqJBJlDfxMoxyVu6w+4/
47VwlWeJlocLw7HeCh+gzij2QuOmCN+E1yEX5HAgXq2vaJ22Z7Mi3bYq2Y6gR7mD
RzUlnr6IbkImnVoKVHmw3DLmUFlF1SKZp4WSHpCCV0xNrtnRZS9b/sGDqJqJbumm
Kq/RycO3LA+F04MFmbiHVPWlpYjB9nK59y5XLYLJ9PMIZSHSL/K8hLtM6Z2Mu55v
46YfmOyMhxZh+fyj8VHInFzU6U9Me1EJcBxGkFh8mbisAAQbmo4271zEtzkEVnwj
PtAFUNpuXXnY0j73GCh8OnaL846o2Gzp3Tnee+KMbVGpzy7pZyF1ap7Nk2FpgI7G
XUBBAR1PkTMPRqXA73vpH2VJGPDgO8JC4C5dtf3agpPbEnlyziAkE77pPU2E3A98
cW70bRf6qB9vPcBcapTFaiX4m6W7ZwZpYNi/3JaE5CEOvDSEM/DjZWC9CSPST6Lc
MjkM7mpNvoB/dS1j0hkjq5lpbDNIxhQn+aGMzJS3JSHCJH8qS4JMSgzwkWlg5brF
RUNpLdU/XYTzJP2GAfzDSIvv/ZTxFAsQLx3dbkZENfMbgD1yVK5eNsJSNHkHK5Gc
gw4mSPR2xHtlHS9ixkTvy3EwVLJHmeGgcsh9Yj2ZjxdgMuhLp5YHUol7tf7pclyx
e1rTbionbXI8vg36/5Zuvs5r9KP+jXbjdPHnZXITdlAMVZU8tFwgbOeuQ1Zt6mLh
JT+VqxOCHHjXOkXa0soGj8mKqF+v0AamkSCQODL5ZaKVegPKW3037gEOxiXHJeVh
msBizW5Tsi8h5uSQ7Dokw9JBxKcZZ0zdI13jZ+TOkfMLJ00yUdEAC96dbE1SvS+w
kgQqOADJJyvn0ZBuCLRSYuyNEkIAIylVZLrnQ58+6E4Of33CbqQIGIxzXETFWbJp
/ZoUC4M/JJgcTKJVuEi+PTvlqBJEoFAPee5x/AgJpSScOk+st7mV4+3WT2zaadOZ
FOPvXzgrSnqSRPOXfuq09IyDFmoiIkxPooSbQHYCQBpnEP+ujjBoJ+qkq7tjfzt0
rpnLwSLzhFBLGnHeA5VX7TUvi8qWLdMRscSd9WpYApWWDnp3jR3GZk/AenLAZUp4
Lgc90hA6ClHwtzbKU2vOQRly57aPAodUExmGvopYdnRsgJcMyxEVaLqESJG+ajn8
ZUTSimlarSqR5UEdiKfY3Smgzlt9i4S4Ykm0O8mnz+y0r5RdZsSALtuIBXRozjlG
ZzXcrfLAcBLgECvXXUrN3e+964Mdp5mR+So5NTGbVxn96ew42nmXPwZJnzJ/+fTM
H1de91FrJQwsRlN1gxBbcE/tDxAJVLNGWgcTYGS4Cp9oCxcvAr+S50ZAg8kUdrVx
d1TiNNwwmwR5e07sh0idKmzxRrg8T24rO/WJdDUO1gYof6NQdYaDmKcRxT9hK6mt
094PsCz4+zhVu5Xe8Wv+S9TXiqf2cK7nHHkxRR+RHKq7GRQbGYihoFtz1/M4qApK
cRTgKLGszBs2gTYNXbY9lN6ronGlIUx1YOuDEKG1dsb6hz70P7Eawf3jvRvtSDTE
gnK7MbevGVidpJCoSBHMW2FOvlIr+pQCPO43ZkdswEoh3QlY9M3nO4WhchRyCRV8
vWPLoz53vGi165NIAatQsK2jA7C2VKzJOi1i7rmib4jdx00f9W6vsukIwnRxQQYa
n5oVgOkt2KsEdoNahNBHJrL70YC2vm/pYqRgDCDwPeO2G+xjcX8BF5r9d86aNSaB
3cP2Uu75KrSsV34bfxI5j5ApvTd5qzbCqYTx+rSZTxom84ow9lcPLi1IE5fcz34u
zPe4ArHMcNtAQDG9J/hkLS0yd31TdT5QSdlbz+UphpVYq+gL9VzBtGJok4EALgh0
iifUNqr44NN9MUhPXflG7dl+YcxBatW4Uer4+fl/N2keWbH9z8SGnUcsMJTseFiI
3WuLxscbs/4VYktPdSC3IkOeZ6TSKwVHuR7lbK4lPxSy5qqF+wMPQpjEEPudpTWT
q5pvrp08MDY53gfTQcD6fgjqAFHYTM/kjhSpsWAajhz0v968zUpFtHWcjE5lDmTf
Yzc24vpuOLgjBJHA2WjE+Z6n6d3GG2Etr4KZUpMbgVs2CpitGK3KOm8AolxEZ1KG
AJ+WVbZakoC/sZ+bCl2ovQjboETEcmP9V7vWcA3Yugt4Oqi3zBiyQ1rTveRgNzsn
E2Nyoil22b2NjwaOSivXJlewiqq/QOcDZwtgE3GF4J9RaHQcWATUe1qT2UeJZKm7
iDDtV+/EtT4PxTCDTBHJNBA8Lhp+bw7KtJA9UWBE8vUgpY5CPYDUoQ/ycKfPvk0l
ZTlWzWP/E18ucd5t+vmxm1DVPVNFN4AOpnT6T1EZiC7fhU3CI50pXgxjNz0q/YnP
/51tt5m7YsmHVryPi3kcZS8AX00kzESLgv9gy537+XQRhRZhPX6YCJ2URpEvbAZ0
rcAorsL9WZMlcqOQZvbn4x2OxfrB0roDDcJDP7utHlCwV2+XcdxsgQIzWvzWMPBQ
LTi5ujnrxK4daMcK2vDAbfH8muEpvM0vpu2+tuDPLf7fQ0j73XxSZ3OEIXtGOtGf
h3U5NhPmfDw0jHbVuzfbfzubpUYbb2juoCiu5o0YiW/G0P867507HrUduwKYgD4t
rrzp2w0aao7Zyh1pLqkizxYvqgp8gifDDTs5bur0pq58rOrdlNVEn1KNram13F3Y
j3dnBtCMVc2cP30NfGpd4i3HQ/zHBUVvCN13t41MwUqOy3wVlbEcsVbhQyAhIsCe
6nwBN1SvS5fQf4r8RXNGx/pM2cTd/ckhL0PQCbw65gJZBFJtqKsRdtTdLjRHId9F
1eJ2aj9xQEfW8vp1m2UXv4N2GRwtiWLlSgLtyr+6FEOkiBN+IvTgjFUio3HECGA/
1jhr36DCMiOUMrEizLDU+Le+sQpuK2o3lc36tR8TJZ8Qdt4Eme0qoY27uaG1Hodz
7cHP2WPhhVyNSF0SHsfyhILH6hXR72n35gV7/ffnSEp7t4pI+11iEkWGuxldRSxT
7dmB8aLQkbo01bK5J3QrF7oBCmYfTJWy/BXr7ofMU/pHB+0KcLfckfvlWCR+zKSi
T2FyYdu6BlwgLtCcjpkPRYX+9YUv/pw/CgGEp64gCjy9Gav4NeZNfusPhgjZlz9o
xWX1F3j+Gek7UinbeHhOIUM9rHxT2nwyPZOK81L+znmntiQU40VlaYLNyZBAlBNY
9x5BGfnRpf++Z5SftrAhc7s0y87KSPotTyY3+D37K7UUlHn9n1oOqrz4NWAyijCa
8ZcbUq4GOMFEe+2uF/bwpJyRbCoyLXQJE0Mj+Aq4D4Ru6STN78tRzFhmFi15qY65
xiU56XH6EpZEqVR4zNwx+x3LBL/3GqTtFETJGdbVPJQYxJsmY3lw74pIY289JQna
SdM4epLy0grMjB7NppstvIzVbRt+yPvFe2p03Ey/YHEzHbfoI5H9/NWnCbSjQn/h
Z2dIZIPUb/AQP6OFXg9iwNy7W6EupHBIrDxuVQmgdwwsb+qvozX5FiSnB1X//O9N
ddu8HkeSF+Z76P2dweSLbpKn+EwHoBw2yZQuyMBpX/JmN/2GfwjKzuan7nptWKbs
edN0nUolmbjbePVdxQme4S+zRn6ZtJwQvVF20KRne7ONBuKUt/78/cDNT3wX90m+
EHcFxh7m+6P2h8AXX77WGg+EDFXzNJuMKSx1FbtomLYgCsp8nlZ+efkTz63/RYwf
ao62NVIYJTjfF1BbcHgsQpaDYqyFt1HO7qLo/LYDR6SWN7Sb0ve5uJEgozIxVKqp
p504AYjUS9M06/9mY7LCFPHjru9U5RlVW+xpK8pTqYjyDUo2+r4AuW3GMTblZTfI
kGXfGnWPq2JUMHO+uruEbXepzQCKq9FK+pCYp3OTlZM9cKJb6REsYqBdNU2fhomr
sVaX0Vk18Hnp9toEKoKWIodhlEVzjNGHszIOP/1QNPkprFRSYrLpXgpu/1DhOMcE
43t+pIXrHHCfy/ArraUhJ5X2M4IUYrmbD7cONpOua4qYbPXDaTMmPX/3Wtfez4AA
Dxk4T7qg9peIFg8mUe+Q5CqHtaXgvXDW5JOETfqS+SUBZ+XRSX3Hi8MKywgFdt4d
Sw6Of2jdcEl5zfU7/8HRILZ6LYyVDfPGBc5BcwdUGpyB+BJxL96aZ5QmVngdpoj1
L7ZN/afk5/WB+CmbMkG1c8X3H/I4ICbpyjIITtgJI+bh2ItMmbg/u3EpajrX1min
ZC/xCPhVYQ+IM8wH/IGzj5TQbV4kB5sEt/ZqrSucQcOn6yVbF1qV8FvipHLmz/IO
X0MnJ4hr6yDsK3WNvds68uDWaqnWM9QoFbSwtBd0PZSNjzwoDwvlCkNAtWVB68Sx
Z/gXLvE62I/cShp6XHuEXH607UrDYAUwjWZ4X22R/5aAM1daLey5RECZ51F4LWde
CxojO/LejMMkEP6414AGaFyf5kfCqXBIc1R0g8L69gmOlMN6Y9X3u2hPtgEmsQ+9
w4/PcQSeOISEJ6Qg2883Kq3MFoURrRelsefrmPkyTntmSklWdFYIaiH5BjDBUTov
e0l3MPfYWsEljjCLbzcGpScAzrvY7jdMq3NaoUUbWpDwyAG3fQHteZgamc3+36KS
OVhrR1zCDsGCg01GS7vhqM78T2BGfaZJ8FACBYtn/f1+NgVGYxynvFuy48VhA6P7
Cqr5ltY5wC0Q1fnirVIIyLdMwbbA2MS/I3FgaJGnwXkTqWztrT2ZfnQeFf489osI
f6GC6YP8bE3GDlicPzifhSKSlI9n7xsTxwMVabL37GmSBeI9yTOAVr2az2t/nfD1
zqJSeY5sxKYJy3glvlcvD6c28DgTiaWRevySN3jmWjLk1ie7ShUiEhsKMxvfUu5x
bgvIBMZBcpqnYH6rwTgbkZqfX828GQsZUlrwmh6TgDILJTIxq4M4NA6z65ooa4ch
a54N++r2RG4HAJYELBw/4BKS6/MD7MOB+wzTMaFL9mdqq3d9esDvTu2+9WXyzpai
2Ti0/szsuzT85iuA3lo6sO1aov+UCtRleSutkVCdbQwk6lCDVdzxX5LafdWXcBEo
U3tMv0be20RDwx+KSdoRUCPve/MoX7bWmdJcIXMz+ElGEoUJnCVKRPkGePQlrIxC
fZi7necA4hEzFYs5FDCm6LU1fqaiw83FqMrnPP7n+6KthAeMcry9JdOYBJrXG0LZ
ctuJRFyqs/QR/4ksqlPEqyEXB/uljS+mbiJCtCGDU712IzSLb6zcAQSybQnAt7AM
YxGHp27H59BowGHe0NCaQqrM5TzDDX/28s6hbvHVA0HVjkfiHEwPsj53iDts7MYG
Xm2Rc6dR3Zw/sB91J9rk3ZlUm5+avF2a8HoiFRstoA7PCvc5vvwcVTAynRwE/dY+
ludYoLmKVLa0xrtfKH+//Bs28HtALxGitEF7uPYy2fZd8eNizv72fwpjMkrnCxqI
AXfRQ36rNLTw4Sq85zpT5dKzKo5okgyFdGygxKB2IzAb6OcudSeIvdmjNyE8LOPE
7koVu8fCG7Jp2iMue1zHT5sebr8NFVAgu8TdGw9v2ltDfo8XLo1gtABr2bqP6Cx1
E9U/9JGVS22CgAMVtswnMLyczNdCe4/LTv6gC0rfRL72C7fLMBg/OSYtxthdodRh
PBP4tYx9AS4KTmSrClZ66mKxnHgPq4pLRymX9Nv8NfCJPGBz58LHo1KLYtYMAwG9
eM9ZiiUSqJuII2nqpH8VhmygOlPT0r9ZxsLaoAZKG37tg5oQ79QugEpvIbSqTwDL
xbR5GxcLBG9SvW5oE1kc1yR2nUS66B8bFKjHBaQsGac5wtgasuPjdEQb+aA/fgmt
RD2IIWQsitgqmK7oiHzhZeqfZfj1a5VzDKQA10jw8WbkYrAxQroeCmHtuqVEtQED
1BhVkTYoPVUJShM1KIpNHvfD8xm5l3glb+qH7M1VSvv0VDGdQKxcvZj43AoRPd+B
wOFX/pXG9s0fMl+GjUVDjnyqDnRyv96j0RYAVclCQlktaPFVRxwHK0jeibRpGsH6
MkuGqJBkocpuF7PYV2cecAC6kbkIAiaf+zG00bDnW+lszVPDqN3ntIu+XkRi7aew
+zm+yVwCIRNWy+Zzgm6XLpd4ObZXq7UCajV37n/lfPMCFkYX0t2LpecyzCoPJM6J
zf90hURIzrv0k9tQ9san0sloXc04TuxHGl2N5Bgrg3HPepyOBlEONXWaZGLNo1+w
41A3SyHTBoWFrPKqz3ug6Rh+I9MapIYBxYnzHuWFWvxDSqSyZniiAiFCaKSdbcfU
iB8Ue6OmSGQPMb/0n5NgjatVjUt9CLzKiICe6Q4Gg1dzBhqeguM6Me1wp8qeXCnh
z5Xw0jpBY5BVEVx1XAv7nvdeaBin58tQs9L4tZDhGq08kPga5jgoocbUHSciEGtf
PzVuOWWhyMvX0S+l6T2zgIWMbLYoA5n07xBZtJF13S6EyAKrQz29vE06rddrOK2J
u2lB/+TPhGZse3iBlZCnAKnjUmn7NwyImVQ9kUgKLGANIARFg9X5MlVNpAEi/G6q
SNcIldUW+wt9lMMlCmr0JYQi+oJ+vCxRFF/XjeLChf9fI1+V7bBuCX8I5vOPHKmT
jxa5O8UsecqChUTU4FbKtS8QmNjbQ3DdnAMClGJHMYfVbU0PR1T1AI3acJINM2xV
qxhDqfvo9IV7Kavd7LrRPrbhmjpi8jgwGY9nKbzRzAFBHxxOfjorqgz1HdzEGFXm
dsXx9qsoE/emObXNTxh8XkSxUOndFAA1Elc1p6mfFWr429Ryn6Ptk2mRCWX7izpp
8o/22ikJCyyMT74Yh+pBIRAY/jisz8BbR5uROoRxFD1XSAsi923gzpqawo2U7NN6
P6vBSKPRaguVBcyXB4hKvkY6ibEcBmq36UwL+qJ/pUXC3pKYmP4QT6Ou79BzZahi
dMyHbThGnkI7HYWWAZ7wZBoiq7Rnq0nKfEnn6J/uU0OxcdcL37N+JDhHf0ww40e/
Lv+7uBe5VzyvUilGKb8rA0eL4CTSemr2XkU4GCKBswdcxdsIImsKUEkDYBBp8y/O
+W/iPAIyFbg5bY9QILQKCFMp2yyzwHfsrbA+msUkp6n80tKZ5/lNrzAZKpxEvvSD
+ewA5wZwjJHBNjw4h4WOzJE0ffKIzeFd34eZem7TL9G3ezjng2AkRMam4WZT3P7v
Im/iPaX2fithc5QPAY+jlJZgug9dTz1Jgkr6oAmcYAZk/eutbTZe23L5iQCQVAGs
peL/+xPMoVKc2PE1yvsM3BIyDT6MZrudWnDtetrbv8Sb1BKdDplxfvpVjWN6K038
L6mJvsLD9QtRr0gv75d4yAkbm7VXf6Sg1MRBgjSBnBeCL5uJRWMn4DxaXLAHuTkh
BR88Te5qSj96VUR1s6MtH2czmBlD9gUsBDTEEyDiWu9AhsD4h1JdP6XXyFrXo5HW
Htcm1rGN9WYAp2/mgTX3FaMzYYAyuiiBx1zfGGZAKl15rJ5XMMhjGVM/km069uiG
Mx9xboXPHhR+P8lrM5z7n5uxAGc+VftKNZyK2jsfuex2grwbFKvK2DhLmelViENc
0ZFit+i5X/a38HIFrgCX8nN/VZdyre3zhzNjHg4AQeyQ7RkXOyRxSINguEAf/Hka
eJ+vqv7qLi9MboOmLhcPwSLoiCHslDCbGFH+agCvMWdR67r55gBu7iEy9PMcRntq
lZQrvEAWOdBfApkoL0sczwYLAUI4i/tVqXjvwIZaYCK0OD67ZEb3QpQIyTVWxV2w
1+WUn43TCd2OFSn4LaV46OsoVLV7L49ZWwKy53wh8kfdPtViptHM2z2rgeVKqhUg
/5VTpIOizJTuSA9aEgkqGH1ZUlJULYiNvpxVH8/KcgZLKbKhzSQVj/Fdr1KZHsjT
cL42TbrSXgawRPRxLnketZOYk1wc6VntNI1egLP8JaO3EtDqNrSDpkQquC+j4h0Q
/tb8FFncZTMNTCipXJGeGM+qmB1Ag15yfn0x0ORB5ZsvG5El12zj8x8umVSBAvS1
Yg2aZ91d1iGA6+Nhveybo+AHw/PNl/psMFLtPNR0S11fPKLE8654XKJDcS64eQiV
jSqbxAZK4SL/Ij0CM2oYlpQdSQ+/uVRm6TF+THS0AcvDCVQ5EPAycwhOsjwhyG6E
8gHh0BgT4pXc2LGL5Yf6vNHkfwXOYpw0g5/jlq6I0EMIlXxNRfp5OWV62MQ+kKA9
MZFKeIso4aWzVva71OdO2klj61PMAFT9RrCN9TkgWstktX5Gi7hxtfX65QpH3Fa9
N2s++eVopnpGfkG0OfSqqbmwk72tSxlJeENHofpEfnbzZGKmb6dz6K061KUACdFx
GlNxv5QrNZunFdvfdjklw6oq4SVJeu0+d1YyIB4E+AAhIJLniHbf8IInwmVCrxwl
VgGRr94yMofOghSXyYIILZrv6ydEm7ie5nIJjpBTvZWJvCYO/eNtGFDVFdkuj0ZJ
NdIeRyQU3EwBTBVlMVsYJbx5cRuh4c9s3tAlnCgveuoB8tDkOoj2pclJGG10vt2N
ing/hLyJHM8IFnzwYogo4rm1wDRvmikJLfVkaksbESCRGJ4SCYE8Vee9ii9QB3EY
X+DzSO0Gs2Ep6/XmbNK2NodcBsdTNK9J8HlSHltw5li5tFSoXrJWDJctyIZ07X5m
Al0CpdZPxlJO94QRC0B+7MZo2Lk82rUsuSajsaqRHjz1fbQEqfP7vFb716VbGXh8
BM6FxAf/Od+7txt8j1yehDImv4gECAmVPA1+fQvYtxwkYZYOSh+2Z+8YeIemfK9a
MHdXyGg8LpUuf+MLtAgpTl+e2HsoB1J/wIcbxC6LxPFy2vxizIhLPHFWkEZMVwtX
QEYNetJ2WeZYcIDKBGxFNzX6RPeTp9cQRpG66YQYzdszQ/v7Z2V4EVszpt7cTOpT
vg4vSsbm3QD2fLBA+uiKBsQErdW5CRWyKLZ8VpMybVYx7Y2rIKqvXJlQgv59Rhke
OUoFkGoj9IY9idZ4652u9e71t0mJLTrgxEgl7Wbyh5WIfxhxA16lO6XGVmhqWKWX
ljjuo8G1eGOVeHdi1Q/oTncaZ5ZZ1mxLkIt3H+eqKfk2SXFhI++1xiDvGxtkgkri
9+3paek52OHDAbcw0PpRjCgJKw+0JpAD6/o70MkHybbr4xK0BWCSNcv0wdZ/i2T0
2yt9GyxJosuvnjCCg1A2r4ABCKhwlBWEy/UXcqaVn99tUA5koC+3b6Xs/aO5PhPS
PAu8Vorv0jsedisa/jLdAuwU2PXu6a1h95whnZP7I+98U5ne0FL5MpqJ5Hh3CNSx
frBWZsDk0jpaPXuPcpGpNs9wVNNMic2oVqJNDmWCwY7Ze3okNwf6f9mOtq8S8gPd
WRJJpVPnk5zDPYirHfs1O1bI4a67m9lbR8CSmXxgKaIMeSyngauYNLUfmjLHweHo
0voRLm80W6Th5/SwteSqYVopq0AKfd6j+VFJTVG9D2qZKCVUQ/shEDYdpv/3SeKZ
38qBCfCQR1Fm86xOUsEcisHDvGNS5fetZoUcAYqH2DTHOlOSz/gwyKU036f2FZDp
80A7EvEVSqISPYyRgEhtvpzvHr1r5N637YdYmCW0RsgbFR5xPXK7Sbc+M8nS9QBE
v+ErKYBzUuh+mKX1wYU3ZFVNNDPp86FaluPTESEKFK5AzAZAtP5FGqcujtfEosYT
3ra0tMOVp6IyiWED7BpEWa0Wvh5mU3U0ap/SUcbkyzqCVrzSg2HUlX/LK1ULEt/c
qvKTCnFghMSJG0HZjHvWItq0Uha2KaX/Pc6cSczfoyxODwB5itUEh17EgcytZqbX
ehyrsuRAHh0ghnfliGyMifeNZn0I5A9Gr63MerGUUmdKnvT2MgYM9PTlBLg/iNUj
qS8yRCK+2ZN0fFG2KABQloa9dtvcnS2Es6zh47qRHCxVJTaFbwOxpoVzSpVAN3hQ
NVkCBr6JcUgXz26axie1Ei/Fqjt6aIHOTepNLewCRv2uidfxcTRuHf2FJibsy8hk
rhM+JT14DdB9cs2b1tvxnYGasWIp1z/hf9tJEvQc+PrkMVNZmXvZ77tVJ53wrSqV
fKTL0xWpmvLgyxLms19A3tnkoyOaVmyzMktHpI7HiGMscG5lZJiswdoVSxCl9kFT
WA7GNBErtt3wC2t91Q1lSQ87GFoiv19SEN5FHEMdrYLr70j9p73jvFOh8ur3mGS7
OMUpCWwiTbhDuLGPvKSe54QEpLvhdXpAn612HQ/lTH2K1HIWe7mFuzE+npsLj1fJ
yWFHKAZNe2T183w0WnzQ4TUIb3yMMT0G0y6eD3Md0S2PKplgrX1l2uBSffyn9da5
hlXI2OQRCJ3qqEE8BT2stLVqkswe4W9duj7gAKfLSq4eCnY2N4NZwXdSJu6CrCJc
AsWUdfjJ/ex5/O3milQaKU92ck8IDK7UyofozVW1ESwO1NY+HUnImhqD4/0+lyZe
3gDgYHQB58sAW46hf5SY2sLAyIozGbgg8QfDvL9+/mDBbZ+9fTlc/rhg5G+Wqg/D
W1dXapHpVx6DhJv3hY+NmSdRAcmXwtak0KSR9pCcKWfG9nVKogG7OJH7TLpxB0OD
aN+TMHOpTJfgsgAwinLwTGgwHSbrpA0yQ0o84qDjcsJxBMKAml81ZQqQTR66tfwW
lgiPWUGC19bG5XMZc/ZLde65wgyMLbrD0N/KbXR1Y163pM+eE66oonJ8DSdlaIWo
lLj9muLPQWPuE9rjWaFVnlyI8nC8BbjoG/VJHzXH5bXHV3PZNqQFsoyCOausY5HN
+yG1WFUsTfKwIuODPhShluElsth0ZUjlqWaLVrafkOUPZyjXjmY8Sp/Bw7YGGMzI
1sXuBurjpMWKcIZv8Wd2l5WvNNE4oj6xWzIrKLqBBdLr9CW+JSDTMSYL55QCJbu+
kSndhTvwzNkKmOivB1tf0GMFdeFadgrejKNmDeQmVclhyN9OFnbcwbrKR2qFT7HN
pHdLN/74JW47/bAFMUz0WxJUADaCa5ovcr0GCqWfqoq5CX6cIs64ZVarI2RYVS4l
qfvYusBCHU8g0wJn1lJRKFvpVRuXZKcbr9vb9BdEvhaHeI6aVSzZ6XkvlJ1p6ytz
8DEAHuEM/L0ix+KmjxXC+9tTJ5a7FLoXh+q0rtcvxiKbSwfgY/tUMqBsguhgWNR7
OXOEPc4g9jLYeHhWd/ExRAVc+lHp1lUKdoH0c87T+PND9NIlmJHEL+DduilM1GKW
PCSFL6+QouSBnHHmiP73xo7ftMe+FyvCFdTDkNvjyRpTH0hD3YC5S/wGWbwutdo1
PFfHgS6P61Md65+v0SYche6UNmGVxiNwTAgYccIiEmx239uAv2tiHFjeej7aSO3B
R9pjd0nFFRn05rPdieEPndC3n9ONnMRqOlU9NoprDGLYoVj/86pY2yh857Sb9RiP
VfqeiFcwAvNZGXI8P0ZNA5uWR3TTkxRrOPWGRsGOy5zIoOsaEJLf2chyt1ps3a2t
+5jaMwC9Ke0g2AUkdjj6Eez7ElUwLyYfuFmSHVqSL6qufj7ryI2Thbu6pBDCGVwB
KntyB7UQJH1Ga4+GnWYTE5AbYpFLHTWRF3o0ufGnamjxeA+CwGbsz/9GhvRPjRMz
bb7+i3bcue0AXPX+dQ8vH43digJoMyoZEVQNwyezWvqhGmdOGgSxrmJuiASmA48T
6ksmxWEtWPa8fvjP7hJG2l26MfmpJCav3UWrRRx/93ivqXlodqChEw5LQ69p8Qt8
ufkT8ATqSWi89gPQtcUXx9fr+awcfb+SUU7VPA7as2clZqAQJOgw3ikNZbdKQDQC
78MVXuobs0PcAphfaxa77x2YhjtlYJSIlIeeOKe0u0I6eED6rNH3pFki0xmsKDdA
Qp2Mhek/MtZieKiVl/0QFpi8AKnJTcT6gSnZ5j2xWqy6J7SEYu9NTcwkYdOfw54g
SsNkWfwCu/R/JwPX7+y6ZQEEDdTImiXBw8RfJC0bEyBw6JEvKUsEsINoRmZubsNr
a/D4DK6TOhQZKpppsB7QnjiY+CYdV1chP0IUcCPfj9Hr8jfGO9fdp/Tbzuwka9p+
a3FrvjF1aeQwRfn4Ql4D4uGGuUexOSucKS9ArTAlOrt+Xnwz45BADMocMrJdHOZz
8lXq0E495CJbQbfmr5ILODLUzS4hviC+EubcPJB5WiiraVv7Q5l2kydvmjVNqJsT
JGDcLvzhGoQQEeK1qnvw3EG90Df/1Nq4szS9LUFYPL/619a6H4fVzDLRO5mLDmNe
lk28i53tGtCJQ4L3QS6PebmRPlEKx3RNJm7waqOtE6qplzXER/Lk47yqszERJQXS
aXNOuQUeu7FatrsIQoEwudrWpRr6eCXRRRo7YfgoqE/1Y8Qqh6WzNd1RrpguEf+E
gI72ddu0X6zCpXljyy4t4hZ+yFXwhFMbaqpYNwVNJ2aEx5yK1uIo4NueORJycfpO
s85EROPMvxjzDquEYgMj2fi0uVWMT6aVRyL7lXKkXyO6delX1ldhUC7s+goJLCqv
w7EDSAxl2pCNmxBtaLBrVQHndVpzXZX1YPC3UkAkTMeBNx0uFowQH94RzldYSByf
lam+2w2OdHqF+TLWmUAPyby8BwR0LZ4m7VsPAOCHen3ErbljJyNBp1IeG7KV3o10
YTXr89I8KDdjzBapEISHHRwhr5YGQE7qn7qJzUpHbVhWr6T7PCjTjOrcJo8MYUyD
SNVvuPfHvvNKUSDELQ17dYUnnJadLq7uRwGE8gYzPCSuBt3+3wxIAFx1uaz1m9NC
pKQK4rYywJRyPcjV6dYCSXihM0tY1gmZ3xDCdtbuOHsD760hE15em/ISmPucOlc+
dxoi9ztZ8lP23AnASGTmISCCVXHSY5WgyVLwrieUMGz/1n775OpTuxnpZy0OjyIh
Yb2l90w/ockvR6iUlq3v1uhKw2Wjjztfj8qMe2tAC84ie9XntEfr4jemMzyKJhpt
HDrnz3ESIn9ZF7Ivbg5f0rRmQrFwrdJVRKOJjuvgq2FA1zr/MUrlQ4B1AhJ46VBP
Duk0vlQRl1XtfOnt3vBidNuLBeZIKWST8/FemreK98YlbX5FZKbSNBwKB1cDXvKf
mCQWaX2GfSWiDbX1/SnNWx6FqDgKaZ38VrBXJxwY5ia5y2IoxjD1A8jF/RTOKcAw
0PUbmWoFLwcr83/PDEDda9WNr9UcyhI4u1rXYBsPSPsK8enJcLS40vz9hE7HeMdz
hBW0yglNyZTkJ6QBi14W8qypZPpdjoyJYVQWjan4LvUMo/XWPa3OtZWwGI6mQKvY
3cLeTy15bYOXETGZiSk4zLjm36uS1FRCSt9A+IX+xREEEX5RMdRX0m1UaVEzs8ki
TVOwnQ1Fs0uH0kO0AdbXx5imxX/MRkSLrCDMLQhZrLpNrMQbs7u6N1qvQx2TB6P8
Dsxe3/MQIqFVibN3tmgFItlhD1/yfXGJ2wxG2eeV4/NcHDn1uMu5DoQEHmgGcjlh
hiPNltnvN7/LWJWk8MmZti2eBuKiRiQ2muLQP8SkU6qli8kYfr24STbSsxsvNgB6
Bg1umivouC9E+qq6J3n4pUD1m+7EZ0XMNKXqoa6OHFBEo6cVuagEMkojEguX9DNQ
FKi9BZ/Id/bawuuImT/Lj/yGXX8fUe/EkXrSjzC2rHKRRuYonEtXIs18nPiFhfjR
OxuM8Z8G3cUCDvfbAGqYdWBpdgctjUj++EduSh0pPjv3Q7ZCXHOfiwIeglapA8kH
sB4wc1eO9PQHhVBy0kc9sYcsbw+PI0Xcy2rY4gUmU20TDEaqFBpNLp9jiXqbJyGX
xcDL9KKiUnnvB3hpmEMDqdKX6reWdVp1SC/HClOejc8b1qhdecF0rQNYCvLlzs40
pZTPsM40enAcUz3GVIaE26qeF1C2lBhoJ9yH2vITbJ/+CCrDydjSk+Loy9VL4Jfj
JLOJZUfYlXln8mIdOnkGHOIjG99Ca1MyMOYPIR4X6DGvzaFgWfyCtJGqhEhmnteE
5JtgTjdj1YXXMn2/s3ibr9Nk4N6aPq79UIPWYKjJdNmRw3j7fIUw4UUxySij7xg9
t0YpqZO/L9DpJdoC8dNbN8r/0DcjYIKUGb6d+jw1S//5sVl03hhNFmRCecKgpjn9
9AWETf7RSWT+70DjZ7R36mmYAUkRenBiJ0DRq64b1whwbb/vyGXA26VsdW22Q56E
4kHPrUgSKGL/DzF8JFKYJuh6WckaI9N7tQcEhlY7Zxji9OpvxnB69VILcEXvwg3c
7SxZEthMEur73t8Glm5cs5CitW1FYeLxpxFUUl2n220boquiR0QknKf22j0fvCeQ
PSt4SEqDLPpvbhM8GfrSppYcsc1mgKeq0ICcb9KHqE+os3HCbPQgq4xK4qgk/F1M
TGR5htXSC+gADSfm+FPsByL9wjc3YVVPVwDTSWhjE5aLVO/Sp8aKgivuuLMXjUK6
t9JXAzisDDHVYWN57tyLWeM23xEywJg4hDQXbQA2qNXEUbqt5m9miSXc4r91yJEH
6kZSFbKK5F5qtzG6lYxtLaxSb2ZvWZsRKr7usv95cO1CWqmtJc57wt1HVb/7Qdwp
GbEAT+YNHQ0CRIy0D9XZ2Q9wkP8X1izeGxZBUgoVaf8HPf+KA71/C5NgKB5E8wFF
xFjW8fm/gDyrwBMMeNrmg0ZVeQqUkw02CSqrYukOFNJmzwLM9M4TMusR+yuGIK9Z
F+iDih65Ubid/2Jc9vfUJhY7dvWMlzpGdL07iMYOwDY4oqWnolaVeHCSQVYtX4xt
VewgAUE/Z3kzePoLLXHZOCSScOO6zZQ75e8T934To56rIvdzCRpvn+JE+kUkTZE9
VmjITey+7p2lD35CFhiHJePxBYmKMQI/cCmQWyJSQ+/tG+QSLeznTYltv35X6cVi
nk66LlcFS36uRcRCfcm5vTNbc6OAI/Q6tIGARSbPP0aZnUSwRv1NiZ+qq9UyS0NB
yS3eraYgcaolqYtUnKan42jZcmBa7BdKncusnMObx0PsfjPpGz1Y+7yTZVI9qSme
z1werrc3CUV0mu4CTVxuYoiKfHmYYTGAaBqnjr3LraK7UMsZkQJop+wpI+p1Lspj
EY9x6jOgsAAo4MAwwoesLpAlslcpMsxYfc1t3LYaA9D6X1an8/AE6u++9tIWPU6W
I3r+FFClrSpxwVehscuuJyPtLe0eI5kxR2gEkr1+kZxP8pipPpgJwnZOmHq8+3LH
OST0YaD7/pPemlXqQ6FurWvql/jCGiQAmBL5sEwqrLIC4vGNFWfo5OOt3tHwz87s
JO3xAbbV/2AtQCJA7byY3F5ZTY5DbA92hkNNWIB8sfZ6zbKLPZ8icvgeZtq26nVG
Uc5Fl5AXvYt1vSgFNWNpOXvbIGLqFqWG9yXQT0s+frZwnobhCRxe33UTE+hRLZi2
1MNNM9jIjM9wgkpJZ3kuJdH7ovddlMTsOyTbbsDqe8EVqbXk1qZQnQplqEKh12n7
etfSAywEKnT7Szu6bMqd8e1AlMg5XJvZUd0UmURx40BQpNGpNRmSt5SxqslEfAm3
9nRSCHszBhPbSh6G0Z48cnO7jIpTGnXtmV91w6MTEzM7H08XVHd3uOKtiEXXyL/J
7QarplzR3m+hmCivyQs1IeWg8cAPAlr9wTgjTkKzufJTPiNcE0Ym4T8rnI7LW2g7
f3rayxeEOWnRh6gmM/zKxqN39nZSznl+crN8U/DuhCLcsj2mGNxyEHGu5X8PF4jL
aXERPpKpo4Wlv8LL2OfIZHwqfB/+WukMCk+Fl9pO5u6+4/93Fb5R1+4Ljuz1lOR0
Ff9+XG0yoytTc9+i6AnKlQ==
`protect end_protected
