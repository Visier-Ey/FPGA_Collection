-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "N-2017.12-SP2-4 -- Oct 23, 2018"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
kqhi6Nft/qc/psb1OEWjEgSiLndDe1Ve6ZQROGu+Kx5SVsBzWqqicnmuqC9Yfi/x
olhBFIodKItpJuZVa4RFuS7X0sZXnSccvIwbM2Cvz58ROXRDccE3NEjQxnsa76pn
tToNlq7wft+9IpNwYOuHGWjxAN8WSUlpYMcqnZyTL2M=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 10048)
`protect data_block
zGds92QJeqbzxm+Hwt/Fcx82H553VkizfTQ/iDs9KsA1yfwrvD+2RnRr/e/hgAaS
ljmqTBMceFS215eL0Ht8+fdW+Fdib/adGgtM/6Vh/2Hft2ovgK09JV56WIYFpOuV
maYkSkdbfEBwYDi6RcDk5uW5Kh4mBu+wb3HSpm1ZIJGW2DXpTrvIAcTjUiB+U4Yw
uxxrwzN6zuoH7oZmAq8PtAu2NGkr6re+UpBdLf0D0mhLkxuvZ81FtHdz7KkltU1B
3+AkH8okV3iNVv7qtcFbx86nq74av7XDTEkvY8rTPO17+Q1bdHh6f+kPGkoIcoDG
TszQ2ST65c3KEvaw4AzhIw/pAeFJzV2xDhNPtmL28Kg5/6uDZrbhJzI8T185EJGq
zve9i2+vYb92wxVUI39iNmjIudBNFJFD2o5sx82KXACYl4QpmwOF/Cx/mHx5oQuM
XwS0SP/7EgE6gLaapUueMuwlJr5HpZUIZxh72IBTGuEtALbXHQjxWQvrZxqWrV7/
mIov6GTXBH4B1b8iSbCyHY4By7sYIei0AXmcxBaVn+byOgAlqYyxPcWtTPVEsEnn
V796CbLyq6yrytfOAMsV9gulDX7k5xpLzz2nSKHiy7BOVFqZGnl3KUXPqZzPqn0b
X2q7DGckgWaHAk1nKNl+16YizKwOcmSeUOKAHLSkzM9BRrZ3t60uo5ofJStFzKXa
v6gDVqlOovNTsk49NspDGCgbwL/lBM66MYEMW0FxFtPQY8sHLBZgi8yrn7m4zgYr
/Pd/be2NaX6iW5sEaDg8mmFlD3Ysl5tMZOLzYQZu5rJElRgkKd5CPazMLCWoYaB/
3McFruHyuwLYaoeLMCeyz5tbAF7SrrMlXz6Jb+0Ty1y9SEn6d4J0jp33cmgadT8J
WpxMBW1iy1zOUR5QyNJxp/nSWir7j4WPS0X4r71teczOYZ6fvIVKoiUs8AjazOq+
TaENR456JyxXHz9sMx8uRyrDk9L0ASYsK47WDRjzZzBIGje66jdR9oEsAMUY579v
k31MVQ9dH1dGxdTWLAZwSKO0pATv68ZQCuHVEW13DIYpS/t526clhRrsAUHtF35m
l85LeEEcBIb64UhDhZ2gJz6JTZ7vbVrIq25hhy+bPWsHONemmkUlOy8ielWNIl5O
TCYX6m0sm0drV0QkUwVNlwsuMzB/7UUM3kJfvAwO3L5VU5AW/E2dodM3AO/hZ81G
jbuvcFMvxIelUMvlGsSMYLKbyOZ0ushN8jGhLi/BSsmqYU2s25+hqkXmsr/EJkRy
9kSYnPJK6Y7VYr+UJqpehisCx92DyOaU+JfT5xM11jSPhQyCXDaGMEAxaxzyPY0M
DLfmIE2qXfXiJLXGu9rpAnAWHmynDQlvRvV0HaxxPwU6ywmS8OhBuPINowpMJmN4
1AgYoxO61Yd84eJmatqQKs//eRoNHIf9jW3znk0sfE4RHJLqJVdHKPcr9k0ybsA3
B5h2+yI79Azjqbm027IMsFy33yPYE+aXujNUMwMlQFtBgfHrT0Fl5MAGHmtx69Wi
qjr1Y+ZaPZpIEDz0exccbacQ/cIcSGiKUlygjWxDqP6RCfnPaG+SYPvvsv9VMs2J
k2BfCzNbNMzpAjMc85VzjdP8FS28CU+6wJQBAE0ybvM/P1FIXJkjSZN0vnShdQTT
sybQewL+E7rs00+PCvGLjEG+I0yVCiFbFCUdVeiGnI7yRPJfI5KPcsjPIqKICKrm
u+HxfuBigrUa4VyDKsu38VulE0leAV0bNkBOd4iSZV5ZfIvZR/rQTbPzayys2M9c
if9XdVhYBQhtqy9dgyzH8c6tHiy0N40uDwpdPAU6AgzH8z+XhGsNN1rv+zhlVl2b
zedy0KQtCvEZcW3pmj46YRlowW/G0mrX5bOk2aIKwDMbDoY+hDIz1SUTooqeKBYT
ie7io/vAE8pyuSQnFy1nXsDiaPPq3dYsSy/+76Wx0DR9EI9A201bwkoWMBqmSGua
4v5MFNC/c8wTKEdT7RItfCFaeDOz9hpnHrT62aImqQu0R/pKoIsm6HOMbq3Ou/cj
wAadv39zoJYgFqnAs8rAdnG3Pqk9VdsoIPJZNy1zRMamiq4uWEE0BDB5FoxhX6q4
+ilIrMS+aLqlpVqJ9R7PqMIZAzOwzU0Yfq/ojW2NlYvKIyt1O8gy0hhvY1fDRnd1
lHfpDyHUg9Mxf9zDTJ7wSFKIieBqpI+mK13fnvw5EmXa+gc7fYiYEEU+D7QxMvB+
6cr5Cpue+iDbKv6zHuhjcm9Qye7Zgr7hBDX5cRl/9j8DLjN1HsABaVd3TISjXJWw
pMLxvvpJMX0ZYdHyA6YDiNFUqJ/SFq89BvG4lknu8JCJA3zHtDS7SV1u5/R5+3qc
5ayDbfcEkEXFMiCa2mrKfRXlUlSPIjxcCZiEevKNQbNLAB6QMBL0A7spfY5HdT1A
4Imlj7+C/E3sX/5MnNcCIhYBVe+zz7hKpxeWkxGq5B4j7nrLf+IliMFBToKfqmAX
ahSj6hOJpcZv4N0NBsWRMopnJW90VLQT0TaUwzhWOBmzT2XRqD2++xvf64zgGZ6X
RGw62Prw0H5z1uxpLH5XZWY/NQ8RevqOtuccIVaYVVJJWIvxxu7gfkSJYI4ZshRY
czMRH8Ioot99plKkxjPRvu7Zs5FluzD94xG7mVwRJ3bRK50dYgI1LyIG1jbjpCdC
K1uiE1ABVSy/NZf7EuRK6vF+ZDfb4OKGDEXS8NUMqg5x5/a87OEiTcj72tkHPmBy
B3PYWUHhP9KyRiTogqZOmyru+RDL+6QfW/26XNnf/Sy/Q5dXKC1yU1Sw13zVsSUs
EOOSD92Jp158A8Z/jICnuPv8FD1MsTRg2GX0PtBm6+6uI32yIj7esrGepYFE8+Mc
F2imX05KxpuoGeiBsCnob/gTHnNpeRmS9ffAhPkBIUNmZONoQTgBdlM3PX90YaZj
blS86TJD3qwxN+SxjZpS+GPlA8FPgla09GhpziUcOG2oL+I5TSEqnbat0KQKVM3B
0f7raYYxDfmYSUiIpe9OIdih6vcwODDRMNH5joBIxp4Y3HQ0cD57r7adJnOjcXU2
+JKY7SEFpg0Zp5jLWxKR4M+hTpEY7lrRnOay2nGgX38Y2PorQmdwgLg0xgEIu3Zt
yqSFXNxeqTuW+/fRPJX7P8qhkcZUka8MYBIJMqvebKQl6wgxCZCY5qSNX6dlM8c4
xFSPJjfeZJ65YMhoxUIwFp5wqP8av/cbH6dPUB5jk5se5GY5UL9BrguSvtklVgpP
2jnPhAReuXbNHHUWw7RwCkJJSR8OjwkVOM/TO9H8ZaoSjE24RIL4DH0aJIa/cvFH
aXFpaxaUfQWWk7X+E4zx+LljyaqMIHzK2EtgvdU8+HtyK7Ddw6+9WqOr8a8bZGnt
ClpVQwjguRFz84WqWKB3WMaA8gwRzSE22ePcMRFd+9PaT/lsC5bvjD1E39544oFl
t0V60iMK+WC6dMOWd64/Uyo3G8EsghuMoG4NTr8k4A0WveFH8FdxbnI3Zk8/yB+X
Ew8LwtPdLEbS4tMVXHQ5UyzDWsNUP6sHZNFhQkhtBZTSI3WW9z84VIZ7DhXry8kk
JwQVGpOv7eC2QaBBk+EUOZe/hd+pltdEj2IyWxFglm9ilmnPV1Afkyw6Oo5+LM61
FrdeJ0cKPi3BsaW0Lwtja3hEvEPZ3zyPGm/KKpSVxLaXecYEvvLwZngurl6/AFVd
b6/vTPy/KvgWYyBkr0sNOTF27/h/cZOcpwA8wA9EmvswTK0SUkhTkf2f3wsWMARL
6qVB94/NYOJeaAAOOJpwcSgW6Q6Lpj82aMwaM/vHwURQOmveLEsKotjUdtnQQfvS
6LTz7yk3uO0BxvZibW2i3VjIhLI0lvHpDXpLtLyJPysBxM+NG/oLwanIF1BmIG44
Qv+T7h9aOqk4HuGtC/L5joq51+mIVk4L6blA5Ftxfy+pNq9R9VkzIl+xwGe68NJM
tovXMZ1qzFV7CM3gZ3LNvHYHBHA+5kq2t2cOoqibCpSDWNzGbkV2I5/tJvOzaIu5
hupD7H7kjWCX6JJv5aJSVvgPTAzxCd3Az8ES+1Nbkyct+YWgTFniqj3etBdR5h9Z
GXc7M2lCWjQS48u1IItZTPubY2VHBosm1fsiW0w1WnuOXHXVqrsSDBWacG3JtxQw
myFnuLCFtSCgphdbhNfgpknt1zhWPFbiVol+NevyV2Lwrc6ZIQax5TFNeYtf/HIK
FsOhwhHNPodNTGD39huyX/DirkBYE3ju/YqvT7V+skO88viHs8suGN9owf7ikR9c
ToPjCMCRRjdEOHzTTbOJnmku2802sUo2HLhJ59PHM7Xt6P5GrlwC/CNiBlPcRuik
szufSFKNOa2jG6VEbVBd+4TGXN8eNhd83oNrY8SlODwqyf6zX2C3k8q67awaNLlJ
nwFMQxLIEvT8PlrpoaRdQGOys++JKcJhzHzZVf16UTZUxlnGOuwKjH5h5OPJ/yMM
qpnb737PmN81ntdk285CNLHx6FoDttJkx8ZXNbKgqvmGghaJE9gtPrY5uwdKYvzg
JGVLyqAmHhH3wj4cVos3GPlXNUl7kUaNl3ZSOS1HhsEbI69X77rFDXVFQRTKvX4l
ufBYXjAhEY5vCSM5CR2vp7N3JBT1ENbR9aR/YF5fdrjok9hNdH8JSStGMShd0v+T
SR+liCDXbAVFU+DP1c0npGVwgW8KKd5OG+32AmNlq/RdAN5zVjqg2ILlekButWQm
FyE9JHtVrMy/q/lnXWgnH1ps+cnQphWd2T8g9FjIjLxO+1YZ0116Csa3kloF1ipO
xpoLVxUhcCGnMso0B4WDjWWN4EzcFSAwUAuDstWfoVjHIlJDPiI4cYtVVIpbMlag
BO8nU0THVWIEXwcHioi+RuZ+DgI9MSf4V/kQT0aQ3b90uoWdU/Y24FGpPMTWniYG
shpKX9/Vz4Jt+BjsJU9OIYjiEvS27nr/Z0+bmldKOoz1MqjxQvFzGLl4LdbrDI/1
Y0AUo8Hdg79TDE0eNM/ycPGD/F3NjV+CyxNpJau785cuV4/jSCD/72u+T3uL5o27
vxIhlD/Y5r0wywn0zv+cywjqdP0dR/Y5q83YiOLkiI6t4RE6icmKleCFpuAWLA62
tHAApIH6n4xzPwMcuL9bZhJvOA2OnrNgrBEVbBnsOpr2vRAkzQFCERXXvhdawmKS
+Hg3rsDWIfE/BotxlSCYLVpZxLthHIA25ZegkR1S8tZt28Y8EKzuusNqX87yIoke
mMUuL42Um+ldy4gyB0LYBwuwWVXMsC246hUEtD11AKO2zC7Ttv9L1WyXCwZ4gGvC
AymUiLvwUmvAWhLewJTJSo97nGAcHjzi9dpGynIGRSoIdba0wc+kkrKlqc7mYC5w
rgn8X8gjTt4ktW5DFx9XAniZ8h+5+dqc9y7G+mZojJ2R2PQH3E4DoC9lbYVDF7Cp
WCRoNdDoE4S1fXWSCgrkmKsJ4/bxbVhdVdY7ZHlre+tZbYN2xJGPsA58m5poUodD
QNwd6rsq6V6Qe50TqI9u3GLOhxfcgg1Zu3H+4XcvsoZr2Rr5tp0X29b3JJAbIMC6
b2PoIgzFbnON2pSxz1dOIufYGxynAti0TqRxEgZ/8fUCBVH2QgX822tgB05TXzxo
g6AzVBPFzntFKCqJyM1JFjVmVIigIJllakCNhescH9Z0K3qt/tHuXe9lnA05NBOa
04xvsYlxMo0mi+rqx1/7XJ/suU7G9/tk3FIsSJQipKEh5b1QgmKiTDQWjjqyRHpR
29asm+6zaK/P38NCub8XY1Eu3w8b0ZBta8hduHOulE3kwqZHMUtkXRd5aLF1Sb4C
O48vgvzXp689/Fs87Of3GoYRwrHbJDePuAi63FSCMhjGgEOxDWmTo9Y9m1wLqSX/
1rETzSUMKH6KZnHlAWV9LMrqLN8eZvjVf7LkynkL8pisZs0XqtBc97meWOcKMI2j
gUulSKMUuSgkRKjmEkcl9UkHEUjNP9R8VKqLxDVLZLLwQIBEVV5pWioS8M+iNW3K
0XBEWtR8YAz9DR3Ex3S1HirjZ8tCcND/OkB+dIHV3/qrXBOyV3lQGnt0PJ62RIeM
w+8J4gwHSdKirT6esOLm0bOGBtMd/X07xVSY9CljAaIuyT4WxVbSrKhvboMQHn2L
ixTsuJVKeZ77ek8OdtUgffGj2vMtggLBFurT6gYqFiVd44aAoSnBOcZFdRQLxdNt
P84X6LChTg2dOzEZC97bZYJkfCEWvvw+tOeJemTgblc11pXOR2UUNif/oglG/YvU
VcZ0qZ3VQF7GzOafjlTrQZhVqTE+9Siy00thyrtmU8BuYC36j1MVJre3essgre34
4vHkCzk7cS6ZKXTZetfoUwXUOohch9k5/7uF3FFowZcBnwV1CwLwL70XaToQzjE/
8n58sW2sb6VLkBtdLCV2f6zMrmjv4eID8xWO//rfIrN/aagALgy950QER+szbJRj
EwI2zgsgM1aDYNY+pD0ZAgpzTP/NmUNHfyEAibIiy5AQI2bbKiDhKDfeS1RWqH00
IPL7plFNuvTbkFJMe+Q4lMmbPw/NbD/RNct2WdoFqcMG+qA6s8rIWMcQfypbJOFD
N904ypIZrtSyTLEmvi4Q/jTnb9PztIAnB3daaAIb3ptVt/4iAgwvzz4Nr/qsoBbc
UbGgQGAKLIi+MI/xiBymH4QF6zowIqJiDuQ/3u8V2MRGHZRyvol3EH0lEGCA77Cm
jivr/W/KUc6YlCkAQxqPxm99uTP3xPPLsV3UGadNdZJnSlhlLR28x0BdG6eNzlyd
SdnOv1TJnz1G7847RWTmCCYxGiMXdBbR769g/8M48eGgDr1CYa362GtABAxUuA3k
pe7sHS6hXVzprjWCH19brTqDhiv9oyQQ3iLlQNgI5y/leZaIsycr9e7Fmy23O+Jv
hPoj7RDYG5rthOSAqvhDwCoutRnPLUDf06U4oafbaIN0j7R5vuCZ4JFHz1pGgoV5
HC5gln4pUkrdU5fUjusmUgnknfXbJVc7OfhscAuYR2o1w0Akq3YOzbbhVxaF9u9Q
02mMGAOPM7uvLr44DEkbGBd/k+oMGHrOwuyE6Clm4+zSAJxQ4vgNUN31qkxVEDlo
t1I4DqJ9S1KT3FlHl+w+n3VXvPOLFXqfk7vEk0CwORyTzGs+vJsg9X8/bBPpTCj9
nJiMO6nHjdsG9JZyDaXdNgUSFq1+CjxYrsnfasIPf3IHxPfVMCBlLzUy57fe4qbY
xXVaOGhKKRfTlCwMF5gKLLMFuvfcfep24L0hgAsUCY7AxfwradMtVM1oKnus4G+D
oDKXfwLWvl5nkYbTnnetMHyI9FXZcOcRts/14cJrPutzmOoT5xm4U/pPMH244uRv
XcBFnmgEgWQCVf1FVI2ibMzYIe7zZOa8MZRq6iIo1dQqwbithhvHtFiybS0pyJkx
5Mpe2ZTTLXOaSGu6nkJzrmqApn19uLg/QwDG19SdPsvN1yOZFt9ygtKntKObjcG9
qo92n+LMREpgrhkB8huF7TweDH463HoUYy8i1kCaqY3eIeUF46uMhdjC2KVT8EJH
+z3iqw5RTtqp6F2xmXuB1MxLnc1Padm57Wms8mw3TCCuOUXlgpKJHNYU8gcUJ1m1
zT3g5YkkdHhQD9fIe0+J+vdaU244QIRs2MQ9eyIqbfCe5znK7UasjNDGh9vJ+pPf
qQ9VauPfJhZ2bzsuF8fm5D4wVwAcSSpVl5h/q112mJH/sjJnwMBRBJ3lK0RcD9HR
qg8hOaXZigHbrTUjKfR8FFOxeEA5SMJ7pe5hmtLxH0Y9dJTtKt6w85pS5P+W4Y4/
fYHSwIZyY1Rza//6/6D6ZVX3lDxxMma0Fum2V7oGI/vofgWmTzZByIvQJaqGsfEE
AMyvPbxqNJAQMiJVkeyCu3rNcQ5JWNrwR5PSpwovzzDINj4QKtJIydWaZolbSHpp
IHRnQFKTjQjynFdONZ+0i0QjsVBMG7I7fD4lI7dXcyBQrj3qnvcthdbYD4rxlSvu
bMtFm4005Lw5LJMTeUtp4tiCG6tJ/kVex7bH9hpWx+Er8WlcNrWrTSZMsFt6dV5o
uxZtlfVVta1kCoW2A1V0iTsmcUmFURenZ2UPvgkB3J1qJhrN7McE2uO3K2A1WpRO
aWh4hj31YGwo4YyaPyx4oRPE+te8i8lAAYlCZl/ht+fu0ZOEhgxO+l4QUOfNRdgv
CJ0X4nxBMrZyKzrMzR7n2UtE+HggAm3PEr6GntypkyI8JewedoxAJOrxjCG25mQz
PCtZGjaFMVn+CteNE2mj23yc+OYVXmsuANq+t7uB+loQZACnpK+BLAn3C1pzUxGf
4poDYCm8zwni7M7VDKjholcR1bjj7trTOnEzJ0CXPOlOPoqkmQvJ4vZPVBSRSPdy
TNbbwN/SoXSpOYKonnVk2GYMIkS2/60+7s2iHpGooLW1hAPo9YbuFiuoO80KXHJz
U9FYNYyJjdsY4KVwLNuDSVIPSD6zdt9jme6foHz5NwOW72wl20FUZ89Zw6wUVQsE
o7EyG3u3d9P1hogpF9fMOGgrB9KKVseEDnIo2KXeXs+6LqlM6QOe+rXuAcTTlg3O
NtvwBx7hZSTyVfOYz6FjeLFj4KXUauTnYorD7uNfeBYAOFRub4NMUjrixBtekdp1
gp60eFa7MbxSXuH836m7nxcOiyav51TF/Zg30ywmZuftde74jdM5zaCnBrmY+TPe
rKib1/cwb9mzsLGnL+/uEYX4Dh3pzPbLrKvkNWLnokgU8Zflb5gcyROlRYuCrIW8
EEBsImIJrb4dEZgA1amZXCjLdAJeBhuyORMPTCAmqj7HSkk1MIHdX5LDzcWCVgL9
n2NoilGr51qoD+Zh6V6RuphXMduepn/lwIiX007YzdwI53jEYDExGwdYXzvUEynt
jlsrrjKwAsnE+RMQ6vlfwVswRPV1tFPWzrSNcXBKT5t+wW/Uam13DW8Jl4r4ibjh
D9854EjgqZWUKSzdM4ktsaUnYqgqep47+x+r0G1Oy/rJ5iVixxWaJYny5Qk9DBUv
v2FirUvwqXc0osQodrtBR8ujWHJOGZFoD6medvXEUBOk/9++wH7j9Bh6E1yXZ0F0
8MODOfFamC4PO62urSZ+pYw34mX/fgUf2a1vkaoARgn8CvYPVxM5J/LFHJOeML1H
Wjcp6FIzsSqe6/TcWv5fNCvwnJOW9shL4MXVoPV6cfh9aQlhZmBUmh1CxpWZoDN9
3bKXdpaCafiZBw5+Mh9fc9J3eI2DdEgmWD5MEdTS8QfmcIW7Kw/+RjS9drqFHeQx
CySHdp6S2JLlW9P7QGSsEwGYEo+jIBpyBi+vAgMkPnSRc97VlDADc7MKm1BUhMKb
0OOOxxo6U/q1Qzr3uDP6qw+iT6/p3VDUUDgsyjFFbc0Y2YKzx94AtTcUFCLiC2+F
BiV0Inh0y/j7ADHeEzC/q9YY6lVktI/zdozShIeUvs8e0LXJzEwHVBwCxx2zLN+Y
X+RVo2sf/eq0wRR30abd+j86giAEOiW7vUEdKvaYXkAE2JRskHDyjHieLypxBkYQ
NIC1mfSUmL6fkUb76tEdJzDGwOAmPrT9wjtOMxEmvwMcdCv6Ij+s283GV9QdlyAN
rlEOP8HUOqxLCjJcRIwTSQt3SkwpTEFYXITCZOUGVpvJbc6PzMxCvwgtGgIaZ0O2
uoUXgeajsl976ywVhikdqyGknCF0g8Rvw2ECjybpFWPnafKKFVjM5KqYzmPoRhYY
GSfI8tYxGwZ+blDVqarJtyJ5t1I3/nyNZa2ymQZ8B7lkXIB4WIeKMdEAdnJ99vvu
7moESheYKsqKlyji4Cchuxsx7T9K25rgfke0fg+UlJka6wATkv3CEVihgrvehouL
IRpf5kvu/BOb/kpOrQx2qTzK8egpDSFpWrxip37GcW0ahVQWTxjK8Df0nQ/wMZbW
CVsD7vgj5Hvx5hsE0edTH3OJPabUHxRMH4NHclItmjYrm1LzyM0rYvaLvUpZlrOu
W0aYNy7vgn9KIwTjFkdc2Y5WwjhUojL3aX+a7i4vm1enHhH0CtxVQvf7gYmCrPUT
awHXxHhJAotOQ+nePy0uw+R1V0PUVfhItL/TrOpqUojHH7xuERPZzwWVxtntLu7r
EjQab3pBKVNvFjo+4pu+1kUi5uhJoNKiP98y4nhIT6bWl3Q06BJjalVC2Ixi2XHj
ciSqDkHl7nCQh47ZAh0CrprlJReaMpTBYn90FxdNEL1OKFXpEhBFpf2uVBmeE5tF
yDUTGJVL78kuQjC2GlsdXblXg/oLXrd2imBLAMAzoj3zMQw0IN7GmJ2hHQW+Hl9O
vPwXY0iwUe9V2XT0AZld4NmmiF+k5RlnIKrtKrn6lgcNOB4cQaSB8bYBhJkFz/3X
DxDyip7IRPyYOIigFbF5pzesmYSGZtjYAuYmGDqwwL+j9T9jihAjKqZfSSYulzxC
6fFBXzX/2mg9ya2SVAvjCsoH8PyMjehuaylAFQfBHxabKkMCY8bzgF9JC1R9KT3J
TAkwU5JwdjD9uRg9ogMx1bPLGJXeDaS4zwlun7UUDFDkICA37PvuqQ4Dyo4NxN9c
HnS4CnYAdfMW5MnAgHaVTcPR85mFaXvMVz8nLjaRYiJp40zV4zQMgDVNRBb+IcQF
EA4/9hnhxt8yNdxZyfeoibOKb9PQqWKRSZbexaHTWvkX/l18813ncd3cqtNdKrFC
ByywXZYRWwjKGYbqVZAXNXPUXHgjNbRB5N0yvLm6kRVbfdiLmHf/sEAuJvhHlUFf
BkLBtqcNRMNejlGOsf17E6r0ufH0QT+lXiZO5+gBuwlJfUUDWtxcacW0saEl+i9R
o2EKGkdnHhCjyhsVd848sEPJ/GSOuiYMRsor5ZkcKHNTi7VBmvre9poRu9Rn8Cf/
4/PC6M6m/qrXdlNBgl+UIYFO8b8hr/LytbRgDE1OcuRJ/BzD2JnBXUUfdzx2j265
KOy7TEb4S91S08zicdkFx5BAagYpwlKB1IEXLzRQMqB7zCyGGaTpa71CABcF2+uw
r65830j6jBeyXdIkNvzIPLiukifClRaEreL82EIAQcbG7H3BDSyAgeOeI+gQCK4F
wP/62fVn1F1v4fMipxAdYJ1jLGBCE6+eFg44+rVZIrHjLnwRiKtO4hpz1jnozjnn
Kz6gMuRizK5rs06RRexj26e/4JVoN/Rr4mx2dXL1eLaJ0SGoFdc0VrzymO1S0NbX
KbdCDJllrRz36rhpcM2aBEEuzUPLvoBpT3q/EkyK2x3xGgIbGXGIpM7i0Fqwgw+B
3Q7tUhI86r/vO0/LM7DhrINkoXJ18BM196+xZ68Sb873lKL2SPZMGGOBxnbABTJs
BDraNP9DPKLUOPu5zJd+dYpnBASalq+pTo5UhvHIs1QuhRzt/WSDFvijbk9iEYPZ
cu/IhgT8slsvtda21+o9Ns0rIUF7+3+N/9jmr7SUYU3/5OWI5JOF0g0JN3zvWJtE
nXyq8kxPjc60fb235oJTDA62K2GiU5bDg0c6sVq1rowaUpbau30u5XaDidCj1yeV
akJdNiMaHD5rBIViOq0OH4z3y1DcOgrv95c89H8rEzKalhhKpoLEx/zvrD4zs2cL
YAiOqdn7E/akN84jkBXCsgk9DsjKFeJbt10jPHMDyB2RBEaWyOGkiqXAtRila+5O
gEKu007n3aU7uyonc4vW0C1hLnpBaNTiqGQ1KnxsJrwMS1aVKaJLGGBviYdId+Ct
TMNlzZnHSljSeT5VxyV7CHuYBYQCVd0JdHfy6wLe2yBDpt+dA9nTYQe6xKrUTgjX
VcRP1OKNYWAC3IPnvbb8bQvqHe7BqC0xByv2HIkIFvyglW+hSfSAkVmUL1c8VZOT
lC0WV1DeO+du1cTuPw6gcajuMxWvR+Ka8c7IvCQsL7Piqh4NqkpZYfMSDEr4QBd6
j7BjwrzaJMBi22vkeAJxPLvW87aANWXrrIcTFF4hki3ra5OHnX1V9OC/OGIaFqcZ
ACFs52zs1R6W8Po/xFH4Dq1Hyy7dTRoR1m9VYzeFHUbfsVw+boaZ+oMB2k7Va9F4
L4S3/4nSVI+uD8NYfCP2NxzH2dd+02WBiVu+nC1ucw1m0nkh7DrHrlEL+NcXqfS/
ZqhLehmtn5n93ZCKV/4GaOcNQ5NTmz+KIkCBlru+0tCinrkPzEdvCzRO/2kN8d/H
f8OOZqCPJRrmmwoYQE9N3JsWt2DzB+CsExthRZ2897YtWpwKGCSTbqp65cslPhqh
IvNchfOH0TEphQ61u5WHcZSEvSmjXAHGhGxbrayk5o7gCPDCWy7RYUAtagbGsGvM
L4jfZJ1Y5wznFvNTzk0B0/1FTATebnuBClYIYssNMX1Bac3HXpiRWan5S49grId/
AEc8+dkOLdxejGpF9IbTAPiaAzaiE1CjMmFtUXkCmTJqsfqN40XYWWdZSFgwIpLs
dhbYUX4Rw46VQ5G+++rjDbmCChq/0zKcRvI/AVfUkrfrcz/gSP38m0NYCtua6S1h
SybydyG8SLJxwRRR4ACMpnWjgtQHfx9EvhKvhtCfLfOzZJgjDI9muR+VGxbdTEMp
xqBzRdu1frhMMNgx5MV4Q74ubyxvnInAxUXi69u0n908ZYpNZhWSZFlY6DNBfl0M
XDoWNLl1utXL/x6uobwba2+gkyCBTpoOdg33wdW3T/tIkfDCqXA8CMzjdyX0m3cZ
CCKlWt6MHgfDQY9+urqk8b0srr/jWxfS+eDaA/3B0gT3ZTEylTlmseDowvVUpjTD
rUauH8n9bYuo6u+dd/Sh88mmhUYAJJKmkXIDGtzOCmpX4q1dJdL0Xj8b3YuPfwy1
8vwoaI250dD5wJ2pP8Tu8t/YHYy0pxWTmzLFxP57A3SBTDMaBHYceqBxY2DlCkpU
LqbkJdjdgcKZ7hcTG2t8gZGuwEkMTsm2g1re4lrMUXPR8k94BrToRkJyzvheYJ0Q
tWdiUzN5itB3v3FiXImIqyYUWoyuwB+GzXDN2MqnMFYdppHB1PfO7X0m14Ii1Edb
yqmqXSJetyLYCmqutaeAGpEVqBZiN+783JEEpIqM/R4tC3ipwdyOx8rFQuXrMcob
9uep77JkYfrxmCha37j8Owg76tPydDNTGvjjbjTpC9C2McBKufaLMh5u3DWCinLL
JUT5k+qDseaUwbxvDSwLoFd88sxn1b0RCDXu45wK9LeAmrueyTOBT9WPqTPks07L
BujUfjDXzWNisSzQDfIi25m69Ld6za8UMWXdzGq+gmyqw2zmmNVQYnS22K5lIVV+
qHs4/CmBNkAO8hbDT8f3NrJmfw8KIODTCORvDkJQs0qyl/M9wBHp7DcUOS0FEoAZ
q6mKszCXgSYAZTn3hHhNSSBF5I//iw1lKj0Sk0G9fMQnOqzxOpxZ0/nFEdkIlDTw
oQphrACVPEvHVyVeN8098Q==
`protect end_protected
