-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "N-2017.12-SP2-4 -- Oct 23, 2018"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
GxuZCaZZl9D/Ikd6M6dd1o5NEHn7wxEkKX1I40P9GCl8gTqYHlYkJgOWlNYqxR0f
gWeAtvhuVu1Ulr1BntjYueTrvNg4sTTYh+uX//7E1IugI4EI/572wPYy4ozMtS6p
TWnthKEb6r9m9tz03a60pBWIGB9RiTDX/yBmlLCUf4k=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 18320)
`protect data_block
WpXGY1yOVEPLe4UhJxR+3E6t1EzEKxxWU4kHnhR8+5hSDsTyJhgrf6yErx2JqGsg
fwMe2RiafimiLH1yCg1eLOEYPS5liHDylpWOO4BTJcppV54neMxxujYC18XpAjLA
DwSAVszGmvWtVSUFNXkMV23s8lq590D18Y4SfgYRFXxXoB07LNlsPuIqdJuEj3vD
8kPmpvvqlxw1bnjvMCvrHLRZsJ1u+ssB5JCMviEiuXynA6hA4DfQeAOc+gBjSlrM
Iwh0gfJiYt1/toWl4lGeJnqejfmV+0gdVzXcbSkqND1x5fjE8zWVBfYhBxSitJ3Z
YluuZAACg/1Lu+s7EzOn4BcOKh37yVrEGnqgb+tFqzzQ2GjVX2mkCPezmXX+Jr6n
lboLbfZ3Os1TggFAi703KIW9shYOjz2I6x8HJomQtd0cGu8e6g2be1r53UFMp9/d
x9LbAhuYkpeLBru8S+EP9bpzf3MuHVAlM7ukc5kNVm4XdmtvKVgaq9sabBaNQuif
4b0I8jm030Owtp/QfZqR0ejqJxRpQcgTXP2lc/z6XUXf5ZFX1rDzQhCcMlqv1ZJn
g6yBcCqzQFxsCBwRAiNcGhFaDOxQ2DvoQVeeEYeIdxEiLx83dPv8yDaSlkIf88GF
K6M4bimxom83TDtAuuEOHr4N42xhET+FnxMpXqNMWavqPfL9shaFWM0LS1+auw85
AMgflb7CybA8BdMiI7vUUG0AIktM7f7+ZRYiOIMPPjalenkwxEuOmhGzPu483leW
9MFKLd0No3T93GWtTEpyO1hHyxoRkQPWzqQ/0gs1q3UPO/jnngFie77M0gir1rs1
tn2+5elTFeWhrSnlkWFqQN+2ODaKY+rwZEy3Ky13wKOw94LOLotXwLEhkEfvrioO
UBzd+ZHUcHX5alVZ4bvkk/zNZ8wrn7AtCD2/pelQj8vr6Czwk0Y8+nc4nJA3I+WP
UhYge7bzpaQl4VdTXW3TS4bwtH2m1VnNKxL4EX4mOWtgaQGmm4sHlWyfRcL810jB
F1O9EbWyKlNz2MCYuGcKXvvqAowFUCO3LjFl2EtcxltjgyzBUgdcHEVR+C1Eahbl
2XtpQf6agK0wo+actbH0mEeS3/L1OJtwyozoA9Do/WqsXiZyjORIt8TBl03KzSnd
dX/h3rChKmA9r0XJ6Kjpitynl9poE0kwkw+Zkl1I5K38CcusX77OdAXSBM29EHjF
ebgmnvRGGe/TMk7xycKNa11RDeSCJ69mCw66PQL5jTLqMW3l/Jq1TnWolbSq4Zyb
SmEVoeomp5pcpzC/tSDfUX99KP9USy/g9EP7YhyIBVbuUOw7mzbO/5RaNaoNDGTv
SqV454j9+fmY5xzmOAo8y/+jIwy/2JCVNApgULZEHwvI2v2xrgvGHcOKZBcJ3J+Y
QqQFq6hfb1t/nOYcOel+lTpV3zIjDKzi9y35awKRcQZuGnW55QxBb/PQt+VJ3k6M
U383ho7iYALuUKjnG0c6/1AUuGqhfM81z539rdwGnA0pEMU1sbvcS1BIIMnpj4zP
7GfY/4katWAozGJqy85aYvaml+vVOfskzIiEyWvFNtHawoLU4Dvg2m4dzXAvmShm
MVXCFKsZGbb5QEsFrrS1k0STix2Qvj5kb1lStY6/0KPaxT1QMy4jVyifDeF9MBvh
1dmytCC9Is85y5kqhU7SMxXo+cFFwRDrZZA6QUbCxHcWNTN2GqI8/8bWiDLFFaJd
LqcYGnW5C46+kycLfADO7uKHPYTVhnRJQlQ0lzAbskRDjMrFqjmoegcHfZ2KYxby
DxDyJbvOrnwh3q0REN2Xz6gkRYVpOaYt1zkiP7cM2kpaH8pi1fhnGzzN+2xT1oA5
+NLrQCqoyjgqTX71nTkQedurHyPe3UqKr5CNg1got3CIZ3JereazDNEdTCECFTL6
OF6N5t4Wocc4R2foElrKpjv8EAg/o0YVREm9ybUptAFbo6ISOUTySVkORjC5hOCw
1Do+zIXy1jr3JsYiMYUOC11HVfpvz97k3kwQjOgKOjdEeKOJIkvi5Ky0qvLqc+y6
I1h3qE92ag7L7tAoVpr5zgssekPfqScyPd63NNgD9WU1V5jImd4jjb+/UuVGeLeS
N0d6cKI+FrehW5lJEr8Y8QMHtHnzNYYY+yqIMwh9k8+L1sXKtn5EMDsxaGgpaw+Z
uJ2ECzKQUOiLRm0lsgb9m4nA3d1VBLLE7WxuyE7y6sMbBwALfW5r27EMiA67lPoJ
NPJQc8LzKineIXk/4szmn69XXE6UvE/oW5US3hZ1V9U0YtSbwWsgNXWLxBcYISQm
hZiac4b1QvXjX/47DBo/dMk9tlUSUq3u8dX7SCHXri7OJj6QXgCICZBZIfe2MTyt
90N85Y5ovypQyLSrI6UdaHTDznDTsRSrTD31By0bX6EQacsOXrazd1dJYwlIj7Ua
ynTQuLZmn6UIvF1QEu1i6NEcdyMr3uk1hHXTeMzCkGkknxDyZD5IVrK16XC5vtlE
Zq2aZpBHZkuBnaEnBNbCjouTbPaBVIpiYDYEjNZ8YG0LT6c4YhDENYFUcx0cXkZC
8gTMwLsuKPgnWu4sDx5zzuR9O4vn4eOUWq3B+HX3/F4nLZNZcDQy/kYXdz0UKIJN
/7rf1qIt4jdtAu5t1P3wcHa6x1NloMgDe1G3IYUW4us3ephLuYnu9RWblP/UjLaq
tJ3QyMbIYXmNk43u4qSBX2WcBhAh83jQcOPeWfgKh1w0HUwakxI4/PXp3xNieHeJ
Vvz3nxJt9+dum9gr72tTr16nWm3pDvfw/unqYpt+VLrrOun4DMJ66oyUJm8CWNz4
swAGOHg3WFNwABcB7tB2IC3pKQpMycLhAL6bC8lceo47OQT29f4ca8gNoFShW+SG
0fGvzhXjSYaCBo5Gc1aX/loNY3V01sQAJ4C/Hx8LzQnWyQH1wFFu67+VXUBMVga7
9XltBWny45ID3Q/MEOF01AnatgoRt9L03rxRw0mrD/XlTRKQmcB0RTX9/l1ioRZv
JMzSFOQyDoTuC1sS3zy4ADuFaNrjBrUvPoZUVwVohMEzr0Qi77CPonOUMOU7WIBD
8o0aUNwIdUhuy7LB+wDCAtiFIQEPYIDEt+Fb89eTHHcSaECKzXSC5Qa6ET6S8EQu
dOgQ00gV0yLYiyYIMb0XPr2gRWvUTrnZBzt6ru07dw/l4USvokVAT8xpPgzeNPWu
1YiaQRKbEzGyImWK5RM8pwWUCA+37MWxiU3CU7mbq3Y79a9P3IfZNl2rZImU9wgj
0ED8NWXWiae3m6RajdahiEJDE3ucCjZh/HmfGd/T8Ml559p8BKJg1u7xyVWJrPYL
ZNfaaBofQwHXR/XGYd46lNWoerHlnfaS3YK4L84+vWwlRbgiqUg6H459497DXLkU
kusQsuRYyyZb9Eetrnq+K0Yhs/35D9fClZx9rp2X1vnDU6LwwN+HOffbG4qUz7/e
fAzAWpOxe8hhDbX2Zr9P1isE2CDFFJth+6O/yudO7kMDsePpo6LnfUE06TVNsZVH
6G65KjZ6fEmOg81/U6G4qC9C0U7/L4r9JxIwKt9jSQ2bkmWeSwF4BGMOLooIAncv
kmGqlnIkFaX8iAlcEJQ5/VyfRBWH7tixThD92ckyaPAxlZuzBiQYRNRjIfO9D/29
mfVB5xwsubBzpLUWe5HpMMpCVZB5w1qc4eiEl1/4H309VqTaFaGn0clzcck+pY2W
p3lISwl//lMxMb4DFVuZ2csuTuYPE0shQZEyaBOZjPSv2CphQSVFG71akSRhPRN9
oTsG00L1eB8CuGwYs752EYiAIna/W8uKxwNo8kBVXxo51omrjYeypSEMgKkRYzih
fXNMooA12xnSAIzMlLIgcDj/jxRDx+xREyKSFi9n7Sj8MqxuxM0GFlfRzT3GZtLh
w6lG6c9lCpuM9r7MVhDRJH3zZ41MjkC5apa8TwTGckNzljrdK4HfpNJQr1QGIGRG
lbIlmSB8eCTg85DTmDaYLprrm7WFVb/+bTiGurwOiIfhdp4gHXDLnEhbtO4ryM6/
FpOkTH+kvU5lop2FzVNCNKUybAGv9g/t4ZvHnfq9Cv7b3CKzO9oEPILcWr9YfIN1
e3wZOb7y8M4WCycix0Qs2dxyT1tbhzKtLR2p+soCs4isPcS/Kqig+TC5XmAXDlLr
5k0m+0e0jQtKb7/riEcOeZuB2hM7ggQj2Flh/LO2ouPCcvsISptDy06nPHc3udrJ
N+5SuG8s4B6mYb+vekB8U/XnxYyu6cD0cHqjNm48C9K0JAH2MmimBQMVXOJhdL0o
Z56Cfs9zPb9eNNggawsB/Tt0fGrj/7npeRClGtgZNY01KmtwSREb6wiW0wEwtE1P
4nozod54Y5lNYzTtPI3/OI3YaLrmvAB1r7W/D2BEZPOJeWKA3sfjNhohLlGhMagn
d3LQWLZ6v8Dfm7/bK3ntvolq75OPZ3W8q36ImQQaVZgaMN0EmfWRfbSJSyqTnzIF
xZxc7uI4l0k0NTSIZoBQcwo6hLDECut0QMp8DbCTNcIn9BsGg62vp9G669cZalY5
Iqp3rN+py6b/FXpUrmOBbLyxmRDZrhKvSK33FhHIt3HqGoFjlrCL0TZaQ1c43d/U
aiado6XfTW+qi1mkDVRP8UzwbtI3AuI6eTMGhbJpDmTYVW3/8UnZPRW7iANDmyhX
HWk5HQsaDOHmXF6a54laX39wjn9WcB8oeNggWDtkFCL5tZHVkSymIp+FRlfO/0rZ
gykaYeZAqnwouVX+op2tJQx7Os/7LRXv0gHILzlvRqDHrydc1fddEKdgIRpG6vBL
o9Xi/kW5t4T8S+9AKZ8IajKoCn6qjYPuxNalXRae8/KRyXn/j4cOirOySYSBRIQq
PJk+IKfVGIYVI4BJLYFcD6lebJRB5x9CUpXt9nAJdtbcsEiezwhK9+j8R3jBHsmk
WHiRWRzPJLjgtJ74N6Kx+/v55OPvCxdmA6ek9HRjGOi6gW0GBzHKgEinkqapXncT
RLI0izp2POk+aHTt/k7PQdk37v7ddDBlh/QhZr4o2oqs1Vv1ZeJVbn8+I643Siu7
lHZKmn6sCyapyJ46N8RiG+o7dil/LSYC/WUwrjcZNKReKLkIWvOPBVzybb2abPfJ
UjBokOSd4kXaB1ggvZJCUR3nwRYDTdU57rtbGds297oPnewrKH4D+TV162LRmU0B
+mNpUl7nmWrHQniahHfcDY2qHIeBrCgbtnVyYipbIPVoqdoOifAQA/vrsa4BJOvT
LN41hiHynV/OHkb6GG2SN9+OchP64vvQhVfB2GYOK1aQvKyod6k9/H0seRy/cV2b
8OG3jFd/v5aR5yHER3EWDRfPlKmYxCj5QVdWIDTBzWJ090sFFFH0Jh/y6ZCW1m9y
+SQt0G6sQ9Uwbm+/yEnbeL5ssvyBK0+ejZ8hgXLLCT7uxMWVqZGa9ifJIVCKS0Br
kyJYjr0Q+mzelr0K+dupvp8Zjl/NarNl/GQKoikJQnNBXh+yKqHVLcegLSX1yheg
k743trX6Kl4ihAZWN16RQiNNDInaCI+IKQcuMn1jeKw/VEHnrwIGJCzn83Gv5hua
81aDWVozdMC2GJH1hb6c1NHAnZ3JFDH2a4lTWwkRiMTCPz9NO0bEcAvw8VuseO+8
XrmxcHErzFwlG8BX7yjwfZnuRvdJ79RmFhfh/VO7FDqleMprZbfKyneoXPm1Mu65
9XVrhTGWLfwGcJCqAecGWbr2SVR9/0R3d1jna8IpcjHXj/Nlz/3PhJOySgfnu2xc
FLP8zV+HJVo4t7mk1TC5gKGluWRbiUILq3SN++2oTkSHYgdpytvbHIEM3Wgft/Q+
qJ2LbqvzpiYxvBdyRw1mi0mPTJHGWHE7tle4xaz5XfeCfXxNkjqEzPcdwwUxWbd6
P5SJM2wW4TGVbRDAW5OYN3RffFjZrZPvY+tsAvpw30tQfFsWwgfyxSW2mGbJMhFV
cuMlIO/FdRcjorSLossEVX5+KRl1EaWCgvptBYfEVkM6hr4pd7whN7O2+ShH3kJJ
o+/vRyae0PjuapmdlXTDt5NZtboRywnFN97UUyQhKMsrF41fr751lQ5lKP68ejw3
/ek/8FhQnxUm/Ruft/dwlpK+AtAmNtaUcYopD3l2ts0sVzx7Ln1/usXJOu2whkC8
H1T1Q9dtCxakwvDKqh0mnOn2x3i6Q5IQ0ML8IKPjwyigD500WEx2TocRtLtlVJfW
kaJDL84J1kZIAsUslbgX11lr/nhYXwvrQhnnMjIWPIPHw/hijURMHvfaqrac5sGT
YeKpPZ78BxGd6W3FqlZIkg0m03Oe+Ha9Q+oGmsiUs5KtNUZANPMy6gXEHgI2agpk
W+RpPIUbz21WpCiFje8/U4cUa2dwOMOJTMqRy+NSLcAR1W2FqpqPXqyqMktsz2Up
NoC6BfdAMm4nz4w0G+taijmUCCFfbav6PXAlxa2VrI2UK4ovLeJwQbyhj5XLp0a3
DeJdIYbAAfl+Pzqqs18FrtZG+PmXE9BMtB0fK/ft9fCXv2z826e0O8T3Pot69hmA
zsWpGl55ORpI6CK6XtWHcch15LBO2JOFB9WdqAAa6ju+pKt036PolZe2xOhTJF58
AhT+QwqnIHo28NqYrCKCIvYm+WQbGp/amkaJT+gIwEIY/xpxW9+kXcKxA+vUMCSo
Ga7LIYpCHji1Xoy8X+OrQ9FtCXKKrQ2AT91DJRL2qGw6Wys0MGTLDf1g8vMIsc6t
oXJeKKLqhulcKk3OB1uyy7k7hi/noUu4WlZPCTx/gOVgklCOxmnE9OlWXLC9iTEL
/Ym4buzgXPZDkvbkEJltJpZQFZk2pxwe6i6B7xvMj6G0KjdSMjo2VC5fcZRcTfgb
gen0KzM9SCU8ZzxxskwsIb33YC1ZlmgqTSEF8BanVb0rXWNYkhfvR2GTjQISwmfe
DdL6NGgNcnwCDKblR2EItElm/sNbvpiZW6kw89rNuG77niHaHjEx5sihAALvExoE
EjCkwzaIvT1OBx+o2jR5GeVdVZykXCrR/MzeEeXKiWi4s2YxvyLRwncan3p9Enp8
53YpoP5iqzdH3PA2OC36I1BdTzCBWdMqbR0GX2QAU1Zs49FIEjP3+o3ns2vDZeTn
RKA2YX7T5FpDWyLv/mP/hG7MX7gvUEgdcCKlW/ueSkzbuoWBdkhTl7ymMMmvPPrB
yCbK8iJ129w/xYMsF+F5v7GUMMl3AJCgRkI7OuO1YI98aLlWUEyllOillcR/ugTB
CPE8SFCvPhmSLSL3zaG3lw//aKq8LdtoK2TB8UIRwxebcWYdPjZHKnbTnTdFSRuc
5gOVip8sl8fEGCJ2MpBFSVBbazmHgpHTQH2GEWkquwI95ZzjccAmqeaP5Rhw8LS7
qevAe+ZGpfHgPuA+e/ix+nKZKv/Q0UXLk+KmCUpFhQHlK4wwzx+IlfavERrvQ3M4
QVFNxTIuiO4DVKnJaYNmWYrLO5bXhhf4S5JVF8Ao9UHwawjT8OaufEWDoAxhz+sO
N4IcYybXofEQTJM9ky00fAblPTycXQKiunQm4/u2OronRcgoqqAf9ecEsP3JoGiY
W1QH/AMUTEk0yAPhk1xZBaTx+ICalPDvoRLPes8Ix12KCbM+sY16scCGRXjQLvlQ
ZWqDc6W93OxqNaltKNNteje610W59neEGNBj0mSbzvLgE6uVwyMgpb8mF6Y68tZ4
GzSg73Ciozq2F9UIUza60Dpc+96o/hzfJDzqMYiiVPJRcTV9pAVyNVraBRj9/Tq7
DWVbeeuijsFxw+fA2Y4+7b+q+bkMVaQfYonY4dB/LG9A5B4S4f11c2ULYcikcVsq
1Uud0234Z57l4E3nq1FHtlx9yDaOSXLww+QumHBqqHEe/sbvNVXRX1XDuv3tncwA
yr7Y0TUIMrhQBJkG03q+w7ya/zZTStvj8wxG6ZMtupqpTByoc2U8M6P1+WGLWpfR
PXsWvoYkCzLAVzWU0eUW9OaF+b+oFOyHEk/Q2f2M55v8gcu0PYSQjzpkWHVm6s3+
/KWmhPdSMUSmz9BrKajnkynCGRRZwotJBhclTILga2r2vGEvlIYeyl88C/9UzG0m
ibEpJG/tarTYMb4RpH4WgNi5shBa3ZPpKG6+WW8HzSy4vsz6txNX4Sk8GI4lgQu2
Q91uNtff90I9dPpC15+EKecUbKlQXGyHinYpGWn6ZI/n0pMG/+v36i/FgP14wu5B
O8+FYQYec0qQWN34XEzD8L/HC0LXDqbnQkc9ba1PQdNVOdS1/A8HG4eu4y/wXevb
tLPsHQYAtjMFqRrrulmNFkPOR+OzGXAgD1XT99l2EVnxZbF0HoWWs10Cm7hgPGOx
TTn1qfCBQeEKiR77GmnpsFD6CIPrHtM3ET5mHvV9rTQ7JC0xhMjKrYohFRz6QgAZ
HrMy58KGvpiVSJGllV9yreEpTnp1pDhq2ydZCqklyggBA5D/aWM0Dao2I14RMLPY
x8P4xrBtuKTKzWkViacOTlOSgNYq70tbDB7xfK1RCQ0/UaYWWNja8xOMAD4hrLQ6
F8w8z9c4ZEkuNvYcxf6icOSgLlV33pokkVC4ONKh9ynTI9Nt6PNl6fvTeTSdn59o
S45GXCqvdLy/rB+UatuLme1AxIxgR1CQwjoQYvABYDIIED9KO6Q9r9XoSdnsyjRq
aflm9OXiAspSUBmrhN4hq1zwurZTfiyfYaoQvuLtmYyZMge92h4QqkQSgyOUbCSN
SeyCzIKWDPt4aZ5ZZnFXviyFlKFHGbfhB3vL7TDskIzqdOwmkj6UrI1OxpxbB9U6
pSTnXR6d5llYJgT+0rMO/p7IImm48nhVzoMaP+HlPkynAiGJIiO65XDGvgRjyOFX
Q0HDZ6nbn2bWXKpgVJVEYrOZakG6Oh1s+0WV0k1MngEhOyD/LSglGP9+LuHL4cB7
+udu6lxPxe0hmpjdOdm5TJZ2uVpIriNVczhfaaM7FTNYhVSLjLRDMhjlmDdQVbF3
Q148/Gotg8ei7gZMghaYTtKfPqaWXvOgla3RhMektPvYhFkCgF/dsDmwxlt26t5h
kxTDLmo5bm9dejwhPDViWHUFAYwB1dIrYhzHSlxRgBkjD+UTiCQ1YZ+WoXbwO+cb
/+D7Es53THJhf14gY4YLwcjo6aSvigphrd0jSaaGonMJQs9LboNyLfmaqYQ+dPGS
d8vAX21M1YJGL74cklZB7wLc5LC9mxPVHLwauWydG1xKx++y95+v+94DFGOUp9IO
EHWMwJX5E2/bNap5hpiuiaRAFFUNlTPNh99NMSrP1kKYOZP2yE1Loc6jmn6G/oif
GRfyLY+R4SYP9m7XkF7IJRSwJ9EAyOQa6a9alWhTy5VZvnpzMjABNq7Jrkp3wB/d
4vzT2BEEzZPRIcvhQ5HZ+HsJRxcv2MO0QOqWi8HClOzFcKwBwdzHyt5hWas5ivo4
Aa+wTeONUzSxs+2NqIvVgTKZAMWSdONgPeGaIUKinHlg3zlT7lkjasN31nBLlZEB
5+Wa2eCga6F8BIYvcUmc4qnwRtERy7WohxbY+EG38cRJQiR5VReuElgBe0i/0SQ8
/Hdi36q8Gmg3m5xfJad/1wzmHPTR3bdtfTSRwZiHyvjWlU3a1xVGhAjNLeEz5lDC
xwD4RoP9oOvMUuCMsTWHqSbMNnZUOLgQBkMM/AKuU+On8RYeSsWFpYeWZtOVR2dZ
dJ1G11geSgLXsn9N13zN04Xkh0oZvoPRwmDrxz+HmnyCoxqqtGpncwVjlrS4Eng0
t+sI3wyjnM/LUfLK3NB2IV8xsv4Ho1a9VRv6L16wppU1Uac25lQ8IvrCEGTdVBrk
G3D6ozl7SvGDi59yCZ7o14XQlGCUSjSOuFsqFivkjEEbTURXutQSfzMssWz/2c3L
axkjiMzrv7hXo2Jk6fOdFSkG2GVAtSq1MsWXMBm79RKp7M8U/toEFxGkhQf5bYGX
8WWPTX9QUpICyIW09Ek8qPL0yPFBA+ZFLyQCRYWli9Pf7pwXgrlMsjoZgvmvjy9J
V30X9pZhCZdCM8evZBLCH7YkQKfOmVHQMstQ8hBJx+vRnZEWHNLOwqRkkuWllEv5
CJsbA50xvJBkdgMgeBOmLnefHTcPsR0wd8Wn8NiKGQ2qiy3Gn63eb5GU88e7bbHb
B3pNvY97p8R9X4q3xa4Rsh+6la/cFcRt0ey1uunsu4rIZ9x910dH9iWpugm8ZTxM
+aFEb1FjRNLTRn0CG3LOaQlzZdvDU6WdD7J6A6mk8l5tlon8AznUnvsc/jciL6vb
vNpdStULZshbU0jOxjnQt6UDWl6kSZkKHsAfG9JMxboLokahZePa/DGnbBHaWSRx
FWCDczIoMCwTSDwILqA8+myvzPggsdkwNGWvDXfoDKkzWjBVbHiMOrftwse11TN7
ca2OYLcbMHOQicaZXdzrtFKVFuzZh+iFcWX1X81+du1bmcf2o8DBaJKOtPto/Zmv
yblePNkKTtmw1RRYX0BDsWOvFvjFYIRWZdU7f8X6legfv9RVu+mVed8fat+8Kmrt
WlCuavGQdk5f9o8tOFQHDMWCyZYxnueDoF+oF4qtqV3buiHwizSMnz+nNqcSHD5Y
KwAw3GVrcwRpvZuI3iwCEU4JnOOIkTEMtpegD52SeUSnJOf+BxPG8HJmnpXGJFxo
WKZvWPHIdT1RGXNF3NI6fn6I+e/Nb5jXEH2O/ssfUMj5BzhUPUoadqPHjNF8UKhj
/cTgBF6Xp/+m5KxOUOTwm7mjTAmZ8NzATBoNdS/3+MLxw8wSsWB0WjTFRV+FPVWn
DU0SuxTwPk+te6J8dA6MDXX/ntk3WZwnR2NRwvkQfdQh70ZybnMaTC2cPfgOsj3J
yPnJhicyVjNp08/9omZh6D3GnqqFbOwE5fItTk6ogcjWgFeAwlR2r8rGOgZFsziI
MtrKADeoz6QR6LltmhL4Cujkk09GAm51VjmJji4apmmPx/0sNNoXdabFo40dBbXl
HDpCYodAlKAIB2uMe6nhBUEnAakGdWZRU4bjV7uEwWOcLORJ/J3gjy5b+4IGItsJ
9BCRqF/sH0YM/E/7ZXqp7+4QNTpN6Mhg75R+fRjJX3u3H6rBbUWlLEaTGXU5iyUE
j+CiCM2dBjlgliSXUfHzubCesMX/lANXe2wWZUgehtR+YjkVcfLTlOT0QzE5CZWk
ivBdEBQ6XRsLBy89TZVtKtsjfnkrDoSY3Vy7UxqTeSPEviIn8GJdmiOxcMkUXRM6
qd7upM+frBtYhgKpFxqHEfWUlGgJalZGh6CPFXrgNL9U+84n9xtK3xqlm4mJDlDQ
ZEwiUkQSR7lnrefJ+i1QFpOyqptMqoQDk84zLOcGsd1B07obpCTuWS6YHpOBDzkT
HtIVhYwGBE/rPCom234pQn0KjRPFBB9ir/8nZkV0z5DFWI/K3Sf/jpLAPBF+D0X1
JH/maf+3eIzdskwU1C1PMQOaNOrC6Z58KO8t9qnbFe+lo5UV6EzNpSkJcbfv/ltY
TwxQe5JUCSrH0gqAPZsBEWaYAiCwIQorCEU8fvwFGwjSs6cKE0MIlttNYEJmroOd
PHOuQKPJFfj8jJnaDxSnNwbi3kq2mYhMMo12YQ1nYlGrLsLvhSE4TV1B4tLkQ/4D
FqZo910C67l6Onuhgk02eUwlGwFNN6dgJ6p9TtRmP+BrpepPCpN0eAav00jok/nI
GkOrWQPjM2QojQK+fbHfaEy7GKGrOwBDScSMsIEKNgAFQxtv67VfJMlnRW2J+Oam
Y+2Gbd7bpKULrWeJcoHTuu4d8XmcNxyjfwcO+POos3y9vM8buLnRrT3RWJI/1Jp5
5nH0OnoQ58A8nusUpJ4H/88PRka0MlQCPZ/VYxM81LkJ6GEhvQ8LoS/vgkjeLxzk
EsX6Ng1/1gC8EKTIkAKnH0iiL9R1Ma5TWwjC8ph3sOov352q4NZCPs/0LHsXh5by
9lYCJ6eodWmTDdHe+vNTljf4+WoDnyJSvXBASEUyRjUdLuglB/VhhPRi3Jffp89T
XAl1AQRAPBwgRmfJe56PZ5EpqEfaJKUOubxsTBJ6PO/3A02gK5D2vZetxXzGAOvD
oL+dcztdtqbn3YXtr3frPf6xVrDR8glSRqHYHOdAXkYbLFyBiFFS3ZyxiXOG2//7
nZKsBbCZn7c2iaajxpQHWXUk1AmJqX5IZWei/KIJfX8CM83RVtLatKeqVdiDv8s0
5lbi/zM6zm7yqzOCRS5OL1XqZfikRVJFV0x/BfIQFNKOGmNTNXEU71mWQs0gYpyV
k1DOa1TPoAujW+Bl4jN+pg9MutPeOldBzkHmMa0gW5R0vviZ1MVWmNoozYH7y+1G
a9Ph060IwyDWf5hOhD1rKX1mB/G/xuJECY320c4/ISP8ONB5lKEqTbJBgQBpsrHF
5ibFFtFcIaW1g9Z2Qxpbu4qYYgoe73Qf9kJQOi/C4R2pYR1fVAUKMsZ55kV4hUV2
fGclIbsoTVJYHgI5lQxQDuKgDsKFEYrjMIPSgX7w/12wCJADHfAHbIEp1bemUxsM
rxU40j8UJw0+gtTE/vuL5H398k7pVfIsfMVmkpQBdNU/ryVvnKHOoJnMtSgZBh7k
hpDCWyhHItiWzaDiagfxIblcMtIspDqSRqSQ7dD6jPfCQz+LJzMvflbQgM5Ejtvz
rfQmToxTW8HEjjehexrosRXUVjNwTb8GsbjimSioa5qSWxMa39yPU/U0Gt2vAf6D
F4Hs9txJNYjOTEUer5n+COaoa+FShGNk5W4upfvgkc1Rlp7Ia9U9D6IPA7c1kulo
BGzM3Lg71VaSfbh8sbUyhj8wBFWo6dOm36mz1thappHuATOSvlVc3FHq1xVkK2TH
v4IZ+shQxLzW4FxD2AGQ+x5gDwh8Q5AZWQl+571MXOp4aoNjf0cxtZ3qFAq52Q5B
kllCtgrP9f7wv7rbzhM4eCbrXMEE9WPla2ZAvANXxVcyK/WuZ/TYpDRIU7GiyiB1
4fNB12XPo8qnCZWfJhRi2vjX3wPHo4d5ywCNTk/Ifd8JgP3nqfvpSlas4dEGtMIe
3z9PyQT0RQ8ysoitOb3mfU94NMAWMGgtL+b/njorUopib81NH3wzZiiZGbMoNPCW
oftIbHSZKmwDEliMH0Xb49Dw2bMOLa9rA6+SjlQM2/WdSrbYFieUX7SL/HUrlPL7
kjXAlqzCezh4m1I4Top/1m8ulne6IfWx/Bg/riUPQJuisjBowJIpDiiU+zQEpn4b
NgGC9PZDbN1MFK1m5fTxypNejBnTlvsD/twbp0uCojT5tiNAyQMz6cX2Lm8ZND9T
GfieapdclH4YDY+Ny8O/Rpsvv/Jv52s7zCidf/Nw+zzXvEFSAxARX364+p4XERz2
PwmvhyVjY3vOvi/phPDx4XMrlvtWRSMYKjb3xkBNTlQX4VOTbt0dulVXvDly5/XL
1kxSsJwOqYWPjDS0RaShBrqdS016sZDZjwco17cAsQmOzqXlDa3SsnvP87I0owsO
MO0WXbp2ALA4h+1oUlIwP0SL9uKjOBjDPVjgtvw23JmGoXwVu/sClfW8pDKGWCEJ
UXHrwgfPx5o2hkMNSqQuabszmw+qgN1QITWEzeVtQQUCttTHep2GApJANJzj3vf8
S8tp0jQcyOpGVyjsacm8X8Y/+bNmjKKj9O4/BnlrZtvH9Q2RM0eXYJsLQGFbQNot
3hYESqiUkw+aLMgfTChWfLFPLqoLvn6NKwzKMnyoEkCidOK8QHCAbzoKKvSMQCBP
yrIcx6tQrnKAb9sqOBVu39LJDwbpZta73SOTFJMJbagxkvpkkj1Mcy8qAX97HXdJ
fqb/3c0OkB1EzBEU4VN5FJLB+wYgY/CjBzmr1UVHhmE73HpemgqUgLv8AN1TVPgq
zt1wyOAWIgjvWJajtr6mA/ZtrkWvwUXv7oX41XpjHKN9KxrRzdy+tiQfX5vSlVsn
Dn0ymx+DUyjqyiMt0/mLuKrOVVGqXtXZN1J52PHAme3XlClSr/iQfcEOHcpf+YQZ
/3Xv3F2lBnUyU8S7YGwrzRSOPGP2du9C00eGbJfHEHsdcTMLW6fRJ+QBtYqOm88p
bhAgSddQ+UH2chMH3UCeyQdAqxgIibRvZa2BOimBVCCxdXJKR1suxPXkKSSeBP9a
BzPqIigXgrCVMcBc9qUjB3k81HLfe0n57N+Y6Zxv+YdCKH4+MAny7+H2ruN6FV/X
oh1gzR38uWeHVL6tjnXTv3++rGGLVUXjfPxXVpR4axCd3nlLXj7voIl/CswoIgnh
o2+kNrMTkW8sYtjUQvjFcSId7H3P0iiZOBfMGpgxZ9l94+AofMSWlQVKk4dbHxIa
lD6xKmwmJ8YF81qG90ZY8NyWqeUJTaeFryf13B5jVmDNN6VpgRyPVff5XU7GsJMy
QdDE8fUXkHUKWPT4Dd3vzmP9kdxiZ6ClCi6L9XVvAdPOzoBwhBHvVR3kNVE17nW0
KW0Hsn1hPnxNoejcKkO1dWPFvvoHlUp7tooiv+EPoumZVg7KFAYWw3+ZwEtwexbq
Fb6CF8nuSQ047Wo0DSxCUcS3sKvw/X59YRSeazuvYDlMGIxAEGrzlCENp3lHPDSE
BTkBiKcDmFKbYXtji8K1a1HzhrcAHLcGRe2CW0aP9w8J6+NHxBL2ySi6WccyL5UF
pJWfLmBlWbaWAKcY7chUGZ6d0vSV+16pEgFEEUU221yro5ZmDI2lM9Wx+JRJX03M
tQZGYXDl1h0yKeTjjPDoAvbQuHm3fIEW/ikgzCKoCavlliGSUUPHRQe/Vuq+nUvF
ZvefwH2PpIJPSV0wQpvAjA3tLZ7GKdcK2qlggsV0NN1Gov3Dysyq4U/Ubv8qeBnO
bjwt58zLN7OaMXs/qzfzypCGJHTcaeWlzMYVT1KNfOuP0RmaZlS5TH95L9qt2Y7G
D0oeZWo6BBZtPyAW4NgI8yTCLCDc4R1I183cePntEfk3kfwCq/7UP8K5dJXpgbNW
jQ/j2Hjt5JxDnJZXVFU1UFXK7RSfgXHQugmM8VVtAQxafehH1vmn11okzZ3ZUeBi
TH5zcU7Erj9m+ghcDzJ/rTWBdQSyhRoRViONtkQ2dINl3Fuviaq9QypvfA5/L8Tj
oRxNW1RUjBsbmQ8P8Kg63x6Epf2gN/OwUNQ1M7Xq/gCB6nsyP/ehU1l/YAu2yFxp
PllEyakP0+i9c2gC5l3on6gO42FK4wJydRwH2026QoOaIXOmaYQVvBD0Ce3h7596
1Fj211grvnD/LEEqTqL2xKgFNvjcNzH+WAZboe32DiHzeCMH7Yu2XaU0+d5lt8id
2lOQNRk1m2M68IE/NtBMtxf+zTi+iMU1N4uXaoq9j2InfZqT2UloLgNZd9vHyBvJ
Cdt9Tcb5rYRY+CNCBrXPZ4eM+h7U5jaIFWC3tFZa52utzK6lgW2DFlAJHd2wmNRd
O/n3paM6/Vwxcv5NByDE+vkDAKZgxSc8a/vKyNAKMMQWdHgDpCvAkfTbMUIM6CLv
WEwrReIoIE4+BeUWS7F/LbG3sBVfV+AO65RLRMqsmYahLSwChSxXABIjQrV8PBJT
gpw0re6fxHAbl0woMs5D9tLVS0hihU+j6UEw9Hk5YHcWXyqqRbg3YxJMeNtOZGqr
T3NxrNM7d6ONf5UQIKow5DtDMkkgx6HxQ+aMaYyIdiLvJ5HTSijtYpvB+Ri7gLhL
vUn3+PBm0R3QLx8hiXLkbnc0rmIZRns9MeockoH0Z5Lv6XM72DNROAxTBVQSbPLP
Jc5JwQwge8OeGEh3+vRzYmprRszMrWmF7UwokPJtCCkzyibzelI+6kxxPSyQAYEp
5yqgHHHl5rSXX4p8T9ydrL8v6jtaFtfSxKVPhsTkqlV+zelq5KdU2qzPc95cT7Sb
5q/YuWkOA2KVzUhprBGAYNMQlwrewij4+NZn2chRcBhA6mYlAF68t/lqqNGYk3jX
6EgRMOeJSegFxp/g/Ghlfa9COF5bR4YhZIfeaQ497Fbk3JHvIEFo+yoWjBWsAz5P
jzh4/uOsNAIiKmtrhSlYPMq/on9tQFcZGt9kBGFX53E4HPBjr/kS6qIbtZcUmvOH
lELYiwgBE2/iyb73An7oaP1n8gIJ9pTiiNpSWsP1jqHWnCjjpO+oBz5Y7NQmexAt
WOUY/eaLq8TBYtJmVjHcfTWKbt0OQyu1bk6nxAmbY0af7VIz1VafKr0+cvtQuBqO
Ib47waQSqnG9g/f84J/I1SRvCYEheYzLEX+6mdE6Cw1IQBtPuH+m3cah4AAyHq7o
fu89bDIlkL8T3Mn1G9ovL3cpjTANzmaSnjSN/G52RTNnwCjawCFt7BxbE5HIvcfN
P2RefJ67Ri0P++K7R4Hy5s4nE2FeRnG6iCWITtUO5a34PGk/xCqH+xHThhgfY2Y2
DXjawh193wP8QgKxtTPYUJXAzq5H70LMwnMyZ6gtF9D2YVzdK5YzeCxJjouxUMrr
Y0k+txBN+rEqZQJRQRgcphup/mczdlbq0/vTTc2rti6PZDlMTHOkj4YAZeHeqQO0
uV8hvWiY4DDWyRjSo+b9AFkubf1MPmsxIsHwN5W7jNHeQ3TM2WONbkv5nNCP0j+C
ZsPFX7hzsgC8PMRh/3Bk88grzDFsKTf2oeyO3X2oBYZOkGJOwEofo8TEKqOqqLZv
U0hg8WNA9bjC6gZQ9Jf0QprRJynDN7io4pjOzaCirtobfJmciEJXvjAXI88QUb8L
KG547vucPPi+kirsIaOEOGm7uY1ENaWevO8ComI0wsdS+6NH2quFCkSyom6JEYiE
IeNaqTcUqGbxWXzP2Kt6OMZsKTPZPbRrFMBW4w2fOgbZqyZtdrRk9AkZPmQ7JiiV
OFk+tEgPXNJ9AsiRoERkjSwqNGHltgACcTSO/uC0qqRnpH8/Z8rfSqPCFf92yxlq
18r+gxoy/i/6YFOVdnq/CuKP8tXuRomcJyExRDzesE8nkGQClXjQVRBt+5TqxBWZ
g+t65s9oxrQs55TexpK6udBPJ0r5AzIMZozxuKYJSEmYnDW0H1J1ly4xl5CEBRuk
2KeL/VGc8D35EHtMqp+OOfXDiYuF+nPkxWrasShmCD6XKHOdNxcPjLlRr88L7n+6
0vh6+vfuLYxmRsM8DKeuomeU5yfN8Ol1HLw9Q5EakGO/0ZGc/K0IlkCXIUFWJtsC
sO6wr+jc9nZ0BZFjz6+jPXh6UCbRARTglHt9dpL/3xTN0VxDNEi/wFv9mn6Nv2xv
7Ra7vTUm5xU4lRrkE7g919b4L7m8FJ3TNtOKhcYZlfmmUNsLRC3dSD4EXwEEoWkn
mxIFbtMKkllCWqC1ALZnz2204bOOodC8O2uPY6+ZmvBgQmirj+zRXeVq7Pw+97H3
WaEDCqdXBzwnyCl10/AMr9+AtrN2KWbLvBv2/r7QkRLEnNqd9n8GHH4vklStyp8d
0m8dhWegyChxTp4HhmKIb9xsdyGMOn0z9W87afoI3c4c4/Kk+30+qhWKgvQSZrSF
QP4AdqAYxKQnil6W+vR6Wn5hqAjakyD0OYONSaszNZEYCMfEHkCXI/gaWnKBw15n
kowzBkUFSmq3Vx/CHIeg5qjvhH9/1UpOPE1GynEzCFaJQjCswW0IWI2yPg6X15dA
iNJZmy0rRTzc022PoKW78mmDakR0Sndky5fiiN8Zo89Xpg4wtjWptatxFKSntHcN
gAoi8qlRoigdS7Lp5+Jd7vne6aiUg+BuLGO+K8Z0B7ZTyLR//4c8Y7kNB3y+Jx+r
tA5AOpEf1hLFGbapP0POVIcoylzBdLdZv2dFV3JpG9fDXDktisGrgwa8zStN/ZTk
fhQw29I7QZGM697WDVLiQyJ3duOfZugwmKbbNA1pW/ARr+RzyChZFT7YDCvQ92Vs
g9ladq4fhNCGLhmHZ9QyVsrZbm6mRgwuJ2EMDspDe3V9Ja5FAiHQvqviq+YY0fDk
8cPyvUz2FDZyclmTsgWbTm5QaIh/a7mIKCwHM7EqhHtbEOQhst7GLmz5LWgAGRWJ
/65HLazzeh6Ujl0sMgRyH/USox9Z1wvat1qu3irxAhls0gH+CgY7x1i1fXYGBDzy
PpcMq2h6AcyC4xAByRoHbOj/p4hbtjtFAbKeEVuIbpCycnThJ+m4V7zXdILqmsqj
rmSZEmOclFSAEiewU/dpX1cXJwnh6tRRUB6lmMLuB+f1rgzdoXe9djhA4QOWWwGm
631MmBvqPFfrF3mvhjEqVJnfIiJHLPuwFdrczGNdbrhaksNFfbUb1jtMVpJFQ6yj
OXMxTxsmhxGuIRE88Znc9SoXYwiWrlKrYY2WA2QdXxcLywIaM2Bg1mQFv4iEdpYs
2udRQN8Eg98cAWk4N+X2Y88p0GucnmuwLDxdNB+t4SqS099wAaLuCzP/fILGOvOQ
7cM2WzRbgHjLKTe6WH50EeeacNLVOCSHVibnE7/8rR7YZLY9vXJ6K/WEmBsuukZX
JyFzRFkaihh8ly8Qpdf/mb0s/ApGGJ6hoM+vkxCpKLs/LKDsRlXJOoguVeYWJnQj
/DcN0fxpMpc9TId5T+A/66m4YyatYQKDofwu+C2oIorcflh8uBPONrMVQX/zLaY1
XZ8v0eJucuOos7Yjn69DyS3PhZ+mPVB6atYV716qjR7/74fun9umck9qNK3hkNvF
lcC3cIlE+YFnZb+NtCtobie/NRQhXl8r4X0kKs2XbsseciT4pnnNbo9HtFYBazoI
GwR5eFZbFaTTQp2snJ1LYOQ8Lv0+lNKRcThRdJ8qJTDvCeM9d4Rtb363H+l1Av+G
bZ0oxuWXoJXtOKmhD4jlxb1YukrmdCIUhY9zDqsTu8Xwa173xDAQmd3TyotlcAwN
vsWCLCOnHoSirOIebXGrJSbY+A7gD2oL/roipEW9xxikbrt3bnRwtpXGOuRccDeu
gGLf5y6jyQrl22ZnjbgVgrnTJY/Yl4rBfGPya0naz1rqujgHrUPyBfsAj1HmkvPW
e1AcHdoaO2G01X23PgwPyKxsLpGXfTKPeKKFSh+m60GKiZF+Dxk7PDxoSwEli/D9
q4gBDAZvndZZZ0fPFdxttf36NYyRprEFujbXPoUTLgG9w6aol/2IIp39p2zSqe+c
pf98rvcZbI+0lGYxcEsU3JH+qKvuYcZyfm7sHrfycV3ydE7jD25iF25zd++/wAPm
vlEXjmzrO09N15sSe1JQ0Ywa536yfwnRyYyIk8WHsJzPF3oICcjW0ULhyU7rO1Uc
XxsJ0Y78WgaYL5xIiA3u3SBzFJqNp0GwStbrfatVheP5T8v3ZdZ0Yo0hrsLWPIpa
+Sx8cXfj2KNHbNNS0s+/zoYJWR27lb9tz0xpDTkAmzCtuiH29L3wduN0pmybjPvG
25KxhBJCEyjFolYozXTojMLa7NzhA5/NC9g427v/SIUPlqUt1IGXqv1oYs7kbzn/
4qNqerII850We2rqg75DSKIc/5eUnFImoSsn6oF/iNQkcxVLs3aRs3lqauR5gBSJ
+wRPRSLQiRcB1TgERoDwpWX6YtWzDoWR2bcF+l+YiuUeYd92xCoKej7xn7vgwPQS
wk0IGUD1IZ9FvmXDP/XoIHOQ47P+BH9mGjnzGqSsnxTAGCCmRT+QcPmZmiJfuQ26
5ZWZOjEvtt8b7OWfQgA70PS41G8mDhRfFkSkX9deb6T/BMkyX8v8nXRQnCi3koVE
T39WVxgB2WzCWi+55cDDIs/PHqYlrues8NXc0GwVV4lIhHMkMZbEUuarERs9d1pk
jxez8oEp/jxkyNRkyp+FmzOOmgE+kFpaxRvfjjmAhFZRys195YGmLzxI743BeZm/
D6UoQtbxkyGz7JITpHxncf2oBr12/M3aMImJvNFWKeQARXqOx3VLfPFcA8g6I5as
i338gcZAwdqCLUQH2hcI/Kaz9D6vxvG3sOCXYBYI1jryR0gbL6RKuTqeuaSSS/fX
IY9D1SJY7t/Gd5zTYdPPOuwSfPZGMcXAirvcqB0G5r4J/K3qQSyVl7TZfesTo4wk
GSIaEsMnaJzO6HKzoakHz3Z1JJ8CjglxiZkpuoA1DQy7sHbU311Cva9OOgGq5373
j8f74eyXeUVXTw6xZgzMyfQMz8PWraq8alobrpPeguVn7d+YzHQ2KjYubmaojyH5
gsnGV0mf+osdRV8YP0pfhUQLkzl1aLTG8bXucYSblQ2I+u1G9AOpd0M1CySKyi9l
LKaW42Adc93dwfDxkxFZrlsdjmwe72cZSG3ycwJqgo6U8rUHWn8H5kO4sk3Clr/E
R/hlg7cuFuq1Qcbc3iuwZcP4Drt67e4LbFzsS/WdxclvoWpnGXtjs/xsxzvnCWJO
o3ve1E9uE7VmXYkRleKrnjdOQ9Zsw1pW/OHIYXwB27tA22Ac/38srZcGRjXDKnAI
J6kREtYDwTgQlsL8++Vak7+DJoR9+c7YAZNrx363Boum1Gh3THUX78FuQ0oWygS2
0OuRw9Qv9RBRsDhRiIJWdbL/UQdjcr2v4RIELhvA4rlxfU1i2htEIlsjZFxdK1Ao
HybsKKZcz46n6hzVkBpYsDQEk5ajodI73npIOj3buAJI7WPbPrZcHrxaWIM4Kk3x
vlXMBkKp77LvfcAbqqekv+/v6jyfs5+5vawPUYxoXHfua9pT8oxsvPnHIE7bJgNb
cbFFwJUjmEuEKjWTvTC+YS4qV9L+O+VUjPuGk2E1aRHeEuUQNLP84uBDIy1+bgZz
EUbzhiqcu3NbtLxl1pNHWnb4c3ftW0pBnyOgnWth7ABuXKRrFF4ocfSb44HUcjmY
WbTaDuxkBY2gsO//vZcA0ZGikm4cpXAyS8mGxh/Lv+YiKeX5+Pc3IyT3CfGYbk6o
0bRv3aY7vfTBiJb+aVn3yOXkstFJysXVh3/H5JHuKmgGcWZWaQVbXsRGILK66kpg
xOqN9bh0dSRB997t8p8G5abn8AAYmRJEkGe5hw2sVc51Ujk9zuAvTistz6yqoDK7
ufNjyzi/vPCJW5hMiqibz0aDmT1Uvdb83tDC2oc4V1fxON7zjL9bmqh8PU+hudxl
9L04QhbY+L6me2pplaNnAlbFKJ06Ffabt+eW0An36WQmjF8++2Zv/PXqnywIVZqb
1VZkwwghxlNvz9d9rUN6GzXIPgtvcWuYfn8VC7on0SeNbGSJJEo2ObansttJyvgH
sToLkeBfiD9P6AfFk+8Y0mQmwalmKKNUT2LtLeky9aa2X5gL2I/vCAuLZZmNblWf
WGIPnVrlSizgCooHo3nCOpKMcDZcgPhP5h/MBnc39+O013vKn12Tox/5Ip1X7cGk
rIWRaM3xcYIXiWD6h7jObzBd5miz+yV2tKoJ8GXjDKNxkdYEqw1BVCzyjrw3gy7K
haykDDKtNnWNJuDuSGvlm/MXMNLAOBJOxkECyLybpR6GsbqOj9Gbx8ImE9K8Vg+K
0f2lyLb8IaYnrkbenrsptK2NRvIWPC0gQDjXj1h7lnJrve6guqbXl+/8W9Q4cebk
VxKFFNdaEHceS5/+h69DO6/DPQUGRRE35DTkIWBz9gzq7uCgoEvoBKM9oGKKrpzw
cXL8sNz8bI4mW5i44vWun46q4hP/URbjXFcQYjyiz32H8j/YHtWUNzXNalg9o9a4
QJmlLqrk38gRVDn2EiNYZafNIFefq1JI/tpacK+hhfaM5XA9sklmoG7cqdrSDoTB
y5cEqblz0kiAIyKrwhrqJIxy2NHDdc5bPO2/ohkjKFV1G1L2oY/KAhIUNgrZWPac
QZv17phuoNrZyhQUUnlI95dEclqfPsJnkOdtu2CrB8QBai8he2RtedKYod6ELc+H
4BLw0bWq6yBHyt2tHtoOuadzPkOzsOYbkX/CkT2WCB1l1Un1V7VlLW0VEtViaEwB
CYbeD7rib/UqBOB084eWD5z60YOcxbhszU5HBrUxDopgA96Fsnjs3TNVT+kooIA3
u5zjdNYqXRNoqrI+sG2LtxWEi+OakGL6SmS0Ftcbf7wFHDxiZjfzjqUwSzAcEc2p
cNHxQqf00FAnDA4v5j3L5Mm0T3+FOMbEbwax6v5E5D9+5COcSfAnwj8CWXX+NWer
buA0cci3to4gp8Cq1cFZKX8o3X4eDrKenqB9CuwBJ/IJU1pet7Ut5+aqHD3xUD8R
lwkBFi/Iwg9vkXCfxTXu325i16W9lG8qngpfFS2WNNTSZGK3sHiL+GHxJa4me9yk
NlxAxhLTa8RcKA8jaMYJhNadBEybeuBHgSJ9pA+3Z4px0LRMv9ndwZxBTlN32YLc
y2hAcWptaN9bzoPCVHmtpnhGYtNFTXnhexNbQe2HS88TReej2GotADOT6/Ffvfdj
Ha6eOdfXJpiJEKX2Ox/vCPNM1P0Fi9ix3sJuM/p10VwodrnD7aqqgCc5wFicGR3X
qIPOHq+Y8s71b5f218CTt2+CEfQ91/4IVcCtTTWE/QffK9jFtOuVB7uRj1NecOBl
oGWD9rvq5zR656O8EKDNtriczmRRKeoSgWetYezr7JI/Mi+CsiBjevUTLNo6Omoo
jEdQ8XZ6JPwLc8wjK14PsxI/LFMBAnIg8XYLUjDA9X75D/eDxTDrpbPMlzCfyTx6
q+u0bbmRIrn7Cy5HHcVqtdBPLQZbf8YeZwB9lq7o441ceCukMTmYFIAjZbTopavx
9sObmAJlUF5shaiZwHM4miYqNHS6hu1X9SmVNTSfWdViJwSx//estXnmxDAOp+dF
anihUsjx8QBR9sBlNvbv4sd38YvIhaSY2dxWxAyInTEWqOdJ44gYNCLUYsPugzNS
PYRLYUuMACiCnmWlYBcBssEPlPWZhRFpkQF5esmOjgVActK4eWo6BsxHPJMRRest
mEyLUuZrSDap7piJIEI/OtXLpRbs5QWBMZ+u+PWD4P4l9sHz9Pid32z0HOWIHAYO
mLjyEACbojKw8pTm4gsw3EB1JMj5XmPDd2ishSyUphw1Oji9cN21sc7WPrQX85ki
76mHfmJOqx5U+7wGF6j9bDJxS1OFwVe3IpaEYfBvbZkeEZ/RvdHEs9JERpB6Krgt
+t24dN3k9MygYRaDDmLSNaUOU3ML/BPU2sdcWup1VHV4M8dTq/f8QLYpZ6pi+QNi
Naq9+mSCK2DhWlKnFd8lUt6yjAvl+5xVrHQzDSXuwaUMlfIiyMwSixz2gtPgBhRJ
lsafdb6CU8WTsN53byjjQYYu97h+KDsbYQxNYpCZ9aU7QH/eiCECI9az/t5Gto4w
y8x+WH/aGOX1P2nnIc8CEWUDvVDweJwV9+bQlBffuiANASNbgUAd2t1RKuaPdo7w
YdBqzOd/M7IWVhHNl3rhSB6fxYhiM+ChR7sSIRUF/j8hriBEeEs48OipNOG3n1x3
eG1BD78zpYWPBMh7rkotBJfzZYDvNjJYt+Zai9sXvWLTfHUc3r1NfpUuxz1vXLuY
ZT6aFb/3PVkqnWkSXnPTfv4M4zWh2n50ewYG7CEHzVWp9I2DbgShOhr/VnYKXIuH
AJcNeLyktdjVlBqPtx9WiLCZYS7efT/67ikp5HEaHUB5PlByB9ISPlSMb4cRGdmu
vwFOpiF3hxWnFhb7uPX02kNbiaR5fz//e0xP1TW5PmBkugkyyHzFn2woryjdxiSE
hiBqEBRlh9owkzMVKz8c2piwuwv5R/k1K8Yx5qSNYlkhSoZu6E0LCMlwY6gU1D4j
/CfUmJ7Frp5xhsnlsYusn0vlXVNo1DeagdDkyCJRBrXxd3f6pIkidZ+MQnWRI/x1
DwIBLkLsVQ5GqIq9jE8ha/xJulrpYOUTWht1OOxQ3JB3SoL8hvpIrb+u4qI88ojm
2gDTVNpbgC60A5Ruqgcv8KNyqXUFznqpxcwGy5/oCsx68nNI3PzZfoqZYMq0ZU7p
Q4CtFc4NAK7ta44dNRDx1fhcbmQ7zgt0WiOZCC5xI9P2FsMdiaKSaESmidiaIT4q
BoWQF3CzV3BjehwfpTFAXaRTJ0y9nAydKYpNEqYUx/n0JwIFMI9KPWQOIXlI7azl
qP1JDmm8qbUiO0nO7IjFYYCX6TZ/EkrXsV+rC2HcJIH26PyKNF/T1Y6s+KWVpl1a
Q828EuzwlUoUnnBQ9it2JFmZQsxs5vx0FZvw8Xsjxy53QZhOWaUGGdr2BGGisS4J
hJOEnvOx/jtVnOgylusaVFgPG6cT48Hzh40UUai72eVc/YCBmGoTWCENwnbM+7Vn
EYcrvZN5t/5U+z52Cva/Zl2S/GHGp4vbuPuOQ5xcK0bUdeMQq/zsXFAMUNxHyerP
zbkTNI+lHPUGUedNxgcv3hOdHMcak9VSQJvs/UCeXXId9VYQnT3O4e65xLBzXL3e
0piFKYZVqQ0JauoaNCNAmOJ/7PxKokGqLKxCtqFWnK3alKwjs33IWF4wjwM6fWtx
UIlE3xqG2QZ3L1x7NuSE8Ykl7ACjS0LhfLok3x/59A/73JHRjTDnTjmDsuflMG/6
UEuqLHxoyXVlOmpCScLu8uRncw/rUJ0vig2gc7wiaXItn+vlJdACUbHhYbpVmHpp
E2Vi1d8Nu12mNwATnYJcXn2g7PXwD4kDOKxCJoE8KIc=
`protect end_protected
