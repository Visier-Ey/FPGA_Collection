-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
xYQWuoK0TIFC7sfirknB6WWhSqWE8DSVkp8z/L/s2xMTOFP5HcpNdln0OdG6HrAyeDQXMHLeh94u
p/MBLdhdUbAllauc0WF1waGv0A2EUEfMowgR78oEK4zYApWu6M7OkEnuZCoqcDAYQPiRVUuOOae/
/j+Y9yIfV/knzqNxfcTP7nrUC3g2p3X335IVZbaLC1yOogRkOa7BVBQ4PKIXJeZd9gIvoqtXgEJ5
7KlZ0axbFQkbyx6YvpgueCX23Y+FIN91ms6tvhgYTue/najl8463cWO6fZbDr9+2F8pbQDYo4rrX
OFHfGa2x23rDRj+ekuD5WcNqlhFQfjVBd6hfYw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 34720)
`protect data_block
P15DVi5bbPibjtEzMPypY/VI9YU+trBy5oLzBc4E8ucVbNe+ciEFQd4oA6Uf4qq5Y3rnqVIDrzIS
l3JhqMHixUrPiKxxbJmmOjMghqMJzO+3tKXwXc4dzlbvenEDcsUDQO0UY6FEiC4TB3jxxgZGAOth
A8WBh4ucjjiSYBLTq06pFYodXQ5nVF/znKtDciiLkHxqCDwp3lmY85Ou5LJHGEd0+czb6bOXlk8d
iUhPRVh69fjf+NKT1iPrSWPXp0KCS6j3wfV/VhtYmnWYMzGtcMiUMsh+TTjQKQCLN63Fw+FOUNsI
utxNitapIM1To3h15F2kL4GMfYsE1wE716OZfDeg2p87nqmv5jb3BRUv++j4gbnGz/vGdKG2GQsU
svVPslh//sdm6Pi7jwdawxB4kesFWhpp2KdUwm5erSrX0Kk6DCs95uEpZEpDLLQDtEZ0pG8UdM29
bR1LcWwOiYT0JIAJ7RJ6SyZHjUVB6VG4Zsz8UDts6qslGQzBCsAJFC+0Qq3rYLARRz/BKd550usU
HvZrcyeK0Lsjp0UQiieXU23rjL1YoCTAb8Ok24+yYOaNYNrwMKiSBjyH2Ns7yO6pzZD/nXEQUCdC
x+dp7fY6fz9DZ+/oXfxFTFBh4QBj4JhzmZ74pnROgScQ1q1X7tAwc5wCEOFCIsMeIaAKWVwMfn9T
w6ZuBNiGDXKVF3c7YU5fgWy3ENFhWGFJ3TnvT0Gbw2dW0LcrkTVC6XLOPNgsKHPDdF020dVrvv8m
LMp4xZlcxFLHRRAguTBPECRelffy69vP59vZS/Ar2mJhUgc6E56634nrCQ4wuUhg4E3nN4FYKa1y
3gAzinGS0a5rL8nzGYzTe7TDfE5QoDM7WUdwOJ5vfOrZjNJbmxOpyFfWKiACIw6MH2tYeD6Bsp3Q
bH80zc8S3IhSZ8J50JWyz2DbpQQio3/7vB5RJaSpU7S+ZtHRBYcV7wg7WxVFkE3PElJndkPQ44v+
ioL3wwvD7BaK7lTeLn9SCjAHzJL/BDWkcQYe0cMmreRRLuCIrS6NOAQ8pFRVrpJRUSgID+4V0TlH
COdd4B6UMWErL9sNXcYAN/ewoAoKHSiPCg2o6M2A5gxYGeH0t0Lu1hWuoVN1ZIBcYGMq1gVhMMWc
OuR8jOxzKXyWEu/Ug02lGTGjjztAaclRy8rGfs9tvQIIJQPLPfBwWWrJkiJL2YcILmHAWfBR9tbM
A7aUN+3KiFeFMMsB1akXtH1W5E9c//BdvsvKHA1WmXVWT9HEOWkPhR8bQKaleUoHdgHNt2AqZGFD
Gt4t0REh8HWThy6EciutYDLibgZ3IPoPKWFydaT3qwByO4aldwIRAFj/4U/hW14CehmtgYHy9J89
Ks7yZ3MSACEp5V5a6eEU1ZibjTDcXhlZycEWuotnsYO7Fw6aL5NTELmWP0MpIP4VTdwrVQqEWCt9
5DRQWnOSoSiVfrBM3TbDCaFzrF5CPP9aPSSA0WwhEGSzge5Tb2J+5kXekqyckebTbuX7K/25dGx/
BxlBia4cIcEntynrZwZdZw1S+9FHm3imEpoEWCNTU8U7kL6ncp3FNIE4uzb1uFaPoLigO4tp5Kic
Yiwk4ZoF2MQ7NWjq5bTS9C70AGJSBJ9zueg0kuscZhT7rguaaLB4nUXn8f0AHeZA3apcqn/OI3RU
3TcrJVXGS/bNfw4ufmyYciY0uYADKMf7IGeeX7zsvg1KLjCwm+IqSocCJSGYhSd4VV71CgxzwCbB
wIOyynlnGmlYEgmDKl+DGE6v1jTaN5AdyIkoAitI29oPPYiybCVj6tYBiiVSsPhh2INX/O2eIMdp
eP4QFuEL/t1kXlMecLTkrlnVVspHVKQLRKjZAXv5xOY2xUIV34eNIn4fXOs3xKQCN11kBQEib8Ax
p7oCf1yjhyEElj0ftE3ajI6ly+Awl+TfsD35dZQg/t3sm73FTtPhMhd7chWqqC/Kp+O2Abzmt+VR
oRZckcNCbALhiIWiylupNN1u8T+gLKD4/5SCOhLHWcP2DEWcTT4UTH5PRBln7hWA5FOsObQNqxon
c5lqMNeAVGye9zvYkohU/Rpl/oDxjsVBoGGVcIcWkGdnza98CqmEDi/Q4NTFM9j3AabMw6EhHeY4
ZmSH6QHYW5ZkA71lzoRpzo41VxYI8ykwZBEMRY8rW5j2nayiiZzQ8Cuvkbv715QefRqLLUYrh8Kp
+O80ylPXOJMO23TzUUcz2sTkhtTQceMndJrXrbMlOl7/0ZcInQXD0xAoBP3Qb/46HfxVHzhbDL36
qUg1V4XvZtsnwMfXuokBdL7GPSf7hrSW6v1lU8xM/IbOYGGI5Z3am7KoOKXg/p/wAic3oXZSDWhY
NEwaDCV88wPuiFQYmuAEpEAva+u2YJ83lzJFmZyWZvoEWEjBREfXUMsc1ssPaA2Yvc0rkGDC1git
4xUcLjPFE1bqfM5IBR3uDOyrpbNdzQi2+9cmCUSw+9H4TIDiwhsHmXSZY5usIybaVqtNeE7dglk0
SOgjCATAfDqhsSPREMaGqRYbJ5xGX9JW+quEn0j8pCw1u8GCTcjvrPiDJbniSrRkIuUCrjmGXpF5
KT15VCG35ZnMcDBbsxTIJha1kzurEHJdLC9jUHozau+8EStPPrjGr8JH5VpcWk1+UYtUNX3QiOo5
ntaYKnjJ1xftsE0+vCxNkS5kYh+vBHnjPcnuMLNMkP5tplSR0Lhrh0DworFs9ebsEdDLu7GzhmEM
B2+DQcMS5tHF64KA0XecKbdoSAbCOPPUXqYKOt93Cveh+sDtivG/LpOIl5rq3MwDYlpVvpFa405r
t1xS9/Um8RUAi7+jDv59T1ItXJmsrthisbv6wzKxj9MGOnKAvXWUKYxDgxAaZy1iry8H2msWCHVd
iMQaJy5JWRgnw/Y0mDUDeBdFG7t0pmGdxdtJ/q6+JKxRr8hy7+V2ECvktPslJOlYRQKvr2hSfCpO
oJlpjFmB2pea/kmLWz3NbLWo2IlciM4VahshODoFhoJIa1mtp3ecCsqNu+PoNrYPxcy1lG5vVCAf
5TFfuiEFmJEpvlT90oICOnB8/kyM/moeZaFM9mGYDep/5kms1zICOO+EjbXeGMnPUg2vldniUOj2
Bh4xgJjzjOpnqb9Nf43XAEtO6RCo7BnrSg+7wR7Nd1MSUkmZ9X1HbweE31mNeSDfwaylYV9Dwkub
XFarU0eW3ts9x8dOaX9Yp9tL/eQwrvLhQ2tVFbPu9tX2TeIwbqdItf7X/E88g57ZPOu/6q3Xzg13
UXViVtZTOk8FFne2dcUBhITImIADcEsOJFfxGOW4Al3jyX5ENG74Dk+qWOylgpRmd6N1suTgayf7
0m56fjFJcFQiqomU0xasOXXhKevfa1OGt2T/HrHcbbXv6IvAxOC0WTtxHpnL7rHgEfYGLIkeE9QB
3Px7EtcYHypFSDhDVCJcQfgTKKN4tdblJhzPoHYe42T2JsVTBO5ng5OfTrk1KITz0HueHZ1CGqZr
VBs693EpTXy15bFK0/8mxmR97IAw+ndlWDD8owyW58Co2GUi4eHoim2Xg+LBwEIsC7NMudlKMcgU
oV0T5RZ9ZaOnUnlBxbvU077GxL1dLTTDoGZj4S0oxBJJPjvBmLJOe6F9sLflZm+2oMEn9JEoXNqI
uv1EMEwevSN+zcgDvQFJp4x/6tzpC9hDZK69D12EVSXdb4mAYofa4qdz7wcFCWyIMO39FL+7wQft
+hrexMNnJTnwlUVE+zuQ2sehxanCqNXEYQ9wUWr/344y7HUtPV8H1BxtdCIRQGnwY/pmGC9h6Oue
xoVDEmprZNQEW8vE5zP6sWXo+iIVNX7lW5YfsjvkmoNUxIu9cgWJmGs8LNU/mi5WuJjOboj6hXul
ZiSrIX6h2mfS1quO/GnCWQju+31zl3Cr3FZij7UWt74C59GTOTEVNfyeL1+iYm7QrttuoARSSZoD
F6EN+fSTvfyhHOyjfFsb6PBkoz3cIS0Ixxbl2l5bDZwGFigDK5X9GXavnOYLL9EDHraY0ycoccs5
gfak0HgN5BxE7Bjdq8nw1ZinqCDjyO9SmG0LYWTChsjFzKMl4Pfgqdl3L1+JhqkCwIDwyKuvHtmI
5VqiQQrV2W6VTWW/wezM/fiDqI+2MWrFofNYO4kVmFcx/TKjmT7XU8+i5xYn32TZxVFnXykRHIkx
cmhfPRDatmFSoObHmYOYZFKDx0l9mab3EKR9qRbgalts/IEZ+Jyi5/tXCxkrD3pitegdcsbP8DT4
/s+5I8Z2UaVigdF1LfG7JcU8TXB1GgXNj/IUTc+9tUKuvThEWmBAeeEv9ZMPpvLgfG/aDU3oIU0Y
n3rAFbAKiNE2DlWa13fOq1/0s+55ev4VshCFpsDHZNPgnUh5owA2fLS99vsLiF0A3v+qUCjx11Y/
5dxsf5l89sem2sWaGZslx5ZJZIF/CLB03dlKiuehSCz9P9Zkf3LP1esx+FRbpcSi7n8PCoMpSfS/
BE7UQBJfGHkoS6XQQ7Xgf4P7ZI+IQ4Ift0kODof7c/IQXwKuEH+qDIz2656els01D4JoU2i9uV4z
Uq89Jg3AgjFW9Zh8Mz8Ocyk0JlLUrfsDCA0WqGFAjMGE9QPEcIa4xVsidLe3PLm/lVtARHb9IZZS
adxSwxyl77qkg1jBs6zPdRM4ZxH+NeZTFUaPrz4vL+nWAk79mdgcAgvqzdSQXDtnonOBBDGwvoC3
df3WJmrilGe4NHJuPGZNvPsilLSQrWhnwpvtQ3zBtFD7Jwoc3Bg7wUUyPr18y7TX9kG78RFjWBWX
A1F7DCLD4y7803KgSfAJxcuSCbDDMpOHkdTWyN8p9S7W+atnI1EDYrGwmxoDINhSg0+ktCwkXmXZ
XnprLwcw51SeBrda17SVMU7ZM3rgo3AnM/KyPXW1iDvx3bfo7zm6Qq5A74oQP98Zez3WHFS6ynIm
HqLZJgk8jclWLZBhrdNmekgVr99dEHz81QvFdDsVWSjYwPX2KHofkiq9ddT/h5O+vp4gi62Ga3Pu
iS0imwQnZPh53D9xEffK7cBnniZp9JYiZ79ZfaBJF8//QufiLVsAvf4Kqeh/IWOkWhb77oKyehMS
8B10OZ0jJeQCQZaL/Kelzg9zfD6ZU4v9FGI24Do8yWkjdjC3tFqOOJ1RgZ051VjoS64o+UtGF8qp
yuLuxMivUnF4/OA22almfgSWvwx3uCQeOR9fRFUJaLR+/IWD+0I5N2AqWCx7PHzxgtWUpGCtJE7v
cu4BpOrrqcHGE/R56gq1qT3t28Lw0dzeAKp7gNOGivC+ZXOlo2IBn1I/8gFUDMvcIHRyKY3fElIF
UWg9ulKrDzZkUPfMRvVH1m13niZsBcsSg6Q6iACbtNkhbMWJclrK3gcbiv/SLNmEnOVYWkAfquGP
OBQagrZpWi0Rgjo1blMwljlhianOoIepUy1az2ZeQcEENFFyRQME6hhTtLRnsdihBIWS5tHNoEks
3nMWQ++DL9mV/2+OOthh52eqPt2sAcVIu6uhQN14yE9eezq10wYgicgcjH1rsQzGC4WMqmBPAOSC
jZiYs8PFMcGyS5Fp3N+DVmUlL8ExuS/UU+dLi+otrq+slk42eKI6wOS5po8itm0/4Iilm593Gf8b
ERmktlyq0dsLhnSFNRojBxLj1Of2e01zrEH67Wx8+h6D/cyV4KA5pq/ca1/GSpCTPc4PCsTmd9v6
ARPFYWpzIIWwESZksEHDPOoTuRW6lwLpCtQ7w2Cz5Ss7ij7iMIB1uENEQxklpT43ftCqL7E6sD7g
Dr77URp6ifR7YUj5T6YgL4SZnwtxoNKhZveA6XFn70qQpyaBOKswlI/P2kwPqXtAcPl3QYqkqT1D
q2rNPHuquT0FMR2uGoG/nmiETAln8BweqIXKfKK/YCSiV0ShcpAp+/0Sxd0bZkftYExKQwR/O47O
A4WH0GtBxthQXERfJVCt10gyNuCEdFdIiPVgFEQbX6otcgj7PET5PiGBpPTIn0Z7O5Z6x4GhRKl6
oXzEOBKTE58tVl/B//MJn5OYjp45vKB2Wk9+THjXK4ZbAqlptqm+qk/3c/lFbqdqn2QpXySPRAoJ
n9whxEufTDPY6Ef7MDoqsR5B7q0q7MYyOwLPO5wQqOUccVe6vVZzlhvhap+D/nZDSXEU/aLdo0Zn
Y8wIkNCYggJCPS6v7AqhQQvt55TrtP9+F+to/M70/KH3f15tJDzkCePORwDf1El6tucPqeEebaVi
Mc/2SFzpSGhhfj7B4kI/eLHellPpRjhfu3s0DtAlk83DaUbJsAEZOSg3ThIhRYyEP789Splpo3Gg
FhhJFdlBkMEheDvYZGo2iEvJMonpuiCrct0/vEe5qGqwNv4Ba8uldWOdvuLhBfuJHy0RDbEel7Px
JcO4w0PPnrnBuxivcZHQwLWmC6ReeVXW3KgFnldaGUAWWqyvkpDc6JeSiDpAYiNlL8b23JbIc9v/
a3V0gkrnMTMLwAihSC5PBtvrfsdTnv4V93l4rV569H5qotzOtibvrtABSlJGqn4MZleUbT8u92Yr
aQiC//zuXMzCY5fADpP7lefC7N+jtwWR20MCU2eeTbgmulVed4hl6U70bJZ6JwMrdGAzlUtoiwkB
MugTdrAllXqKb6Ppohnifsl5iD7LoK4A8DHKTO3JIb8pjF26CVQGudS8U5gp7tykdz31qn7yvb0h
AMYoqG57TJhvYcyVBCtcQCNuykILGJRq35OsQrHN4Jiq7DpZ+8S3KcmyE3kTZLQ9tWplr4Ktqt4N
Wy9Be/C7syGfp6CfZ4rTNGGpBqCuqYjcZBvaUpuTmPLKRBbKCHsTvSiK1CpKYH2Wxrt0Sr/Isew3
u+zuNXu9LFKtRuI47fvHdnxwjzxgLxxdzIXDdz4YEOhK2tgGF2SRkshOLbk4gM1aC9/5Yp7knots
u1hedc5X2iWlTS0xZv3ypZl4ijaeM/RFTTcc3XPdJI8sx4+mH3QaIR1SrPC9ErWG1aDt8/iiMGkA
HuvrohJkQrwM5Arn0zBY4SGhorg/xghI754E/psYqFIbE/etvEKy8Vy/3+wHUgmAQd6pPVH5i92j
P1/me4fE44H1RVXvw+ii0dtQ4xOwITbEhkBog7MkhZ6wy54T8eLLDGJ5IuIxVeucAVWdKzq62Tgx
usXsz5IKt6wawG0+eAUrTZKhmt28vMBVWVmsjULZwFlkUoLHNvi2RV3U5agXx8/7FiYdDUalovNm
Srb//mb8ywXsEk15DxPfRVPjjIVK3u6wjLhlAh7I3Q6RtJIcUFtNFosoD4wwp+SxHmstvhJ1URQW
hbDD5QOE8G/hngyRsSeBDxiAlefrAZkfHaLC3m8hhIyecb/L1p4HAr2Rq4TWiiINFOMdOXh1Qdso
xdTezbTrn3ST0ktTupKKzE9ZHEZQd5tkkDMqaP6Z5NIXthqxz+09KTxz7yVOlwOTFiHK089/yacr
0cryn+AVBNhRcpypD8c09s8HHHBgHnOnMzUgrevlxCoTT0xQPAn+O931VQGDCEdbL1jOLvVwig5L
BHC3kvIK6gas2NhjS9bA9temgdX35hhEjB2jdk29lW/qPCGFyzovEytHVJ7i2bNS/LGJA7vd3C9h
BLRkerWRAirbcj8SVRaK+F1Tb92s24mYUqo1+s6d99FJNQqOr4sZ8r4QqqHEkODEFeebzGSZWYqG
ahlFb++3ton41VRYp1/Kmr+zDErBLpSsnz5k/opLUbd1qzTScTHE1Y2DS81cYSlSe8Bcg1UcEO0e
rLq0rTxfM/Vw5WYNc65A1cq0kU9yO+JwVBAvMu3PFwF7viXH9VXcQfqvjZZIeYCq59fGdcLyMlHm
01Dm3gAeJVCCyyGtrSAf96e58pUEsIGN8egBIc4AOgJsGHyRUg1nOl/cuGNZ92Lrc83+xuQGlbQi
AarNjkhvGNE6Z/ssN1jp+Y6no2/ouw376tjrJ7M7S++EIaKoLdrsJ5gD64048tycruJVfawDeS78
ac9dvmoPsW3Z1HOOPJd8Pl3ikulIFf2tPJs9ZRpC+mi5BSKe+tWNLncraTYcep0O8VoBbl0jFgQ6
GIBlbgUnBQQ7H5jprnKKK0dK5N5gqMZWavcNrY3q08F82zPx2VX5WDz1zWoN28M5l6t/jCxxX716
KrxdYD9DIqlC7cvPmsAUCfD4jtzGu/YCZW8U6U93BmcKLld3+Ew1SJCmlQOxde/t+RKowCP7TuLm
ao5mM3AwUcNI0O2aN/HAM2TNf3QcBIw1272uzPSpIyTEvjiY5VKzhKuj+t/vi79fMaLZHWge9yPe
qwFCRdkJy3vVgMobIHAYUy/xiC9DXxNIT2zPkrmw54IEw/YXzx0+N6J+EzeLI/nxHlid/I5Ico4Q
q3RaLC7+oufmyp8dTd0bLhznW0rBtg/fekWiBV2l/rnI5HwBROHWX5n2eYBdoPEAYZWArWaHt7K+
lInBPYb7bMWz69ML9WKb/KpttR6WQCPdZo3b6N3NoWbFAjjlJQSVk6zx6qhYyqncx3BhXBdetZIn
5/c15Z6QYk6Yzk1Cn2/OtC0kvPP03WHs8OTl+kOnw1OxeIBGuY7SIpZg+2syP6U/fTbqyVi1sw9q
zZHlx1jYgOdMjcT/J7XErkNoX2o1bIp36ja1mMV0RWAoDeD66oVP/Xt5ju4liapT/sOf8aBzRqOP
VCgZylm3Haq/LoO53Ol8VtdjVZ2sUd+UL7v8qE+o3jes8OJvBDYWNZiaJEBFO8eCGrLU8mslEbSy
nOWtVBMIovXUHQP6pmu/D6p3gpQlHzzxZ8lFeCzzBrGQ35UTmyxlGo5eU336ehmLCMN+P8fhkaX+
RHSSFy6XRbBwhftTyJ2p8Wceo8Wne7x64nS1HygpwG3oYZYj7eFhnb7LetFC4oiTGbjIgJTR3Twe
/LbXJkPxzzcYOnYrIHcWsvFOkTRg7ibL7OyWc/R75z/jNv0+Yk1dD/Wp4Patd/wA+/gXJ2c1qHfO
zOlFtEEhrPlxbSTz5pzgl/PzsU0E9QjoXu3+4q+Af/SEHK4izpW0YSJWJkw2QieICUb8cWF0DFKT
wy2XHjf4+CvW9swSBdGwXn6OICSfhIRXzK5V3yO6YmW91hwkqzpMn37rtGcFDeN/5erEZ6mADSKo
tN6oJ/Gdy2UaJsatkc6Q0g5Ci5TJbnBl7GsdstQFKlCjhfZ3ST/zNo6xDT8A4x+CCpAQQ0FddzkM
EId0MsVgjS15cg4i2rOz+AtfOuuD6LzPuvhpPi2kfX84inbJXtd8GyO5jmZMewONvXs2w+YgbFQc
inehUfvis4LXE2/i+qYfjV4HWLHIycS3OWPtcCoBaDUkfz8VUCSR9eOqU0WkzctvEzelzSrXAXPn
KJOrAD2h1AoRdkOCDvk836frRfv9gPH5GdvJMAuaGg1o48vsPEeHW5g/4+CbuRFnuznEH5JhBinf
1ic5zj3XYhN4uHNZTA+diO7plgOqTGqThxBWi59fb7Rp1yEcpdDOAxZEWnrJaOtvR1N9VYBfXJHe
j46NulZJgcXbVHbbcAvR/QjdBh4oy3Mp4cfCMgEhwv5sMinbyo1YeUci3a/HRIk3IuI8S7ShjXkX
E53SNp/zwcqsSiSAjVu7DFXq+VZCDlSRHwh6TLBPQrNM+gJsIQKf5+17zev9kuvKa0U6QIX35kJ9
/nuUr26Jnc0vDL+RdtkepBiK86w8qv7ZuqmA5UC481TY1aqnoa91Q5y9k4b9q7wyTht/yYt6+h/P
8UlNkenXKgg2IYwGiOJdLjwdd5UVj8EPDd+Z+WakV/fL41ez2DHtfjYKeTqVHgbVbELKOjj+lwqc
C7Kd30jm3E9UUwZ/Lq6KiESVSC7ACjhbWKoZyPFcu4nYwajXRNsK8+nLrUuJdAXJa8uvfhA+/XS2
HoYayH42Q7lzHw6zp6DpgoQ/Kzfw+BVLoGYeSG8JB+o4kMisT1DxD/BcqXjUr16c+LK5iItqvj6u
rBpEcsVLhB7cfrzz2Mk/b8UDJoH/FSFP8Fi8fFQkkLcZedbE2yAD0mbOndRRPo7X548z2zlvRDeJ
L5JuWgWQrrYVbjNJ+noDBP/QxIaBLHfecGPd2YXj/ozz8p88U94PKMSpvb7r0cdbwMbaYDYjaGLr
jOVYUApqSMD9+fHRtCjOEe1LYXpWfUcOOLiIYUwZlgWjUy4zLNzy8IneBXiuyh3iNAmSP2UTR17m
l+8+mtQBzda7u3g5kRLekOfSgZCXg9UQGsYvcCwlQT3+k7qkIZvObFP3bN+hocWW7j619/8U6ZWs
LNoobJMJpjA5zHXO3D7oCoBZxJCAJR5j/18vjiORxNbnq8VZXj1ZYO1d0GD0zTaDIZ9qS6X+dzhF
T31a8VdV9IzFCbolbORgf/kYAfLKBCq5AcR8kswRchm5EZHlgQJx44F1/VgoarpmQEbcAUvIf8oo
8GqhFJsmigbNMWzlmrEmqTQ+GZnBhNY/X+ojUwYvXx23HPsduMDmZZzxe0AcaF4hzW5H9fnKNN+Z
W82Qs9R7+/RiLmgg0Jrtj16+efmxS+xNodxAxVdj/RPwygyh+pGMiWbTfLhddrj0rBcsuNwdcHQi
oE9SfWWr2vziW6RTCxO2aOtK4cXPwTMLc0bUtoDx6/oKQBL/TCG1+KQbuylRSewQ6cfXeZ7Qj/PM
dbqI2AHKLhTovnhnloYGmRRwYHIP7PDlY0l1XJ9gZpFFGl6dNaVkJ3lne0w3NQjogYMEqGPDn9uy
xBCUorS6FgfCWdkJMxX25Gt8R3k17e1vUU4qAoBjEtmWhZtXeK6s2ClKkUS/34Dd+0ldpPimWo6r
mlb4Jvs0X6XnCIjqeMf4sOvsl59f/8bxeOw1jOKZIX7rCzbyWX+n8C6uew566NoJXoEzuJwUrOmK
iT7t4SfzeTJ2RUp8tvL45Fh3WGJgpusTr4nAuUI1fnJJjguAwxy4nK/t9YDUlcPt7byRUurXzSFz
vvM+0hIqHJnpuzbcfwKl+IDfG6ZpClEpMRsm4rTgOQc3Bz0ruiSTqzo7UOguqHS+lRrS+Nhst0yj
oEVwyQB882aIsn7NdEAYh7ODUX6r0ACB4Bn/TfjEtOZK1wgH8jrCmsJYkKrVd+Q1DqzJRhhU1TRI
TVEnTDO6WHnLW0+lZ1D3+6ZTWFvRdTnlveletzh4CfEp10wt8ogB8hwI1a0aZX0xG7cxMAvPWJfP
Y+vn8QGIdsNvEJblsKhY8Hy/H6ep/FkIJTiNRgpdHWGqJTRhApoPN8DVkwgPlcDuGsPRSjktY8g3
YN2iiB5Gp5pNNMcmuemMbDZZs6AH9P5BI6l5unagRZ3mNPso52h4x83/jvdvDlDgDtm/pUhtVC1s
Sa4NY9lNU/5ZJtdO9nq5od0LxNKp5TqiQwL2NjdlM6DxpJUUO01WBSDfSgLEg7jD+jDS0RrQWs78
UVdNO2kCqiqoUdU1+pmr5dBGAW78WiuyPPF2X3VA9ekz/VGib5rstmsxjXYlDfHYwGYjDuS2Svs3
pj7H4cQsXLOMKrq7oY6DiwA0IluR692xZt4C+aopTOZIuA4USagUriENsi+G0wCbFBW0/t06DLqx
9/1pvy5TcrdFazHwIaDtED3RxWSL8JGsp3OcJghI208PiddoNF8mRrAiT66+Q4gnBR1chdljBgNo
Yf6DpdzdKjNEIsW4VjVFUqXRKw1DdXbpwlj7UAGRGGIkh49Ypog+Lxpe7scuRcCWOKd+X3j8V73d
TW4qwfLjCWEM1zavI/pVpjU6UTbuOSPBouT9dTLrB90dR/LyJFKVrNtXsaCHsixZffGdNK8t0N8l
oYi2bP4cC1XUqhT9NNBbsc0i4nICUEte5C9tdyWxJn/idpMPsbMPwqxLmy9OmOBhOqxRfuk3aiIG
6XO/Bif28neW0gaL44kl3UFIkSf3vy85xSDz4BrcemDG600C1VbhRyYprI4wv+8SHcaZhyndAzfw
CuVEZRxltn4+rgv76SEdifXDhrpMRgeNQ/GWdwXadfUooUerqK6MlEvDABPvBacmlj/0jluJp+CO
q5uXQefslV4qwI/TbQ/IK0cLb5ccJVlIBM2VqpIj6+KLOc6nV0xfEGLrFNoID3qapUKOxE9/EgVr
KOF77ZXek3t+pLtU6tkstK8M6RtfPXRUdtAhC3mHRm6Z8b2g8RpZwKqXNcOCbqMK+6lxkki22WS9
pLIfRaSN0zcDZlaXSCFoIIZf72t7DS7YEtg5g9RJHNVMkJp0mJzbabI0X28FX7224GggsV8jjnSb
KGhfPhvOwB+EHUuxC3Fb7MZTl639aTfQgSTPtuPRKa20AXf0JFsRXDXoB3/o1+vkV67NF5pIW07j
YHsgKKtWsMlLa8mvhonu+juT/l/FDg8XUZz7uAcVf2oq7iYXrBLXtNimlsuDPxfKP/arfsIadEZu
PA++WnePcGgmyqlTmgFUmIdRCBLuO3vsH5a6QLUBo9GqWDoYK5vjpBfql0YLV/o92clYGyGU3cGV
xvxJYVTfM9uuLok5CNvjsZKA4jR7sZIHDnA+PmSuDjOlg3FmXRx1wYEGm+uiMd2BDmvAZuwYHkWM
ig7+oE6wTQPu7fGVnRS3WrTkebV3jw38/EpbPxShAIXUGEKTzQPtHTIBbAPfmyrRxp2/k0TLI2I4
MMhGClYvb7ssirt+FOZy5iBtjyy0nUrpiNQekuZbR7cAXq0CBPnJ4OC/s9QVjz1d7vyOzTmQMk6X
LRYd/UZERCrOH5cDXEIat/q+7KuT2Z1ijAYcvIvo+xsUyXXAw3AYA7Ss1nJcTl+/rSYsOPvxA61p
LEu3pAVdHjqUiVDgfIGIPPExgzB7IIJZ7mQFwTTF/k4O/K/kKC87KCqbI9NnIHo8n0ECRItI752g
nKMPOqThUI1ciIPKN5j2iAAtbFDvDtbDM/wx+K3zwxn6Yxgd9maQ+cqju/WXmiAvNjnDHSJ2uml9
ik+65pzbw+qpRmpJI94Wh4lYeH9+qp/vt66mKsB1rkkou2MFl7N88TxI6i4IAtYFwOEB3y+RQ7wM
ZxkbUcSy5hlQB7P7NZDbb9ecpzmZIvbLqMlgMIfvEUpQQEp9+N3d6Rpbls/cNfHqIpuUsJs7tqbT
gpcGD8ajBtMtQVFMBPc/QLOQXg7pEczpV+T7KbLZUDacIbyIAVM1XSeSgOnZjOe/YHkrWENi6nmD
9Y7wwEYbeTpIDYUjxps6NdTz4T1XC7oELCPDrKcUc7AvzKG+8bpWGH2ibrj4QTDkmbmkuiaOmFKe
Oj/LP7cWwcdN/mM7ZG4nU6kWFu1AYw6dPgaiEJll7IXuXPNIMI+egAKE0i1Lae2qkn2it0te7eIS
oudMOhTWWfwjjTNGpQJLocfCVGebaiBHLXUnxeF1IqZgFpaBsZHn3tlPk/frSUtNgdHISPwFX/Y5
g7FxTTuFcv24Jbx0xGAmFIrFZVMBoQy3hVYxoHLLX5dKulNvUG1UnvIvnEfYflQy+ikAMU23D0T9
Z0u6hPbSw8WXZsCOOXiNX26aKxl9r0rMkqv+Z2pKyF3h8XuXV0XKEYwU6bp7qmU9aw+K927ZAM/z
8WljATaiBTfTxKlcznsA6lZBjHEYFuAzgmCtm9NgQ620bZ1B2BbvSnmjjOn08CSBqN4mykPScaEk
8IdfXQ5wDIw67eVk8Li6SrbmL/fR3wTF+VwI55kx+oN5fLPtk+3q2I9ZKnPlHOuKfAdz+y7djFBO
xDVqOMHUFCV8u0yf6oulmTH0sKw3MGKSVKpDkHuQ+4o7xJ5G2mmI4ne1me3Gd1zgZbed9m3kVIQl
NnPUjpyCawLVNz2ZGOkumQvVL8F9cIYCQurxB7vFqBlnSVXlDiFbWta2edZ2v6mrbbX3rI9c5AaR
VneT064bF7BJgYzx6tIPlUwWEBoS6l14qfRMJAEni5cBOyUVg2La3BxksEj+Wus85HWNCAFnoDJ/
Xk9XV7XoRN8kgM7BRZL2ZjmuPgg3kXpt+2o13POwrV3CzzDMMPPquKx6kTT1QruNiuyixqAHhY11
yOIeE6iSK9WM78rRcYziiW8ejmMzpcTGmDz78roygLT2PdEuQQ6MCBqVvbzfGFIQpLnHXv3Y5/mT
6trPZhznrSgikRSyx8a1hat2ON4S0PI88SJDdqWSUrbTzRWvHWxCslDhe+T9huS7aQ+G5lfctRt5
Xd8n6p+dHmcHwMrGSteGE/G8dEkDk7oJbE+bm2gdV0kK1lhqhjH9uug4Y0wBbhvxYpDMd88sP7ch
iD4jULcCoSg8vgDv97xS+hi0SSADIjPVj1y1SsnRQ3ZeSp7yu6tzW/7eBCrgHbwPDeEWTwB/xcBA
U+t9VSVN4Hi0uR8qgUij8ICM/rUESpJYRRyhdwHwYcm3mxJeUzcHRgXoCmnxrx5SQHz31OgaZdSx
KuLu9f9nkYB7kWfB+sBVsQxGa8nn1KlwfjcJpzGgU+AQNVIUIFvNvR+FbhvtxafgdNrkbFXJLoCI
JP7N637d/rr6wSPUs0MNa4vLDV3Lsp4NjXCQMG/uN1LlG95tphWyAG80F5w3JdsNWVu1sWGdq/ot
Dh04j3tqXAwgrLalhCSsUuIoYY0ZtzLLGY5Vx0Dr7wuVGlFjblchj2oEDV18w0PMzv+ZX+Artaiz
0p9MpQUo6b9fW/yfxXI9/T6rY3ZWQ4y1B6qdvdacPdURYpZw2AmrZlfD467btrHq9SxAxTrEIjQw
BSrMke6rQxbdhytrI8sSTnYg5g8uPz9aMDT9NJ3Ga7K51APZYwdDrvm39lOVfp7elUYnB12hUZG7
jRFEEiDHuVQ9a1NA2gcbPj6CvJ9bXQWjvXQ2bPSQEND/akU2qUxY40EeHCtEeHPTGwNBGLrrURm6
y7qLNZyhcJMvcPljbyEY7O5q/tjVh2lJZ7/DpgXBiMKod5DFkcOY7vHdd8t1opaCLel00IkkpH0N
iDj3YD+HDMVIV01BT2ucDZaZKtW4x79sbrrvrPKH478tj/6kS9QctXTQnQAUOFIG4wQkzMEId+2T
OuPLStUUCw6cOd+18dbp/u7Vm7/bK9BbBaJk6pyZ3R0u3aFPTxp15/TExsKqUSFozhNHBsb/tmYZ
jIVGxzhUx6nRJ/WdCx0n7gtV+iIh/SyYBKiXWehWJPNtWnGHt9iBiMLRKECtGDMcWuLCT5QsWebx
SE2FqU8zxM8pKoVHEhjcNVE12TExBk+w8QNhdCpFBk9l73SwrKXv6R1+TPWygjBI5Mt81ULwDjJL
ig9Ju/F8Gl5lXTSth7v0oXq9K3NHOzSsvARyWcOnmpdEH0Lzrh1f9ThR7InZp4mKpz0vfNeGhMPY
ihGMEFeKptTD2mn8zKscBtRPuk8Ts37XIDh88TrhK+DgDUsm/WWCTLxl8iRIAykbE71IfKLW+aYx
3sLeBAU/rstQ2kn8qbotPkE6iX6dUjEfYVsMjXyixpl6Sig70JU6XSf+ooJYK9p4VNeemzMfGnGS
GJEZYv4V3J6JZTGlFA2e66O+t+/6It3gw6jqqTu/I2V5dgBW+AonYFsuBLIYWVC+USuTWUgSzgOk
E5wbkkZVZhPw1f+d2U6ihJfEfPE4LT6+W30NL0ZlGs2shS35dUfvv06XVuwxs85oPpDrlsII2QEe
Nb8LiqPbLL6riIr/jcfn6OOE45Y1QkUNTl/fRV5CVzJRdIrV0WTeVzBdJeR1GFG+6umi/HWHsca+
q01N08KL9XYdP1MOSWA+LFk51x3GSsYRj7iM4hM3lJ7sZvsk192rGTjJxKZYLsRzLFgMuOulGrtW
k5qn1ZsUiwSouFXPRB2MV/v6UxA+6ZfC6LAq8jaNaaJ+yDkCLpu4WKcoH6bkrQ478GXUk9ZW+n91
QXS1ZUWG/UBaL7NvAVG4xIW4EOiM04SrjW7WNubnUdPX3wcKNfeeme2C22Agpyy6Ypk3xbamcQ3x
lzCn38Tc1jEkXv9lZXqWDP4pPhxY61rb4PlTaHFuAVYfrCiI3NaLMJ9HelIPLiDQfF54xwGUmaPc
/0blPFkTqYKW+4J3NdfcgD20OP58qmWtWh9xuyTNG2fVS8AcM7f4nzu4vnwSFdUNl0TMMSpkUTDr
LBgrlU4yhvAbatzU07MaGV0slGwfhi/YNg1MizF/DLkYBICHWgC7DbtbT0/7XmR/pdvTCvmRhtsT
Gta11YJbsJuf7RVofTRney0NpMrOcbN08u4+AhezV/7OB5KJIOkDlB1sb3V/dKTCragSM3DMyMZG
oN52STuTsWCxApGhASe/BkUmzRY8rU+P+DE/spKfs6GNVfB0jVbd5YjcV+eawfFN55pE6bNpdzgN
fj1Cb5ZQvvqnN2jtqHv9wEOR03fibi4E6G+YQhesco5XeZBGGCde2+PzIxENQ64TO95JVN8t/+c4
TFUbDo8GC2vVJOYEYhB9HiuqktChxTBNUfpyu8YEBUZhNrPxa1WZlfnPmvAVt20bCvdWEAPF5Ihu
Rjz0DOCup98JmVGfgEuMKJnuZ2hczDBcCbFz9KNFvpJTyakRVX8SuQSKYzO4ehvGtpcs0D6u7x/8
RjdjU6BAhAhZ9pn9e5+k+l3FAq1VyHVazVa3lcoW/Ks3pHURX9R6mh3/n9+8AUr5OrjXRvPvdG9Y
9zTkQW5P6+9GCcl7vCRombqOoHOYJHsHTNzXjF59IvGHS1DiM6vRSofJJlgyO/Bd8sn2/LoRMUkS
vuFtFZy6wWgCzlgHCNHhT4U9PRGv/KBVrEuWfLkbvZzB1B5kN8u/DQkXTU0R713GnQhayY6BvLYK
ubHxZZ3mOLBAf88GMNrtszTAl5jCvcsCFhfCRWOB0Gz9nHHsuYRWEDCY993mbtJMbW53mbhBqeq8
FPKlVcJbaJk3H1zx4lXm2sm/TIhyn2nolU+4Pm8Mh5BXyx/Iw3DfAES3M+pQosQZj049Nny55pPc
EKM+4mW2wMVxy1iLZBm1BT6t5Y+Ohu88uCJtKx+kfcsl4pVvGjBbunP2JI80GgFEpBCgQoS90JXv
KHXfdaHeldvvUqn9hTb4OkDMDZHPZS/0fkE+l0sE2H9TIw8zP9jJ4XV/Wal0CbUz0GNEoGAFiv7N
sap2V/DUhy+lk4oBW7CxeRBdUDFPQQ2n0hIts/YWDCu0ya2eq936ztlrkJzC9+n84Xt5ns6q/bXK
UN894A5SYSVfW1gk5BPMbeFDNAtiv7i32qIxGzsdI7Hmm5g4vXkbN5rnAgBryrKzlBLuOs//6AnU
s3y8s13q31WA176mnyivaQ554fxVrchw10jllhXx3uzVHz2PWIo9xE5MphAn7mJdKIFrCXGZJ4Ap
5Qtzy2/Te4M95GCZ4ZcFqgcTh0U2JGCFxDUP02I3bcwhCm2L/0UGINKI79e1ltQjoGA87NBxr0by
5L+0yLZlJzCFqKmJW8K9rS9SbwJeKGgINQt5Ivc8DAjstmra4hxOysbpmR7by4dsF258b/ZhEu+3
mUEOsh28cJxrle6u05UgiZ28fMCFRnAYnBNnj0OSIdTXIfp6JYCl70V47y964F0VYxUvhjPgNDtk
OVKi7VuGO/G43haA9qeV6sdswYOJNe3MK046AbHUQqnG6hHRys07TRycojPljDnC6CHS7zSv0PWb
6uUKqKgYzEsA+q0daoJlUKcZwder5N4pzMSb/YnPDcbOCo/jLwXA6GT+eL5S1XYOAGkXznPtq8/h
TF349yoxDjrJ3t4XDVpRxzgZhWwdoMrPf2vQgn4CQawMGOkdDKwnn43VLPj2OyPU6cnPgChK05Dm
wzGqzbq1V8wCpxrr+ajQDeFJI1Rd8g/ILCN/ILOE7oU55Y0nhCnZA1ajdURxhHOuQ2QWC5ncYnnm
Fd2qzaFILrhri190Gu16nShH202GTV4tDvpTGuU8umIt5YH3KCs1pMrb7eTdTQHt/O40vIjcLJg8
U2ED9QhpwNsNaOpdGRSqdB26lcCOiK0mpksErrsFZC44KLtaoS5nD/DI6TOvqE3JaSVYSjXXFDAM
7K27cohmwDKMCF0lf+pgseCq7wTw+/XmqubVEF8UILBx+ReT8rTUjG/3rhye95xw1+frKjWAybdB
AdINF72eFh0hyrD+5Ih4CNv9fM30wYLrKuf1AeTp4d9S/nnxLEF0RVf+JZphsvuYgH5CfmgsAhUh
0/2wPMBL7rzcSfy3wmGMRnJLxYxJwQWCS1qnw/pUq75to8lnaxuHeq5icDEJ+euH1gqF/rvSly3W
3wBSfpZPCDd85+9ewrfXEFWdffuMqTQbJ6USltE9f+hMQYBwHnRSzwPErCgwOurIH+SZryJGybQW
UB14KZIgQ8IMaBpgiWATl9QeQX4jhQI4qdo16yARhlUM3OITuwjAOjrv93vLLAYKfZClaIsjrAlT
h+zN2svHNNAUWdjDmcy7Whe2Jh/iIEsKOpoBRBTdSgcz7R7NGcIQZHF9Rb1elgFBHIcN/eNGqeOz
texoqWNShcybfnL+m6+rys9wVy4swqE5fYJpWcuunm7WalR/5fCSyOBd3zxNzo5lJXN+Eeoi4Vue
cfahcRyMZinItQaGu5cwj6iWtzLqEP1ZlwJljsz78bd8BwtTpdYJlXl4Wg4kZ6Kp2o6vuiZIvlAG
IS9Ln9NlUNCYGp6ki3baoryNHNMrUqbsjfbRwAqRoYupuvMjaxFSqMEkF3+lcBS+IgCzHSjElSnG
rfuVJe/rz6A7m3jiEHBcq98Qsm/7XJYW7Iwkij7EspCIATlPwQHHfnJCdqTtkDXWBYfsf9od5HcK
gdUuJIW1PqGdqw6zGLhVYbcOK8imL7F475HLO0nx6AvDk93TqTW3xXeJG+UcFTwPszAD/aQH5iVx
rknHDy8/uPIbTeQW8bVy98+VJZ282zU8VFeLMUYfigPl8GTzAe0faXBA9CJktWKyjP5ixF9DaZBz
qPZled/7AIW0JGQZF3jKNqKIt/F9Ml9Z3QiWtYvKXzFvpOOPfzAFw8jVv4D18y5kLRrhmrbcgMsy
8Q2uieP1DN2lRC/IWNiJaT8hqJvIdV6iJlThg8pLaG1/m+Fvqun9Gh/CD9pI1R9kq5tcV77UNvJL
+/78QVFA55etqGYpXNg8nRp8ZCeJH+R+oIIbCmgyTF/20WBB4ej0E4MQzpqWk2gFe46gWzAA9TeZ
n52h65F9mg+a9ERvPhl5iusK2kqKxb2G46u/F+vP46+LaJP7o59ho4VlBNOyDTjki/EBm2xbOciq
Lisomk3J4uumOQuIU0qQAVgrh4zBy5VasJ035q3GUbRmhxHna1uu2N/kPxoY6qYDOmSSnt3eiXQ5
rta3PM1ez0P5y1Ekzm/teBTgI6Z2r8xNHQT0HOx1PRTMAK8KdUm2w7b3/5SfHOQV0iVKTUBvU9Nk
m6TTKoDRntNKsRDvRIYHWTPZPeF87epRBdXm3XoieP42PT7lLXG9kIOuoGFdVhq94HpToQXgexXC
Y0vZa4PUgafx7uG9bR6O4AM/LSuOApXA43bQkLG1gxkf9d4ZlKN93SDWp4KLLQrzE9EbKDYZR3nF
id2forEjWgXBx56GJkkFuCaOOeoEtisG3IxohMyysuyajmFRxXdkWzneiqOdmWFTufOafY2yQuYz
upwTOBcn7sRrezSqsLaRzyNnROugKEC3+nWP4CSrxUzxZLQwzwQyBoP2LJIIuqoMGlGMvu6QKzOd
qaSiCSi6lCKbrBHN+sey1ljE7ET1/RPOiAf3jFnBkSBKbJNmsE8IpUM5idX4R07k9MtcS/EaD2VZ
gbCyDr9qizyNkK1vnH/z81DQOEFSaZ76xBPD1pak3cAC21FJ0FHfZ/UIydZ0qYoP4hfOtWvygz6W
8zK0UPl+npbAnCWbpyyaT/j8/hTA1ThdbCfufQEsowA739Q4qysbCN3NL66gvsaA3JJ569rwNfAK
C+qmrky/iiOLADZ9mW1HVIna2dkCcIr8rtxazauvtUOjd53g9i6bkDUQ1a6cRI/83PyFGdcyR5my
8YO5zKswW+ZntMA3kWpnzM60ixamMtx4Wz4WXDD64HZVKm5HY0h1DTousubU2jOGIMWsqrAwOSqx
6pslk8woMabqMkQHzVmhYoiwfyOmM94wqkc0AXBz0AyMDgQbyEufeuwSbepxJhaOMGD3vedDryrn
wEdKSQHyprZ+NqP2y1RLE0AsQjoAmBcLW5RPyFN+KymK/n7+XMEmNyzxRtLmkrgr1q/gWoFz9/GH
7GDzSvEdt26de5KQbPHbbmx9wL5WgQFkngdvrvTgBfHLjFsEqp6L2HOzkMPk/brVC1Y9JPJTDn74
2gMHVvfcPuxgvfIUdQAOFXuqkSKX/EU1aS3pT/KDEcUjmhg/EwZvMvQhmhjFOTv+NNElKLo2t/dx
fVdeROY5u6ymSupCpD3kQjv0cMoiGoMfabrAovdjZdQYbOGm3lvocpzfI4GGDwAYw9zAkWT9vGj2
k+GoZimTcGX9pD/H7OhswfM2dph53cEFzayIO6R/RIJFl/I2mrIQQh+lZPYSzhI9f+d8kjyr4X0c
KfAoI9o2z15EWnZmH5i7fooPkIfFErDetx0xTW5SEoWdHgHU3mJLcdDwbqFZHgU78B6jAN93/qmL
wgvbRgRGtnn8CHMjJlaF6agyw+SwGaoIQpgGBeoBvCU0abyZwAvSxYKeh/g3GBMPBPDZsQ4491du
O/5TgaVKGq3RTKuJTVpk6Qns1BUOSR+iUgb1eHWC3RqgarTzgwhVnO22vYntWSIAvkaU8Ogv43+A
UkITNzOzJLKQgoJTttr/fYUrIbDebpsxdowvo4mH1wsUeHmTQ0TD0gMDaSULJ60e86fxeD4qraka
HlYk3zlydzJxivWPyjfF8rl+jz6F0p0YL0HD7KgpE+Wu0L8RrDxHBuqVIT8beca3ceHNRv0vVF87
siZNK3nWREDQo91UVHoGqcRlg4PD6kLnAgN6mEa/f0Tet4PuYRxuuM86/1tFQezf7nG4rgRvmgvq
JYuvk2RGqX/v6yeuqYznyz78xZCjnNpFRz6f3I6pAZQa4rtOErwC+wnl5fPTK4/Kl/seaSPEgvvz
p7RbPRrp9/jSf3x0npnQCHr1eo7ZL6bDIZD4efS6gCtyT8H5rJ6QHvSzDWqmEXoQCAT5Hn98sQuB
QCpOs81SvqCm1gucu+p6jBq+o405HiO9/vPkA1tnqUtD0noVEFtaCKnnFO961IhppJQLMuG6DVKg
54VxvpzahJimaSQYmkCNhnSsOSmR0jexkUG9ebu60ACDiB/GSx6jq04rbufakB5BpAdWfAgG6ZVC
zWbnO+cj5Nf2Ixp5ryXU1fcFaIlvkcXfLTiLR0uZTbpJpbq2w2YHFgF3fOhDyTVrIO9RDUo4NgPY
gYW3OgFWmFMyK5q7mPc3jmq55mXQT5yOLcX1IGdWJHDgA3X+n5pqN+OujFshpFbbP0DkIZb8gsnw
XGkNDx7WJfiw9akp3M0o5qVe1E6n3L1osaH71O+5FNOQ+hIzJSdDoAO23PEiRf3lYv5KUY+UMiVM
t0wIcqVuMl5b/+rXUQ9/EdGB8ZcuyPPOaTkz//spg51EnuAaHZAmJSCTGt7HNDeF03Fyz0dL6wvu
yURS1TX2b7FrPRVVp9MNBR76f0n0vxXxd3qwtzYPXbbBiXPYLlIINGQyL7YHt3sb/Vz6BPK6+AXB
ee7PHChctr9gUOpG/VhXImQS9PXo2hmmlqTCeOuBrxG0jBZVt0nCHuh6XusSGsY/z2hVjc7Y4oRt
mVfnj7iVZYcZUatgWoXOKOYV4frHpW6quh7Aa+v4x1WRYffrAnMA7zWyC5tGXUTUse/JMEFs5H46
6ZlftObl6zLjcxDXTkONC4J/3fzpoxtbl0FXy5Q8zCvzc7rhhvCjx3Pu/QzebHhvaGgCuNVmcWZ0
wuvmSkoo3aIz//6d6yDIeleidyebVa3b7b8WTmNCoBvCQWasONx09V1N7VN2bCw0Qf26RgOvL9UR
royhuwjygd6+Oyx/1ZgaTEWjCmFbE2qzqEoyPMzoJ+tFDMMtWTz85ipEWVhjqkcVB2Mlt8v3oCmz
1Jvw0H5hiVMOJNJjEGxBCwB2F6UdzZOlpvapQ0aB3x9syc+UPANtxW0ihv/jVsk2phDQ7Tj3+U0t
bCL8VYETAs2rf9RwD8Apwa03rv0vD/orBGrY0x7nVYKPOmdSU81Ybt3EbtP4FQn7+JI004EDXgbJ
5cu+1z8TosEf/WDSlyuKcnxd8o85cBC/630du9JgsWqubS2XdqtZc7GVKg7iMTY8p2TbtbxsGTO/
TmJ856lu8pjbmqVmUfYkhUE1L8F/IVqvdo0Q3OD0H+TexG7og7F3joX1J9wVXWCU07TNW/jlnwTI
7AcEtagrq3b9+C7LJi7UM1UmQEuuExot/jJ9XhXU8w/Zt7ziWpkD6foArnZUkPduJGOLrdzVTJCE
XpKgmm/jlcmbABIcCGl33tCcBXMFjsSA9T+Z2rY4ijh6HoxV72onfzwXL12kLy0yoeAhcHF58OcF
LOksSspe7oXGZOITCg02RGj8WaRwUx05hZRPzMXHdTFbi057Meq4Jfb3xBy7Uql8SwddR77vFP/k
x6V1++wzvGxRKj6lPNfeEK2ZItbTCaW2SE9G0dWrKM1g9oE9knudEykG2CbcprnIEg6wekzgb4uV
LvmkWnB+tAi7XOxl6PKiY4sEKVQUIMV5oZ83V3qaCQo3rYA2VgbfqflYasj2QtlQfBkOiZERSAjg
gfE4Ehl4GeOWQv+Gg3iRhSpTwzZDrnbd6qA+sXK2ZDJAOC6sqI08K7Tfvg7zi5U88iJSoONk+cOr
HrS6C7d3bbKweBpMP7ypWEMrumWvnj4bebmmjeQFx0wmgOMe4obFGgglXVfmM4YVGUcVFPeKy4ug
J653HhJmUN3AN+JI04wtc/hTG7gYrNvF6XiZQV2eXcdc+8W3a2ekkRHCpOf0Qtq3/qHz6tozHwqj
zcxMf5CDrkb7qLiEnPUa7ihAkjSqnfwI09f6PwDBFk/ZtV1Qw3No1/YTONsa89iGuyHVBeTlmw6v
Vi7kLPN2pn10P2JF8ZAGBG9l2Mlu4Opfiia80L7Es4cQD0E52HTbNEC87JB7KWHdrGygdo1Z/ao6
tCB72g41+sG0NNPcoJln3dOfsrLrXN/H73miri2Gnnj27EK5yiPCIly1lrYrtqV+s2L/mj2LrYcZ
XSIX3POPCixNGyYzKU5xQRPmUNvjHpUEJXp0dQ/2xcP1gK179VT2CDbMN5+bSsC3VLJnkyw6rbmY
wsCHxYgX5A8DVLLF96D/WVDm0f/CkA9SRCJ4+a+xLteZxW8boM1rfhVqxe3Nat9J5LnYuJVwJ8Qt
MuxFQh2b4rUg1rjT2giR+p/a/atcEPc+wzC468+qjwp8jJaTDwe26DUvYB1TngAiE/IuCLonCFKZ
BF89TXr7BrMHEGp+q2Hz5cc+CaWVSMYszULxzZhrsjmzaikLFVrfWUIXo7Ovh8MFQ+lRwIjIfL/P
1AId3mow7gkaPXYAhcg4Kjodhpasxy6t3lupyCmVkAuWpWvi+odhivguuVWFl1c4yKDrZUKm9dIT
ROSUfB5YZ8kBlJ205Ds66iwBJG2lH2N1JAyxl1dkBvGOM1lUprPn7R/OeO5XHWKsyXtP9MlXQelR
9I2wUktk1dgwVSpBWS1RXPJXll047ufK6sUxDl/jGG+ndbd/r2XmBZpe+nJLc3l48cuBMuUGuBJn
U7cIwQI+71/mS0nxO9NbZHdSJ5fB1zB2tRSglprTC0yECpGk6A9wyuxQHHrE1pr6C1saQOZNpQHZ
InGCbJOIYZh01lfdFJgtKg1ZWEssV20AxE9E49IcNPFqmiqp8okKrPoJhlpZyCuBpDQlvknU1twD
v02gR6uRe9yfS/5MSPP5GSe+TbpbzG5Z4t9VXb9ZsIQkcQVIfQW2LNybbaNWvnMJfnr7HPFtCDna
Gl7yD8mi2Wok7knU+bNyRWXAt8FRJR1IerrTGjuqOB5nmyTzmboF8CPvbP+I97ON7QSFW6SsO5FL
Qq9XZ45Fvk0F5KLPSBOj02kB9SBHaexy49mpzgylwp21KPmhJ6/RkCTwCwbjJsaGH3UCzxAzP4pG
cOVhywAw946uqyL5ntXz+OdK3XATPMpyQlNvyKkyI4hgMfbS45GmNB0Z9HFork5Y3uJ85oDQdE7F
4Z2C6jreEeh0KRkh/WyVODzejFk7sqXRrgS6KmqP19v4QANiApkx78KTq8QQc6LLfH9f05pvA8xa
t+f0Wipoq4hJLYIdCE/uzdUWFva8kXcedUQL3D/eC/DfuHnfqVBOnJZeAYo3M4X4N4/I+uHED3gv
B/9U+oXBlgl36pvWQ3uK6WdA42Ty4k+mryUskjRESZrb7ez2PbqHTRsBbni5o6yYoIlyNXG8ueZA
ONIruzFwWmj/sVwEEkt5F6+IkBT71B1rhDuGMI97duZoco5as1FvbQWu1V8i90ZCaTxuw7i2651L
/d44YV24gwOMvK4DAmhoqL0f96MrRR36xwvAW6F/6oLaRxf38zxIyZxF1CvjP5U7PknH/tMttSeF
iWYlD9E3MEBsG+7Ta9eC8lzvgDrjlPUlmkbulDZeRsK5wlK+Pn3V72RDfEXc0ZQGs/DtXS1HR3qv
sguysHrS1Yqsc8mn0ktMDAFMtt4ss+K9d9/yQRS3HlAs3rEmJdoUgFMAfEG4iBXiZjCte1FDbkyP
oisBKSf/B7zQNSNKcgFlL9NJHI/MgVZ4Wti8xniH7AlqyMAhf1Fy429Ev1XIJ4KWl6t+xrgtQAQO
z96PiUQh1X4T3jyuzytnHMz+RzWfVOZkL1dxhYl6MNEeMv+Zlq/6USBwn1Nu0IsWM2OhgGsGKKfj
KswmwdayK5bFFArBtJVDoDuPkRjt9Ny3IbeHz0gUgeYggGUBGdRtFjXxhO8HB0J3UNZHOWMp30Gf
NqQQoiRUIZcmv1KGwJ6l2jxcz277IUOPpYEBhw/MCQsCZjNtCRXFjizg71VV8h5mD+W1GQDz3dhm
jjaK0jCklvAbiYNqHVEFpfwqAaWrspLCmzXGqK4XYilVC3tMuhYKw4pEOClyStPSK2AmLyU8AHd0
kMIgrE8+/7AYhEQ2ZHr5tZRwDzqTwGmDLlDBf/q3OCRIFRu0zOp7MxnuCDicAVD77Ni77hWPiYQt
DwpiZaVwPcTo5t5Sj88KlsENgFr4mcKoNh9CGZ0F8kulF5BYnGQHIuCQVQwFGhsfyMg4dAxAK3yd
s94Vie04GBXQ3XsavQYtqaMQ8N56G9B414rKfTRmjlePVnXkwGHGm+4VGzRoKRUyOWNqaA/vjDdI
1+pbPKZfeV0gGnFN6wI+Ul1vz9u1nI7VcoO2AjKvw7iskPBxj8X0hWbPmpqLf7eiXXhArbkdGsgX
1cP/KyaNJNK0+s2Ir3GernHWxAyPoXyRWqLTTirxQhfAfj+YQA3n121eri0kN0G0hNPSfATg6SRn
ksIEIxyOkqS60WAaSdmmbI/GxD1IjsPPu/0i27N31n3QoeOn0QSrNvVw491o056O8nRG+nhccfCe
NH2XrmNwRRu9ZjvFroJ1kQkPZku1DpFSsB+laJTFFKZrC1V+3Y4sUq9339/VGlPoWf81JtDAPrt9
xBUbGpJ/QBYmuwsTTxHcMacJfC9xMOxqLJEquL0lw1s5Z9UdE/K628MUKov6ADM2kT+IPZSV6KX9
f9rxq4pKYMEguc/ttXvWaMlzG17rq1VlheKdrg3xLLwUhhxCidlxfyQrufPnPub3G5O8i+zpAy6A
gj1jblseP7bEj0Tg4txDxS18LYTLJnUXvocxL6hjZHHNHdxGKRG7SjowbZtC+KrtDnO3n6XQatJE
BO1eWVgN9jUqfOlpOybstXLpjmr9+Xz/FxRMyurzuJYetWd4pKJLJjOhJEoeQzCdp7NQYNaRUVwR
uwRaG/gEn1AVstDJO83iHP7Fyg/WNOYUcNi7XnLpRoARF4hTrqWBNKXEyHE5XfexZjiyqooinWAr
omUP4eiLL4nMSfarGDc4Q6rArcyPLiDy1xNnCdq96XH9QFSsATV94zcLD+g4MZ5NSxI/Iub3FyRG
CTbKLB9oBIVbnx9MIzfTyMgTHaEbDRfQ2+QmDACB5U8Hd9jnJI7P579Wp8zVXS8ULloP4u6Z0kf1
h8nsHJ3dyso2hQcJ2iuPmgfWjZFAJUGODvMoR6DSrpRE57xf0T1TMnuJO67kppK5GiPke5qlr/Ac
TVn6weMtlnutKXlUp3qjbdW6ne8ogEAP7brEIfqlME+gNqczkT2k9Xy4pKRl3D4YmPkl2vVv4ZP7
sYoGL1qL2WhNFiKsgU7fN+mn0PYwbj9GupvEZ8LgiT8tnATXPIXLVH25TNqGoLFmGm1cy2/L5XAF
gSw6hZCVYeuMDNYvxrfSck0DPvi6Oo0y/RtMKiK8IRp7cB2/fmmIXQGpmLqnQ5Th5mgpfO9hOAxw
8QvqfVklyuxeMe0YdJ9+pnNzCbagBkw4ljv5vARxNQZ2hT3syhAl2h/D0UF0Rlkt4atpwFfEb1QT
cVLRfJlozBE1kmR2oCI+dI4GgPLdeG9OFY9gy0AQyaH45RSoN/oqCBanx/n2pC1d8rZ4p6tar0lj
Wa1HLU+X4oaLVGwAfODuujqS55H0BNxKLNz01Ju0+CTvZMWvHfvk3+gXtf+Ajavu8NVw4irZLXxy
Z9Y8k/tmL0w0gQuQyUAKrxngns23WADsq6f6NLd4MWvtu/6x8koACUvprT1jxTj+64X7RmnUz9L8
SLmkNvdtpFGYa3wPhjd8k3k1cApNnOSjr0n6UqWRBCviCbEePcWRJh9zku02ZGPitYSCJhqBs6AW
Ud4Fm+GkUVt2MfSXJOirtRkRmdWR1AdN4UbELAXenmS29bcb+OZyHWF+96YxWzREEkP+8xaSdnJC
oL/9gaeNuMuTjaXgBGpvR9SWotSC53rfnHwPYl2RaFcq7/gi4uuvWkYR8qrkV6aERSeyAtxJYLbG
0xB9a3jXRDOQCYHVnKFwG/x8PsGtv1nuEnrNUun50oDJHox8dRCJhZxTgf28Yk3cfS+JhFtDSqOl
BFbdA1W3m+1cAYy3eEewKb4ew+PojriOzfnVNTcrohOWGxMISjSLwql4tytDf57aI/uzpeewYZHS
6o3dlzG1vH31vWR77NdeVCfV+L2qHi70/XK2u7gBRhky6/lWY8tQ4rRHnsQ9REfmN21oeq61Bq12
DZcC5Fv14uwy1T6U9MmXn5yQ5Y4gLbRT+xg0z3tUfyoNerS7zZ3YPCC8KuA8O9qaywFV8k8cFk6n
N8wuCBp3bQrHvA4XrAO12rYA8CXHHYdPx65x7jxD8b1y7ddpIm/ZheXbUqWQajFuAVI6YUTfyuRt
MqW8+GIlKYcrt34ByRPuZoiNsj1xOofUx3BArzoV1bWxVCYqbuSh+H0vpLPEbLmpwvxFZnKUEgU1
SYIm+f4LJd90IeXe+dnl90ieK8Jx1PdhSVi9gIkdiU8gqCwHvplgUxXPROGaD+aOVHAR/f410Whz
F+Zg+uMEkPeah5gV89p382snli4GuswI1UYu6ulEqHO3Zp+og7AFtK/oqZ1hXOUQTxrdtZERtQgk
tgnhGtINmk2YLe0DcoMevBAWMlUS6Ml57ZOjj3oVyglRtZfs+r+DwwNnB6G3VvH6D6zSHSOIXM34
SdTyGwyB1/PIoTpF7VMgnT/Fc+DtxnNrSrNbmuZdfwN7iDiMr/aDbfnVR/NKMsPkG4VRpd2Ms4OX
Y9emE/NM0orbXRFfTbRe0fYMy9z6mPLmfgf7aa+BOTNExl9u6I8poge/6BEa+VQXzDOTyz0IM6j2
73G9xisTtBATGVsqeb9PZvp13vI1A9rooF78wcUjLTT8bjfOKnX23tfFooSShXOTUCcFZusKVxgj
0PsgiwzeKjfbAs3/b1CDKtHpz0ICe/VfWbSN3kLLcRfmBmdq4iAfKzBPm24WNf223vP/16RFlrbn
P0g50JHp+/7+LhzzPklUYZ/cJhjT0egKjGgwO8Aj4+//3YHrVHDqIIA4ZS0azC+k/jsS3fxpB5aS
PgERZECMqrgux7mmPrFwVZqkjvtIQREuXasmJtsA4lm3ijn3iGS5za9AL7LzaGR0/msl74jBe9Fd
JZCVsgOavdlVHKvVi8tPFO2gEDnaIDvePfQp9iRFRMBRVGQ8mdFv1KNFcwXaBxeBmWp3Z7J0h5jO
PF3qGRiwqAuOF9MFaMmTAlQG+IhPP8Yw+vmpvcAyuozdQ+bSNGdNzrxfLgd25kDWN/gG4ndOHhge
g6fHXF3XayOLh5lZR3BgkFTZvq5Q8izxm3VrsAb1VpIYhgA9Q6JbAWJtlLGq8ocbLJyqOwbIXSzj
xXan05RufcVmDQEhGEc7TvxP8kfwkaa/KUyDTZ4O3XWU1mqkAwOUk3m/v7t476NNFLqHeWao3rij
UuM4Bf7TivcjTkjQiZSTtm9H3q8habyxxaNSwmRx9+Kvt+FJYJ4wf7U55Fmpb9L92oTK9BQ4QeOP
YSaGL/YUyMPTko/9XkUoRCw1ARWzssT90Eaq+PSheX6KJKGMtiPpnEm7W0dr8ZjfO72mySkT1+YE
gSKYbpkisNfb4V9R6lYuOsWP77JiXAL6Q3aJaRabWXti4BKf+QtNsOOMabHRgT+I9yX5ULzNfJ7P
fj8yGGXyWWqurMNbydX79iHTRjCtqPlvE0UL/1pmHXmFbgbUHb26twFmed/L2Qb+yFsbyOnYP4UZ
t60IoRN8bxywFppMmU6/jXXJCP/yw55g835+cQwrxmH7v0pkwyQDHcTgnEf3zhpSxvz7OjRqOIEs
aUq80RZ16nFXaQydlwksoQvQIj9qvKuYmrbWv7FeX6uAToTaGPyiVYZPX/eHn9nAU7nu+PAWXSW8
iXF7f4fmMKmg8qBzxg3wRdmT1uLbJSwRo4tNLYygmstWnqwNCWqhGoBMMqnw1oKohffSEHJ1X9QH
zzabx/63V2od59mj8HwHcHCqsWld+a49894zhHh40ZK/po8L31nxdhk9LLG6tnYPiiXczpNsxQFa
mNMw/kMQ2CUR6jMuuvuLChaWQSRKtkQyM+66TSjMElC1JArtkYREWC+hadlSt0EHUIPb+htHkif/
VmlXUCkCal78JLxKYMDAr1h44NX4cZxz3XcsycSKQCkXhN/WWqUGLQJyUn5JjH0AGSyU6G/LjJrI
QP5uuv7tafa28nX2y1+fa6USslFPvE+3ifNU3L2oCzXzMGgGK+q9puQXl8Gnnh+NNPCJ3WbiFOaG
xUKMzdvnh7vAbqh6nksyYmUPklvpSV2mZ45Y8HcHH4l4JojXaFRbomvAyuqlxRby705KvGj/Vdyv
+dzC2HyfxaUvjh8dIhCFdBNthKvqFeqv6+vy8eVnxkad0DSjyw9g3QR2NV7aF0D1JE1iJ4ptXrAx
4P96uj5p/JgWZKTosZnSP69t95ExLeSYQF94H61TPGca7kKsqdLR6Ph4TYdn4QGmB4Rv23WofLFZ
a79cWBCDkBrSlqT9rqPuYVPovuoBKvTHVLZoTBUPKSdpdEsW24Hg4dGMSOJ+cLLDs6Fpf4iCj/xj
XcpTXEwGomfCRflXZheKW3jgC9DpRIw5wA7EFTO0qh24xc1+HPa+Vhxp0ET1BivXjd0bmYfIiWb3
IJHeD+LAokFWVRk7EoJWJYdMJAqtTjJtKvQR1zjBR6FLi9qlxnJyOKUVC1s9d8ebaYaR/2HX0dKm
7IZs05pyqVd11i+NVWpDjTZEpmiquMlQizJl/VQY34xxH1khb3cCvCvJqxqq/dgxHnM6EcSJqeyS
8UXtbiCXOdjK/cP7mi2OqlgqM+LCxXvuevZLM+DZiqLWhkb9Xal0DyRXF4SpSzbtg9o9lw+NToK8
bft/meIzb48h78V8AZ6kj/vB1c7YeGoa9dQDcPuYd/XwLXBuFyXadUbdzGbrWM53FKI1p8p5Mr/Q
6dQKjBigDkoOX3ieRgFPHCGB0MCf0EMxPLVIV8vGuxUigNhg7MvoOqMMBFi/3YEmTp3fbdlCASfR
xJjpohBlav0y2iFjQX5+1WTW4WLvyB+nuqWMIKxvO5AQ8xG0bHX0Iihh7Iy8AO5RcWMIuSqSGCvP
AMg0+0ymC48Yw5nsqbbZU3plfNb/xC3U9bVM8yq6y6FK2p3JHJ6b6AbIeqU02S97T80CYZWFW2SJ
u64ZldeXr6fqsXBcQQFT95hZUNFaJOIISKRIqXfCUbQLFGNUJLlpGl3I1LaNzF0IgB3//ZFEPv19
I/UWzGDMucJTrR0MjcaDV2oVZXdfqGj2SBsvkPdaph9nkz5ESPE3yQ+7DkKnTxZrCYssCoYy2zue
d3LR4x4XwCyYk4LLOL4mOsRtExp/AYsza7qWvveqYczJpp38MT+v0eq9niVj3pexMDk8+2trvcsX
UzvmCujuVfdTmUB4ZVJiKVkZWuksHyJIcBfsIHQWDYibD4h1qQVOhtRMXWkt8SlMPvfbhL0xL2wW
hTiOSxIxM8jZfesynXmFuwPKiV/2OP+W/Z465kgJFTW6LuIfHb5+nWutSw0f5JlhL3L0typQ4rSb
wunpljfCazG5MdNjp0g8lYPlUv2Ewu6/CrtH6m/4bAV3Zg9zk0jPbQ6U58J+7/qdtQ+j4HyXYp02
cEu/F1G7OntYKfgsffOC0zca/hvAmOlRP+7/SSdEaB/uQjgV3xV8h9aC6pjiUwFGTLkEoZx02Mnq
mgCxHxaxClNMdgyukww8Yf2Qt+CTOL7ZhCT1GD9lnODKts4EmQWRkmLdqFZsmxF4mneGkGgMYQfm
HhXBUKyfcgEl4JP7Tm+OKOXmLg2nItBzq0uIE9j0BLozqsK37Zp5TV6lJY9ALSKsX8b8Pv18eTGE
TNp0HDL7R2i8Rjb6OQOogzSldBYiJw8Y3IOnNXuGLcV9l7NicVJfugvpzpuNuQMnXcZpTbU0yQfe
eE/hX95lmNvTyQNevRXoLeljRxapsvUbsbBOPa5MXuorI4LxiInXPZjxabzjQ0GCdoodmG4BOnQB
YIHuMVoTrxetnRqYU6T6ylxOYgWGRvlXlvZ8rlbsdg7if+q59aOhpFmELG/uvYhaMRdSHsj1RTrJ
iOJe4gTb6pIOCwTYENCN5sbpA1Tc32I3cLFZHFJoA6L5muqee1dZXzxtkBKgBv9YJ6cPu2Amxo7N
CifeQLLz7M4YvrNlpvki+L6Plk1HbiPVlr4+0vYcR+PAULf0ZGhnR/MOAaoqXY0dn7USWLpwOiBm
f2HmmACCLEf5dvEIO8UmXaC8NsUNDZACW/nYq27/zRJbKwLjSfpfb4Fd9GzlsROrwLP9MXKHT9sN
TsnOICsZAXQYH3mBQS2juLntMibmgVLZq11Ah+cYlSReWgeRkAK/i1crk/jaLjGGiQYHL5nvb2Ym
aCYITxZe1lQefr55jvRzUNnz/C50kjxfWRmtStIbpRAMo3NPvlL5/kbGM7SXBTOf1NjBN0OGeGEF
at4mudxa2sSipUHIaD1x0Wlap7Yx13xssipRkfEEtRESJwBFtN5eRjWvckYYY0MrKjQpbGut7eoE
lE8ht9HnsyG+7wq3XHv2g+VTMI8Qz2blUxQ/8PMas669mDiuJfLX/oSLY2jII3lT6OygYSMzQHaE
CBNJ+AbD8/K9amc+9RilRlSC7qR1vHMzoUEB/779GyXOkd0e7DmobRa2Ooi/CmNptyDQzlroOwii
N4qcoiCbyRbRErYCc3PeqdueXO0wEXudluKa/6zRExLJxCRhv90lBgS0zOvtHVht5BKi7aa40P1H
r6an+vXZBctyueU9ZtqyYval+Joe+aybggcrl0C/IUivP2sruxxHmfK/A3w9y/PgHEac2+MZQjIn
YFcULRkIeWZE8Gg+F0KmphDrxXR+f9QJPY1vXAyyOW68ABm19Uaq76wzjpbc4nieP4SWiOe4jRZA
QUj5ozbY7A1SucJiol3OjhAA2jeBJ7RfhawMF3i4+IelDYhmlqRUxn//bPDyE5L6JYPXdgQT2Nwo
LHMTfHTXC8lspGBLn6OOzVbWdBk4fqygWykUufMd/YqvONTMeHtIiW9XSvQxum/dNpo1t0ykeek0
2nbXHMbXErwnY/Ys9aMJ9osJDtfrk5j0Z4Ws3dyWPR1guyUUqFzuPGZDNhjgfzyxKHRXLXr7syid
SEotUy+2fcIDZrRFymtaI7Oj9VWtTriLebauXghyrzFn1MTYugLss1w+oK5tjDlZ4KzPSCrjqDat
07T9TQDjqzKjfeZGlo3ICqYnZDg+9FBXqaIjpE+nys9JglJ9hudOul6lTri6WW8K8boCgliUVik8
9r3fhzUO7fb3fvWoTwjX7C+N0k0y+NKwdfULjQee+vxuLZXcXOCez9MoFmzc9hrHa8uwhDQJwtOJ
heNc7zXbNZ8Lp+wQXrmGWloEmeJoeeC3+MqMgN5aUAPUTUI1NuNzdi7ZvDjWVfaQytYDvoq4Ib2G
Z2T4B14HwYa+1Ylv/3fzJzB+QBUMaaweLmSO94Pzxq5U6MnvrOP/4wO6CdMcoPS0jSiOlUd4SHin
aBlEF3MVVV83tdndAry4O+ioAfQ3/csoEWgaIaton2Nta0rGx2YVfdHxPntl9mVUmprsVER+Ih28
mq0kf2ucwJF+er2D4gJs8QuhzJOaPFkgwlIaDWGoIsX9B+th1VoEnpDB6ILpAptOAgfP70TfPpWU
f4fnCbwspSWDCHtolLeDPgdoPvolYXLeGiomEg69QsaNkE3p5gnXnHV5MsT6OX++4WCEO8JIXda/
5tdDeVNpz+i6a1ITRY4P6GChRr4wnRShXPnakyVWNpk6EUbzezn7a+WsLHoVl+7u4O1lOHHBEbxy
oiI9A3FkbJGh7KttoWjywsa9B4iCJl9KVWe5ipvsOcZJaMvFPRpcoQxFc3mXlGPFRORrcuwS011O
DbZ4ZyhkpD7UUSvC1XRZ4OYp4QRk1QMmmXhAcWcg/jvLlJv/etCGigZfj7DHAIaCZ6D8O7cqADzv
UAIvUHWd4uWMFYfeIXnxraF8ZB7dyLr75jdU5gbgr9hXrRGFXHmtEhNTGKzybadAtAJUA6s3GlWa
yloGOT/RxKxZeMUNRpxO4DuaKCoFfiLpFDEStS/VuZtCxePihkTe5aSq5+uUKoc688uGa3BzF/z/
pMetURUN3P1xkXKdOLgxy/TKJgxFAfyUnCQPqAmRQEMXHTu4FB0f5Ho/vAxJWObQOBeuYErd6Ily
z2KKn5OaetdIztHLUAY2Hxdm/Gdsie9doWxhi5PW99Rk3XuoIrVDQlf5GmM8uiEa/BO8M/oUEdD6
RcZs6xiz53oMeYNYranwZXvX6I37+ZnwWCMKYlMCnZfvEOR8azolHj1ABHo3uRf6VncB6XNeLZ8W
1qT/DQbBYqASyIoH457Z0NL6Z+ImWf71tmnXinajZaWMJq78SYoJmTeYkVB91t/XyaSdYq23WjLw
/UUwST4lHuP79BAhwrQhKCuViq+23iTyVwqhKMnAM/tIByI3dMGbB+GzBZ7D3D3ZHEgShR6V6TCU
uDat9Y9/+cOKrbsf8p9zHM3C/i5BKHeZ8FgLWfWPMAXjekmGN+Jxv/40MQZDJyReZ7oFdokosRc5
FqGL9hBUIrOlVhN1ieoI+YOms6U4VTCnDdBk7fbJ6o5N4lqTv+53fMLApZGXhK3SQE0XlGGq0+pl
Zy2BYRiNBEY1lycj4DPGzirFEVD6nPmHJX8XMiv7YMSSrRp2KSCp5JW3kBS/4p0D1f6lvTnGNu/t
zh4aDoLOQB0Qie4KiAUaTUZDT1Porv7B1H7w2sJJSIGcOMtawGjWpd8hoadH7UFbAw6o48cUPzz/
5rjVbGTMvthMj7Pap6jG16H3wNRFO7w4GDt02K2KDcTxTLCo4mF/oUhWAa4JisV7xPrOx6z/akI5
YUD1riFU7Gjs2vupKveck19u39KkHkfBLu8tmFwZrRio8ugqxpUO4ZGtYH3qjqOB5EEndMJVYyIE
XUpeZm4JnHLFSrQFfNQ2Nuo7Lfw4XxmmBiv+ZDPKUmoB/Q1k2zF1CAwy1+Sjrirdbi6TF+MS8r2D
xWKKuzyUGKuvKs7VGKwzKAAOCfhddow+EuyPWUKIbSc511bvpwHn4MH3xVWys/WybMXb/lWPn6Cq
o1y3cYF+eurZD/RRZRyKRdZvPozaHVyGFmAzV/OxZihVm6tljbIVvmIgJqxN9BQ+yi6+FirbjxtN
NupokKOq222GluevW26huLSFFx2wFHSTXCVrqn/NlCaQ9H3i11kX62MbzRIvMurZI4KnJtHfNgyc
3LI1BiF/Mqp8NTFQ9cheubh/WM9uTXQgY3tm+xBcZJhq3vFqSvGeePoHZwm4mh5M3v+/9Yx7z7fW
sa/W7vXEhbCUHDmzqbBxD6Q/u9sMudI4MYm5c903cF0cgPtoyhPjSnM36BnWR2icef+OLSD7l1q1
6MGkjRMW0gHpURea3+R2g4GD6FqjY8ODHD1EvHBkN6BCVPuPJRMDSuncS6L52aNZicd4ld7vGmp5
WX0sRqlJHYg8BV9JA5Bhh7GZo/IjcSGbBag7IQMqT5SIX7BkjIWMLEI5zJ9PmZiBZXA0cVVPe3xE
ZEcAOZQap2xxJLlrPZ15B7Yz9MqRRgYjXSUIupX8fhqfikxw6sbe5H1Jk6F1ArCrJLdvtj58ap7K
ENKro2YRN/W77cuCHHejGBcSZgQtPhr51h2WiLVzIGSVyctoRumyWs1UMfLDgmXPSMKxTUdniQxF
tZ+reFXoKYbT9pcQ8J1sA9sS6VtRnLPG82M+ndBlYKFmev6vrOccEw0fFYExTiif4CXX830jscNF
6n/R6KxgMh5Yz18/yo3vtTvQVaCT5bofKjQJuOus2J7Iu9jibMqFdJtoDhupYuuo0inWp0XV8zw9
CsgRE1LdFS4ynMecJg+fhSNxDL8XwmmygO3OYLUFLxYoW3tufq1WlaAH3eon/Gf3FTBIN/2e3H6o
nin4/c2zsO4WZNq4/hYbLPLdtn8sYWXnEOU6pGSR7/P5+YvjQHg09UvqsEZX/qR4I5y54O3vIovS
qj0nWhSgKGdUNKG75f4ZlYgvWzByEF+QshpRUkoZliSGel2sBD2ZzfAQhQc0Jl0G6Wsf4oV+shlE
icCJcuNUatkNzXZX9uFWyJB5rFZj4Ww/JkEV50Kvy3R+QPBaKorWUZ6vSoK+i9yZFc1Hv3LbHClN
CUBRrKIvpJyE4n1v1i/SNhm0sUftp2D5lsQYL+HfFf2D0V7GHMkIaadMG20Ca5HZ8J+UJmT4LHfv
mDEb4gy9LORwMUYSzzneCW39CBkNNIJqfGdA1nU/MA1U4DXdq6jPXxy4aQfZhPcaR81hOvQ6yxvV
fQVV77Ha0hqf2iDJubgrRypFr/Bk5HJ4pU7FG0BdtvkvU1UgmA/xRUbbKj0k/g3UDHCXU9KPp/MY
gqGkGmxJ+G76fsB81Tq4DMmRQAY6CaMgYleMxr0YCuXgKOKOZJfwn+vhKSw4o2mytQTHe8Ry94mT
CiRvOA2mmZ/vZ/EUOEIfRlokXzqv2Ho2S42JVfwWOwOEja/G1g82AoMSmcjtjmc1xbv0uMEJv1WN
fdFDKWnywtjtuWR2+TAFPR7vwJatdNIbL3p+768yUWEwgADIOUmycHBHZ8P2ijGKjwe9pEqxvlgn
CZoJ77cv01PtTEs6QoegPV+vxXmbK/1DziIDx4dOcwVr/SI4FlM1t9Bmux6vq50iFtxcvxOo8XDp
qS0ofsQrMLIVXyebq0E9udbIqa+Dee4DjmkvV/qOgF7jj0rPDwC4Jhkk1BILprfpkmyzx1yNxdEt
K5/O03uBEPY5HCxD2VBen3vsjOroHMwc4ly/ZB8hbnj3yzr7ZWgSnHaD9AG6v6cCP1oGgVRM3+SC
IHLPJp7+UGXoldkvWsZWy/1VSu6C1rIt/rAOVIiiZ2FDnkoKgHe7B5qQoss9vtdQvmqfrVgWfEzu
r2Bx6JwQ7NfyCR7ucqzRzx2XSqWOZIcr33BplgwlRSw+2DTbXDNdyofVYucar/GFp0CrDXKHqe0r
Pv/0djf7XBnYvy2FyTsAaayPFf24Ubn/jQqfCLWpCavJ/Om1Xfevm/BOSV0CiKTe/ctQljc2ZUoR
tho4FJmm7DVsnDFjTg2Q7LsASCy77hgBImMrMGiy+76qDeLaE0HH//7m5VzJdApF/9Wza4Nux6Eu
cL/ACzNSmh2lklK+1yuxuX8VkFUkjM//NDCzXxcUKLUl3jzMbrJ5DuGYHN6ruAWEn6S5kqnafBL+
KXWdhxkvrpx552EO+hjaiAtxCra6QCN/kYMmk2qZPkuF5cFv9ScWo0tK62zkAjL31KML1e/CKGAq
YXovrWMP6HfsOyCWSx21bfqyU9V46fFWJjPi5YE9UPoE4KnKB0dEfVQxA9W8atAki3bofB/XecqE
Z7xHl511P/2vecIjSy7zzZ3ctIJl0RmGixmndFrpWgjwK3czMp7bUhx9At+0vrFkmlXnrioxgRb5
Uystsr3/wOjf5Ea8PqHk+jz0IpXNqr3n6oLyasJ+A708MqVL3smwxA29YYBsYzMpWBpz/DkaUQqa
rZZPW7VWRd0CWQEEyJnkoAwU02uOWpCq9hP5uc2EEEKslwT+NEU7kpRU4ollUDGeFBmpKaHuyZo9
0wK0iGQuY0HSIL1zgrRFDtAVWWpvDLj5HyqPIJvBHZ+DqPgq/fpY0TAskdeqa9NIEWHgi5+Qn0OU
pvbFUJsxZ7jQA+ShyTCJgO1Q3lxRY0I7tqzNU0BL71jFLVINJ/v4OrXllCM9bXUoYM0ADVVOUH9e
2hyu/MVzFAZBZ0YdQtHHN/Bni5Pv4ZfA2r/+DsPfpxnQC+u8HUP9tzhVI349DwBsrwJeRqk8FrqY
G+BkG0T2ullgssFP0nmI5t0UvTra4wF1YL/ka5JAGjH0pPX2asn3pKVquoideVsuy7Zv29w4qrDF
6zz932sYONt5p4oUvQFeKFhXrTxnwEfrwgAWkCaHX6388fk0j4wbm90AsnvqfYDvs4Q9joq0XjS8
+8K/+3PMubr9hE7MaODLUJm5SXoOWTCezNMND2GC2FsQyr9DKKlEfyo0EtLzAO8V+GmAG9+yPaM0
bVkGWER22ZBCMw8B8W+RoiOZ+Xg7U0/WIsnMPIr3VKj9cUdXD5mCmCLVt5nzZksqB9v3DB3/RtGC
vteHvhpx9bFhrvg35WpepO8aa31jRHqm0cV+78FSSZfOEeA5edxrxCARl4B5UQynwIZdpUusvoj5
98QCjFxL5idzVVucpeWjTiiQtIm0xb7mAnP+VcZE82QAAceXYjIbXhunC3CvNzdNOpUhbknI6YiN
yZhaF45DvspZyvaTDY01My+9f57pUKp8C2jc8LwlW89JZwuEG5Pjv5jla7l51T1xtLhnTUilvgXQ
wkRwP+zT+xEXlC9m69WmGjsyW0Fo/VgAPSSIsiQc0fQC2VzH54uym7XjnHhN5WNcHyI9NN087sDi
maBHniiIfP1WStQjxSkF3zldkKuyOqd6fUDKtYS3/ZpsfgRafz9UxituLfzgicogGTMMXF3q+Wmu
wY8o8GMZJJBXDOIiPiOQ4Rkg3G74tPK3pkQFIgepa9RlxQFHAPtdzo9u87G5XzB+5tpYHk/K2NXF
iTIv5bBhxwwhK9mAYbi2vsAoHY6ZscSYMHUnGkkfvcQt8UpWlGquXqHsE940akLLPZ6RLocd4PqH
+p2O8MK5ePt9wtuCsxJ20I4c/p96LPNYKPzFWikKbOTREo6oGIvdREbpx9HdTFm2DiHOxpl2A3xT
Tx2Uc07FEvrfUIeK2afWijGQKpBWptjAOdnuYJPFjIrWpGPak4eTQStyL/s36Cc2BgdxqtIdeoYj
NAATFxUaCGaWedrj+SI+EjuBEJ68osD+ACrdgCdIF/5FtwPpZ6D6EEsXYuTCRgURw8AmzBwTc66T
lnvaeE5h3DBqHolXWxzPy5SUzRuwM4KpGgLbWsfA0S2TXnUofcm0rLNqDPNoxg7q03mW2+4wMOHj
nqAPfCr8bZugw/zDBdDKJRxsPPQrY4PnYKq63SCFCHXEUnNt1P+1/1CIGNpfI6K0AI06S+2LDB2i
ye2sf0mtwcWcF45OgK/q2qWCTXfOktx2cxscW3CVd6vMogT7btZ+AOac58PaoLonKks81nm8i16p
xEYNsIT0uFgGVTNISu/vUqz2+KhxUIPOFkKdPPEI43Z1EaKrO+GDYM/Jc4cfsSQ+ROaubvI4rsWQ
/UziJctaPR28PA/PTkpAvgeIZCkjJRPiAcM+BaDQ++esVH8jWaWseww3yegc2mdF8yMNg2MEqXdP
Qpn+hMMnQ/WiBeLMvolewPixbPdQsYGDUrHyVrDXCFYPMNiKMV9oZgMNW75lIRtCdo7YDGOkS1xI
2PwTKar58T81cpdS90Lb2PJFpCcpDfgtPVDs0lgGjzfRnDtSZp0buF25KFBERIiR0iQ7GiwIL+uZ
cDVTLPnDr+9sa4LaFAREnip0YbIGv3HWu3gWOyEzuqj87JZRXTzjAdk1h21NZt97LYlMoX9Bykr3
MQFg+OZnGaYu/xB8Q4gAT34bR0EICR3gv/nNbWlwh/KLoxgtuCM2RI2f8QoMb+T2h0RRup1w/x5K
yUww02fEHbOWJcNUGbE2DmpoKJN8J3sEikXjBljxW0o2z5/sbzCFvsPp1/rU85zUsQ+zdI14Mzsu
uHcVRl9+gv6iKxQJ3cyQ7XC4PehWRLksiU2JzSnV80R9fu2ZY7IcCKaH5bypSXmkzl3z+tkaf/12
ao7BshZQHt6w1lX9epwJJkyLS3Bdl8Kx0aO+gcOqoWfSyprvl/ZaiTstizj6fDh0tB41IrSA2Ppd
Xq45Ds1BylXhZzlOYzBIHGi2oDIbjq8NOm7wOIq7AcpHgNUbVK7jhs7MT41/6hwd3pLHEVlTqQZx
21kpeRaX4GJ2xxBDojNDrGVzq3BzihA7pEeeqqgY6UwqgtlLl6AU6178IdqZ4OrvhoYCRl508N6l
ygNDO0/ixH65CPEGiBHC8lMOgnGx4DWjYBR8zR3TOcN0zgxQ0xUI9dkFTPE102QvjxXlghdWo0zO
2LLQaLRRGF4BLAF2WYRuZugMJGMdosRmyQ5jIVUOahAhjejWQRoLGeGFdjCEXzaR9PQJNhMgZz4K
pFe4GanJ7WW0cGRkw2TDVSZBRtI1SU3K9hYKiMnFRte1cuW967Xp1IirdscHWUjZlwFNmqCPPdVH
jH4qYrRtLfXb+TIq9PMU+CFORoQkZPA8QjiwpybIev/WfgSIYVEjmwEBVT4GL3MVYM+LodIccjfi
dO6e6ASOEa4NbCbAYMif/w3GTwMOWpuDI/VFUJvX+ujI3tz6EE1VVhQAEJWW2QYwlQEHsoY7ZYNh
hCUhB59v7QpxC6RpaBClRz2GwWinSE7hxbRZ10Wx/bJ1mGLxNo5/m9p+VAhTsiQfjJ7/jfoA4qsU
dgs/ppVKP5x+kziJdjmJJhKZ1vLdWZPqgde+f5c6BQbB8eNWm77yN88AOP3xQ1VYa/KkZ7F8pQHL
+91JxjqyP121PN/ER0o/X9o4MSQ78kAbhC+kK4Czk1DWmA79Lp5LWchS8GzkBbDT6Bm+Fm+pFcwi
X1TywdiIUXe2SFIwk0venC/1+o57bv5CWWLakSCsYxyHgEmD5rRDxmUmeZnqyM/ryYjHERL8cyEh
S8puTu3OEpvQ8a5OvUAXwC/st/fzhS+UifmHT5MuXYwOJG1PaB13lZDGb6i9zLX3RAensrjEHjHD
u3nfLnkWWcPkXAIpYShO5lxxlIiIFivrt20m71Fcu2GmRT9Dz9C1xq34DHzk9dhniwwe3NrUkuNv
1SJBxZN9mqsFhl0EPn1dOLOmmBLyK+nTjmljKQ6QF2D07IS+x5xi3PB/kFy1hSBI7gNLAZC8attr
r5xxjj8L+y7FQq4IIfZEg6ygLld4Y1WQJrLJNT5Wy/jkArfbnpsFEeBt7uOVtqvaC3to3ld31JiT
wLB+9NG4oZ+bwvYyiM6a+Lye6E1a9sFuch1Xo3ruUb52QJlcGnLLgejCKgfys3omWQdTTyXlizZ3
MHEHj5AsxRTth6kTTQnAp0VYQeIe3UBJXZiD5o8zfdMnvhM1PpQZQHxY41/Upjd0/6CMEZfqwIVh
wDcbKX6oQ74zhEZb+1n+yCviIbUGPugSJN0Mh+12EWtu2RmL5Gdzq81ymHbB1w5FFL+iKnCHLZo0
vvXL6Nwxb05V5jE2aGIoBGInXC8gSJnJDHYJnCBvTQI/o6Hv2Mk2Zfk12HC3t4xREiZNm4NIikvT
gg2aIQxmgt/4Ja9Uqk4kBDQKWBO+oytoFGgKwdPKtN91HV9kJxbfpQI+3y3d4mznhINciiS0bf1P
yEbta9TPyP7HziKMjJknvKWbrRfhhNPyIPyUpGGRgcXnraTRKW632ieV5IDyIYZVbXRilbaw3IBr
l3chPmh4P58Z4yqPcJZsb6I1NMaembfw7o1EeZMbX7/lB8vzGYgt7RpMU8fPiOSK9NjFCRFDifbO
PgGQ7jDsXdV/JOfLj5PzetiXZheOZKmAFGIEAg+/2SyYNfA8kemfOeHNDjEl7nOUWism4Cu3MHtH
EGtwwGDR5IHhTwbFhvHvJeQSPWeaEbDRurWKBEY1ABh3A0NAXhPaQjMGmuiafeixZi5qsheiSzwK
aj7l/+eHJfUYvauv94CIEMYDdgdPvkC7t87fdrRwDS+KH1j38mNFE7RacFeOYIX5iu4FB1UWk3Pz
I0c9fH4amUC3C7TwZjm4Hlq/TE7kBftOrFtcgozuasZr19eA3IewmREo452VjmcmXt8c9Z1DngLo
j+vxJ/sSBlKGaeFeqtVxiBDrVOKSc8reI3x14+SWOR29EQBNZiPKVy/sFYoBmGwXm96yY7nG6kuD
emCxda1i7Or/pL95r6dDyfIMeOC3HzatZDwPaVmcio1Oib/LKijcWU56zt+ZgcG8hD8el1CDMHs9
19eXyHmx1TYgGjfWrXyIx7ul6TnWJlaBV2xbd5jVmFeqxdPexdygh7uQEOp7/U7J5aWUG4tX32ZX
lj1F4VMPzte68KTtOtwpbVxlYnvr5ri2NHava49wa+DO3hS7KZGbL+tUn4NOCQyVdH2hyA5Uw73C
fKWTuGUVDDSTHk52bSinoS7zYKOknzKlnJ5ipoiy5k90GzOdaNyZElInbJoK6SSva18c4vKemEU5
tu5pFB7rW/KEDMy/bfUjEAazKah1h1iVgTnpaC2uuvl4g/vdYaKforR659xwHM39Ph53ILHAO1jH
7n6twIODrEQqfrQLwVASjNkEz4S3zwaFa7k1t4M58+gGLzCeNHGnFHfXSMRYpFylPlYfxHaOcAK0
uUwgDSR97V+kAO4JE1on7ekr3exX8UODrR3RYrUolXvqygy3nW80ICPEzlDXcaz3+jAtsNY+ByK2
K9nu5GI9To+TSkeo11TohA9oBD8LlbgClQX9FU4EPYrMTi1jd430LDj6i8wUmt4in4l/8S16P7Fj
XS2qMJWUWKn7N08Gvh2/87TrR5wlVyYKujnk2PKTl+F2O08eGdc41f3auIEUVNiI54mmsG86Mauh
4GovbLlWdscBb6kNRlx1mPzZsA9S9NlNEUZvW0UT6+KBFapGP+LWpsCXmkqWvMgf1FeeRxrAv6Nl
IGFeQB9Uy7fyRRlr/B2bGsBVvwavcf3S7Gqrkd0a6X9smENnaz0W/Z7Kb4q5sSBUxqYlf3EXhau8
/zVHQbNTfiMcp1e0ACe0rljdBuEgdPPI0tmAt8D4yMJgNyjCaeP4lAtXuHn4+g5VvDtgNRH/JgY4
RV7EGtA5gzX9j6+WYY1/oL4scVAbzjawKuviRZn1PPFE1sbpJ5xdekkLBbCPtU9kyAAb5T8h8jgQ
Wmq4exsMXdHf3lvDO4207xXBjE1sgnt+RnhVG5jSd5eTmuxEC8W2PwhrJRppP3w2QY5FJ65Y2IoY
hAPGN0eT/1dEKoKdcvZ50VklJ4uV/WQiPC1rIvnGgwqv6XO6CZg++1IRdTTRQeenS/LmyoSk+3XS
AvJXUj0dPb14T+TE/KPgY+Ri3b7XGFmZ8qVEWICRuJ0khsMoMIoLWEqCEX4S0q57DPp5McL4XjBX
XaNimAZhA/4Qo1XuKQVPPtf1I4l9N7J/RewTkbVChtej2hC5XLo+sK0qxATc9jxygeaPLLbp+W66
hgQw2XuleAj2mocC2b7IywjevW2n015W8gmxFZ15OPDH4+3+U6RFhFQtD22Rx6zkniLUD9cCVP7Y
+exqf4ZSivfsZ4eqOK/Qen99R3ERn+gutIpLlrfeJfYMKD79z3ASOYm7scRTtNMec+oPmGKroD2S
vyCMohHFKs/D6zzv7SZKS5CWxAiP6W4JP/eFw25l1iiPVaDfiBeCXJE7xdNsln5CdySBBYDWGSDF
dJhqK+TdyWcBqS1fG4VUApPR8kI6z0sXNgBFlYOVVsHuXbBjjOfswb5jC26TH8vqB5DpBukHIWGB
kugkrqD3Q+lwjrALASotEeafw+SNxfvn8XJHmfXPQ+jOZyVNlz8p1/KR8A+0XUweI9eX7ZnRv6L5
DdLZawudVPei5bQdf7qEalHaan+Yg6RgHIS80uraAAHfjeKkv6ZsSkSSI+gDdMDY5IXyLy0gtpqG
LPibdRsLSIYlqNu7OttGUEC37Z2mG9/iEQ5AVdWEdrrhARjFliVV32CYgt/k0q6CghLyRZi2xkpj
f4WwnXaDyNcphIZr1zN5Ve7QQATSOzth/8PL6g/7EKP8F7QVXkjquvMfwR2yuA8C1RIsJ0gyTUMi
szXJLL6DBVQ/Pj0WmqI8NnrCIivVHPt5jaicw0u+61kTNtHRLczPZ/8+I7Vnf202ujCPROaPZdRl
ytp0YVoDZIned4+eFa97KWZIgabTraPnbbp2dX7qFKOWHZm8oNliHFAFAdx5u/tcyZVrU9QxR6+p
jEQmhglJ3TPLOmF1wTrSid718/nAzHE8UtokxPxeqaSvyIQT58U7HE21660b+42PowCYm5QFVk7h
2R5nHLGpoTfQ8cFRiD3aYAm8A2+gzJzObfDYfO3ejcMYXdpdW3HWM9DnYyTf0vDDHjaiKms4/cnM
hR6PA1G+qyFOcx9Iy6Y9c1sWECvrAjgmqqBFTnhf4LeWSyGJZMZRL+1wvWGCB2tBlAu8xnT6t/JA
2WfMFG9KXgCk0XfHvALvhUC8wMZPNvy6P4YuBKO8ILEeZ3uiBNd5bC1h0SppHolYz7TxHx6M6Irp
SMb4SQOkQcporDWNPhFP0PUAfDtaORv9exOkWpX2psQXe3EUspxpHYrN8T7ORkelkOcy13RFHwn2
jO2JEN4lVsAQcjiKanr6DBrdBjf39O2JUwP/iEfC13VXgaZax+rSyIcs6lgN8zJGckzhnTmUv6ZQ
OZXi9IW5YYc2UyEAoDCcB/7u414EbdfYEdeErfG1/kSjQc3szQgKTVRS8dLIbhSLwXY2+UtA/4wG
B6p/seD+XHxs2Q20PYAwaq12DIwHTEd15T+UBg2jqD8jmBoIpQXaQUIyvYtq8TVw5+iz2BMUwZkB
Kpv6OnwsJ0J/IaO5SpfTT4aEeh6/KAKTgrMDa44cr8SduW1jeRiXhj5WyBY+9+o9GxNb2mmjMqxt
d64GWmIXtc1XgHtK6v2t/4t8sSMNLWsQFk3okgwdSmo0TChx8mqQVN9RwjRt7TxuJWnUCFFFr7ne
XP3Bx8PUxeOmZn6eqe9qPpkYT/nTaZoUFglk9SejgzEY4leeCivm2fOc63TXp3rWR35BajxxFsVZ
qqh5Q09yBJUQCCOe5sCOwr09LJwH4sRSIQ0hKsPOF9pt2ROPWHX1uzE8y5p8RBPGDmBsRUCuxXwu
vKXDv9m0Wmz6HMvMBnLCpa6JnZusAZ74jmN1vu6vtleQxuLoeqHSP8w5cbJCFXAywi1zpW7lzqiu
tcIixlKtrtmzgztANOKTm8OquLXPOEWplIh9qvyYazZVaJRtQQEKkPCYmoq1MZCeDYcvZMmTo7sN
9CEHjvTM+vBNECodf7nwDvkBNzapyghOgqWwdKJ9UpcdTawgBrm1rzPfV8v1iFLJlJOzERnRKdhO
x1ccw48lX2S3iIaplDy4U0lkajl+WdbvNZ96YEczu/Lh5nmtVg1aIiY9JXN7u/cXhi3xofV3OGUV
msgFJOmKbvjQmgcmZxMXCL+LTDxK4PXXBTvd9d/837JX7nVi51Qwmx2l/mBEHtP4QFqArJDnAhVS
XV2u9Bpd0pnqoO83HZiHKdRDWhdc8rleQoQs3RF5PixFvIZdkeK21iIRBPIbZCzaAnML03ZKWvW0
iEROSLEVUQ7iMqlW1IK7K5MeSuEkH1ZIapuaDTQ/PZ24QeASkw9FT8y0MFlhmljLXEBaBrt//Ufg
rNH9KuRxILbNBlazvjM6L3yAcYzo24cLmb95VZg6pWFwIET9lUWSFRYOPxdSLinHYU65sUUJfr3e
/WBuhw0obsKPwRgAyd1B4APhWSJbMcZ3r3G4Y5NYRquYKxzXGVz84CMqhjYZyx8y7STbCjvGOwMD
n/QYeKcPg0JKHdKvSd+K/e1qqkbuQreXcoirwjULCiKRKiygkKwNVPogPAU5qakmOOE5//gI2J7h
MIAUesNY7hKbUMt30kYcB7eBhO5+ltShzAuTkDv1N6eR3rx+aKanokic9MtrzX2Oh48Ziu0ys4HA
mttzy9tl0GIXeh0+7fAH3xuDK+AMb8lisH1JuooxkAHF88LYORndnfdzJosWUVuzhgzQTk9yCZgJ
W0aQw5AV/ttvafKbwzfPjypdio3NfOcHMxTQa0AHsj4hJGmOv0m90Mr1+S1pp5vraeMrg5v9a1Q3
7UhljjhdSi16BGXQzoy0iwJZK94lL+UregmduoDU/eROJwf8t0g1QqjHnUsrbQBI//f3Kiv4xmKp
JMCXaOBjLrlGhgdZc/Fdbrg0Xyx87Y7L1mBEoAthkhOj5cfxm/cN3sL9Mcn2FyWI7S2XZzICkJcg
IGVmnQzh9qMXTarN6h+bsPgImThAswldkneEZDeWw4sudV+7o2fF5Udnn8LB4O5nk9CZUjTNueyu
6ZaW1PE0qvgVUSiSmVpVoHofzLNWlVXqdwoTuARIa8t+KMTBk25/xNI2cOLsF9OQ5BW40c0/S+9H
9eCnx9xioeWnsDpS4Xt8mqrokxRYPBo/XxIVigB7cg9W5CS6RSpVT+ytzGKoMnWjzfGMCSuu/k9e
QAG5kC/OVq7Sd2hitfPe45IfsIHFzFuLxr1gr2RBuXhP283p/u5ocV/RY8dg+ZvAm1cWj1ndbnO5
UpvLcTebkOkR3xnWMNUHiBhB61vP0RgGQMXWlmZ+3ZJc6ZyXAC1DpS7/N5eL+ZoJucxzwz8GhEWU
0y8Z7BPrg1RpXySx4+E6R0I5hHxPY7PmDnWj+xdu8QMN6I/4qo/2fQy04Cp9VIBgoUHXeDTPzT0x
7vnJPyZlC8aOfcvbzwMABEaNHgOLnTUcP2AWYCJ1zERx/mK1ximeexIeawXVADLESWkyqvMhMDgT
A09D9MOC+Qf5ti7UQ4G5zv/SJmdD6wAG5cjgRrLqPLD/y6h5h78bZGtaqN3h574xS8QIMc4Frgu5
McGPxNhD6Thnvhv6dzIZkTq5ksrjzxItTIOKqJpHJsEdPee87cOPELqIML4XtqYQhWC118kAbtuU
uwA5gTMfp6HIcyAn7ihLvqHIjdVwMn2rFRQd1s2LuCjRZqAVpATJ82o+gEKbFgLQoKWkbwuEVTmb
BskrzRkoxQumupeqBWUVwDd8Flvb6G+4xajRnW+x5owBi6DSY5MCajUcdO0jiIBGPYAGGmzz3SVH
ubnwnAQPoIrmczr/XfNCSK8USSYFMacCUT/02yMJBtDx54O4VfoM29YI88y0IQNuHNOlg2oStMLk
FASkvUIV5OcjzcVnoFourOJvg7mRrlnjsD5iCk36P4gZr8UjqWoGg1jguSef/Yqi5T1mKLri56/J
DpWvWx7/qbIfyiXAVrHte9n8g300rsLNlc70urRHBbq5z4smP4NA45CerBca6lzG653IR0iqjbJw
3s/7YfSd1lCLKRSpHPwEO5ANLS27NYbEQ9Rh35tSwBpERFUgVufyQttSM8/cWL3aOCif1PxI+t42
qbKo9DCnPlisMGDD5IohUe4c8udgjpVXkEF2Sf3SZR6S4mm1RbJKMfjvYY2eSVviA1jTu262wuby
7ZojpzouTQrX8yXgdcQQZNYPOJ921NPEDjd2KGDJtvXevEVQjunO8aqDTjXF2RxFCIFp6t3UT3J+
zmzHjki2U01rvwM8SgC2NgbJ9ePSMb5FHb95e1+uDwG6Ie7TOnfv7q/Fgeq8SdaLb0mQHc9Qzw4y
lD0eNfArDg==
`protect end_protected
