-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
1hjwzOmAACX56mZRafyXBXC0wbY5gdp4rK9Fn0vsPwnV9r7Te1Fhm8SrCYQb0fXveeVzgQ7UQHN8
+iXaUtO1jPtPfv2gXQdvCVbkrKBxjNxiPRamT3iQKwapCMDf2Jsf3lT6fsrR2PDEMWau2PKkPn+w
/8c7bHOZLiwAbBfquIkBlvs29c/2LdWtOO3yQLiE7+FF7M3dRzRG0/350iX7Cu9uxueZ8WRttJUw
CWvooN3N4I7KRYGdTYiRU4TdeKw5cHjjqV6iLxi8JUoYS/at02kWljfldQt9nsi/mAS1+JYl9a2i
UpDgMMuEjM6mwHRApWqR7uA1bM7ndyZlEpgZYA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13056)
`protect data_block
6uJGEaZDuzECDkcgcI/WpbmLGFLSQISWLFo8+WjlxlkEZQchT/Mb8gKKq5Z5pyAcIVCLQzkMSSvc
0Dr0iOf98WRcVdBjQ4PHd3k389kEoB51OquGJ/ZSheJqZxTNcCaJkiPnmKQuiGWqDnEiT9mByP4d
IlXkbjO5Xi/V0gf+gSeeNQYaort/xM/0vBytQl+9RVsGf6+cGpFXvj5VD5LvYLKt177xbtHTV24k
PlrK3plHDnJKlEEg8NP68u00hlPFpdBB6dwaxsjHURGT0jFhtYAM5UEBun9DxVQqj32f8pP0IY/W
LB4dGt8BXpy8v4u7mT/o+w1HWOI5+hCq5NoGY7kEXHFwjzE+xSFr/0ePKum4/NLKaBftZ7CyAmyY
4GVAoy/gwwqYNrre1P/sicdbznCFLapIke73sp81zIa2fJbXcpm9SpaWt5tJQJtYICLUcVYuIPQa
hwjEnU1e606QzrutgqfiUrHvcC7BSdFhqNf/awesAvl8S8cF2pSGST3erVz10yWIUmMU91q3QqWF
ORYlESFyJ7SAkqGeUEiVE93BWQhAno0nbdgTN418jVkB+QW4olBSPxJc45h32SiKbsvdcAqXUQQI
5L8O/RzxHIv6oa/ksl4RDLIP+qh6R/vCycMokJhnQGIwEpsQV0bp29wuQuxkR0tdmLCqiUvy5CTz
ninGbJ0hKGB8DEXrlkmsrux5mnJ7AfCGHUPWQGdkUW6QXh0O6Q3GRGuOWgdMu3Jt5hb/QtYhyOb2
PXStfh3FHV7BzUYYyFYBYvo0dlpfDTLr90oJxIjx8glz0wAYqytmsZcMt6VQNKvjIVmCRcIwai2e
0rDNRNVlAZJE6LS200ITIEKSdAqi39phCQDgqSRpwVPO4SQHpH7WE9ogpxCkmOYJCEVdwfeS+sZF
y6ifpHmirz7Jc+HjTgs1uMDSiD6xoWUPlN16eRPrmrk3dfxtg4wAuVLlySAqyPOHIiqQWYjdv387
XxwHARPMsA5uci72tUpFRWu4qfcW+zNUk/3nFN0CEedroXeJaMY04ZNQ6tDKwU/9Ix/cjZ89noBz
60YFj8wPv7Ns1/n56WBMOlBNqrODrJQSCxAGEIdRQfDOPn375a6IXjK1q5t04rWmC+2YmOoLFCCa
Djffrk8KPKXnhNw5K2kBCrqBgMg4pnX4M0XWrJ3Fw37G/4oLZI+g1kCNGwzwUvcChK7QYeJy454d
5lO8faYX6VzV61MJE1wq/DxE3c0OUR/ntC9XAQ0/2A448RLbDsIdxOm2Ids1nmF15lGgHrC0lQ0I
uZqKS/9cM55l2ewYvKGixgOuyRjbmuMvyWGnnzCsATtNXoldkvv/y7P+5yWaapntKTjzkNRB+rDZ
64FOB0irmBF0eALuyAjbLjaviIq226FBfyZ7mdYSEt1/N9YXJYKOy43KK7l/138viIzCPqp171H+
/hTXcsQNk/Q+z97yr0h10ppnjyaDI6zInFvIy1SiR6EgVuS1qJiKB7jezd9umFA/niyC/VICCbFf
VZ9/IbgXUL5S+/YWUPvR53aNxyejLMJTjXA4J2Ktjt6u9s98CRCbHNZHsIVXC3aTp4N+0braymfP
18fhJpi7pSyGaczT8AjaYf2tE/2PY/MEl7F2L9YYxZNNK86fxN+b9LPYxEOrMvCCOKJNhSUjLZag
tuZEF/uz74MZN4ym9AnrkP10x6lBxxANS7TU1wrweFb1jve1c5AXrgXeEC2ovqExfpiZp0SbCAcD
Ii+X2T0l4JQpg+5dSO00cTlV4OhohHT+u8jUQCT1UYDixojRBkYTBrf9AEUdf61ddaY2yTP6j0t3
52oItBPZZHnJ8bKpZ+shGsZv816hKqIBjCfHUEeYGzo0+EvKpHpeowiDXA5T/p+VwrMGpVU2KsLm
gDJChQvN/QN+KHptMwLcX0Nt3gIb8s3tQQ8lodT4Hj0b3I8QcrR/taysZIPdDirwTYokwMIjFhGR
CNuFKgtyyUlnE3fc1nsWTXB+wpSoo2dCsPvj8SjWtMu6OwBMaCUugXpfK4L1RqT0ufD9yvkjaq1q
GL4MOMc6F1if+/7EsZr4q68wDKz1RKF1wEZ9ssAV4iG4GhIXkFstI179hNbmy1AzD18ge9cMGEMo
XReN4iXIqQL3WRdy5u4Isnejm5mKIP4ABNPLfmUY6T/Rmv5fCUsCslBcGVedvPiCHbEoV9kmC62h
Q055H/leSqNkrKAuY/TCm2suoQ1HcmVaaQEZJ5y30yk6CCTbOdslHSowPA1x9OckNedOS8ONXjuH
FG9mpCC+ZuRNYtLtMp50TF+udVgfeaWb/33SVthcQPj0zq+97zxEYGWpAbJ6R6cRzWVErtIJSJvu
E+GNiHfCzHff+JKs+9w3MjR/PGYyRb+XS9PfYxYzh1atxOtpEJ+Rk8g9pHq+W3oIaU7cT3j9Nyk7
O431TpJUXZOkwa7V5VkIkE1TeIygVyYxyRLKNyWHOKFBXbHrWNsXNN3dsH6raE3HwBoVOmJkhVii
/mlVDhMIeML+845RW5XN9xm//8vTSUz1dXoHvqYnjL84AiNQx7Czbnbpewqg3hBN+K/dLRDd7G8j
zw5+tgRlinxV+KV8usi89EVGv54f0QmF38IhojJWlH86bPV9xPoTNmu1Z74FbgG21/aTpvksDPdK
arVRkhBt21bRgY70o9me2QcMt0Nll7UdSBC98NPaO0C0HC6wNExrk54n79P0rRHMoF/0mHLHgpnC
UQfysTrfZKzUpJRKURLw68PQjZnUIzSZKLzyKOe7V83aR5VcqNqh6BbE3TY/xCGWn5shj8EWl9dR
5Esvm/ui8yY85BoPhMYG/Vty/8vRPyaEXSJ22GKTVaaLE3CD0fOc/PsxVT0SabR8vWdzeZY+dbkJ
FMDbT2MOnE1/kc+ED2i/5lJPtagp4IcrVOHQsoECHDGgALu09XOXbUfggDxLNC9DggzPtMPgLHog
07B0CvLi++ga8fI83G5NyEeHv1jtzMy1VvjYeWOzcEokZ4v4+jWPOX0gd+t8T0nGan3+pBPD2nY3
9Gg154klthzTLak7fmzmQW8XQfvUMuX6jCTGWeyy8KWLzzmHgGvTLHSfpwMIJ6mfDJY3NFNbnqOq
0gfkJ4A3prY0d+S/JMpWRDj4r/g8rEupO6VV8PD4xzjXxDY6T0h8dwmWIqptOZj8Rht0SBGNzgUL
8thLkRjUwKbLxqI8w84KoPWATcLBxX3PfMFhEgGidqjo0p8hhCjECoYDO3McsC2HjCDT4w08n1km
3Wel6ijYsDsmtksc43RWdFt+1EqEmLTc3s/74686jtwSgKj+59WnmSNCNh77hHCR0DI+/8I2QBq6
1xUp5m7qI+901Al9fruMCzI80Gcdsc5rowUMN/DZ2lyuspL5YNdC4YN9koMJaUL4YjYM+x/vD8mK
WtkTuYbQKOWaD3sdPIBirbL/UCSuwMvaj5ED9TfSgPC6D9idboe0rf850qLBIrce72SjwjMjMA0S
KDQUJPGo4Vs/FxEpmnSDUWQK8xL2f7PzcUzSrOMXNfByo7PiNZcfcrVTV49tPo8N/EHnyUHOugGF
ySbU8osR9mQH/w7fCPuDeRVbhmIdTIlo6W5PUuYZH+3QPIhiN9I0D50fhQXCVPTQz3y5cuS64zVD
5BDQgAQcIOamIgzJOfKp/9HIyolT+att96Soxq29CPuA+H2czYjq97RL9KDsLbzpbJL0OEQWmq1o
g4xadgwMZvTqyiDfSChcTU/TaB9bHcsGSAuZQEepmMoi/TSnTJfV5BuCYFRM6Ms3D4g9Ezzp1Uzv
q8bWpKZlg9pEaNl0oim91DCyH57xg349lBWHU/cbwSpabwH9agMtGMFqROVlS38+m9ifdmxoRMu/
5Ze4ryt1nlD8mAsiAgkOduo1tuSBrb8cM9kwuGX7M9i/+m92IHIJDcJMOg4DWh7xjLu4B85xZOey
x1bH9rfZGL9JlNkuW9MwV3DXKmorL7861z9tCW4gmvex0mgOT5d9FACDefmTBt/KD6bRZszzRtHC
Bb4ckmd5YBXpkTVObtM13aYjkKoNjBC+bcApIMSuF8bADJuJd7HP1TihZ1eK2CaJIA58uRDSrXXe
jZKNgpZDEWl4Un54PYOURJl5Z1nxV+CctKpKCu7EvxDQrMku5vqOeOrcWDiZcZYZUxdqNI+UX0+d
csL3KglvyYca9x2DO/Sqga0691z3NXSlaHlB2DuqHx2UPQfIdH19fZNdPnw1IhQDvcdDoo5J/rsR
ISFhxmuFuNJkBvNvSg6ojZQPiE56keVe8LgTSkIkPWt6gCjeRY3pkNrQyW0u3nbUnvxSRG1+fsKz
UUYy8OmC6c/4bAg7pBo+oxobDDUZtmBZKl/tcE38UnN/altUp9po9KvQJ4Lnwa44+RF1Or7zv6It
bBEM+7Hz8FRStI+uwql9NWU/FZOLFtZK7XWzKW848e6hTVRocF9DiM0qSI3NWBhGyBKqwgUFTMdL
DEpwKJ07TKJ92at0duPLQB1W49UoTgPAO/xGijb30zzP/kR8n9QCi+XMWGxUnzLS7FLilKMaZfDm
woWl3WcqU9r1Uog79HtwH9QsxoBbJHPobU67fyXjsBkQErGfdCwA1WzIkofG9Vu08pLghV35kBsb
T0jria10ZuadD+l5xISeTmh51BJdLtGzq3McDy1liYMHaVIrLRJcNFG1CnPl06uIL0ZbV7B8ZLUq
dydfHgl14Wp0mMgkkyIirdoJ+DHh2MJTMHpmisaygmylucZJxXrywL4zP4x8o8zycBc4Czkr/+xe
Z5jVh7HxF9gUEwX1a3OaehW4tNLKa7q/h0anjwMUxIAfVUH5WB5DkJ3Zre/iulWL7kRLa/2AK6cF
f8snhqRtM7hZoAIjW0/8oibwDmjtfvpnEyvmaQvWe3j8UjtDxMHuk9iwKaQs73H8UkQtQCmw9MLd
wivhJM/UxyazFK99zqql9nQSsV9AkgMTPF5+Ip/1YxdbqA+/+GNFt9IpfqkIJ1iXyYVZ3hgKtJJU
eEydkN7R1uWvrZQNMrnXiwWxClnDwH8UGKJVajkBDTvYLVpbasvzLmNekPhQ6NFN/Xf16MtheEDy
oHEsczpQAJgeebnHGOV7Nogydl5roJ7tjzhE7iS4dtKIcjo7Au/Ays4N2TEvOm+wJqg81naUFBKP
H6Ula0TM4VLaffyb4vw+5Bi5dxMUnLF1+w8vu9E90rmALZkQ6yI2+c8Fdfzsl6xWLd3HCRFBOh5S
AopHZ74wx77fSVi6Fb3wBjfFObBjTUG7scUZaK0U/O4RfR5+AM6mt+zBfd4KgdasTwCGkGmfdf6O
lEAb0oh7TOKrczwQLaW4J6xNRyCbzA+wkJ0HnEhqiFE1g6aNMoSRfO7FWhbo1//OoZrzXFJvpFLg
bPFDTDR5fB5ND6qMmROezGPL3EQ60drpL19KEJ2AT3Sl4hTUaJA6hAXG+VZUENl1CNeYOtErOOcr
W0i2zT1maj9kHg+9JnZ64yCOrCMksU+QdG7wdoqNy9B5OLDJl5tuAfBoEw9Bmwsl2i2WBPJ+HTc4
+78EZWTuG5hxk+nwO95l/3snRiLx1YaM2Zcg3SLC59g+eMfl971VliVaRYqmc08P4jFUI/9kl53k
I73SAmAwB4l0oDZrl29KfZO/1JF7GMKzLfaYn3j56BKYi+GYwf8iiUF/Gyf6IVnyDhsqEPVn5xwf
qd0hwk51ps16ZFudDxAx/1wCSpuTDA8XHaXhynijq7n9nzJnUX4DkD/Ln7I+xRtCkGICRVT9W/a0
r/6u+x3Msbd4kX6gpPDbittvbboT50V4kydDzAGf1X9QjdbzOlH++dHKmz1PrbZm8KvEXV9WARv0
iZ1Jb2xuwudq50sLH5/V/JpHbcC0dPo+0mBR7Y6dVtiCfpD/KzTJJwJ254xUAAnToUkyu8lFydHc
bbbtUYhfyMkSpm9DclQYzQUtQc2DFQ57J+xNyOW/dH3GocKvE/yKcDTEtQOJ06e2AgCgk3rhrgjy
HvEC6bMiACKWNCRFca0CS7YDdwi6nItMkR6N8I4En66LYqGQtExft4YxB3dOJMmExHknVkWzI1FE
GZSX6lYQDxSV1VZJalXvRqCScZHMHnjS1D0PzbnBz9//KjrTOK4D1QYPlCpWW9W9StULHjgWiQ2c
jFwp7c+yi941tHpkDQ/CLTvWVRStpb7Jei+76aYHJf3KobXSaSUqIB9xe+h9r9LlffHNMVpTlxwa
sYzpwdDwCQDzhq8wLtXeqkSDSQkFG7VGeunkFunVuIA5CQGDcvYFshipUujg52egTpIlCnJS37bI
uvzYpfSeGr4ozPOgC3433jS86FPzoMQLjDTwzOgENuqip+g5g8SnlVqzofRRtrHreXVu8unXLcTg
IT4acndjY8qUW4ktjE9Gbv1/CdzOrGk1OY1yzdageYQW39VD1h5BISzp3nA29tvdZ7vYZ/zYpkLI
ziM7ecu21JAybNcnB9dVP9+bStf+gzr/YEj83wBdFyuta2dUgx0J5cF0Kyr0Kn4vW9hFRLbsgQJp
TfqwbiDWCHnlS0L0wZPhJwRn104RmT3rGXJ6c9BZ1N38mY8afZjJ9WDN5tYGiAEKG44e5c4PksEr
sblA/1f5zlrU21/nuJ1l+Ik5abaXIHQVCgVsNZreQ/YxDhOj9kzDGRzo/M2n861w7qGTjWlqipJP
acSJwXMDEW9DsFRoYwjoN0JHTJIX7+BURc6otRYKmmfOoXo7Q1i/QeNAwynVc/FHkdx3T97R3Xdy
aGhl9OY755XWQqbKJFdSLoWxW5KSzAC1wzHOLrNdxOWEOYgDMD5H6Nvg9WDAMC1Oa8GtMivRDT9G
BX15EU0OOOorW1RgVt8GBUx/Cl/6kvQFdttCCUcmrF0DpgSbYj3JLr2Tro7Ig84DZ/xzGstPfsNf
+2QE6NGRAu23IQVQXV5D3fG3hZ5ocRAhv1jQjHwxwwMhTCfrfmeSFEiooNPs8XcvzuInH6bGMoC1
NNhy4qqcH1cejaAxa8AVURDpTSrYbtozHTYqFOKnhvoFxCBkvWtWTTwfF1SaXMziaebAUa+ofG1U
sb6+LdBJ25UjDHhNOB01TEeZeC5jN2pjFM47LPM8Av+jmJSBg0zzEGdD6pH8JJc3+d0lhlfcSwGC
23R7Xzp6LU/lN0LshrzEf+XMK98bX4hGXQ7j/yxFD05IRF42FhHFrUXPG4LXKYvKCHE9chjO3faw
hTbmmF2zW969fiOhaKGHwB3UFkz1gPcdVO7zG7pOTeucBfDnrh5/zKzEan36X2uzO4CVIJsGzJqo
cgza/DXB9B8lujWWaEUdLkeog9RfQ4ClzjOBgMHZC9/LSsSxFoS4cwx4mCvFQXhHfciyyZ4MOdGu
KAe3NK6p7Ny0aZiQCPGvuJFn5NZs3dKFvaXOJnjR37afF+flithcDRk/G5d4AcvBeF4eoaTzVd8d
5RjzMv7sW13UjPndJ3JNsdorZ8zB1kFDpAjdsXmgpVeJYyKV1MB19b32Du3wnmAB8P7qyc0o4TvK
QeIiY82RW0nI+I61eXL4bAyXJwcfJIkUsZ46Qs9Is+YiD9lFui2UG0EDQ4EqRLItFjBwzJZBjhjS
WsYZ51GitEXmULxsHZWrez5LySSHZgR88uNWaVXmaZ+w54CvZJWCIY+V2j844ZL6hJQ79oI4aynS
BvGDidBDnbHrK8tM7vFU5Yrm9X8wQsHubfYIUKYy1Zn79cjTZ1/jqR9HbFQ1crxxCibRqEEm71gg
jyH/Oq/AUFnOP3JX17cSwJNK6BtoJfsCWVKjpKTdvs8gmPwzUhsbBH+IwsFIEXmEmnYjNNB9cn1b
TbcDcDW5xOGEvrJt2zbQ+fnMpCRZdXMBTXrMHOnpsbxy07vmxfpOsithsMrby536sKnm+J0oiS2e
3ejBH4WfSsWcDKf6XbbzVlMYvK5h1pX3X6V4HUVy3t6tB0CGCj5Ao9bwTl0hxq7gtBLOV2TaT26n
qlvb6DxQY8o0BySgaHV+xtO2e10EURz2rvfv8J9yJx7j2mA8M4ywqq+I8DjmAuwbqfAVV5Uprlsc
/pHo+nUEYV49vkCTAK/Dj1jb+O9mJtLVIoKiM0iTgDET4Mi+oP/0kbK8jPcAXBLv6gaz+uwLUUoq
61KNybefB1Ghx5PbvZSfRixesIRDm2Nr6zcetTI/Dlg08gqJmH8d8wdk76enryGpDjjqZRyDKWxC
4BJnpIulkAnlAqt0sE1vckscfKjK+llFCLJBaNQ3iTJhelCoOKcnQoKZfftjxa4Y4mSZ1x9Kw0bc
6SahEwQd78ncNOmsFOMjyE5EzigpBEEMRBE+8ZD6TNi1ubMvbaQEFHTKR1VJpPsadQEPIUaruywd
p4O59zpJFaheix4hNSbpIhh26X8GYqvxWMHjdHsEfViK1x+Nh5YTShNm15nPUhmfghSc0CQ6sxKE
jOlrL15+GLzXw37bdQzPYh4pKq0Rq/+iRnyQBtyVmSZBZxYk8eNbzAk9sGOz160nkqZafeAHzzr0
940aQ3cnS944Es/UO8Vs3VS9HlR5mNugcmKEGo40Yo48nG2jSeSE6XCNKKPJJ2/07KBEwoDEf+87
F24r7q+wXZy4i+G2JwoYRL8mbjvlx/IfvYjMTdPX1NzMuKSFG9NzimPafL4o581r43yML7RCAG6n
ff7Imv1igTwNFgQJstnOExKczzcXz5X36VB25T8xLEl8p1ykuQlmvu6QxSccLxCoi8hwoz9H5G1A
ysLTe6MjVVmneHwoHmU5XQNMf0Gvzl/G9jCDICXt0RexR2vspFWoErCmpbYZ6mmdmKKAdbAFqWcS
/B0uV00DKJhq1DiRTSWkDrShm4TSXV7azxUNgq3oj//UfYlyp9TysvA6nP1cI9sw6PSMw3eYoT00
7D9C5YuboaP0wRpIc3idaaelZWOmYnkAC18xdic/0pV0jYB94hkYXCu26Fn/lsjM/RY19M0V5tyr
yMONrDA0chYYExKywPYJZAJeGKmS4Qbslfod4C7tZpDjG1qO7zPhxB4oDKSOrflc/nt+s4xR5sfU
6VNcxGBgroz8zUfnQSs6PM/+eInVXE8iqrIRIRnlprH+eCW35n4XuoPi2LtCa9ipdxPhnJ9JUE9R
2hoQwmooYdyrCEL6RFanHlzSroTXtLTe8/0iahpKaYELaNT5sjI3euDd/Y9qeo69OEJNCuksDcTV
zzmO86uw/m1WrthUVJ9BbIdLfBLV8m7dg/IF9TWoK3i6YuqMJG7GXk/PgbUXV+XKBBrE3MdxhhKD
t2vIgylCXebNagwZ0uB3vAb25AvgtXVwud8+hBDENPtmQlhHHpNGM7jnrpX57giFJBAlBFX69EJ6
32HAtThMaRqwn/thdeXdvCjFVoyl9v8SdmqPc3vuAV9KxwAofOGMLo40WmZwoqxuoHn9B1/ZEUvB
Ct7eXx93HPMgDOfo+ZN1XNd+vSfrcl0TscpHeaiKzAY5d4paAEJ4BM2PKsHpxk47jNRarL2AyVYY
Mx6BEReWwNcNYKW3RMlz40QVP8Ilm8xIfvbRHW0KN9dYg0032FZSqnyJB4J8r8njshm2s2Hf/KYr
VVhBq+bpjx8citPB6mcubLJTs8UbMTKgY3FliGZsUqQ1ZQzywY3spDVe7xpYzo85rb5GAgRv0Fpf
vzGYSaK1damQLEKG/Y2Z1hGGXJlLEaL5vXZjiSRoIE5RUZqjeuvox+nO0HrV5g78+5Hp5jHLMdHO
Vn/KwF5RUwusAy0fcTd69JWulHJzgbr6Nj1Sfqzu5AHEEfRN7rQM1o+I1ymdGRh3Vqh2yZmUmb64
bW7hO3mJ0CYrudMXEQ0voo4DAhEnsdVpIzZEtdwkoepQHNTLdVQlESvSwV5Jk1nPxFrv4qEFXihT
AtLTyoVwVzMEBBD9Chob6a91uYRilbYC94NXWQoT+7dVnOa4YOfysE6Aa5FZ3DVkbrKBYM2rL0R1
5VaRTwmFFACRSYZa4ADNKnT5YQGoP5OGFGGnE1PGxmbcL/hssayDWs/VSKe1FhL+y93ZojYZDJIb
DR8S4cxMpRcrfoJdWECR3c4UIUm5htq6LwbJWclBIZz1Cf469MwPZ5wyTcOLAYHGex45LyAfBzKH
mzTRN0wVsOa3tnvIu4NmEwZAqAQRnqu3fx5SbSZpcB39LMDP/0niTk4+fWHOWOnxCixIFdFKrBSD
43Fn4F0w1MeMHQf8zqbdySiX7zBDpFPkOLsqTlcYrpWa8Nzv9VO2et8r+U02xHR14dvcqk1RSqXy
NVervwl8+TotwVVH/0wHLww/4wP1Mw4fsxCjNDnw9xCDQuEhEmidazwIOYgZxEZBZVhr/1PUmJMW
KlHxRzHtGRLhtKsw6AvBUo4xCZD6C6NSBbERWuR0q43GVf8zUIdF2nI6GgyelN9VoY8iTFf4BPrH
GuQbooRmDLq0bvzMjcXqY+a4mwh/W4mAGWG51LcG6P9iFnqo8+NsiPe1mTlDfrr3BXp8gmUU5TB/
IfNLVl4uygPgsmvVqEFnB8FSXOlyas2ewQm4Ay4fALuHsVpOdhABUPvvmoSbNVks9zklXvh+J67S
dsKHh6yQsoJc19WWY4O2l7pVeeOleEIO71DdhnHExe/PY713yAun/AZTxdz1Wtx6jJZ5eCxcmjx2
XSBrv/cNe+3Jpw1qIXNBw4H41mH1FWFQa/J5jZIsphvrhjWDyvNeUwiYFwynISAsit2MrynwIEDR
8EWpIkrvmWCY9+8BQ6PCCXhYby1bWOKHOBkG8fahRbwsfIrTJpkwtlnAtNj8Ez+4QHI8odwSpdx7
lLBchJgsjnOeRZ5KgskL6J8683u51G1vfSmS7ZQ9QPSBibAf+LGdzvDuKC/+50dfzid5crrC3YX3
uyvlzsJeic90ccALBk1sgkCwrFk1/2Yc5ky5VHd8UE2UwMtYdrtZWmBDtoTqVtgkgNTL9lQBPYq8
54a0md6uMl4+TU/KTmVAyquwLJi/Hl1dJjsBmG8M0FOLivrcRm3lzbam8dCjKmR8NlYGkdbsczi2
3i0QQMn8y1uu201EreTZp7RuorhiikHG7LUvU247DeCSjzYjHV5qBvThMpdm4yY3VpEpG9/pzKcy
ZMkvdNniu33030dmPTZLojNJHj4iVunznenIQ5Og1XstQL/JRO7KSUFH9mGwA72huYVZV3DrHPqZ
85p2vy3r3AtkHNrQgxCsvAJm2SbWVXqyNkkA8bidkPJOqlgjfuJxNEQh0ilnXUPRRzRsSezNYVb3
W35GAgirscZIGoHuiX04RqNiV5GGW8QIp7pagEQFduwFwpYv2W6HQ+coWYKHqQOQ4cvNIkKBmJ0D
1RCeOtKw0SJ2p9uKxuy5jtyzugbAmFGWN4j8oeOX+l3C2SL/LbHXGM+CbIczuPHom9qVZ8bHOdXI
ss5jHc+Q6KcZnSXNJaj3xfsO1Yv+6W8E3uidY5Zlz/jNhQhd3UGXjObEvDcX1KfQNoxmbGpVP/fs
WlabhlLzBmDyn53j5Za5UYWDrlrfWtvS1IwgppnfaNH1ViceO6ktj1u6rinL35gZLzqbEfVMmu/k
Y+kThUSRht4aF/936+gg6tIZ4+CFitN77Hij7IEwOL16fULBZ3/tbIk6U+rJr0/kWgtmX1aKS08S
igeBg17dw+4cTyqmVL3T2BXqHt8NU9fXibapsJk6JfQgmP9aRwVOdZRdf0ZuIOXFBoeI3LJnd+nr
JPFu58JRQfq4HlKtC3fiE3fvlb5VNudhPg6CBBTYrGLY5Vgt62Q2p79OcnoV7i6mUoxtNcHznlXm
ZAfRskA5YORGRqvk7x+60ZxT4PRv4CScXDhuo7Ck/6E6/G3XZXALb2J2gED2c2/j6VkTyW0/LHok
dq5ykaNa4Pq5T239eEUqZu+7rNuRq7NMFKHCbxJ13AjntRV6GSnRCNUsoa6sDYpvxyna7OQzCSrt
MLoAULaW3STU3mlz/eiqYLy4T59KIqo3/62NZFr18jqGovEcRNabQdDvcmtdA07tIHSEvevx9CYO
Fs/f62MNO08VKkeaJAD7Gh6JxajXaVN1e+s3zcA/zmVB393pua1vbMxx0ir2fosV0CWgWJEm4CbS
of9TV1X42Qk7QsQDMZod68mzwLqK6jprd+KbP4H8TwshMznQ2Tm8z3Fa6hdaBFAP1F3vKeaWdtXa
HDlxEHUB9CQ/HDwOhYNNOQ5bBcXdwVPuTHgAq2fKIVma6QfVEuutI1E8DfvmhTW8wBbw4uZlbc+M
/x91o7rd1itmFQwJIhJQUg4N+FM6nksCiY96dC/cMifhcSHZ0vrRuNdNPQNHveb0u8bkHYmm0Upf
TeifO1XBZWBVox73C1IyeuqpGdMQ4HXvC7dYjP3SIKxwfWN+yPQI3d3KEx1/phkpd9FQKl/U89CF
anScAFIF+IStZ4rD4OxqAqaaBzMqQ5EPXBxtQXjLS4eNTiOSBns3zOmcJMK1mV+1WhXZ1G2o4eh8
EgRufhAcHyI3jj46HjMEytWRN0RHPhyv0sgHIZMMUf49x1EBE+cbEGYAPEW2/BouxUSWKN+ZNo4M
3pT6JM9psdajt5TATKd8fHM57MLp989+AxvENgaJauL8mEDzwkWk/n7Fmpj6MT49iMLsOXmC5NBw
yfE4MKiqviCN/L6G5juBzQJ0na6uipRRcWkALatqbPSyykSo6dyvX863ZxQ53wHFrO/+oPYustVZ
aVjYh4oQE8S+Qj9KePDRghWoLwabQ83y/V/H/ALFvacakzj7WqkA4IBkfHUE+23F0ASrpjbKGFIl
hZSvGILJ4YLHEaKzpnXj0Ggu7+OJJees4kTnsNanf3ui5rYfIqGRoxn3bpLlGUPy9TLldGb0YkM7
aOX8IIoGGlPYIWcziSZu6jQvSnsk41fHyR36ifRN6syHSvPCQMdZPiQXJqWWfFHvd/HbpH+74wwS
uv5rh6A1Ua1CKHza3LQ8EbADBPOg4BApOG4WOYmV3r3l9H+zD4LQsXggH94R1ei9ntU28IH985FN
nmrJcEi3SqquqtjurRPTGa5zuhv+L3Wd6BVMmuehrqp8jWvm6VW+grkq8b0SdrSFSfdEDiiqX8WD
FcqiYua+ftxKOpP1JKN5XWCUUPXWgYnN4z3b4SgdWwbSLbhyRrK4JCbqZfRIpJ50TU1IfpK5a1hn
vROXdO1CLYu+MTulF1arGCRLyne0T8+KP/mYsK5rgL4i9wiLMxUlkkQ0fUzRfQVvyOyaHoe9CnkE
m6WhjzSp9DMKkBfLnT7CPUbZWA5S+HsolRg4/CovKS9qoXfi6wHfNmCdTCO3c1kQ/qvkXlmkr4uJ
CofxNgnVQa1BZsNjlUvGoBHY39U1aj0Sd8jRU5DgQJYoKlxRB0+DEPCBx35Z0jBynKYA0Tp06/bI
Hl0xk+6y9qz6L8xlL6OKUlNvg3qXRmEGQJ6dek+DtOAvBPO7mIxuB62H/0ea1guA2AtW8khKohF5
1hRuCxYEqHjOf3oYXBFcY6t69/+hfoWVKft0nCwjusD2EAEkvJo1xrFP2rX2fcWiwqtJLXRSrtsw
IfL+H4G+JYgccbKAfrvrNSrLU084K0YBHZd9/8JAg0TEe44Ety/eDbgvt3OFwlWhnZSupBejoiTW
0lcvazMs5pRJSsLcNL8H3LHAMuiCJUT6p6gdLTfQCEGcCLiHm8AV5+pEJkyDAO2T3+FI6hhYKlQk
d64nvVM0rHyv7RKzuzQyQVS7IAnfuD8kVNu5qhkQuxLQc99SPNcCM5dEYz8yxJmhXTBm2ASpaXU1
HT2Ll3bz70PbURLrQSmVdG8HbWOHNRcNashQenxMXmxZCOP4Gb1Q+Yhkn5kfjWKotnVdHW4DBtbJ
X1hhTZ8wiwMWCI/zehvCuuRkdy+aAUOeWcxB6z4oe6OB7c0QWFuZ1T9avSwe6e6olhusoFiQanYE
HZh1uhRY9BfSW8uWtNc0Hz2xov3cNQoKmvxXRPOVfyTKjgJJh5h8NvowuNL7VGa8KGF5/s5SiO7x
SHk1klLVuYTcA6e9NVFsX4ltSup9ty1sWxJKWC8D8wmQrciaFIvLgz+z6RcSdAzRwN756L99mMRw
NrdQnO2B2fA0/6K7WzatJ4vzdUHiLV9hMh7XkFxmSRSKuHeJaA2uCrpLNO7Ssq5pLBO/PmdOFvRV
QMezPRUL++XbASFtT4wdcs8LyBnNRoneIKRz7qkfLuS4iruUPzycwPvBjT4iRR2aUpkDVtQ2CADD
pVuB5l7U8+lyFFvzEwOhVs4fFqcH+29YAxFVd3ihmw8Vfh1gE8LbidVxfuvHhbeuBQK0hYFb68FR
ZO7meXCO7XnkREgIdadSgjfh/pq8+OBh1l/Z16DyVvvegHhaKlhM9xAkZQd8C8DEQj3gl0/Lstua
/AFVTdWu3FbDoBiPQ4c1dXuSESU7uRDWZsn6QAT5MxITjw9EusUf2qAPjWLmxuoJgo1NiYWnQ2Ea
mSk1AVJ0ed4hjzB8cnqcL2ajbx9VU/oqMQg/kxlw+lm6mlB8ToF5M6VOTLSVVg5BvCThPYVOZbcf
+zD8hqZMt71dBzKOlk0WLPbry6gGm3pXlTUnJ2VX8i2Hozlka0LXkR7OpvCg8bJNhwiJiS2ENlpG
yIa9mBC0Ski4D4uq+OfAewita63ed2xDDKeIEQ5ivvP6w7WqZUlOonR5upd1bM0ryj1V3sqJY2xR
15Oe/xBb9rqpCYlyt1ahMr4k9ENlNH5ys2WJCMQUJYQC+fXnNgcidna6whKWL5WAU0Y3/IH+2JO+
pswElk80eX4WhxwpfT1mZVjek/HpE80rDoskfquCeXjK18IDOGQ9hhmYogg0awQ1cKCW9ZdeuBJ4
sAKE5rCUTPmdMXs+yNGwjH04eTb0Bj/0PSwZwu1+hIhEnRsRgBQuvJtvFb+5W+UNT3dU4G3pOh4z
uYUL2Pbb7skVDtvp8ZTqtmyrNAN/S7SpeCM9yogl+8oqy+coDRg9fDSUqMgPiwQJjcYpy5uw5YIj
kNqEKoFyNIzOl/CWlHrWV84DLhnKPo/cc2Lfqj15ciPw9KaRQhuXr3qbyXfCsqB07QiIMiaDRJJ2
RoI+wSYk4Cx4aRN8r/YOQp1nO31R99izVwJ3v7UsQh/8+k+1KZCQgpeTQMJC+9cPvQTpyEB3IX/6
RA5eya4WnCTNoozzIzgD4Y2DLOMI/Ia5Jfh1eyn8AJRuNHuNJIEf28X2JjM309ent4t6Q6YTk7+g
g+MSUMyOTXnFusNGLcZTC3W/RR2m7qMjogp9ASDQTWEep05pMEAkYsKTr80Mc04cu+kcmyLpUTrX
AIwp+DntOcBOH9HLSvHF2XQ0Ln0xFaWO1b2SNZVUY5pEVWlN17ySPeVdOyvALxeF3kPmiDOKVkjR
GMSKUjgY8rz8cK8t57PDh17AHrbS9sLoFamDsFqT+4n2C/UUT4wkY1E4wD5UAkOzdIeujA6bFSFO
wbOEmc062s8qkOGRrbTZ8IZntgWseYo2huZCArOKMkPNgtdK6LzKGjevQEf1+6xwIS+Tq5ZdP49D
DPsu/LUxcizsjN4sXB3YU/eVMMRHG+h4DCDXzYMuLvaGR3KoGZR6AJjg4rQO2o8M9sXdn7GWfJ8r
usFiecx7o6piPpk415DnlkIGhUwJAQ9ICzziRU6Uk15XlNs/nQ9Nc93Qcg7A2TwT4PPx6+DstDyc
imrkWN+DzcHrQEVV4zObIxh6A+eN0K0WNyCxk8e5Th0xQYNYOS4RQr1OH3Afb7TPPnh9qlO6M8Xp
HYNX5PedKGk4rMNkJgx9ryCMIoH0saVwZTxWf0kA6N08jJgI3W4k9d22rUI7CvtupqNwWLvWsu5C
Q6uyz+T0EGDuhyl2EkSnGZXfF/+pCLLtE1NcrjJHVysBvPBNyPGLHD0zclQf+eyhRaBOwmj6QiVk
EzenT50CLdn/qAsOyxf6YZ6jDTEGF35rDO0OlcOCc1KgeGrmGeU2UKPsSKdP+ul6vVsm/lbmA/iE
4uI683dY24EzCsKQdswGOlhps6c9H9OSOHE+7vQyR5saXkY5Kde9SYZcRB1mzT28A9DIfi8pBvvj
clNj57wTtNjZKsh8oYzR66HLJscS+8K3S+WxiKiuoirivdvtEqzPuaCnPbae08MPxsESL4OVAGaL
k+xc2hRbXCPwYH9tAXmATGh+dPkK3hoSgTHKqCEranF4cxfMJDT+g2U9lVqrcJUgaKkh1sDDe8le
OXuWYgnjy1xWfkpMl62NauRlwP+hLdK4j/sQkrntcxsoghruCpzlI5Vx97k4A7kqomwn3GGuYfws
ge/5KS9644DU/PgOlr/M/9pevnl1+jvMyDxSVUU7cdDC+zHdZFohixT8qdAd7N/5/BkVhoiBAun7
cUrAfJrGvE4r1ztCHjqQAMWhKZVVYuefK66ZUrQd3o0xfRFCL+xNUnSYejhP+I2uNdtSQaFsP7B2
/1cWujYbtrz1JdYq3KRgCRQl02exA5Tvncqx0p8P4gXB+TQrqJ9kXzUmvwZHKPN12soCQJJBAdjK
psCoy8ZBVhw/S30TzwNVNofRqrVrarHZg5lAwTr3p3LemcVdebSJ66pTwMz316GBOrhvyp6vf76Q
AJrwCZmCiIA4q6qwAYQBglll6NgS9HTGujo0yFcgn+RJbur4LItpCYGTFJkEMBIpf+s0map+SJMH
FRV5IvH1fFriY7sP6fQVkeXA6IYysKsXDID4AtOQA/lzy3ouUMp4JVlizM89SeVjTUil6XLYfRRB
RgqAQoSemu8GcOcJm1x4jcCiWpaHW/7Mp/9LcdMbv4YelhAUBxI6lHsVLiNvwxRHQBtwI2pY6zhl
IXj5zXZ/rE+NmbhL80MJDEfZaMzuBr/5hPF3uBtSnVYkakQEx1t/6oU9rmpvaT3YMXsALQk5CklV
3tX8X+ZF/EdJFVNyuSXddGltMaLaVLGMG4CoTXjtEdV+5aPJbUxooYnTWFG7BzQJdj1sIBUrIS87
3o0zi9biGNiqW+nUqCYrKslOTH+q7Qoy2EwnBW3NAQ/KIxclGceaNskgNSyLnoYl3KMxSJrrnrpJ
fZUhvs2PblO9FkjptSIx9aouEzZtxFgJv1/5fAXhFR6ZoOaBVtpbng7QOl+rnpbmWZAG+OFqavSG
rJ1+7pbZcGD8fY8b4fy213j31M5xw9SFBcZs/eG1vSm3qWsQLeRV8VZziz0uY7KAEJJ8YYaWhIf5
xtqodWc4a9O8mayr2K8XUuX7vBuQLHs6PX/MA3bYt9S6+9ylPG0x4Tg/rw+Du7GzrGYGjfPzGlgo
eJky37kWhI03surhfiWG0vo1yQfWe9Q6IGaa7YNR4GWw/pqs4JNSzeW14InN3XSNssgxuFCLsyHP
KF4TN34mwAYxdNVzH7RsQrB3E+ruy9CX69DK2vjlHfUzdyTKMchJ/0NeC6Ucx7wvgJVq4WzTvC2s
vzvK
`protect end_protected
