-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
--pragma protect begin_protected
--pragma protect encrypt_agent="NCPROTECT"
--pragma protect encrypt_agent_info="Encrypted using API"
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
--pragma protect key_method=RSA
--pragma protect key_block
iai5J/kHVByyOy3+5vPvLoZ0LXMBJ/PqMZAJlQV+MVnhf1qQb3baiAifX/VD9iE5
ZBiVQ5G/K5M1Qrj0hxOWeIt5AU9xpm9I/WPVJG2RMiFyyyEI7b43se4JWSQOsCe5
DAfWYdK9F0aHpq6EITop9QQE3BzlVrAnGoY15EBN4kSLgk7emcXkXCmxouWnDJa9
p5iztnSEVC5d5Ia9nuNNy8d/XpO73fDhG/Eufty8zpoFznCKKb1+6dsdiML272sy
39otdFopEZ/iZ7j2PvpC3hhGLG8o0n47oNLz9pYIXrCex2u7UX4zzNHQXVpSwubS
VjD1TEtZU6B/Keof9ygyog==
--pragma protect end_key_block
--pragma protect digest_block
EmAslxSDEyKKpFu20uDPDlywbjg=
--pragma protect end_digest_block
--pragma protect data_block
uLlOu6xW0RmPqIiAnjLAwFgBAgff2FCYuBUvyMiUT+BLpSKv41pvrcoXvbPGi2lC
Ucp3hI/3T1elBu/cXeX3YuKRvFq4cK9XOuaJwJ4yxX1okHxTEBQNxrrHJkjIYsit
TxsKOgJyBv1LCN32o3/dVh2r+56E9c5bEeYP/wxXn4p7u83jP+Wy6cZv+3raA9cY
2eb4teJp6r8ebqW2/3+OsyYwwE3BxeljyAP4IzIN0eVMrcV/T/inV7lKmnbN/B84
zlfYF9nPTdl8Dt3bqT278OI8IYfnFYarh8L02Mqzz2mH7W9TpDdX8+ehW9nb+kFp
7rooNp3OwXElMr4lp6FRkCGuoAiZ7BH0O5OmJNQEiQYhPPInIcBXy5Jb+OBujw2u
jmEpkY3sSZz2/IYRZ3akyPtHTAx7viwNV0ysntG2o4P2M8ed1gEdRaGoUlWPRhqA
6UOO0cNlbE7//aJuz91Gaiy7HZCfvdqbGF7rjHDKK/T08nkT29dQK4dGYIEC7SRl
k+BwSz63yKXTk3b8RuscTdyTKOxou1ptpsu3vvgcLZ2jd1sxLKbShcB9KexM5lDT
di5sV8ClGH8Pvk+RHd7mg1pHXLGjJ2VxHNOJociSL9vz8eGNewyxDxXDxtu60I0c
r84dlrE7s9VOpUeqXhQ2acz/sXksTTdde1aClPZQxcpUoDWWlXghds08IhM9UiQD
vf56/IpufLq7imXVJ1bobqM5YT9LCXnPRsrYDf3eCI/1frhRxrh1RTVEm9s7AdN+
y5mTT1ZCdeWpE1C2e5IAryd88w0Ff6dCh2iNfFsG012MmS8xoiCjMtlXL5Gsinjh
DbANm/od5qwFb5wK7LbjRofxt9DKABtx1rc728ftXZiIx5/F8DJ9HU4HoewDsjWK
de+dnmWo/3sh4hbH75DeIHtd1TB9o9FY8OMiVczT6PReWemxIfiQ+ZHNwmvF0ArD
pm2LMjhZpoFVYlYEB4My4F3i11r6Z14PH3SV+N4MpHkfNYG42o26csPbpsn8FWUR
2o21wIE1V8e6pCRJnfx6cP4pVnTfc0g7PHL2vibiH2eM5U92eSZlDIpSehKsVctp
2R7RT65bSpXaMuPchMZ+WO4cgzp2Kng3w/HKvT4T1twjSMNCtEZ0yxGFS5Y6nv65
31nAUKmAA0aP7vTXVd9pjcWAPPOylOmODXAE4UGd7+nsZrxSmleZkIPyRMbsLwaY
lAGhE6mnfA6iPc3pwWj6KTxMDhhPU5T0wUGEUmX3x34hIAxGugvkbgFzQaU9U+nY
RpTrLQG6mr/z/VpxYmeKhJt6l57bxznM3lCDN+GXdzo4Y4HGxJTo3SMcnNmBjpHC
mQcWjvAHIo2IxDZQkMUiRKuAuJOacr66G+NlKJbfZQ//phV2i+QWFHVJwJ6FY1oZ
h9iiihbY69ArPETig0sUC5jeqlYizK2Q14RqeNE+VG8ne0hXTCYHG57oswCTi31N
/9uPk8ysXJBP1zodaF8xEr/4mW1gR4UddIj2GW9JFrdvvxFEvL98CkTujDPUkOqR
TU4o32McXqd7n7NwR3JPTivj+8mFKwsStrv4HK/PSz24QmG/Hpt34d2zoA2nQL9n
Kr/MqolmfUdX6J0AzIBvCB0nt+hSZCTrfm4T9rvTOZKLdy+u4eDSmmnRcxihiWRW
YcNwhFcQb6EUtsU6IYcIy7dS/cdYtCqaVdjtOIfDvMZVqwAtllmpxZ0Q6m/0IDJD
/TZlAiG2J8lIL8ZLbxray5H7Twpj72hxMknzk5C0qojzb95GjqIDrWDJkk449yU7
RYwcCAadmU8E/yJoowp0gB/IaDf3JuLUztmja6+HHJvkaMMOKyCV5o4vOL0rbcf3
FrhZAO+MSp78VxNRr9lcLLClEfLBOPTGoK4sPWeRt6gH5tn2rGql1OyTGuOFSvS2
lD/dc0emU+Z0iKf5MbyXNFZD74uw7COmUqLOALrjPgQDXoXZ31E64WPPfpPCyVL2
PY+SOiRuhxF2CQJ/D5MQRfUh3slbQqH5Yu8GiU7RFfO/3LrkkHJQ4f1F/xTDBr8F
aijHQjGAfOiZYyG6SnM5+ZesaiNfKPY2HINZaUbtOz4Gf8X3VRr5JcnuHIpFEXmO
gYZ4vO3BaCpEoyVqbxQIsxxn6Yp8lQx6U/scm7GSpHnmcIZ80icNoOYie8y+njGu
mq2Gx83dzvDL0QJnLk+PLok11nb3pD0Dm5d26B5oOIrIp9GxObtAI3OBd/rEMhJk
po6rhxVgneOCY/gpM2tar4dvNbsalCB8RiLSVqjl/+0zmX0Xu2v1C+9U2phcpl8d
RfTM94WXWiiW0RH8GCm92bZRNH/tiEVRzYDaEPJIhsWd7MtAb640cM2KZ0uPkhRr
lVx4mXToL9e8C8+QHECATXQyXcRFrGTJkPayCiakP7Kt8pZyHpdar356EcpQ3GfO
DFx36yGH2K2wqEz2Jtmw2szryZQ792ZWQT/JTlWdFX0Tkp2cgR+G6mx6OvmOG8JF
vy59gPihF6RrszJODqhhpNouw+63YvaG9uiytyIqPHr8FmAFz3YxXrGsQGQAuHHA
D51qzhsY9EtslKyJZRJoNfpNI8LW9KFVpoa3QIja8+xDHY8Uf+mb8l21z9oc94SC
aDWZX5S+qiJ2j9myge8JfA5+qG5P0RC74cZAAmMUqit+kFI+4fp8lJNYCroF0O6e
2LBQjs5x5Qoxbk1pgPT17PChRNacvl8XAr98ZGJeXrLKKfWhxxoR1/uuKjmI27j2
AfX331XA6I/diqIIKlpoGU3pw0g2IBc5KD7Z7AybbbBONuHdWV1fYNAphPgUEbvn
FW9Y+WwrKV3OSqHFXffHS4ggelNaN+hSLdh0suW959DaNFJ6LfFXnL3t6L1oplPp
16y/yYngy6png9b90BZpluSeRE7K8ms7gVeE+nf4L/sy4AaGscGw8W8jDFhFTQtG
kIR7t26OvX+rQebb5cT8UOjYBT+q0VGA8aB0/EJ40bZXw18X9SzO9tmywvQjr7iE
zYYMthzXtAJjPI7HFvAKpAAkufQTm0sdXSluU8+V6l2abkgKnidMUdhk2RcL1LBF
4C5vk4qXxn8Fv1NRoyGjYmOHkws7atbM5J6xyDdwY48DaeMLDJcsDqemRmjuvh9p
aqDF/ib+zWK8BirmkM215B4BMe7gWsmPevYybH/nECbh64KrYeQK8SKwU+L9v3zz
8F9CWEsBBAlw19vnO1Wg+T6xEACId5sQvwlSIBdB2+QCCvop1u7C/Mv3TZXnYcks
4tQmOuxMTsUi9LQbWzFw5lifF9h6KEC85z6JzGFa+OdxSrPF2OZdA6fQe3zL6+E6
RGN0Rdr+//QbqSIqotw/g58iT+V69jjErCoiKqzKmIw2DKv2OShJ4U2DoFSZkPDR
k70R3tavcUwth4Ijg5xC6gaiG6tG8WJ8FJb9cnJNOC2PKCoCi3gJWoJKqWbI2nTn
d6V5LYERzL5XS/WVDbAKVmaMhRNmrR2sYH9fnq2hXUlhkkqLaDzD8+/zBaLFTW8h
zPpH8B1kC/CqfCtsU2mbquwxMKJqlnrIv1fUwteIDldyBd5zCDjTgizBU60k02Nx
IPHACnMoZ3f355AU6L9udrYWb/ureoEtfCbZnAZ5vEBbBq9tuhbrggciEczepIOP
F0AYBpytbdj5C09T1m95CdrkjU505PMfFX/xppafh6Z+lsbffyVmTzLY9XiC/1l7
KzUYCNrnxOf7HXhWwGx+Di+y2eZtSNl1prYME4d1vgrqi3jss260Lnvl/CAWX5d/
YAEelFri8QDKg8WroiWmsJknB4kxxUZLF6YdQWSlWsE5CoDMEdUZ/5lxtebx5JLR
Vf8NAas5dEMDxHA3zW71JAD3K44Hgo8FGwiX+Bt8IM+2E6p/OmdAYjBv95hLRwnv
kDio6JQDKhiIyJS+RyHQdx16EGXe13KZYe1lxtcKxbNHZUpwYnOuUJBEyrC0p8GD
rnuCq8Kt2pUWrBiEoAL2L8THYHY3l7VBhY2kV2qPbHEq3kGCCx+yfZ6yniI4wEF+
/+Ob/ebH+R5r+HMNYK3lsQe6Oiw+WO+AR/k66fCG45LQjhUt7lafEAuOZntSZ3NC
FXQQyH+L2komZcfSMkGV3TCEh+042ge7CVtJiLjJPVTOIHhVsZ/Y/SCrcEi+y95D
DVx3Pad+lIu/AvPXKrg7wc97gllr3G+nRcYGFhlv2XmsnBFpSn6U0G+3qBQQr1Ks
4AkU4x+KMIZ2Iz2dbMoE20qES9iGjM8nmF255BVS7Ie5nSC6+w9u0nJCtblgeg3r
VmUG2oE68FACONKCSdkqsi3meAFcTxQDx39QguJ+26uurC29yWLKGH3dGUSoagBZ
kjhk+bDwGmhYrnOVrJ6d897U+1ZUd9BwLpvtEZI+DCk/OVKHuAK6CbYX4JZUVOkp
a8jXfxhxCnnKI2ZKOdiaflhoMLBVLAEPRarF8gje9qU/PwklxyvanDxpCtJTtKtm
cA9NGGLz0zXKkxbfVdaU27gOwNkWuNEbJ8tu5QEkMgTKWqReGHP5bVhLJ1ZxQ7pn
50Uz8lmY2xwkWnkTHIB2qg6FEsrplQDiS6zg8/LpQZiw+kOUfrLR8ZDAxSWjvrlU
nKZ61FOyt3j9BU0edt9H7+D5Pmg67Ky+aA/XcJsW+5VDJwRNNcUm0dnuSzvbAL2K
QfkVzT8EsNANGGhG5LW6KiT8VpMHXEXlK8bsiIWYphAYO+9lrFsNQQ1VAbjnILKk
TnQ6GsCSQ3fqrLDzoyL+VOjtDzGuu6uk1nfIVSqtQP7DTDuoUFj103U89XnPAMWk
o0PCdXX9j+g3PUaqP5b6TeVHe3ndsrZd1tIC7UcjAPY1FjNoRvLjSwBT39v+a8IB
61KOg0s05M+TYAH7ZSCuIAWYktBDMgTv9jLQ1R8WyMiQR8qEY+IOlG798P6+UZ5Q
LqyoRfGWv6QDSHGQzae3onfJmL+0GRXW5nvLXE3mojOS6Ij9ef0Wz5UJO0VUBQ4h
r4mlqhYgIig7LyDqHcg2qVr4kZo7trHB22OfWwwpM4g/+MYwomWYj03531WP9w/a
ZQWc91UE8UzPR3m9TvzLGgdGbxIlXDizwGADkfkLdlcj9vsyWWJE6iUkxoYcakNv
tAC4HL7w95D/wo02nYomHfev2Ww01pNZdEElkj6L85fe1rfbIsQhtOyTVvfQ6GET
vqZlpefR9GWCjuY359CQBHTq8p2AzNKt0ktx4+RpQSLrzORaYU47FBqpC+7irsuv
ydWvpxISab/6Dl1OsFlI/NiFaxLOzb5dUWY48LJyJFeOruv8zhXkw7uuqgCY38f3
nVpMnC8RNUkWdhuVPzDBcKRhQQYGv4GFK3UpJN1LY8lUpNjxND8AKL5EJdPF7cog
OE+nRJTcg4Iy42P3/dqnwJ8E97JEX808Givv3QxQR/c4W1EO15Sy5s6wecUM4WTn
axpn1WF85bN3sZc9aakkZuygdlrk3bFMazB0iP60zvW612dY41TLzYMLCIdyAGTw
MSjsYHAR7HFTfX3NaDfYbJxy8BvGcYtzwDmscBPACf8SCDrXMDb/pklATIUcvnHL
qWJjWnD0nf46kPCnVnYmfkoqoK0rNT6MH0SPc9jb8KsaLKJYU//4mazSEvRbZJLr
65fvsRU9W1jiuBuCIKkwjZuSirLDAQ3Mru6oQzsdXhuDNlDytmKXHoQYXnDPRxA/
a9q5s33BrSfTw7BCbVHlUvUqcMmdw+pOAJpWZWnJdORgOEpZgYrp1yntwwf4TYEJ
WDxQTJjwRVH3UWRLO10YNSjM8vwd6cSdy/G4OzhDINuZkm35+a3FmaPmHM9CFz/Q
ZQPDqEFJpsT/C4DpysKlpsXsHJui2WhvEa2tLFMeotT535SXpJcKqwUjgTVMOpEY
aByCeU4BmBm92vsUouI3WHY+AdisYWedjsS2/kKPyO4IDnIkmLDvRnkbJJPJtauq
9dLbOulS2rg3Nn5R5204PfEdeLuGmftJjn3Gqr20vUM3s9vAK0cvwTSK18F41fuv
EYhWVJQ41TpgRrWDsPIjunaaH0fitCu9BEnBSTsQomB78IoKpvvzDcHxGOAPcSmv
WVpcM+AedzTuMnKCcvuqFUFJWu3fD+dmty5aBIDmhHnw4iKvQP1W1i5/gKIHeZnU
IuXpWZ9xwmijTeGogJ6f5Zu3EwleqOwqdlsSmDxR4DlRIy51KABRyA2R3tyBa+gP
ZCk+xl2Nba1rqp4CT1zQAKSdTJy6s9APmCIF5XsHllrbgFDBUZBBR0HOtsRdngQx
zwbIzWxy7gGCh+/fA0losZiPzGBt9ZxPUFzoupVin7Zv4FuDpkrKl5cPvKtrb5th
b9A96Wq6PikbtTuOsg4tGleZHLilzN9Gyoqv//fncsUAA0w+WOl+J0qECSbEo6rf
uqyi2y3/24bmuQ5R/B9+S0P9vN+dev/1ivjA0Vrnl8eshbE1JxKdjPtC2fVIvK3w
vNxvVCZL0T2YESFK8AbJ0VtWxcoZgWMQ1mDjmSj4GZeCWdtMskdTAguTvuB+h5uJ
w0VFoRyaHIbop07c61zGIzvDwWeVbXWQ9PPfZ/Gi0anJ8PNNdb4npNkEg0iSGGo7
Ht1DyW+1uFqfcP8mPA1KcY5QE7beesLcc5aU6ulLFbVgyTzqSDgFN9EZHZ8KUeJI
364JehIYja+I7ZXESH/b+MtaKzmaTZPEFV/w8NVqLEQ8IOT+dfpdHct77ci8p17+
TVMH4F3jcB+/dDxSF21IIPupjZl0RVcTXAW8HF3rfaxzsUpLToebwWEo1PCpWwWc
I02+Kype71T2svBqfnK8jJ+Qy1UWRy34tcnofk2fdEVFMOD3/kOPcEruQF7ioOSx
tHtdBOfi+gxmyKBqhTaCZFWwrvGIt9DKXLzDNYH/DTRF/RtSvj9LgJMRLd8C+vFV
Lr4G3dk2oUfiGTIeQGdw1PSQ0ftbE0mbUCFNTP2aVlJgXZt4znWN1pZG2Ouu4SZ3
wMk+PYtLrOwd4mpeAIW/iwnn8JLWXwCITL2GDAnrnDfXgVQkvBekHCm5UdQmRhY0
spziSoLdltFzEVT+ZU2UzNEfH5FMq1LSn4gXhGJ3WCewZ6xl2siBExZa30z1p6K9
eFb8TOvmGtVIOjsPvZ33JOztynrccQzaX6GYrUlW2S/5dH40OiwoPxilWj4HB+e/
pHvdZbthE73NHXFYU1ig6NpBNpiwM9j1ClYVZij54vsjTxahan6Mr7Akr6CfZyz2
YD5CWvoMAFZYf5pThzOhQIApEz7sse2gKCIgkUatNlDnQ6W8xqwgIDceOrML39tQ
7bwx6lyo4e5GBojO6sUSdhBIqAo0z/4aO1+j+vkxHEbMrJxIkLI8Ik0QWgDHRDx6
V1QGEnJnaHSaxEr70r4+yhNk/6g3/y36msriUEDAbsxgWSu3CKgOe2+8lrCcIlYM
x4B+h9vqwXNh6gIhMUGfE/OHO3a9ezEXDtPCRSJrBuixrgKnO+VIvd8t7+gkV8kg
HTjxNDAD/T8zYMEuYJQw08XWUm9Lc83WFe/sQ/lhq7Mq0WacciB+hFFvFKZKzcXk
hh97DsfNlxQZ5scpqrdkaNlDmh4M282BKnoSCAaBW1I4VbUitE5xbSjvOc1YpWXX
b6W2SCHZGb6gEpbXGY7tG0tUyeASTEYowZExFX/7s1LoWF+XkDgbpMVTbfj/S1TB
mWyB3k0ltfTUF3H0KgRKNx75/8uXVUatMbYD9NzSlO/o5i4O/g6jQ4/p5F6dHWsB
QheZ7XOMw9DUfQQIvkubGMpiGDZqo+Qx1xoP0VzBlZNK0MoPlQLRlQgEC7WuUmAy
qinedapSCnMNC6vaJbS+1gbvFqgddAlW08LMKoB2vYDT5TXuN9fHhpNJG9kYrl2L
+fhQ0u9ZdCXQsOnNC05ZEKEQwtVQ7D2MX2+B4PXqizQwmWzBRQHavQ39yLQw3Ytz
B7SINjqDeMxTcvUexMwSEMtgLc4i0J1HaJBkE7ScSR594Y/zxNf2ZFf810unrpAq
5Dfedp5clFN68Cv0u4NamLigkFv/p8FnXQwcYr4yF37rqNC5ihsn5q+LJ58ZGzk4
JzInvG1S8LB5gvwIp3gq5rNGsMrs2nOx6qMVc7mIeECpR85ASFoNi5vW48Ipu8SB
4z9lMPn6MWzjMdeR1e61Gg7qHMMCNZC7HE3zk343tfaDK5XAEx0or0EAyoDsUFQ+
bncQbXPLRdioDTa1KPj86fhgm+vIxMfbQ/z948F6qtPo8i2rCdxnM1p/tJJ4MlIf
OC8Fz0FyPVIa+OmBe64T5dt2U6TRbnEp8rIB+tW9I4CSLK/Z0G4KBSZUb7hrNaI9
OdqVAUtn699ZsbT8aplL3O+K5ImOiIuUbHBLp3gEhXdjVhK8pX0kMTC9hNDQ0kJa
xuiGpWso6CzQ0bqh277amSByPUkFd7XNtYK4YEy7VKQae8h/gm3tv+7ZspB52xYW
P4H6b6GObnHift/lopkbb1juR20kXLkTCfzcVqikQmSc3XLpl0k7dAhybF7P0T+f
axqDLURTi8KXHDHzgyjf4RJtU5XwT5mhq8QATVmPQa2B2kb+IsoBRUlWXETfDqy+
heAV0pSqbqW2kyea45UgmtB9EO4JVMkkYBzac6Q1blEQ4bVvXQtrVUC0Zf7VZ10d
LuYX527mmZhFiOWF9WitcqRYi/mBF2fqhZ1fhn3ESsDAIR9F8g+aBJIwFArPhr0/
xXU8IcM+nJWbzbtM3PbWmWN+pNIIguPdTWi8CJqaI/T+6ecm0c+EbQoOK9F72Vzz
nXNxcKe3DmYTA4hfgUNP8Y6ce5zgmrG9DT88Yk8YJQxM+Q6diXqIAFFScuxF+X5V
E5aLWUr66PkxiT5JyMQ5IRuVLqvBYqhfms8udxQJMBcf8j99PBnK5JK2vN0/3YHl
FPy166nyXcDWwDwCMt4HkEwC3OyalnSQLGR6hxxCDGLqtgYfNBtsL3BTl1RTOyCm
hoa3CvjIsbeaDAPidECU6rsfJt/3op/2XgYnKTGnAo6Z8myjA0EKVDemNhUl6z4y
gKPoT2RgtKgxMq69uU2ap54iF5fWVXzxDnu1zw7yucxuJpJ+hpoFIYpbxUAgBsiL
LGyfRn9xExgQP5skKvcgFslGQ2TqIfv3/d3UFzKm1aUuD1cLCod2zPIYxaTvZxts
Pc7eg0OYDDWOvJRqKKdYC0pUbYxawuX7IvfXz1oJ5Sun1MAMUImPll93V8+blKL+
w0Y3w2tAmhbK2meUAo87rBVTnAmqIoYzl506Yxf7BOSjnU3Ri0S2PGOpqbXrJGac
uFclHP/g0U4LNTO3F5KMklM1ClXGi5eT1nIihwMmfPTcz7CPViPA8TlH7RDAONxr
joEhWUO8513XWSht2RI2TMmfdwGSoykVn6/UZgvpvYGrHcYyRsEUjuVt+rqT5KRg
EJ+CijXDg1Rw0vhMWyQPXYNAYsqtecrElW3505+2cDbRpryOBV0skjlFctBeDFTW
SLUy3teVC7W7GcBdpWZpSvSSiw0tgzc0GjbV4rm2cfeaTVmwDPnNfJdal53Z7BcI
Hfo7dtxPxNHttfRdTb3/Ol4S24gBikL6JpCB6wDPO2lwjKIacZmt4JqCWsLijyTa
+IpYrOfvfbAVA1Nn3fE1pjKroG4LbKk1XcreW2c6E3mnE9fqS27raNilTPNSgFqQ
qZTNuucddxGB2AIBWUR9ZxRQzJ1MLIhJQBi1ETkKkvmmUbKIfMFX2/s6BlX+opEY
66x04E6sd++RqwAVvHEaI7KsXCXEjIsI3ahXXt8GjpA1zX0+B3jmefiPsiPwwzJZ
jRYnhjsO5cjF578jL7D09cKBJOxrRibLCtPa/9W3CVv4pBbda0ZJpDUmI/Lct+km
9cIf2AcyH+4lPtsrIEc0sqvLm2bMrbAtbC6pxC+aiwVDg8ov892FGsuKQc8w5KQc
GNMfsLlGu7USh15hOLJdG6lC+DEDXaJc1s9hJyLV3x2Ud2X92yZM9GLc+1qfZwpJ
DBahU8ePbeVhAA3bN4h16FzcbGjr2N5V/YnPViDmD6PdGfnd8PRysUgKM1nU0Frd
/tQolLTvDCU5xJYnFVARItEeY1AHOJuPbsvVmjrTmeEiy5obTDRkM0XjBdol9sq6
1+cBoEZRXAE5qKlLlYKzeaU6GTQ44NRKoOC4W/D+R3h/XBOLXGGRNOKdwfc1EELw
5ezYTKB7O/lgQ9HeteS2/CxzzLDxMFgKVZPCr0NF1sZqWi+F/vSDXfsXVq35uUwv
hrDd+f8cq3cHZZ6ODCsjPOhOMEJOLwcX6r9pQ6EgI6UaDyWWx5oHPn+rry3E4eQw
2GqkZZ7dgLnTNyfSBj1+VU8EWUis1YZbSC0YS9J7pN5ZnxwkNNkUO3iuGgYJP2O2
yFaiJOipVL5PTLhLjOyvrOJz9feaNDpv5u7K5RSoeXn27d93/c9P6spuDN067aa4
24ew3us8B+fsTxXgHGCOokRsiBH3oVSVNVDK+Ga4N4xxPw7wED71DHYtGRCQMlEp
fMiqgxdmN81cgjLymcVt87ABna90ZvfBuQ8N2Istzha4X0leSVe3f/iL/30s4n0y
umPSecUb4SArsFmg4ke9V79hmU2hHOMI8gWet54BQMdckB8PKZ3je9dNm4euG9Vn
9dZHuzGKwz85qoop2un15ucqfKHuXnT/iz9ufV4l9atmBuD2dx5US3sIonGfgsLX
zs679xEMJLqnok2LzGWyrybVd5VG1CcfJYJpiuZjsU2dsf12xn2l1P8/2dLiHKPr
Rykhm6IXPo7eL5Kbkm3jdwjZqQ1pbr1IMYsJ6cRS6Tic3aHOhhtAWkajAjeBj8Um
z8Czv8hb+Z9ijODKgH2oOW8Mqu4SI4Mu2tr60fuV9pIxK7XsHUbvGj/4qnPjlu5E
bDGnR2Ox82iOW89ctRQzRI7ZAVNiQ0rySr6sBnAYaeb5dkVeQEHSuW5JoA1fFmia
--pragma protect end_data_block
--pragma protect digest_block
RSFHJ6sBWtXSYqRb8H9xpoLF2IE=
--pragma protect end_digest_block
--pragma protect end_protected
