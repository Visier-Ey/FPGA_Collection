-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
--pragma protect begin_protected
--pragma protect encrypt_agent="NCPROTECT"
--pragma protect encrypt_agent_info="Encrypted using API"
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
--pragma protect key_method=RSA
--pragma protect key_block
bfQhH1J6JceopiJ4WMtqD1q4j9JGIzEtWNwXU7BRy3xdvfrDJbqWsIS+DVhYjRYn
SO1nvA0otgV8Ko5uA2FjJwu5HxmdAvIHHp7LWy3wiEk0CcYLLTdYOmoKx66ImBMS
MMg0Wzcgx2Li4vJsPN7uZR+Da319AhNTQHtdIN8C+xKg8eagL32okBRD4Bbpqjqx
jXZ7KNWJkDwAvNKDv7ziK1EmEbML4ehQq9irPYY0+/CLz3jKV4axfKO3RVtalEWb
s718sgkF0ZXQKyoQlMqco0uiFE0U+5h0Pz9wS1oiFsw48U23cPaH8uGGfxCnbzNH
PJNWdhuKLzKi7nFAEVWp5A==
--pragma protect end_key_block
--pragma protect digest_block
cb3UxwzQd+Bn5FA6DVuzPrndCKQ=
--pragma protect end_digest_block
--pragma protect data_block
9QJUVaRIZ9vNn9IIuOP8n6IDFjAuOk5ZohBE/I4OcwqSp5Cfknyj6H4P5t5Zr1tw
qV4E9ktfXsPmRns57K1DFPUncYjrJ2vKbBIAzJm6yl0LH9jT8Rdi0tUWyP9l1hPh
aGy4VN31JclrBktjqEPgXS6n1ez5fgS1VWYjS3VOqfM3+G3nInvU2JrXRz2teu24
DjkdUgX5JzC1tOe7ybUIhF/HokJdi/M6Qi1LbdsZmZjvjd/+j7xkmm+UaRS7JFJZ
9VgW4IYq9KmrDBFmcIpDXSTcx1buf7lWkYI5Bgi2qksQS5Xlhu58+1MRE/iRudfm
z0Y5ATywD/97T6Y/xCItlMUfg5WpKjJor/V3wZ7ju8VfkiRI91GMWJERz0oGH39o
WDJlW3+QKyPbbpJBrDPtP59j6o6TsGCjs2Pql7PDNxBKGU91+T476+uBEyRrbYZA
rPVXoijz+hyXaCZHchBU6bc8VV+hApJdX5vItFXT3nRKMAObuTkTrB0vKPXttmNf
PidZ7zqzB0js+nKZkrvnX2OF82WIJH2tGoJKd9v6ooKXK2mHq6aG3LmYYyY7mdxk
+jiqsnc8LhUnw99LbCOXfxuvaMEGOBrV6cdv/Df5EewWZeIAZrDRr4l+2G2t8mQf
9Yt+TFkhitZJQ0+WzW3zGMiJf/vkC9vAV+QfkcHR6eOvU0VqEHr1Yw14t+VCi9Rf
G0W/d18Ga8q5PF6pDuL5R6JrAa6Nmb/4PgLrDvX1CVmenApzexZa/K/iwiv28Ow1
KJXl2RSV+OUuQ+HdTesXSCT32yKf5YUaqIwgPVGzLSfGMfe8wdNUnhI7JbD+dXPd
REvs2pg5kPtmzEKCdlx0lNUHpsYh1pzet8zXkcmFaJ980Iypric7GZPMHllPnckq
D8B3O0O34uUPYtQm6+YQ4oKbLYGQav159JCzCF+bXwBja+YHWIc9DgNS+2WAmy3Z
O+xyQDWLp94r1lc9mCFdwzWIF8WzWyfEk3lbo3E0zsGhzZo1eA5qZt+Sk3McqGxQ
eDsZeb5bHz3qzwGGkYWR9lmRyyKsQYmuF1KQnnU/F0owpWm/lTlfBFTmlREfSoob
bMLg8utXIT+8QhNhmn9CNDC86IcW09It5GfupXIudD8+R2NRAHwu3byIIDQ46yhf
RBVzTqydw91FvQHIn0KS6NZTYmkcriMlHzgZBPnQaWKeED1t88L9O/NEr1/qhH95
8V6q8HsWIQE9OukcwVCtaBqeYRPs2GDxOZIUKXSL0rlFBZb56EkdT5GVDB3/qGGS
9A1tyLHdZ1TPvD7V9N8Ybw8M+DykWNJJbTh/2NcU6gEeTBpmEQEcVDvsE06rfp8s
YtE75/KRWJCJ79P2RR2mqoZxshFon1yFHoDE+x3iQZuo4eNd43fJ/r4skO/xsdkz
2pJ6FD7yG2XnzO/90/HIs6z/Ys/M/IdQxoGbVj8iWbMj1A21sCQ6Tmyas7q2K8Af
lk2IJk1+od0dNrFu2v+7LWsMD5KOXlC4iiVm3mxq+Xj+yI04SLW3yL7Lv9om8tTk
cQ8a91wGOejkofRtVy2LrfwbS6xYSlrX+KWnl8bNO/Sj2IarnksfMWzX5fOR1XWM
6eUmJxr8qY9raTis02Cqhwym71iIhnHqqaFK3GXmo6p/S169JLnmoVeNsnFOX7fd
WIp13xw8kvXd9wE82DNDUmJThRodnBqOIDXVdi2uCUBN92PU4LexNa+EzWnQiuAR
Kt8uW1gMNxEjWH0lK5TPG0GToYBQWO4nJKV3M1topj2gjpEZ+Wiygr+4A0HBkjhV
L2wzNKgPPI6lt6VFteIfzWbTU8jZPI8TZewwJ7IObVfXsqPUex5AfnZERGOnl/Nm
HXrlz2DccNlqMlDJQigRnNdCr5az5DUAhyJYuxunovyIBmS4FW8S2JlICQcjLZU8
TkAAutgXcz9Xq+vKA2/TyICAIfhe6hbRt6Z7s3MPRFsp9MzfjupERW4AHywq3P6a
GJQJaxu9VgfZRTTuNJkyiwA+Pp3YNDpBy6KW1Bfes1FknOJr2mGmrirNpRRG/A+7
WBRHyj+LwMJTUd7PLvSzp0Mj8FETIFlhMH1lv59CToq+SMqJC8MOGI4BzIn7w47p
1mDINJvK0/WEzO9FoujFnZI5/LXjfIqnUb0gB1SxcNXBmvmv+vbU9xCEJAloMjTd
CzDtOg3Z8g5uTKzg3c8U4fNtBh2SrSNMbb1oUxkJ3+yQie8dSJ7plZPCw+qaVL85
kGd7CaaLiBB2yHQo+ZBgI565XxQvqNF3u2kU6sG8KMxvOrDiylFSC0phYlsoQekB
EihkUGJv8WJyu7eDmQ/TXuTtusFstofGwChQbv3etwJsUEl1mo/HkD2nqsXBayXH
ukDr6i9MMXrcAcr2ZqIdn2X8YOeDmZNTf/C3sK5ll9xXugYU9Flbr30M2QcQ8c8C
mtZZp072UexdjOahwoZvu86guWr4Swg2a9uspp/jhnjOsiQDd7kG6s5WbsRqzUHd
wD6c+2pT2IKQhl38o/VTEtPPnbb9uHbDcN2OwDgdYA2VDSIaygxgxKLhO1nQbXTv
ZBdoqZ2yThq92354Nw3A4N8zRTFh8Tb9qdkD9CeXM6BV2A5olRlc70Lh1s6PQKvY
rOBlyiOQnuyidglddD3Q1AdNfdAnDzqcYLxc51FRPc/aUnJCJi52HiBggJbfji8Y
OMWIt8YVxsrhhFiCJmNBTsclK3qDIQpQ4t0nfxkYvPPw073K753jyAsWpunfJLdC
bTo0War0D44KruYi4x2gwPjI2MmdjsGPLbnlXXz+VCngTZsDSMmKaHlq3sTgRQHd
bzuR9L2nt2iEFtxpiZHWCqC4HPgKDIblcLYnF0ztOUZFd1JDM7Ggn9gvFyT7gnQH
JfRsINtMM/aXQOT8ZNBJ+l7ll3dja/E/sEd5HPwxIRwIg+0iwDzamQV6QiFJ8hVf
in9xOBXyhY0tr0PpiYXJKx9zcyy4DdEQuKAorzotEpbzTs0h/sc2IZpDFHgw/hRe
eCpLD/zD8LKMUKtjF+1V9MaqCQdslyaNe/nin2oNPO6GkmyYHIVBer5T2PNkmE1g
iHNafyMW8b2VdbGIAUbbc/grT0gvVCeU0flGyOytbC4SRWEWt6vF4oE4zkr0SxOJ
KYMAKP4OT4SUskNXiYIgbVFceJo0NqHrPzFXlUG8qJWDzx5mehQ9XPoh4tOdfocN
kFZJGQkxndrHPX0cCC/NRrU/EnLM07CDlWIzu9G1LwBQ2YH2kCgGcp7BUYUoOzFu
hBfFYH98dNeTjgigtr4RP6cLLhE51X/M7skqHjMN58bbIEgbp3o7PBUJzsO3FmlS
bbRd/ON6OmQHqloLZrE34BTuqHeGO/34V/FXgDKgVpwu7mti/ts1yzE0rfD6Zjas
MzvBUJ4AnVshCfjt0EYin78M0L5T6DlYGl5IdrUQWKrfHTofYmW1DLrQzQXkFay4
CRIoR/Z6KZKg8cj/NZpUqQSh8p1v+sM4sBdHSAoUH/C/Q0Hn2Z4gXIfRFniWk65p
Kiwu78CdkkEoas19ChXat1rsCUjsMPLuno3Q9k3mu7xH75RVONENtzgvrsIvQ/j/
PWqHEd0Gm1PQ+Bx48zQIRCI6FbEbwxj7wwYgqqxlNZFm0uLUA61N0vvaalrD4O2p
tlXwYd3i6GWE2hbNnFYTjVgdFMzJuZ8WTAOodxIp8EoUFVdWNfUyOtNm9iVodHYd
JqFtnQtck37GvyBCK4kyYg7UbWjKBDGKkscoHsQKMyLdfjJr4pPHzWI5dpU9YMfl
JCrUhV1CJqtDpn2R2E2YFR1d2Qlt3wVBBQMAI9tbMQHAEKzxuyMW7D2gdu8n+FSa
H+EvBYqOGV6PDUgWg+xsF7FMjJXZEb/X3J7pBAFzejFcT8ndetngep4HLSJWX0tU
b+wPal78p61IgfY8vldL9eCJT0fzLEYmrktcRNFglngDs2XADm0FOokuKrura0YI
Wk0D4t5xNyuVjP/beYHLiCeSVgPsNh/tbjIanFFI2DeDuof4cCAq4qOJOevct1DZ
+0zG082A8TIx9HZ5QEm8xH4+i62mkniCEi3QSb96Aj5KlgxR6uGLjoq+FcoFOegp
jbyfiLchYyFImbFAETT6+V9y+oFLgDLDpVeXtBHDsUnQEi/yKSMqNWz+AxH/wUQc
ZIJgdfuDhUv+cZSw75A17WeeNDiegKSeo1Cq5zsK49CLi/v/N5LevqRfZ/G3zI+3
8gYDy/cadRN5/wlMWktodvFD0hCqoIi9P1NEcENYdvFWXRsrcn6SStM1kbFd5K8A
oDytOxwI1kld/P2QVlSq0Csuf9SNvQiZlvpdb62IsMPYaBBTaymszrFG9zSZq7hp
8EfisKEIEG/m2PW/KQrK6FFTND/L+WZEfu34JiRbD6YGbIBOA5z4SCMV6I21D67i
gTCeT7Z2yw9Wy48uHfyTIW9SZKx4gjpjvCAdePVvTHKjh4KESoPWfXl7clIAdQEG
IYF4tc4fWYP4CR6jWfv7Fy8QWb9n0kuEiFg/PZSQo/D7FpeMCtBywuiukbq1C4hg
Y726pZR0/8qQXLOBNXfPJCWU2VRheABcZ3Bdg5jF5H3aEy7y5xVEdknq+5spiRDo
aTiBZ5riVOnqsDxGV42fjUEZx+jc4VClIytfw6B+35kyWOBlGJPnvvrhZmOn694R
YwU5TMnNBQsEVGmHrH8Nddjz2nD5EGGDLVabXMqzcvO7qeuVf4rCRfoeM3CjHZ55
HrPumFuM7U6hbOCkqhJwS54ypt0D3k0NTQjEHkN4aclxka6h6BdkiUe6e4Apw9v0
5nG7QtJUDDkALqY1BOJUzZbwsxAb/4wsj5gp8QQGI4xa97c/QZCuvvGdAUvUnAAW
EoG33PSTVasaKlU00SUUgOAfZ/9pmMYr0sDOkIDPM/3xfOToSGhUfO62LZC3a+Pp
9fpvvFXDj12IKdtDhw3jZoLJ/nLAKT5thprvcoKwkfx5vsszvHEsVYMEK187Zmjy
Pv2BmelVWQrMblPWnUDW+HuB771+61jVLvxg6nSbDM2FS2yCN4/xbWbetWLTmjRp
qEpjTADj/PFbue9a8hSecDMgE3RW4qLbRXE34Sx4CAXEGERUSYFPgEmmxSqRTqx7
Dd2Tao8JvQ84aIis6W5nF7NB2gnjnn0d6vsahyj55p1+dz+8xbdBgb+3qjys1zBn
rFjbu+dwmRSzUkJmafkmC5mLnuy7KCPETM9vLCiy99r2/NP3crLwHJhLv8ypJEFd
LZRHzn4Vr8t4dgRVvGV0A+j/tFVT6yiI7Iu3G6LPMRHsMmgPk/PE/qaiNf62m+kN
R+e/x/gxljutt4EQu5q5T5nT9WRP3zc+oKFXazeGFs6hdPrPT+pjnfKhp/5jbr8m
db6dzeavbXcdJwwihoPhEXLC7/iad7cZQFUJHixumjRZynuWJT34EYXcfoSHUEAl
iyFp17uVt+Iy5Q2fAZbSr94PDP4l0KDl91RdJ1x6bUP078EPFPOwd9PC8h2BQ83+
mCEe18QrM/ESKhiJIcTH38GXogQiyBAgKPgCmbtasiEAutZ4xo5r6ph4jaD4fkjL
v/pDZREJaQTJdxmlgZEG9aWiBAOMDjJMsBfBvYNvMgZk0fiDQb2wYrVllJMzFG8N
kre4grOIXviAV7qBzOkdwj21zMtDuSIrFHeeTpeaOtwg+7uJjCpB7ybnvpxgJxpj
e+YHGUkNRgG6o6OTr4nIsvnaAeDX/R/nEWp9SQcPFZqmwBe6Ftd6RvArbh4Z7xOV
K4AVeIrmat0D9o39nFHBJSraTHoxCVosCdZUdFIISk4TQJMdklZiTp7MYnyTOGVt
467z77PceEKYk+ERqyYFSfpdPKehR1RA5UihOlIPvPPE/fblCGCkHsf29FxQWMAY
15S2/D6jqpy0m4x86VfJzoqzKjDlx/KLmT2tNXQYPh+DGX/BSbkRZl8rAlK/4NMe
clm+fvJxxOOH/gyi8h13UfckT2Fly87Sa7fK4hGJiPld0mxLvH2g1C8sy7Cg7al/
urxvVu6E5gqksk68w5er2pdvDdOF1927PC0xib1Y+YV9pLgsTdS5UfvHoO4BZuVX
mMHLjkOY47zHGDfE9MzmqzA8le7Jp4Q2b7ngfOWKLVzbz/oz/enXX+aRI/n9zSzq
vXxEt2rcM2MHRez0zkRjINVx3YaDx03xXztM9sg4y3GoBnWyJGnj901AuthU24NW
gS0pUn5UNGjrmwPCCe+xZTPza7UthMcpxCvj55FRzmddr/G3vE7zNS+owf1j1ePc
oMzzk0JrMCvl+tzhEvDN4i+8aVsftUHRej4oGqcS7L7lWC7FBwUtgghDTqHEj9pv
ylj6PY+TL2yjXlgbKNQiSrKYfLlh69OeHynCXp+htXoFjqHwJ8VGrIx940RXhe/b
ryB9pFE6HahMSMniNQyzRmARilV1VSMwgeMnvIsMikBTiXCWw/0MQEM1b239Y6sf
8pB9uGtM6f0Ne6UG7cqgGUc9kxBQwGhPKrnDJHzXtG5yDaiQ/YtSe1AtLOU1ATUI
IIVomMN9YjNfIKgMH/QjYdcwluqdXy/RaP4ne8EQfne+5w7I/hrgjtpZpR4ITK03
W0T1oTd5rBOFZlTpuvJL8HoCsU7CtokLTCkiuxQXSSoOq6BX6eqy+cFRC2WO5DJe
vT0BcCOH91R73ExrSzAhT4jQFFjGQ12iIzEYvvOILaez+Mqofwajd7sZC/s/tqPz
F5uIM6EVf0DEvkAMONp3bm1nlcdrsB5+qgynUub0PjlJ1oIVxv7Z1uQzGCVXSExR
ODUUFlmUA4eb5ouJK2I64EetARzcrz/foTlA55j3hV9LoF3WE0Wgax/r14Y4K1aP
wPa/3d9nkSiveIE8yaMfrShu+0YOzt7E6JA+WH8GUNDMecw2Q4rhoGpGBd2c0Um+
X3YS0Ik1dG65jJvOZucenWHU/D0kLqNOkJIYNhnR3v0NJjaHm7ESMOHZPRgvzGvf
cvN0+VMOEJhFA+K71oPU96wQrQY78z0TR5JC8hiNzcfu83DZuxc5e9FYYxr2oB+z
CS3oHxfi7DfXDeUc6idfLW5Eub2121paUnLIKDFd0uMG26/tj4+OljMOv6vnuher
Q9zHwCKf5Lepoh6m500Xcz8j+kE1WLvl64r3Qy6+D5mVLPf8/t8m44NUxCMo1zPX
xLkChXRoEHjcdTf4DJqWnVpAlV/J/fSzWnOsx1VmYA0teJ6bU+Z1LtJ9brQ0LlMZ
DDvEHV1lQ65JI4DkHlbI0lzSRI0VHMOxtIV4w+5ul6Y3LeeQQI3hUPIO6fvasKe6
lzMgZYLrnDu1j+qHoeapXbNsF9Ty/Esdw0rQs0useIImmPF8cZLmpoB4UE8DV/Tt
zxmY1vzOiIwb1gdbF05ZgtfW7gS10P6SguX3AvtcJO5FlKV+dyqQCa1WYq7lBU48
4elZ1EWtMZJWEBCrqqI7M6IUdCw2YB6Q0mTLH+aegh7PxjRlhQJdqomwgHwT8cD5
HV3y6MrXzpIHJbDApaYHj/APoMrlO+r7ijaQzqkEeJ1Z0vlY51RXKxyjdlMC8H4T
7uJSZtzUaf9OkL3ivjk3sY/jFRX/78IDvZ7xNuYONaygShcuL+uHBXasjGuL7qLu
nOKOfU+AxNIf0SaCy50aRM0+q/Gth+rmKL2nx2MySOz6Y3XWlV3bytDAJjluTKwu
3z698E+q1NFT3hE8pzcg9YYhxZ1h1jPuJGJrQ5wjabAVMdPP/Mp6Wt8g3RRUNMBm
lWoU09qL8+QbJHr0LwISd+Ii7PhK267rdXICGqfu4GjAuizfS1NHSnHa+qnckzhI
oBXYZiKTLR2r1SGhA138bKVvTM2wIysvATK3CuLg2xOMacsmoptGcgpRDFp4E3bb
5fduIYqfHWLf4qUGwOa0ksINlAuRFAPb/uXueku1D0PCtz5iehpXV7BzVRQ1KSxC
gh2AlR+4Vd9mkM5bdlmCCYmGO0heyDtB7gY7pspUXMmQCJrfyM0GAPJduabkcpoH
1Not5uXGExq8NTb/He+0W4U5qbsvjkHP2dlTqSZ7e76u7v9L2KA7JTsWz+nA3D6G
i5H+AZ+MfVog9HdGkFeaAVxlx92udcnIXFB68YQYk96iZdvDtJBlQNgWjiyyqfd/
LipXg8oUmPetIPgETmHiJrA7A6bHMflk6S9GATiyztgX4W+xLeWMTBrbuRqxJp29
Lkx+99p4vOJxstTLWgBHXVy7VZFRQ9JulsV/IwFan94Mi6Lx5kW82jPGcz8AezwR
YAdYqMaimaWXURvjOZDbFy09nh5c0HNPQ8wLN00blIrgZ7M9bQmDQC1udfABNTxJ
kYaaPOP4l9E/9aiaaw9L1H6sKUbVuBs2br+L/yxuZLvpvdeGoRRgUSCN+9BBCd7u
QYh0zo2F+W1newaRNhKJ23MXImLNtxAcqaxJkuVHzGP+3lmwp5ZQuOobE8L2Au8v
i+pliGjVF851MlYuTkP3QT8VQ1tHDPX7WurYKeDnR1WzWHKcLFnbKnl9rtZTTMGG
LvSkm2GP+vJBydBw2vzoLlXPGqBFnnZMykGJZzI9bMCj7fIBwWWeFARJRDlN1D5E
NU8aajtQMpTE4JWZ/hVWbwAwgHL/qinEzfeHrO02G3oMUPcX+UVu/TIvkHL9WUoq
vLUQBS7/WgRmC+MX0+ay62vu5KXFovz2sF7CZ3CYx1PvUy6sowrsegvd+ctSnipg
3opun71457yfI8FAiwix5lH2hZIxAGkE1pZgWoKhwlEe8g+I4X70FR0yk0UgK1do
ivORmsHRgQT3a/ZmF3HqHJJawB4zn0CS0lT9NZD9vhrZwr8F3SpRkYoQVouDyLHD
d33bK18AHhsY8XHbY0s6C/dgA2dsdntqiF4YCekdB5NVppNjdkJJvLX8TGL2Q27u
hy7EdfmfEawy2xKL/n8BriUZ05YoPANdEa5GutQtlMzL82EV6Pd/PJEE8Csyuq0J
RgEn+dAYFW513dDeAJ/+wEIFERR0ryGOWn+K5vkEUca3+Tliz5fwDQG0bZCerFvQ
8mHZmhFfbXPCgItXkVH+e7+i1MOhZUkLKCD6RjK3iQ/hlgoOHKGYD/o4wJwVMsjB
KCt3RpKdUrvwc3B5tgu/H3qmqcaBGGOAOZVIjcZi5WZLh0tRmTPmUkgkizXuIJlv
OWa7VtxuS7OLOaNA55oAYuLz2tN8QHBofxwOOpDBn9/MHdymU/SD8TAvf+EtHzuo
DzoYh9Z0r2/c+0Rqg4TzufjF1bo/9zlDj4GZn+GasU+AqO4bffEBNs4U47rUbJzV
z628hGy+iiKHhz3r94oeh9tZJuZliMAXhSXZbAnZkLcZjrUzviHqTFawqAFaMeZl
i1PRsB9tGWZxveG81d8FhQ6TydgoKs77JrshxSzUCISLC5Pi49M3Gi9RxZoe4LdI
w/5USKSYl54FhEqHnQxSyqb8BXEOP3Jvtsl76Of4MbMRIjLMwzRr8XTJRhEYrbp0
KvDdgakgoLlXLKWdfzuJEFgdMC1bq2VPiZqMb1NE1JOaquBLzPx1Tpj2rtSKHsW0
ZOl1dYrNULAru+CbhFql4KKGtkQAdeF86kGtrV4OHi6Z9LLIObQPM6e7S3meSkwD
JbkrINDFVHRbqr1Jgrolu+bqkO84WHJ0ybvmwPYYqTpO+phJZZHXdjvD6R3gUpgO
2HmmEApqf4G8Weev0r1sCj5nIjptuzSZLMxb0n1QiI63/16DCIX7TcNdKyybT1vU
Kc/kmNPpGWnzmojWLqP6qAL9GUZ/gntsV9FcQC5XRU/ytG7pGLKZ/sobIrToxFyV
qn3HviP7MybZQcdHmPriNgxjY1XNQHQjs8qv5BjBMW3NHwViwQsaomVnW6X7URCA
Ahfa3sC0nkcZNlUdkaHFXt+NdyLQc81jPo7uLUAYgKMt4fIyukNyZPJPFSYYpVua
f9cUAffIubA6EqJHfK5Ndjogc9zgmrSHYLDIg0O43Gjrxdm8irBkQ66CMzk2yB4b
wDUriek5dglIsnVO/2HMmEwkJouKA9AUXL/KW1Nb0BfRhqN58Cy08QlsNtQVodhY
VSnIJxgDNEx+rDbMdM/rfnhAcGptOHVZFD/7vQ4duzRKXqkDxByAyu6v3qxfUNFy
OSZch+BNt5Tz3ga4S2XgYDsap1I54lCPWWcm9P6+v8MLna3zVKBEixoxl0QCoLXQ
iDEJwG7amHMKhVkCks+6DC5p1CUCOljhejgFziKxtfQ/RI9D/6HJcfC7b0bG0T3l
zmKc52Smlhzk7oK3pEcT9iONu2U4mFkC9wTFJQ6s30qSem+wZPMzN5UvkHHYFrRc
GjUeVgwbDqYO+EwdML4keaDhXAdhWeJHYZQ/WX+FD+0RQQdMSieO6Oi6xxDmn0Ji
yBTxUBxOdW9a6LV3Y9FxPeBBO22OdTyq8y1zly2QKOSXxbnvZSM8StE6PPsBxkXd
sWsyehsltpybLwZEtxj/be4HBvkEDNwdApPs3ebz3t5MsTCgmhjkj5xljH2Yyhy0
Jk6iTKdZ3Z1zJIlyKVMoK2vjSoe24kuRsjbPiVUcwfBdHWL229BfRJcR0lBiHuGt
HsbN7ZuBNUtHO+iOMQVshOIu1XgU4L1FfTtA50FGpuclzdUOy63ETdGNpyKCg4XL
8ydSQRBIQDXnbndhfyXdSYNmOrQPfwwTA+bSYUvyWmLbkW0dP74KGeZdJ3j8JE7w
4hUxHldb+UBNar4cnUaN8hi55wGcTE2smk75mPzsy+St2cSA/+dAq+waF6SSuiP2
an5xrCGYHp6C6WECANu9F/fCiCe3KgwfmDs/M0ALXdEu/U7p+Wkc4wvHCvb0tRfF
jPjHq8HvjA3gF0RuXsspJVNCeLe25aLgfTZnW9MHOiYO6MVl8onx2r0h/BOizOUB
PrrMXg6r3xafwnaOtW0Vluk5bw3cEGMbDRNJQtFkUKMY/5FsE+Me43Rpy9WNVpBg
2svEhhpS+MD3XPOyful5XUQQBWXZn1pvpcGfmcSv+N4grIf8Cuticjdf5bvMV7UL
22Zm65qORjUybNLA4y4JVuo8xTupKbnszqDRMWa327RqNPJIZG7LFD/NfPHf3+GK
rRn6V4VQ9KRdAnBQTV6mCUh3ecy2kDZsULUXh9wWJGPab+EWQYSF0p9s41bDAEdf
leNZ0mUE2abRYWh5kqZadAhNhX1eh8VhxbeJWU79nw5LH0lwKmnxhY25/hQMtKvA
56wLabF6lXEJTBDB/T229oM/wvBaKH3b5jZpFdbJcnpMKsZAwqNllOMb0sbLsdqs
/O8ZBfey8oQ+15vxQ2wPj3OZi9FkHXQlzDqjFL+gtXzjR8gFyO4O6i45lw4Xt+Ct
Kc5+SLJSvbwOZSJkap+EFSmcHHpZJ2RmzTdvm80igibY2/w+qrg1Ws/KbSQJa3ss
xmgmZWtFz5R8lioHJ8wwnIOyEfhb6ouC101kLUCE0bxcVCfSHkq3WY0hQqDSJmlH
HR4tHsonqZ9ca71v4aaWvl312SEBmMCFmViOO+KA+IPFcA/R4ZT/uBdqp9y9LFjy
TJ2qSBlQkbl7cLb76dnYY/N9Djc69Si5HFW4Ts6ovtJ6hMBed4a7Bhpbu75p6m+A
4Jj5qkA06W/KB9AK4JZfpxeaT0Z6c5/hCNccvC9SKBcWsqdJTk+KlXyXACGfJoq8
E2SqhN8FX5t1+s4JV4y+/yo04yuxsZttQg+gt8NzMdNfXnu+jB1L1kP/KCNpw/pF
/u0LIGT+oQ7gb5KJSwxw4vlKmwoSNTI1JxqDyG09+2Nwj4uO7YseEqzjGGA1ddNH
62fY2UUECnkrPiCVXv9JswQsuZ0kEpJYKRmCMKn+OgBXhDLxUtE6giedXnJHr1LK
NSnKO1C8gvl/IxG1MOjKuJZ2k4A1TiYL9Za2e6GGlSpE7RIXrwgw3NjPv5g/xU30
mEsCnqe/yNn2d7vLEc9n8tzJZ90bB7qAqmcbnJzvx97a1QMMJl8543tVQ/DFJgxE
gJn4Y7De1mYzuWm8N2qv0BMwr/q7foHyfyTG7vafgF/ghw7iF09KY4rNhX9Sm9rD
LGPukF7uK6GjBgqRiEbm0ElMTonz/pt6aFeI2u9d3C4yt3nVrUrBBFHCp/0wjJFh
m9ccQRKL8ymf91ERWSTo7pscX668m8a9Q6sMCwEOnrZUJlw+YN7WPiBNWO7wQB4E
2MoTKAfkkHj16QjhFLuGIhjE87ttzu++Zr18vr4+hZuY7BgUMpdR06aocOPzC154
xn48TuJWNmXxCftYYx49tQ1lJgPEE0X4IMaOjGyG7rNZ+T7iiWBLgf6Lt+7yreRa
Ghj52Txuo7q7/pzHRWNa+Wkezr8hjC+0b0T1EG2jYQbnxhL8ReZktcqpLP+4xT01
hRwLUUNDdJFQp8ASyY5otyOtsHVxCxPpF+wWs7ZO4qXRlfZl4WgZrqFHkgGU0cIK
LN+zUVBiY8e6Cy8YTj1XBwJqWiKXjJoJEz/lQJXlG/UUCXkTYxtzJOQBw0MhglsR
muSnB5ePYsQvemXvKeqJ3j2uhfiDOTaV2RxXJ26G6TSJz077eB60+aN7OfS8L6DS
fPNLzziRlSElhjwsUqT4MxcuW601Y5nIAR67ypm0NI0fvmKahJy3oRMKuKILYCud
tJN3qQC9d/mS2wAk2cNRhA3r9jKQSXj1btw+7e/Zby8A9DT6MsfX4uonNGQmYl0n
xKJgboa65L3fjfUibc4IEvwwtBO4CM67i7EbNc3bZb19d2n+x0YWwS2/06v6ZoVl
2R7gkTLTgilK1v+y9n9n3fpvC8bC/CrTdIaS1X3LcoC346dQjDA36BTdmKOYAO/4
9IkBRvbhrTvXhSpXZvIaKUhCBGymnvAST+J8RJl2VFoQRA/uMzq6nVfGNm4yk9Kq
pof2RptXrVX6dffs0V6UDR0w67xaZtQGdEjOh0xTl5De2ySeolLiV7KvTjIigPOo
sKl/Ek4ToRGIBFeiwuZF1Ac8J0vvuJWiPay3HjxV+TUfDK6deotlwBd/ZNQZksuz
sIKuTuGPIY0VZgp7WhxJ7pbnZHDzygEZRWobxBuTafVg+LLGZnSyzVx4eKLhtbVq
lxoZtn/fRZ2sojX0ZcwRd/p3igebMK28lqh1iomJ2sHyWPkIl6XfxKCg2tp2NZGe
snLBxXfo4T+ayRseuJ1jh0KirQ4yCvKuUq+Gju252Usp8sUSNCfB5DtaSgXNjYy7
oEb/JjH6Ss113169feDD6mciR5XHg69ZudBsQKVIAqQrx1YYhbfMUMAvWJyGAI9b
GIUcQFCzeirqr3moZzwmnYld8ltQBNt9LdE8HcXdw36WXGiX9popOtj80v2k7Meg
oV+jhTwzmz6DcfFfk8SctZMhb3Z+l/tptTyGiKWFnP1XNn2fSbokwxn5jONrWE88
LbfZXiXPVYnXEQNqWpShPNgwNP8rkmIG/AxcLNo38dRMOjcimhe2Uw0cWbuTtVIs
B7rvwXnXE9F7LBm4UevcMTl/Rzv0qIm3YsfcOp7aVaT0XMOnmaplk40IVw3wwFuS
AljOYAIsHGyHB7ODLM+VcM43nuCsD/tgvM3UfWyiedMMLnybTqzE8oFbpVNsAhbZ
GA6TT130LrSICbkIdjgRpbA+yhwBfjRMDeGKfP03Dz2UGwHYPAIrFM4B0T9RZhAA
QI3ey1I8LLuHTFyg4Nrp53tWmSoeNuOj56X7zFdCqBCXCgS0bkdCjmgNp/agvFde
jpKAzbt+UVezBVzX3zdFlcyvm14XC6iJaIk8KBCwcrBA+TW4Em3Yx2gcRLYj+pD7
DkWpKtymHQkCCwDYbdO1LD6CGBii98vv20MZ7agXCLQZAn9DrfIDYVc3Nmz/OLGU
OC3Tqe6IzxXaxhafD9QeN+sqyyRnV2p/xrp8a6wADT+URN2iXf5J6eg7cYhbidn5
tfaPTEX904MVbJZZuoXin8NOzK8YB4dyWdiSjUJ8eodru1VthqCa7gYmJuuDBILQ
G1fyNe9a8H+GzTFjo4mfpVk5CT5Mz4/r90QiMKUo//IsaxaHtOoqRgj1eLFwPW07
CGf7S8RXe87g3WD9j6tyHwNpXmqHwO14r9xioRVFe58vIhUo6AP2yJulaXifIoGW
aKlrjnPOFxDJJAhf+BbZZUah0mwyP36+OPd/wigsVzEudxCZGMlnNuYpAwz/BpEM
CnD0ancDnAkfGsWutNV5i+Rk3TTALRiIBfbbhhWy+iORjj7q36OsB4cCzqFmKKwf
i6s65bSKkHuNUGFFN9fm6WRbEP+hFVjNLuY+QcelLrgbVT06eM0ECDDK4xrP6B01
A/q3WipoAt5DNT6xaw7GsIzaP4VQQZTyCVeGb9OfHJ6eYHu8CClFrkfQLFuV3azL
YFOklpcd2kbGu0WRtu/vtcb0T/DDEnXGHRDHqtR6iMJY/vBguzsr/UHANjQ9QZ/o
9P1+u3DAIBKFASSCAY68/Be4Qjus/qA1Z8KVM8bXsStSrr2GiPWFEjPhSgywGeE4
n2FZawgKpmtLjH4WrH24uix2qW66R0jdee3hQpJi38rS+S3RfqQlBd2YiCDGfIxM
aaA6oT592nAIa5RdneUKHew9G/hJxSNouSvVlBles+RYw5kgiky8PwdlUIrcMGSA
CFPZn4Cp62bZWf1YApVx9nczDdoYKNkETLuoqhjIpkkWcbtq2R9+XWbFXClEYi20
RQq74QQ7iMxCAo096KxVR5lWl9kZ8pyy7IgNLyotWsNs/LAul034VvUxIKX678Ok
C+R6xsyoO8Ux77Tx3Cwe0njMxegIHw42SWOdIoGl3McE3IP2kIMxk/SxJbclCJOD
kDFfd+s1UaZaJVd+gzTI799WOVeWb2zCsd1kRC41nTgJ7CJcSmx3Iy8WqLuskjHA
YTrYZjqX9U9Y0q/WUoKbIlim31uNlsxQLruFrjiMuOCpQw3stUT9otloaW7utOGL
01BD48M/loZj42h9sWPqR3bAPN+R7qe62GPveaoY+/EI64iVAIbAzuqpG3NBPrSj
OD6yfbxCymdx51vxktcxN02egfVyDBl3kxEAxcIjiTlc2tTR21jkz3q7Qxpd0jXG
Jn5weB8zgU01CC9t0o7kk7dCE9R8zKN4ELV/6hNF+7ZB8Di8VCUqsGUFb5UKowGV
h+mNQnCdkDS9S1h79+KaGdw4Fhk9HwduQ42MykSGviD56wbAUgLMNkEfBpkdwP4B
pk5x4+gCPMp/9bKdw/Vc94pp4oXQNk/v0IdgCcUFODKAhUGasln8D9RTALSJwDEj
f00y9IYRm9rH9m+SCAHQI/hh06uYcg+21Z5TQdR4GpfPcunE8qESck9CwD/lJHCL
P/p9PyBVEA5LlrujPMZFEvbCIIAYa5DAI1tIHSTlMUnWvBVALg43skebmNqLlBze
oq6KQj3opHs0VyA4D7Siuuk2DVkcJpQc/dQ2Gk4bmWj1lttBR+Z4rem+Y9Uv3h+O
uzMMjsB8dpwpBTdR+mrcX+FONPU+wIA282446kqULfCSsQb66wRHyBFpRilyh+kb
FCr4ybX8VDiIxPdpDZVFE2FyQAM4/panKMl9esvzSPM0+KCLqZrs0SLBxLty/p/e
QH4Rnqu3b2WLAX2PzjQq0O2I6saLHsjXVgqRbRQVbHWCQQWimYZBSW1l35lVo5PX
7+K0F3sK0XnCcxKs4jkHXw8P663YviX5jGs8Gi7FoyjyoKAPfT12GLaGlZUMqUMl
XcV2DcKgiMIXA+dybTeNYJaiDA0BS77Ubyj1FeeCwpvhubxAoL46uhIFnaTPo9MB
uxix4bXxq/8Az7onaWy4LE5ULpQ/Zwkse3iOOS8HZ8GweixXlRsQA6sTZ/i4GIDj
retIP/5IdF8OTgCxb+YJlAc9lo8F1xwJ6BtkbqS5FcFAuQbJaEX8VtUlL2+J4MiU
JsXH5ThqO2Y2N9fmuzUHn5fJmHhWGENqIq7of+ZhM8TT73fQFLZPspkEWS7ptMwC
QBB4x0OnTD68JAk22gY0qKcDoj67ofsHPGiQGqrww9W9mUqDjpAkmpdWzCC7n/HV
9k8Ia4BB2Hssqj2l9bjPPZuKjhdelD3vW0SRj45XxK2/0RmeyweFjmS142IUMGqd
1ZGhROORf53muEMU0C25a3bmK+qo3RFK78Ogb+XAV3FMRjnClSKzAb+M9METc6th
GyfUDtIIUXSMYXb67IcvBy9Y3BNBIEW3+9FW4GEZxeJiUKfP7X+uquQ23SPsuJv5
L6mw4Q1r/VnqegD3DpEjSOceazLzA1R9ptF3x6//v0Wd128LdXrKmaV4Td7XOh4r
1qFRA7hthPVxGsIqiT+bBmIhAkW61oCCvf8EgeSUYhPjcme0MOCinADwfAFkpAky
q76mFCVJlb53Fj1mQI33ln1MJ14pqVef2awYpz97ClKKXgUd2YUQFEYNAfFhgqME
9QpdBM5rvIX6Vy0ZCG7TCfInRVjDhKbRnzso1KVzS8CtceIOYJxluyRnoaXuPaAl
5Vzcx6M+GM4M38O67sC78Fur57boGu3HzFBKeZYzz2L1YwxPTOx3zCXh1tmV3c7Q
c4Qb417rntM4B39ARUUiC9lVoOO1PMUt2YNvwe0cdeJzBn6CgKlpmxC8scnzzw5J
a5qsojjm/IqGy6SdeqetBsqsLRYeALTrXy6KCW7+80OfY+106sTlKvsbuGyiIoX7
NIWkL2pIZdIynUY84ktQfnnfe3/wcJi5sSeo0h6V0dnVLu3Hlgp4RzB28DBJobbg
dsAte459SyMFnNDxTyV31EqERGEum4pyi+TnZqj+i86W8kj+kRGnQKfei+KIzE1F
nBcDvr0CCUkUxHQXv0w1ZXaLRdVVShQ467xJi28BlgN9HjvqNvpJ1NMraSCddSFL
LT/FGEzUkJUh7i2qW4QSK+7Il3dp769iM9x/q019UWTIv0Pq/gDeNZnCxO+FJN6Q
o/KZv4iXYS+I/N9EJgaK9RvytloUemLWHNB/OjBu7ZsEEcOqQOLDf+PS1nkgY6fV
fnN/KWma9gW/R+LV4whoTNp9FKRp7G+iFOgJPWRyiT7w3yMr7bd8izam2Z8+ntMO
D3fiUNtK5RxtwvR5DRi4pj1dK7VrMilGsfEKq/lRdtrRmxGzOJ3wbV42rVKWIu1M
bWEzYipvBP9tXJ4kyrmNzI1muFhxMm8jvE46H/Y+AfqBg4saZjygMD79k8VUsbYM
NDk+pjcQHPVmsn5BRExrxpgnlDO92UE+s/KbMHfk78idk3A997fiMAQT/XZGb3S7
RnQh2iBpAE19/8GEmYy25wAQrTihBTqdvKpM+rYZPvdCntlZmyGMxo6itGgVSSQx
Btb/e99K/DbhPsNBtJD3eKOy1fUReVs9HJjuW9VrCo7cx/Kc1NjoPofWyZRcqXdg
3WucuqN/XjMlP2B6r7ormAO6EypwL6w74COe+8WH9ZylksGDITQoUFwJHVW01XHv
2q6DXWmedr0oQsykV9FOiFqOYDdc0A9WqfJM3r1rO3e5efM0O8TV+jOnMZadl7hy
GHgj2wxOvnaXmTfa6Ct30KffLbTiEVS4Pub9vdnaDvgp8IUVzWMyPM+GarSYVvY0
PVGZekLuPEwAlJYFSooIV/o3vLCBPkULTFjXOKMyH746NpEqwIwr4F2PRSeGq/2y
j2ToRKq/6vlQ5a1HQyByKU+bGgyzCRiEUsPm3dzSy4LATMm72aicA8Me6HUM1hki
FTUNu3cLSyEyoqTAY36mX68gB/jshQzy/if2TArM75nWTlu/ATZSiWjB01hIhZzF
PVUOcpG2IbMUx5iqYNSdWM098GQbQDxSl3O3ujpjAs4Wef542mlpVBT97tBKGHrL
GhAa5Wkudp0Jf/4AtXyU1T+yOx1yM8M9n4KD7OcUGcohCYujy31TXFWTgEqz2nrw
zRlJ6/fFZpt3m53D6jft3n+d8sYcvLcikWWoYNZikF9Q4Ka63pQnHMH5+7O4a4UY
IZYpQNDKj/OUlGymq/c/4QmNPhk5zuvL4T5JLrY1IW8IyXn+p+xJroxA8gjIu37T
jhDsVtrdl4zV0HkV2qGoLwvkLgSFgr9b5jllb89PIKrB0lNhbqOgBrwUK1SDHWqP
tJUjKIuDMxaUHpL/Xupz6ksEJc3ekZRK+Fjw/e7rTWUV88cMXXBGLb/tPizXpunl
D84Tmpk0jMku1J63IJhURXM/dlmvX5gLsSxKGbDc+hDJYoEDc7fwbO3N6kCBejoj
pARgzQc7VNMqZ2i9owJ3C/KiXHuscxAXnrC3hipEZgOEpj4uPZTvf5KkLBlmq4Dn
Uga1W53IKBeVdJYFswDRZqBNY9Mk/nBD7Xe7pu1Ea0TCoyALWgggETbWUxve0AVv
y8QisMiQbkVmRo3/wpspA7rLnBKJB90QvYcTPzhfZE3848s4jhPt8xDn4/twKlex
D6BQMyceGn6VgvCKnMQXxIXfueGkQrO636KJ0/xBgyvJ2SayUjahTHTPINYGh901
JYlcoiU7ch3ej+8adqgVebz1nHx/UCf37xqYSEuZPdg12tsOObCoV0btM+gqP4tN
ksBg1GbpIvbVzkAGr19gt/D5fNU22vb36r8ZSP5f41W9828p+EXIH3y0Xfbm1vRo
lNdF5t9uWol2q16eC3NFFRhDnlHMSVAGfv3g3DMtu9aBWZqI+J/8uuLcu55ypfsr
lEoZonpzTqXrM+HdBI/Qeg8JoSQt6FmbzPKW5+i6A+faPjFuRRJYa3NnTvkOl6bb
lvsCvLsKiPcpXYy7whDLxBMG9hYtwGxNE7ZIJmG2HcKQaOB2b9HiKqjIUx5EfwJC
T5TDA5YhCknThpqgE0k/5XU/T630UmGwPM1RvranEuTHYXGt1/ioTK9ZdiD87Yqk
SldSvNQGicVWlGHWQFhcq0YgdQuqeqU6A0lI1FQHqTURNYXSTGqKUNtbtGCKG4zp
Jp3e0eZvSxl6DhbEu0L8zfIa2grYY79+WC4MoFbDK1Fa//PwQsYm/eBAuGO7lqb9
/HaMGTFWRJKRYba5nCisyoUGqPO1gptt6Xb07OSfr7+rD7/3f3vagIQRUikF+0J/
D6A2vy+YLnt0Lcbv/dBFqmABlO2jBQZmTV1Y3SSOL/NROsdEA8Go6v6JEmKalI6/
2gyoBj3EO+lSwJUYBCJjRZscRqDu9C3yBcSalFwL02e93s4O9GmLE9ebIwNq9MXR
x4nPkGryL3ggSRkivOCZ6dDpIcWWo2ASBXJchf0BkNaWBWALZDVH/4/NhevrCIBO
Qk6tOErspb3+H5HweovTdVaedWLhaRN/MbSS3htAsVSkCR96kXOvwi2SWo8Urzqm
wO9zL/cw8fX/dqwcJ38O2Npu5uhU+2X9qWUy7M+86uGQ2Ir7MC9xDDillE9vsd5I
lMdbHD8FbzIwFm94eX6FDXXeLt8IWokYo1wM6l+waZGvc34Bt22O1xiIrMEY6tvb
hFJfwwx2E7yYAwPgQmp/scjzwExEJCobYBQzsxjZpOHaFvUl+dBVd+gbNLURh2wD
XIj+NLupD/id2bo1zxo3u914O5ZGDz0+/yeo4lavQ/wFt117u3Di+UHe4Zdo0rip
Or1IcidlanIi19B+TWtUF3EteHscGFk3vVBooyarI30B3m+8ym4RJrLRbLSLuhgI
sYLQULbswP4xPrFO7aSnQdQGRxSMYmZK19XK4T1rHlJVGj7fB3hs+snMvNp3cdel
ZWJoUK2G2IUpgFkuJEVJt/ToJPDesyYE8Zl9TmLn4Yjl8bXjp35fHxqmw8uajqCh
6Ag0yIuJuQh3/et2m/7/TdFITGvKAEORM57TRLyP8eUf9LitQlcxHFGzTC1nT4wn
zrDqvIt6Q0aR2wbelJ0oyu3A5C9X7wUx0p7MhBqdNWUcZmzq74h493LK0wPCvA6P
Tl1umWCPSK81r98CqbnkEu7pn5IiGd4AhsFhJE4YOF6ZnWY5YKcq0jl33UAJdwIv
at3PQj2IFftYTWwRVBaLZVAuF7MTMmKKQwFXa4BmerIj1It1LXNW69DmwlNkF0um
yppOS2yVgm6X/2B1CcsiPOOTxcrCqYs7nsrSiUHeLC5LcX7xGDaqsPupQKmtIqYG
ekk903MwiXlOQYxugLE10tGG2Je2qSHVeEC9uREuScurFjM9FDPvndq9U8eAtSsu
f0Smkra+qRF3RagIxFB3KKSoyaA2Qo90B+TQ7kmdUmtbp8tSfm6WdFNceOSUiChB
mVHKKCXyw/EmN5dGDhR/tIVShGTsTBrVdvfbIRiJIOL5xHevt4YBmzpF2WAZO9VR
a/RdLCtqRJa5/I/H51o1Jw/VNwbKMayQ4qLEYOebLOOahHt5Z76/huYzfNLnoadI
dnMrOJ5A4OyJLK36vGDlhPx+JMN1GGVgNeytehJeDNUldVfY9B6L3U/rGNf8yafQ
idCp4W+Y72MN3goj17m8WAVAtRVyO1FAtQElZo3g28XkgbP2MciG5UQ7/BJSN7q2
pYyewQwMlNJPlVYCKBzO7C/0W1j5HuuTLsNl9WdsjeiqJZBRSEHhQG+z48RoJIJk
gyPAYxjfhVFMbNtPCYL881OVZjgjIamR7gPPDp0VU3rOn/cig1zy+Y8DZzdMTUNp
FbxC1pZCIhGFQFHx7Zsr6H4gtWOOAvDDpUHNwl4Q/hiO1Z7aIxWtfUxrCFWT3f9M
bioT7dIzcSOku5ytRD9G4C7BVbvxesTsvj7KXjJfjlHPv36PIuQwMLZVpHp3gkg4
LvZ73VpUzcpncen0EV/7T4dAyxyhdlvTRShgVe3WxD6OATkzeNVC9esdzaf7fgDR
RXoEI2Xg0mxHKtIZL1aP2i0R6P9lc5UM75Odgljleq/hvYr/ReMP6CzFVlUHD1m7
mqEe6obsw2Q6iN5jkKzCwynBVMrrlTGVvVVh+/78nFvhCs5LbImSQgCwmLf6L+Yz
qmLiZeViIpxK6Hz2jG2xfp9aVFEFrGSJtwf6vq0hV5etg5ZK1Gc9gX8zwR2dM82o
v5XA9SyC0AsuLnRH8zy8qObcQDEeh8h26q8skOOcI3Gmk/Eba195BKTffVhAuYQ1
hJYWBpukiGzkfMPNqTZLzdX0nLY12A1l0rypLBSlyLxMB8OGgnSePBhtrVtdOZD+
WNs+J/BtNKtz/U/eUA74yUs2DpAEHSmjjXyQbRhQ06NcR12xyU/WVylwX0SKeQeD
JB4ibQR0INOWWRe0dXSpp+2C1h2zjhwWuNhHvMw0eOMXrsOI7+NQfRVbjBLSd7tK
dtKqls3UbvT4M+EULQiWpL7vgK3H8P1eE27NaxUXF+rUlWBRfi7UT1XtR4oyGltt
dLJ+dKCF9boiSoIlNwBej6xcHHn2HX5Ke6aotuWK2fmg95rG/Z22Duq50dtQFMbs
JdR2TsnGKvaSI7AwTfO5IanfZlG9I0f5kyouePiipppP6QflkWgNz/YJx8vrqOYk
Hqgfakrq97WI3LbjUNIAuX0luwAcIAay9BgIMBnfUuq6ielrbZg9oFecR/jOy9za
KgZ1RGsgZdbaA3lwPghl57OSUC7VhKX9ZO6CoviUer8eyhVybPUQVhH09m1lA0tZ
cqIZ4MwDOE2oBx8rME095ExKI1bV0vN2TfoRd2h/TaFgVZv+sbo1Be1kZBuyOXD8
nnc1kuDmW/ZxpAbE+2b9qkuL8vajOVSV0yiQdWRKSsqo5YrkhFB8P66I/QGpOr2M
0CgMDkqtLzt0nwohPbEsdqhZs01EBGkP+oEzVKwAblXoPPKpIrgZDWQNEOBeHFMD
++Zg1t3Me/nXSYkRqCoxK1C3TRmC+QuGKzRqwI6tZXl/BCe+SvYPBfbpCxGxezQm
yLpYGp4uBRK4KL9r7E5l4iVvBwTzBhcsncWUK7t98wyVNDhl2qPaMYyjodylCs4s
PJXfhI2Ol024EMvHrHgjbiIYzoY4DP7V0QKy7DkWVxrCGHtLzaeTiMMG9M+GRYRX
cpCdgG3GgVaEvyRjH33I9jg/2sX6UFcOLhV1Jwsfl2sX8SW8Wn+hLjvzmMO4DVox
bZabZ9mg0qyERmmGmhCoX8iDWwrAZLc/XiWkmmREzVep46mx8RVjbi7U4iXPJr49
59J16kJO1O6HJwrBMlqw0GSIEeWiaiBUYF7fbRkPeT6lW8exyzrCnHoid6Sk9hH5
Qxe1vN1418rvPzrcY+IALA4TViDi28B9OX0D4Z8fQivJoqZ6+mymA+LJvDhfgHJf
4yL/e7PIeSOeowlmwQji8LOUKYh0+urpdvZ932VNrg2boyYKe/MxvN5blNP7EcKo
FmwGMRvv8Djo0Kxc1LhMM7RLrtBQlMv7FPKHiBaUqQea322UO4nLbmXuYDVAob2L
FWy+i+bhRuuXiCj30JmQWXuj9p9Ai6/FPt8FswACVyZgXWlh/lKPCmJitTE4VObh
qquls9Nqxh3ZD2T739q6K7BoSpkWk/GXAAs2sEacwo0xocYs+4eCiknINc66ck/+
s3+e3q8jd9iGDwVTPiRDCwKTqsDXnyvtEq+Psoz3x0Q4JQaqbUgfdCABHA2geWh2
Gbwej9o7sRewKGrUjQ8HjG84asVurRJ9OKsnWD+FWHlOXL91kni24Oveb6wlv77j
q7RlD97xso59ovgecB/7HxhDFX0CpThWn4opU5kvUEuNn1ZQcUB47J3eSwfriAfr
M+pcnn/FcnlPMYGUrpeSpzbMuVDWNsYSXh7AjxYBouz/jyoNMn3jwcm0tBSzh/di
uAnMxUITp2+sin3TDQR4Y10I8eqeZA5Xr/1IKU/YScsjVmM0zMG1yWoJC/QWJtuM
Ivp2YOgZFCJUW0a7Qk0CAdgkcK7uVmsLYBtSIS2sBGem0VSvCpcwulsQF39KQZr7
tGyqRah8xz1IKfaHPwwDpO7HU2mu6bQZ33JGLcjxVk79z1GpDYHPP1+/MTCGYE+b
SopH5cocmiGBxbPu+aATUZNnkFiJLdGFYXudI7SknbnxewuRfhzDEDL71uNBZS37
CAdgwT6gaR3rIB4Hy+ZNh7s31uA9bwlKRdAbiDSSRJCkcwfAsfkKRs2AjDg7AfrI
ob0DO6vVQldL9H3/hvTc1h+ImkNRVfzU9XaFyrYNS5uPHPdY93JVelcpWcBD9V4E
BMJBsYP4mHrvQQmRHdsYWajdVxFc+z7VXpdBHWN2DOjDY+TOB9f/zUoweVu2IhuC
aC5igvW7tr/uR0FGLNebYftCcXsMA5YB0nMdWeG9kb56puYeFhNh7GKyqGCgRwGQ
EiCQmQJ4q7zimGbrIKN5Ebt5AsRblQbDvofnTn5CICvURenV6R9FxyYClJhlHW7W
jKhFvkSvyzahnIcT3uixB+b/BqjVq652Se8IwXahw1D9DQ6lcY99nemaw28+UIxE
1aaTBhu+WF7tisNirDCtZ1PwilM18RBMssMhUhFr1Qxoa+dT/qxl6vZrZ0ExXef9
Ryn/qDuNrW/KNGazDmgwwcBixY2ew9GWomiGtbHzaUfnY3u3/L4ifls01m4VTRJn
5FCS5Vgos82yG750lrkIgeBMGaZ42I8+q9X6FjzbKLfkTg/Km1NQbDF0ljWyVCer
SbAZi3tfAN5eFuOef6qwNpjy8ilQOC4Bg9Y1k0Ts/hITFqH/x1qS2zH8yk3S0cN5
NKSi6GsmYHBxJp9UvfuuLpKtb2AldFJnPN/kTyCZRWzVEvgmR9uYe/zp+LToRAnP
jm2SxGkTNkLjXUVzUTnlwSYiAR0W/JdmSARGPPJobefiGA7vOuhfsUgy+wcAdCkZ
fbBZFWGhp9EowSE2kqBzFMk8RfpKgAa2XUqZa/2EGjXjyTjgPizSVFaERkshwErb
X/dO4cmFb9C81IqRGMzKUGB98HEamD+wYc+FLBEmvwd+R8SHZPMMVSgNUqLgASaf
bIUkBtLZc02hHBWBHU9/TKDcEyhjcQGK6VXWwybzGHEqqBKmK+pzWY0EiowEBuCy
IZQ+3/gWv1dJ/fRldMRtOeb+zNnDCwJHaqNmmJPcKRH1YIAUQx2S3/fnG+EA9hUd
5qfUvCLNAbCro5K7satkgVGYM9Hhu6sREd6oYAYvd1dlW/SOWki5oVWabdQdktNg
KH2xOnZtXLNDE87B8ZeRK04WD2Iltfg2ID/YLNu4dr2MXTwdhBRCL+bPyygnn+GP
qwBZG1ORyFStUXKe0q/6EG8rLhsxuHoE/lV9cllZQbDle3+i+1LHCGrb6o4jZ0yT
e/+KJ7nhDoOb/qrJY236ZXdvV61Mt91/KVp+XJAmYgYNYFSXKDOt9JSjFF01XV4S
9YTY8LAy8LJG8lnl/3O10ilNVil8cwXDs16upW2pz0fpJ7OH/pTbXjrfuRmL2XM2
RiYH7fYOYx+2bgXilLJYNIcrySIpiz/Ihg52HFsBDyCS58a/qNjBxTxYva4K1Ask
VV2aaDywboIO6+ez6UkxqotncgLiw4DgHJWxiSGnCj4dw+i8i22L2GDWLMCAg97U
iGNKI8rnqYmtnrcUjdaHwSYRSr0/1XliKcwpnBkzZGJ5bFbVArG6mRmX2KJNGVSR
D6plqcasLZcfcmT3+RctdmeQ3qbF4bWozis7UahMitASx+cLqvC3R9xgcUxE45Js
HnBV616L+9R1I8vv2WMQ1MK1m/78D8cd1WcysnpBMDSuSwzMZB+QjKfYQCEyqOdu
eDVD+s1hXllliL+q6lQEsZSo5PdQ52FJgC7fKW7JFfymQ/rJOzFZglFjRzEnPD7X
6sgVJsLp5RsNo0E/iq1oeRe1kIpCsdOSxrrUbyyCNXHXyJMnHZ5+Kdf5WLUN1SBq
4EwpL0KKHhI+mFjmvB9X6wkqdaENSdQCpEuvkYHL+w2Xp4Gnzvf1Ybrd7ftuj23n
hBTJ3IavyWeAmTfdf7PhImkKHHjvaDq+ODCE474yogulD4FIxKmmJhqGRyxzi3pV
yN/sZzolPVLkG78g6bk/fDdq+DWaDxO2FcpezZLLrikIFBqRW3DJPlSFnjO13yC4
nCwb05ITwNmfaDAa1WjrFMID3dRh8Kzjr3FVfX6ea3+M6latySxP5Gp6nzjURp1G
LY9q+KMzKBpfq5deOaqaBd6ECJipuJUZT5lSwleSuGZYRrdcgL4Ydm3OG9PNbLP3
6yGqT364W3mjVqKXuxgkNhwDUaahDAwxFC9Aaapb0RvNENhObgAENetz9XjbYy/A
kldbFEZ42REzB5pSS4znDGPvTSyQXjmfi4SuincoSjOc8dF2OrIXNG7pxv88S3QE
CfPSHNRoUBNISH9TQbPfFdeosT7l/rhSmCFlSrp7IpOHammAEca2kyfr97BLEWyB
w9/A9Lzs1Y1ZZzp64kKRmk0QliE7xT6uYWWseVXOrawLevRmJzyYOk1FIS3qBUaj
tppysceJax0ATVoqi0Fx1kG32eGDP6+hHWJMzMNaqusQcnGbvvDkLKMnhLU2yhCB
yR9CdlB1us5H5SfgvVK7mRNbGdVTh6SYTSjLqP1nUyR0/+hNVIiY4iH0VzusWeVW
n1KHeT+XXGB82H1gAv3fVOswHFlLmya3Id36AbTVxmsThSW74PmX+SbVzCIMnxxL
jkoGbBAuNjEulHKFDAa4a1cyEpMFduvZqhfbs+UAZwBNAEUKR3eKecwkj2R6m3J9
gugYBCfWIdeQCGIDtJNvxOSU/zrR9HgjZ0rb+DcgIeWW7Zp79qX/r+/dnMn+EQ0O
lcQrAyOil0lmWVEYD+rO7nT6dENqdRdnWLtRMchY++kKReh1zdOxnvR2Bv8dHFRF
AFKeG8HDkUqbmjq7z79ghrOAndk6dwDsm3TV3aUGYpo89nxODRjg1knGecaZaTAg
HoHl7/rdj6oco+SCJbWwS7LVvy0XZFT9rktycdxSaWFz5+mZZ3eUK2dW3s/+uR7g
CAitWmpH2hC5qwtDcASDjC8cdODUvTbLN4sDdI/nz2OGU74Aoa3CsMitut0Qgjuo
cUS17kahSidSp8+VUhV5rRy8wif5Z7z1zIMsSNjnzdGOAGrhroueg3uEl8ToBEHp
4oXMsgw3ViODSpgimGcCm01HK0d2AOKXsiDA9tKlNg4LP5lJdxQC62Xjp3o590wr
/NGzmBgqW8WSTIFM/+tFSHxco5/pyOm95JMs1Q72nQaywUbKAcFxDsUB5A1npq+t
MOo44aMU6kyvrXnfCcpNvNzoP8XtnufKlqnLxouoePTg1WoPlezkl/jml5oLg6kx
Ow5SOJET0NiB7xTBdTFLIsKn53kxKN2pfMv+LtbDbqN4+am0R0BS6NUMDydoaTiE
wiCZhBTyedASGIXnUO5ZR0GTG3CpHS1etNRs7pp8mXD5T8YECpQ1rRK565FVaD5S
3+mizXiG7CTQC+/DiO8ZOOGejdv7qjUxbtMnp4wIMPELdUOxbdRfopMaKlAwye5M
KZ5AK6yb1iWRzwgkhsUs76COQn+yA0on0NiBd1DtExyQ8uoBkGJKD6j9AG21CoeZ
g+dgBd/b+DQa9QUPb3TNM7zNxy79i0mT28t3P1OnGtyYzNALNB4H1H0lAxjAhvRe
ZZul+XdfXSY9hyPxvUwi/dHrjaOC7hLOHOAcdZaxRVcmAZ4yHQZpJoI+CUyryzAc
BSBBlC5j8SM2F19b18m6Q2rkciMxsxXipXNaHI0yBxijCLXuKi2+XkP3keIcsv+n
YgvJtKhJ5Ko4UyFgvStlPdgHQrPRQCEoDdcdEBVvqQ98hhrWxHRi/vLe48xBn760
trR1vrZZeyspdcBrTn2YBNIWJ4H2pQmrXgEtDLg1wMpAerMpZumAMBpR6rWnQ/xZ
yuK1r1L2wFTaaZRZWkzzYLriSHJ1xeUw2VqMHmItQMCXKMvCKhOv8MpGRSgxriXk
MatI9BRnro2kVenI74fZfawYwyOoLTlazW+lQDgdaq0S759UaXjUZscKF0CmJo5b
cCeO+EGWiBcl/zJ6EtppfeYxDitigLsYKfe5gPstcQKztyl7F8QmCrsqcYCHM0QL
lHMP3r9RaB9SAy/hY0Eg0uodbZDzFoyKY7vg6o9vawNgf/DaIrO7p73RWKJlE6ie
t6GC8kMWyJixv6mfmKevlGNkFDDMDkWsJ3sbp29TiTL7JfcYReKeWUyDPwogqTwG
7PjvLHyuh4IxjbJ+tR3QvstzIdmMZbL+QjL8U3Z7WksnCcnP0Qmb7ixZTjj8ckyo
STBimVpSET6bE/VQoVplfhSH1D7GVfJ67ff3mQF5GPEL5YodxieWl9RxEHw5sejx
iisKd9wJHEoNhXWRTfNldnUGlCpTunRerYXUvXBnYC1xp0mXR5+Ou4ICRbw50aGS
QXoo1iJHV+qJ+RyHxXfEyDXjcIwrEuaKkM2vn4XmfcKDJ28BnpXfHEk5Nbs+fET1
lWnTma911mxW20OWJj9VX7RdT5Y3Tz+AOEV8aabPuV5yktCY2nUWhmQzTJWKe0IK
4Y0f2Er2qtQECdPdF9fdllsXAznx3wQHmtW2lPLMlo+CzQ2PW9BJuhoEpOakwWPJ
UGb6pAH02J6wiwRdU4qZYIXb+PZxyXWl38m73YBOZGdB4ugpM5tF8yTo18HSpJUi
Nifu2QV4fq5mLYekFkqgdk2YCWK3KFJTTTHDI/68hpMzPy4COrSYAswCUb3vrCBN
cjJAA/skBWP3u/xPRZ6zqdaQXdIo9Oqudcqml8E3pHOKe/UG89Z1OkwsYDcXIwf6
5AYUfM3EGtpI6O1TxzZ0IPI8R3mE/r2TyDKs0vm34G0R9R5IRc2yJ2OXvdWHdX/z
BJrys+LAQVoEPOsD6p9peXflxFUgRRtuz3E1kQE/7UPJC8vvUUczxNbz08kdcqIb
aJeCpKALWB9FE4P+NR7On3DN903eE+eSppgVtuZPeF9F7MZsdLcLb3uNPfxuyRah
8gRu8Y1ldevsKmaFpXwf1LoVfYkHQsjg+hkE5n4Rx1FuIhrmAG6QQh49sC+d1Gun
ZDkOYwq2h0nTneMPP64zU7sFqmoF8gEEhXmTQaTmix8yLt1BYe+2lyvlellsH/lh
dSNBdh3OD/W6DLKmn6zjfBf+dNd7yZo0nKV1+H8RSfC1eG1g4nyrH4W0Ict1v6fm
F+Dus6JCeNrd+rSpaIL4IMKTKm3PV5o7N3UVoF0XGOtpAJQu7fII1FWYveXwHB1x
CxBAy/eNheSqeD0V6uOHupPjT0hw+/56Jn03kLz/NyNYjRAvCounhUrbN29b8Q+p
L/Ysm8aSPX1JbCggdZl4EoMs8XFdlDM5DVgveNOlu1M/6ULbrwEhUE3P9fT55C20
mgo4kJlth/Z0uON0iZfDKwbahA4LoskTHfap99sQhoZhyh1VQ/4PCWuuin0wDZip
p80QyWlfWb0BUeS63uP/tR02lFEVPrkyPZqSt/ZyMIyLQmaj5c2kTBISNu6DJljE
uNXfq16ITW2L73EHCSzotzviyh7ROfejO1Qw8Mk12jaN5Qpmzrf/MzAzwXvoTjOH
HQHDnkenzP1R/4ZlKX62ojqQDmFpkmORwIfx7+Q1eLgKvS7BhrRRDV58wrCjWI5I
hwu/yWqgKOIVZTkHEB16aLm5m91pzFKswdc4Kv8YjZc2k+2kQ4djIQqA2qgRrCqS
c/h8JW/o/EBp+4N6v/aZ2yuuB7MfAGfReVPS2SjCyG+TZ9EUv4EOAbQYBBPpSVRH
tRZSHOtin9BjSB0M+x4ZIcH8XRkwPTQbjGjp7MI9X7a44Lwv2aJSYYoxr7Yy+PXN
fx4vd794zDBD7N9F07L3Umq87mv+T6irW9oNkTeCWc4beoQ/MUXE20G3gq5ZUX/z
/QjChCAcN1Yo2nWq3yXMnbn/cszALrtkmROvizKU3N+IPLTx2hCFLlwyFmZJ3mJ4
QgHGwA3oBLakse8NI3YeNszPYkQ5i7UHCCR3zt0DiVn3DHgrO1gBL89FzueimkUp
3rxsyoy+J6Y4bZ7MOyQbRaARnyKp0jFH8ZWnELi45LtqbVWM7odQon1cv+XD0lrP
3IdgXxjQ8q/1EO8/Q7Gl9/kmpDMo6lTEIYaGkOmC8u0K3dtMw7uhdUcjMH0+uthQ
L9TYkI8/AwXNL46DowlwdZYw7YHCOqMOnoJIoN2LUQLovHTnAAud6fOSk2QXD2B5
pjQW/oThrWgZKUIDTsHb1iABWC3E6wABJdEWK/rKIdoddXtYaroztiz7iyOlMqK3
gY6ELiBqOKqajwSKeJ937TdkyqHX4aGrTGvfyQCCcodWk6c8J/1rsZkOFsRhuzzF
B54h8/2ItJFbO4tAbmKyCfno9J+CPNXLGx4nw2H9qGAdQd9nXYfkOQnf9/+MnVHD
EJ0FSXANlmXaDxWe6Nwen802XZijsDtRudFL8uajtkcSJPiMCgrTOHzhnO/LGLha
vzT8bVmS+/K2Kbx9Q/I68uZ6gCnsHh9EMsd9xpDKcRnkzmLs9oUUQwn3gKkzXzmj
om3hLZ3Tt2Mfqev/ffIuY9hocs0Sugr0oWvUG29Z2r+JvjG3G75tQBn/8gOb+bXv
GM8uh6JONa8MhfBu+RI/QgXNAj10krRFL5hSoVMWq5OUT0A0zxW+2ftpww+di9xD
w7XTU7Hpq4WP75aVBICFeFsvCoNqikarH54Oz/GTr2y8kuM8A6XTlvnDN2AyXynz
Xg0e7Rmww71z0s61AV8yeNtPqPwbyFKjXiTjle5SD03yQXX/VmmmP/wzjQBeaIv8
k3Jiqg8SqT5SBIbr288i2NmQ4ddDvOC+F5N/ktRntRNZPESu7t9IUueY+qF2KAZm
rdmxVZA9Cewy1EyJibH/XRuUk4WICzokmhpR/lHuQuzY8gxxlkaXY0m0icDS2fW3
yoJZ6Dob0uqYONhGpFBBEVLoxyKjANCvZDeF5arkFFvaWeKmIlToMqf77ZtvGWlK
UiHEUT6gvDTgA/qQudDesD+gQEgbL+/2fQY8n8B1VRwf+MACAoylHSwtb5zBB6Jv
mBcLW95JQL5WCJsXM3Ly3HPBw8yYxH1lWyCZtb38+MqLpldK7Uv07aPZRnuI3Oe8
vcS+7c+doZpUKSwO8xsm0w0RiKlEVbfjJtQFkL9PhJPg1raMXhUgJ1eOGLsVWrxV
PUAYou7ArR0flMYiKcJH4sb+u0XdnZqRdqemZjcVeYFg5qqbjDDtvgbbbPI2uOYS
kqAzIHKTBGiF+d9iFk97tpjbtGAeAZBnHVb7wuCywwWW/hV8qSO9CHgG6EzvNOmM
ssVO5U64hKZHUFJ+Z7XaYwcwBo44lfXCtnv/nNla9rMEEQa+ZFXxqnUzfsqj9aXQ
gLtIQ03Gl+g/qnOx9iWE/eW9lzqq95S0t8nVKjBz1jHdWPhIdyWERQIvhc6AZqU4
mZSgMM/kwsXKKOheac3DsG15cV5u78XwnM+/yY2faRj4U5akRuCcm5L1xHUtzai4
Gb03+jwsNgNDTWmW3DY0KbjbhkeHRoF7fhsLjmQkCx94cZunQoSEB2vYUn+hNa/S
T5JVgtCmVhYO8BSdjd7bqUEkEM9pAGSi/l6F1lpnHy4A9RKGdrjHLV72UCPK4YaM
fQg1LhV9hcOY8hm0xCalR0s1oBz/A52Mmm+46dK8+rTkT7T61KiqLqmeoMAHsH+L
kB+SD3ADotCl0kt90b1EEzMQJiYsW+udrE20ugatkvGXFAE3R5/eMs5Kr+Z91Bzs
Lxb3dPg9MP1riZfbaUjVNfZAkkxdqQ4P7dE3BFHyohePtJCADLx3+WWVLaz968Yd
sBAeTX7QPzGcg16unX+Jj2rTHKIv0hq3jtXDUNTW3Kc1xvotiDvljLWscO0Bqt18
9D18/2F5KvPAqTT7VsKaGwh/fJ7FpRUujTHCdYg8LUxjKGbw2wLe7JtxGOC45k9X
yf4mWGjiNCU2KetRKK/Nh/trHk8TfJdd6BZUqzDxykmsG6QF1ZMTXCgAaR9nXMGF
CCZbXGr1wWc1oblgN4QfjI7MRUy5SoYHmRebsP97WO94x4PL6PRRcSaE6impUVc9
TR4nLM6B8m6qMxZo+Riot7h18p3GEFeAjFYJMLhP+x+yONDtRLBSX6MFECPzd2tR
OV4bOSmCo4v7J8rrKrP4AwCNmxgN1Xt8OQszCHaoGLZnnNnsC4biC4Qk99deXq8c
taOjNroOXFB11TiSQR9wZufFkFzq48y1SW1ZBVADvPbaqJilW3btOnhmEL0wtyBD
B1FImbRN3n0HUDtwgKtXsaULaA9W40yOfFDWmuxnMiojNHjOJaeGMBaRXiIyry5T
bRn7TYDwm5EaDJb8We4FkmBfHot75N+dKMuKFtyYmz+nQzGMxuRpkmD3Tam57MM9
1/Nq7yYT95YTQp3qZk4xKnQpRhYHC1MWrGKczFQjZ0O0ygR0p6NHz1ILLTHEXvOa
EDX6jr1RkbNCjnfifxoMadzUEHK/UW2ebDlwYfBxVqWAQ/8XvWfoMaQ31uIvoHeD
HMpfrO1A31CKl1yx5dJOTgs3VLVCeI59mPwJDmLBcAezt2yN/CLYm9bgJH61uVGb
N9j1XJrnkK4MM1GlU99nvKoJnEyQT+6Bfrw/akJ8v46DaB3BHZgoChxxelVBuHQx
n28EKIw2yDwZgg13OkHvMoUufI7/ayQb7AV62Rg1pDCKUGcPiSOb7K4qNRlBT31f
bWJGCyvTe06+7eLtYfHClJ8KYxCciXue9r4SFR8ewZdIfzoc79cnr5tZzsUY1Vhm
eo13YXeTJu3UI+7NhY6omtELkdxUT9zzB4toZ5LOVHF8Orbr24tvTluP6J4GMi8p
cu1cDePE/5yQOcTvM4T+/FxjSBwAMpbhIQ5fqDrc6kv/68rPfFX9J8xwuMBXka/x
TxTp7QIJ0LB9ik42eTBvsZdAfj24BN1X2pHGcN7am+6HDAB8Qn1bAHjfOYJqodNy
b5MDvO3XHAD2d/Kw4SjBHO92waxNpHk2Jz/J7qUxMNaQmgoMCaI7A3QyGg4vQDfa
nFMyfKuDD88tBCHRxtNXSJQGYK3nIffcoWlGIBtKTOJpxWBOmh6bldZSDyTpsix9
q4vomeDG6rcADzTzS/dBwUmfsTV6348Rft7KGxKdOGmAGdB/bWkgl7LNm9mC+ULt
Yywq0+VpTEy+uaYj7Ou/SwlEojT4pYEfwIFuBL0EMQOcvnHNkbBTi/6nt/ruPPtV
wKkUxKCZSo/7ywcnfqjNzoUQIu47z9r5yh0s8ZNN4P2bobhAPAAFdZ2Mo+mPpKnS
ee2cXCZ1nNxb9DnREg9bM5cpWnmgJrAXf2i29k/GorYTyNdmlQNGi8E3lQzToK+J
lnoiPYFmogsbijbvAOVQ2aJwqxDRwApEid8iCWK10mwE1D9UxJwOFogozza9yAoX
oAjhpJ1bQtZtTXcYfU6LSfWwdFjDeIXyheSSz4zE5ViGF1kzevV0A5Nk59CvFL/A
BGcIG4o8oGhJ/RFSBTN28lQyEE1b2UgiD9Kvsb8gYfWBTnvExgOoDvtn6dahn7p7
8fS4NhNxFrmRpyweve1qNhBqueWdpz2zJQ3Zte5tLGB3r4H+lVEQEtRi0eBkOxrv
mHCupwf8tPNeExyo5FnZhhNQAvnLtDgxDj2BfCO0t1KVomRb4fL68v9YqQfaBKL5
gf+KnasbifWXUeNrnGg3Kg==
--pragma protect end_data_block
--pragma protect digest_block
HVoexBmKGkBDRxKqM8/60KxzV3k=
--pragma protect end_digest_block
--pragma protect end_protected
