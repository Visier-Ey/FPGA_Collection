// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
1HAvw9+IzWUszk2EB9oB+qy230QXJQez8yQGdjvalFgTdzQI8psX3joBxHxg4dJJ
O0o4e3gs30oGKSx2mxIWyz06MwxGGpQX2zp8k4SblhDYrj5gAQqICnQu4jwP30R2
FBVywVA/QWMG8BJ10YJQ6zgJo94Ni0j/GCZkTdoVv58=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 10864 )
`pragma protect data_block
I2T0D3zJTHfKUwx92Cjk5er6om44RHaT2ZEqPijP8s10hkgC5ARLG1340kuvII+T
5PIvusM/cWEejbb2BcBTngseCIVXnOaY58ARP3dJMeH2/bXhnc9slAvsTCRhIBaK
5LTg+363Kh1l0QWBKU2UHjj/eiB2nOJTCkoY5/PvwZfQCpZbCHJ0rEgfg/Q5EJCl
vjRBiw+P4l5JnqzNxyuGiFVPtf3NxkFZvLr7fjnpM+4TlOBnIfw3F7zdbkc4qDI4
H7v1Yf418pq7xpA9CdhyxR0RGqbT/HAuuucFxASzh83GXX2KQP1phWOStLCKhxNq
jxEhXMKndABBPRfv8vJ3fctF/zk8WdypXVEP1SnEOWcRHhMK7GGXe5VaDA22dMqx
rrNyZxgjVBcPeQOZioUM5uEIHpWyQTY+F6ogwkgzA/n+C4bI7kKnIl3AclAAqLl9
7lNYTQGX9zauArt0dsFV6TCMO6aRrSWtFgtcSBSDkeYK0u5AYT6uhfJXQVQZdRFt
G8ZBUB/BSBauJPaTGb0YMsJUpYfN8O3NZxjG7UmTPOjfDZDp+GUUIx9alrgEWIEf
SkNDlMO2CI9d0pia7uKK1Rs6WV7l38QpLRKMiCLRHCkpZ1ap8PfP7A3Fy9ccmiGK
Mg3GPKNu3QRPpiKO5NxMHzmYU2Caef+Qw30KdIZ50I5ZJXv3Kxz7eV0d4gmITukT
zzGTI/FespcagB0BIAK3RHPjo+O2ODBtQGVJ44D1wQp0UBi6GsXqVuloiEfPT5AU
nlPQer/e4w9AB5fx+pAdVZDqtN6kQKAi4FtODxlcKXM3IJPaA0u7iNunqxNllZ1w
iIzx+AIwFuEx5YclY1KQnq0dOXuuxToDXnQzy6FmH2TfZ1VTIZ/01NY1s2F/gOyc
/GV6wkiIr8gLSQKO5Me488riM1ogBenHeKyfJcfU0aNYEWffTy+tDVSUw6ejCi89
20UUYhQHNAuE1twxRkk9133GqjdinPUaqHKL6ObeZ5HMYXYJe4qu+ErcyHB5zyCZ
9SJ9Gb2Qg6k01Gk7K6DfkBDUx+0BfYvpFeJrOVmxPFaaSHMQ20QI9hzaMgAHmmKP
MO5QJLjdtjEMJWCPKC3diySyXr8rERt+DC038NPk9siU2KNTrgjt5PO8XtOejdxO
9x4KZWmduWFDuXp6gB3srqmZ/B8Gg7glYyl/rlWHJoc+CKVsuhk/TJGceuLhwav9
UGhme4Hv9LJrJeJikO2igD6SsmSXCBLSzV3KEMOvG9kMe8/V2kdHaZNG6uV4FnFZ
aAcduLV61u0n7bh7UEfhtoMcJNWhWfzVUx+xCUOnFZSmP24uKcGGii6i38tmLMyM
Wl/4QZaUNLaGSo9TShBf+Nv/TaIfc4HO7s9UutwX1865ByFq9dak8bR4AsYoitv/
LY7Dr5B18KKO+lVaXIRg8lgCbty0axRa4JfgEd/MseKsrn9MJyc7Uej7GCdPcrwm
9B0uZUN5RTd1WPY4kUaiii0GgQyq49koRNTf4q9+BofTyMVh3c9FhOKHf922CK4P
p8j0HbpoBh1e1nBRRoG+cTvSGCiLeFSjDbkoRwZBWeuyNu3kdbVyURgRGwK7VcGQ
5lMeFLU3IYc4paruNaFWdyJgbCy4UiIiT/LqqsP1gVTz6g1OeW5ZvFOZRvWMCm7f
Ujq2cBRilqFae5ssvRf3rQkg9mudk/LVG0sv7aVrM6zrULSnKwCrAo8tIrtSj90n
wm9CFHn0ypWgWRZI5aoUqfAMqHFixpcERu2UYtuogBiodHPmr3npNx6Xk/s1aNSJ
/dxef27EIPvjEv/RblhS1tQyiNyz358TBsuxuFsFV1IBrNGehNq92YCDM3fVCCi6
p5AMO9pHfK4Eu5moPqv/CrSqgDbzNmr4HeXH7hgRtle1t7VPyPa9rS+b9s0iHJg3
MsL/XsGeDS7AVBReeAF1TboCwXBkmRlz7H5UmbeOx9XFEs3vT8hLPHhyQU2WmdeE
0Zwz7vverx+wA0F854Hc8Hul1hJdZoAcrsj65b3LGSRtqTeDinvkchl2Now/mdmK
gbQ6Fq9vN7TzWveS8eROtPwsRoC+79p0ErdRye/NBVtRzSbkNUU7nFX8G0qwsjmD
1v8SpxkiTiZrl7w7YI44ZJtvnS4pYolOrxP6sUM+fUY11H3mpifRIiQ2wZr2qyf/
caHLL+VB3Rcy7VkNShYgUvChWDZ3ChWXe0JQW7lhalmlktGeUu8FNkq9Ho6M9ZId
Z5hmHW+990lj8p41w2GuyKHBHW6+FGMzuHYZKBNUT3/Z6Vga3uMJ/7djc4GxVRji
ZQxoA0lNSQIGksmEGaItDru5jWjrf9xbnpqjVnyv+dQe9Pez1SGTzSqjk5XpBWMA
gz3ToXOpBfOq5lcK7scTnGQXskaDjKlLulPcqOwsB4jTQty0pfCpvww3SctDkmT2
wsxQukmh5EQTmAyDdAzRGl3jQ0j3TCQ4nmDbs4reBrLnLKh6rwbO4dSxq1G5zAVP
PeuN1nnaYFqZWu+HV29zrubajZdShUT96eT+MNQW2jrgNy4GHBYDRwSNcSM9CYBg
ivtb7XVvW5X6M16bGNb7S0bfLk0xKQT9sSmH11xQXkNgFLQ7Qu5w0FdIL4fhXPSc
i3Ldakgl82HpvIRMH4T9udIAYzcwhmbaC0Z8XvjL7PycNZuCYxYzCwJ0xHtS2EwQ
A/zlB/yBLj7UMYGEhdkIpBOGuUcp/O+6iflch8tDrFx24tQubW31qyJWB/orndX8
2ga2ujO0VKrLUIbo5ZQMrjO0GmqY8pgIaCIXYd8B3ryInaGBzasaFCoaO++sEnZ+
KvMPs6vkwNE6xqPgLuwJLHxzEraAgVndRcETlRlrO6/R2FnRlQKEo5iI1ugCdqaV
1EJAOUPhst/d0vO0XuBxNSvhn9HInQrWNo3I3ebw5JwGo2nF3X0ra6/cnlxXnbi3
rH6nWqBN72XJ6ezvIkOTSOQGt4O4bErgyvzJrZ/7n8cbGjGsSyTQgxcoH9pPagJP
u18uryQqnBUya/QdsCbw0lbV9U8kJu8v+wiebLkUWhwgoftt2wRtkpdv2LkYZx20
7Ix+/8NYFjOPzr2QTQC94FxQ9Ft+SQ4/ODexPtncdbUJY28Eq/wbS5GPn5VLMZG4
leMbAdCLLzczHGmQVFmRHj2D3ku2oR6k2R/2bxy2BZK4AbQXDcvBiwigN7dDg1l/
Xc9ljRd3G7B2CEXDb9/ltf9KeiR0Wrx57rxUYy5+U0x5yxFNLwdqvtf6jhmsdc9c
i1Xpl4yDtnO0AXI3raZCXp54X2iL2oYDh18q+qfZKtc99WTanEA+xVYdEuEwVnEe
bdihlkk3D7Kbx1PxSdz5wFL+c0tijPJ+W+sjZNtwg2YbIqrFc0vun7A+8dqEeJoR
kcCeMlDgz56QJqQKoZLfJ2SWR37qu/F6c6gn0+yHCmL8UXpZPiAHdD5rBscAhJVn
UvtKScQh+M+mw2OVYpTP+1IkApNbzTOlK2BV7NZ3gDZm/VbUnhy4oFzjDil3JwKy
BvbmUbCioA5GnCyAHGHYiOeTW1hEC6HVfwKKHgdimEdatmQSFfQ7omk22QEME3tC
TgQG5kGpVCeM48Ut8m30Ld0kPd7WpPyXdkuiy5YySpGUAYt7bRV27RF59wbltHBF
qGHosAvhGc0x/XHlSNKHYcLruInM8wlmuGDhrPTZFIc237AyI5jfaVVzI3tyRtwi
4t8tT1b5oHzSmkGEdn4xzZiliKAbVmR/l5CVE8T4wYAQNLSELxAjPLIoM5TO6PVa
W/oHdsoxdGEmzGcluVXtJvtoNDlZTx//PrkzRNl6PVk5wNztRrNqrX5x+Y7YrnnE
+7dgCB0/iGZcjqst9gQ77ETkB9YGNuAiXxXQ1Ysd4R3w6Wg8b5YUR579QWD/1Jww
ubo5ngbub8WBQSZYKbJb7Rn9eIyjbZeGJK4JeZWv/8zQmr6Bbnhc+apcte4DKGQ9
54SMnxCkLhktvtfF+PoxGle8Bc54MjiRpT1LzFuIOBWCpZmk4nr/cVI9usnfrQRP
t8cG/UBomX42ea6h8I1ZJo2t+OERuzZFk7iC1zgKqlO9U7nTTpb3JxAfygFmsNZh
9emokv8AfwvC+iflrHfbWqM3hk+hMZR+hLBqTflUb5al6Fjs0NhhjIP1t2f1Yuxi
R72hs4XU+eUmP75FMfYiByOsynKRJPqaFB+91USaRFRUXd54ATlFE6SpPXGb6JVn
6vGfDegUD2BQTMcJtxDOZEQLBrZqkxgezvBn58Mphl0JE6031x/lj7y2Bi0vOYw1
/aY7znA5mzetFk6rHZpe8OqaVgU7WNZMP1km1yD1HFi/AM/zhvd6j92VDyPtp+cY
1ZwRFcEN/4tu9Xlnq04fPBIhFuTYHGnhSHj5bjNQvc/eRc0/Q5i0DN6CY4o873dA
jVqGwFYf0RugOJMcRzSSEFceQ6v8UOVR8AqZdZ0V0MLBm5n0kMSpOC5hEcDaLCcz
Kt1VvuO5vqzvmnynE027Aj8FdS+deAjlD8J6KC1mrmWLF4u3lTptWja7ILzPv0un
tVZL3C8AiffoTxEYh8HfLpeUvcZdUcUeiWyhs19bttv1UgUSXOUPLAXoE2VRk6WD
gQnJ71VgN6pXcRzy3DFpPzodDCrPnf9/uQNPZE4gSt4FHJ7D99I7LZopPbWbruC+
KS3TysIYGPQDJTEkdDny59AWzhGHk5+LfbNtAI7CUx5ShWcOpcQ4gE/tzjoKQLCf
4MBMIrYjui+E7BHYgnrwtxt7ZvxtLSDIDE9JnmjHWFN1WxDbprIJPavbTSnVHiGJ
9Z6fGoLpEE28x4SuTbNuPQGb8GdMT2nD5i6YTkIp90gYEYLVDETNosvnb3aPnhTF
LzAwzDd3NPuzzEo8WyPJpoO0vnHxFF5w/wPnwF9hrZwjp3mUe56S6VG7XxqOGmg0
ReETrtHKecNDOb0D1VCCYzAYqsw2b7SnPru1p6LFsKs2IthjTdOPdT6cjot1wefl
TapKoNwpL2y52jWd1Ur1yYvdZHd1DJ7atcV2l2HZ2OsZho4+2G5lAUTW3YVkI12Z
YfuBM4lDhnsdpC0ducoP6HS5DVmELpjCEp0JsfWMEUIA+d8vUB1puHk6kLlAvFwn
b/Ia5qUu7hVRUHHzHgy7XxeXvfU42Ee8Wgk7U18q5eP5yS3LhVoCSnCuC/TWnrDw
y0tGVY4M2wH4GMlj7VxU96c8cuXK13I9iRvEXjn/dFkjPj17rcWTDAFwOcMAql3E
I17DT5tLKtrGPerjoRmV3JGEZtRpbhlvdq1BaEcMdg8X1QcDa8eg15DN/wCewRKX
LnLEwKzWjb//E61TNXSFLD1N9n585FDz46sWem8X66TF1TrC1BYnQpSPUMSgVDBf
No+7eRh/T9PWYG3nvtj52O6QGjnaY4qgITOyIzXIXZ2kcFaq2AxyuKWvHW/rs18T
G9NH4Aa29qb7QunsDyLrwvlCuhCHo8FbjCyxJ88jxntJ26ixCBGy8UR8DiMo+Fqh
vhrwlLfHLcV/zJOW+78+Cetmw+gty/9UlYvrGk8pYwNVm3vFkf3FqAvtqp8gECi0
0AUOTlXpdeZI2pn5bTiiyUlHWlozaa63Ynb9W5+fzUV41NNWvld2352u+vUprjXI
d2w3mRG7mqvDBeW3eGRI/kOOiSS8hC/rOng/NonDJ6A553/bDIGjm6l62EQveJOp
nlaXLvEIl63kJUh/IalhbU9pDFIWNNTbh1YUE2/FL0qX663N1vTzw9D0LuI+TQ7T
Fj29niq58ZCCNYLx5Osd3HCkW2W9l9LV6bQvmbpooDFtq1XXCchFD1YyZZu+Wd12
KMlfm3aVD2e2ks6eojly/PvBbdoXQlpmORuoWSFwki8WAspMOf14omfrnf7l7+yH
nnUEi9wJFPjG3rBlmnTlYG7c3xPvroP903v8n8LjFb38NmRaE01FH3lJxeLSZ8EP
F2WFknfl5U2rFr0ZfQn1+LqW0y9rlCos+yT9JIz64A0uWGvwOzSoNpVFuYJ5qryE
1GBlfIV16lcF/VavdkrHDQHA0Ia9iRIWE1i0tQgAOuJRr+Ud+lDT8BoC3lz1Ddkf
D7pMMSnm5h2Zg/ZOOwsODN3S3DyPDONehByQ+xKK/oF8iKgk5hzIdWtZP1LbU9BL
BBEJgmjUSu+aLzDXkJ1CLxlA1gGJ5Ph2VxB35L1SjMGVDgrXKic4///TGjhwnogX
E6G6qA9CtrQ7ikVHwIyNwNU+73nNKxtf7BxUzdEhlCmltNRThEmEcaZXdcYZF0Or
5S1nf9nzsFsyesPlnqKq5YXMEi5vtpx9iLDoBG2XzyrnE3bpDDjHREkWmxbQD/k/
P5EFQIAWUZyKc2Ul0bgMeYOd0tTzWKlCt2RGtDymgYeJUApxRhYebZkl6rqITd5w
piQu+jAh4jcC4JEowSKB4kDXXp6RD3I9xmkYHnuLHaFFs1TIIfnYV8zvDkr6Q1lU
e8n01Bzus/BwnuTdk3TWpBRJtsOm3uFyJPi5H7tWD43LXIzEupv8nTKECBIZCVOx
EMtpWzMcpuWTe1XDHj5ZjWvHpIHxwOpHSEjZobcETgiOJcwabZOlSk5iCpCHr2CE
0F4n8pxmJ4Kb3khtsehulBjGcxeeSUz868BGIqCUZ2QnOxBuoMd1RZua+ekHbPaU
hFXwqgIb7MaFRJdMmlXXR2lIYtgXtlI8tfZz/AqYo+k8IJUw6kMiFlVziGx5SRcN
ahJ+EfjQt12v0oubGIZMVRFZvuCuhGJZLANUuLrh7XAesO8pG3kO3U922zgW9K+w
4WD2tZfG+xc7WpXnknZFgTbM4BiQNibohSFPss/JUg0/k/z13uGYaQfx9KViYOGK
9NNSrvEOWsN0LphXK89VsfGT12Zuo1iqOo9gya7EewbiotPBwsNwrcyuxcxRHJVE
HSZNi/Z3smPQUtZ9ZjUmady3Ice6ZakhOx81t+pzb/cB9SS3ss+h6UqOwALYUdr9
GAybA6RXD5Iuk/7uizZ0OId9xxX8JM6t1u5KAqpTvtJD89XsJQ+wZ7FpqwbIh8zn
bSY3RkyyPLutKHZWxbvIaN2ZtqUSLJ7GtwZlhnEg7QOodAc8LMm1PYozvPxy4VEs
kow4H8laOfzoDXRJrNVmJADflUdhU8MzLU9IKZB0C02c5m7QvdIB+DUvo0v9X4Kh
h/1IKzngNT754kb2/vjt3t7xyK8lQ0Rhsn47912PlBSpMDd6o2uK5qKLGwQ82gdd
iagONeeIxdItuAoOvgLraMuigomHgVKQXR7m2vyBSZFJ/d8g8e2Iti9WnvK/oZau
NLS7lB0WwUNBdrlsrfq+05rFXF5r23DhWlGTPMM7RH6zab827MtyEgk04njLgbG9
OXJN9X52Awk8bhBNNM49cebozJc0gqJLp5FaFhpXDqIm8j1JbyiBU0ktO2qGvZv6
1QFJhrLcbmZdreTDRHq6QWl9OKQkThYFMiTNsaQxryLROvzDBUiV8LeN21Vy2s7C
pv4FBy8ePiGVzffmC5+nPGhJ/6DMYQzdGmRNw4XV/dwJ0yYQo4rSpo7bI8eV6YBg
jMTKEy1PAJmxySy4qXK7VGe0OBLMzA4UN9S/rW6hLsHAatUYQ86+ewosofNZn/Dr
0d9QEs3XYOh3UPeJbTObETGzO5dnw2IkApE5wkYtK4O9q0kIpMPXh71l4sJyGzmg
eeejk11zCCIP6AerBwEVoLcqPAS2C2+VhJ935k3gEJhGt5vuxBQbieiABhkRYViD
xsOPFbdc0DK+hNKlV+SoM6aBxR1GMUdv7hv3ZW4znsu+vSmqfgeqZIuiaYevaJgB
ul6Sf2soC/ttNr3ZO4ufmTwbUiDL6DYC/1FqiGUPmo5WJ1CSXksLAMI6yGgFBMul
GDqgH3f285cF+PYoo6zblRztScP+b7dZ/oWerbccr9i7syiwvwJBZ5N+q16ODkIX
YAdrWCMQI6XEWUpY0JMcT2fSwSVk9UUk16Tv5gE7vmEzoW+Pr+j8uXvizTUArBDJ
vMfrGZXbzGBxCtfI74gvOCTaUPrmaYstN6iVxbrHTdWwE5ocfAwavE5yumHbhZAN
Z6BYWo/MFpQYeyN7z5EGcVFGBp7+rjnUS23PaAJMS2Va2CzNuiGS0yLkmyxtJX5C
VIBmzXql6GKvutaRdecUGCkHKACMFXEr4pScCy/pT5RhMEPL845uSa6mO8GVpEv5
7lldJFtXFGgCd6R3zPWJc4KGywfNm0T6w4T0M+9cJaMA0dBRNxbYaShKzrq2ztyo
NicQsw+s7Vzussq3tpoy2BeG3r8VRnTbewXS3mau5dkzvH+dVesc/TqzCl7ixilB
gmjASCceG9TzxaInb3bvGKGsZpZg6qVr/mpRdWpYtRgrvj5QN4nGvyxjnwh4BgJ7
EZFwc9leuDRHPyJhMO9emQylCiAm7/fPphFy21DA5SF5lmUpuTXLv3ZrxYoUhVyh
OlXdC1pdhlr9fde69Ju+YBt5+8vmv7fL6JA8U6jz3jkwU4rMZ4Za0NKFHj0QUEtp
9t3UrxoswNnvCok90RyoNsqC0O7vKEwfmARF9AkmgfcSa2QhQQvXLENu/3i7c2Hn
GOoeRCyddzmRRuJnOK/LuZheFBayiwPDKOvqtPuGBj5XIkzQiOLnxiCyjzuJWKVp
8UO3nBIrvUIQkOA5ekRkP8KIC5BXmu58VI0HNY0VaLll7Tgk5OURENkfaaMyRAM0
AQSh6z8J18n09BoWCjTatATgS1CR5mZqHvfX3/hxVPIjD1L4Tq0Cv2LpQ+1ii7rw
0DWaarLjz8g1TRC6ky7hMF2mwjFqzRGfMpzRV3vcZwOaEOWBu9bRVxikc29tcRLz
f4VqWM4Ivzx8yhJ6RYBgWH1yM/+L2F1xKGXBTXKtieeHbxNsOEwlvvIHQPsaMzxA
Pe6P1fYXQWuvywE8tedFz+SyemnxxI86PuvqrAJWSkRQifWEwDQdQmZhuXPPsCDd
Ah7yHi8f8mfrgIdgOgo3QjnKWhv59s3PGV05kqmHO36Km1d9pWPhFjJirdkmlv+z
oKlTmP+pbDoC5FRU3xT4+1lGzXEWyB8G04T2V0/zUChUt8yn/JhYjdwbiTQYXvq6
2kogK/wwE2XrsUGTTLZAXQmVsBL+Iejk3UiXFZZhsZelQ6Ui8VnXwslcG5z4mIsn
/g3k+Ej8NgBSf+NDrHCuj0RbxGdB+7jNtP0CHAeZ0+Iy5zKDeHkgnJApq3LfB2je
eYRm2AmgVJUQpRSsBAKCbeTPdKrsGWxHw3mhapZ58W7ed/FE2nWgfdne+miE5Hzm
J7/PqbefGntoGCkMHCD3OrBxJIQdiCUS8qE5WOP9gu5loX3wq0PsF7oFLF9ulx2k
scof95vswbvmuRJPIqb8xLb9qLFW9M4KFYnID4bY4rouzbN+orM806lVm+Sq+5OB
nkNT9pbD4O/mXd+3QwmQALybVA1xScXfiFTjFQPOMlW6/M+IDjw57dkNeQhX4knD
9IXZh9Vpn6ZS+Bd7G2LDQ1j5E6v2Rr+JbGR+5yAdAYMaCBbFjTsSJWF6r390KL9R
cK767DEe910SHNo/Q03J3FrO0XDh634LwpSQw7KXJpG9m7Qut4z4YHuZDzy3a0U/
NFvZkdkBBHhdxOzyxZh/8KW4OaEZw3ABwKpeTdJAz4YK/v2sz2RRKUov6ffkNWHX
LtTXiJkSp5LxLMcXm3jW7YDu6s/1Q8fsazQjiGUvfTXG/vR+ZH5dv4VxoAWn7puG
Es5aBbiGXxgbTcncEdvRIZk/AKD7zIKfWlLziP73tZlRT3pJVa7SAF4BvqJIVbk5
qbDjtlzMstspehVllDa8tfwxBolUQJWRnRWKnQrNIcfgGh3fKuVkQ4K1J4JK4Lz/
gZ8QN3pLPtAplqCJexAbUJPVqiM0Gu/fvrLZsAGX6o6x7UhTgOj9GiUuSVX+oNl6
3azuOw39LlwbT92LwDzVSkyOW6YpX8qpmtE0mdN2n1ytHvPvcs/San5IKzFFEk+5
I9NE8D6P3Qc6pQgmkmlfyXIXTaLyrl08WSA5SW69I0Zu8OiG/4zHhiE/ndnmieQX
2WoI2JVNvTjngoPlq4ty2lAhCGarDwT+phBS4hncsl3+UWFY0PrKx3bFCnKfDe+w
EDFJomHBNazkwPfuAUnYJsA2oLSlIwpg1/YyUxtucU/hIW2dRgNiEl+BJi4YFucD
Mo8c20WVON7ObWL5aJpvrtIArndVgart1GOhiKKGN1q2EiGzg79j+r45vodM/hTm
VPDlH0+1lKijbbviXW2v83T7WRdeH4WxtEktzeKLePlzUvSWbPUZmBjcvckf142I
vXKREWgzCAI0srih4bgCXog1akj/uaLcxRx5Kq0NtuDwEKtfBcZv3XxyvZBb3h0l
ooU/XcW7PLGgh2RW80ydomm4v3iYp6SSBScgIo/7UrDXo9Cbzn445+rWoG+FPA9+
LCOp+rC5jZai9RSeiq7MciM2qMuCNk/RqC1kAV6Rnn4IqJVNT0HCvaR0Znq2H/6x
a/yHlHVJjLAuMEvLIzk9as+WmES9ia653wEDtxYIZgatAMnTH7C2QAPjB30J976q
5YuA4CvKetPBstTl9i5zpFdrePceeUOs9+TaXDSTvfz9Bc8153uihWbOGhW8DQdP
LRK3oHkF3ivzrT4JTKUWSmTC7Gl2yalaXxYHOpFTPim1/7/nUv76yctYpfv56gpu
tfH1on8/DQOhteayE1tPk+6+7vuZRWQylKOFlKiUjQstWF7asZfDpwYaTrqENA/h
U/LsFoLvuR0xMklqZKE/gdVUH3X+E2cpBtcvaoIeo8+i3nvDGASJ8T46nXN4+tDS
f2bDysmKMR2FzpCUwyVmud5w+2u1Wutdblcd++qICtZTIgZK2LWFCtfTHKpIilXo
I6tiBtxS5DXRsQn+u1Rop/61Zltqc26oSeIU4F3wLXxU0t0qDABRhK4xCnclCKO+
AsyZ1R6M3OpK7uOIyPeO9s+cd5m+5kgZveu1YvqRMnwGO5yoA/pwE/jGQnFozdxq
OSG+toYQtf7aINtKvJnpRNSehJHbXVn2rqFgVrOWIseR8RFQy+PZmmgIJzCHS7XW
0SVVqQ7Pv9rFQZ4sLwjpPrAZmWBv05NXvC7n9vIOTFigVP60bJANQYWVKVR1kwxz
/nUL/mjtTwGtvhgBGprDE0yrmU7ehHkAqxhfHzdjXPuriqq7b+enDNumV2v4MsXc
O/YMiBSy1aIllN9ys1lJ8uP7FZ2yWrb5VQTBPrXi4HM2d5tQgnFvJti1W7pKpKfY
laec1jmT20LErp1ffuH00xm7+6MImyI5+xF4xobGaT4ah6xJ4aUw7pqC5Xfp6+/D
SjJszi1tQU+FZHY7HTFCQHK6UQw4l0uSlTlFBP31SMjWSgcEW12Fp6lfDxSTPaNB
Pd3QkXToI62FdxVqa/0nyk2Y++b5Y1ttqM/Cl/JzmF73xeccaV3GC84nDeN6x3rR
UpTRS7vyhpsPRe+rZobIMjAJnOsEF2fssypPkRLa7EdBS1Nvu/ELVScSyh5OzydZ
jIn88QVw3TjmsiL5+EhsXzlqHzpVtxLnl8QDtcrtf43T64aXGsegYlV6UjhKNscF
IvlSwpUu7FnqyqmAZtiQgS88S/ZlDr1Oq5o3L4oadtrxnw/NuzD6UKUstfZRMGbQ
ROIXrsJBZJiJEnNANzm5jHqSo9cw05lemwz3rpYCoGm5nDRrpDWxplQUEHIf6EZ6
ExYt1G45tRC3jiC/mo3qanCZ4Eau8MjYoeA6RH/QabGsj5Mn/Dz/8chjp797a+6U
e7XOFdG1FdIIsGg+xTt805j0CnB2mO05lln5/p2jy0kTMbpwTlFN82qbUbdIPOXN
AtmigTPuG9MPjGSuzHoYMCsDofmOg2r9A9jMzqUzFW2xDy24shamnRi6i6/b9n0/
9eJbhP8ueEWR2MshLI1Bny8YihtiuIhh+xFqrgvYd/Ub3duYZMQUHqjZcpbyOqO3
7N3GAAUYBNMCC5cMhKQrrUP9Z1mVvLqdqStRyvmeD0He1Rz2LyiAoiDtAG1edSaW
hTUe234KbNaKbq2FzNRARpUeErvojuIQLIBkhUAdKNCiGmi2cfycxaNo/25mVY9/
fVphh2ACr6ibfEIJrPFOk+Nt/taDeKFqIlUus9A3rs+JOVgYO1bjZT+nPG4AjcMy
EYsgJoJal+UTD+R1DSKoBwzWLbciRhbfx1TOQ7FYEB8sxmP6YoHTGp9Fj3oiufgg
rZpWIl8Mv5lpmLw9ICkHQacfOsc9TtXOMKTC567TWeMxNBnwPI9L9xliz6kSGQHV
jZiUsiJZY5j6BqorLNSuS8vlDpErm1yeVdEs4vI3ZomIJ6fZvjBonxeDPp12YFnp
fhzWjFcq6OhaUw0/r6IEbu9E9ZVVGwpuhWbIMWAvqNLuuuvlcnWsC53LrPU/6z69
FJTk/a8h8emzWscXNoCWcBSMHYdgspaVM5dOO0nuq6YRPZNfvNAqaDeE4QCd7JsV
ItR3xasqr8tJOi2Bcsz4elWDF5ZUx1tcXUcVZN962Z6h9lM29BaFl2WVNl1SaSoU
Fo/WeVC+7rnkknL3OWidR3ZqDjAIIY9tViOtJHWk7TID6P549EdCQD0WjqtwD39S
R3QFI0RbMHDYjgaGeiBfYuwdTZkvg7fDR4PBHlaNPlzeW2McjwbT7kud0CsMbUqv
FbWlpDznGKBSOr5ZKz/nTBuzAjXCCLetG6XXrQwFkrUwUENBiFn28WqFCtqNgj2Y
NE8wqcHIbKYxZie8PWoVm4YcEh/hWFcZJQ66sBtJs/VqOA3UlVjjMY7ZUiJCnx+7
JSghjcM4d6kUHrIUE1NRv4EDJhYumYsLYfAnAlOXbklIEPRJ91wNasLV9BpLlQhp
eK7G10MviWhWP+jCR7DQlk2XRajRLjxw0Rh8XS3/GrvlkMBZ6lNo8iuYRQ1C88kv
/Cff1l+jetS9WMj5VI2O5+5WTYcbPoTlCvZTRwuv/3iUoWkk1RoawSgWdV3XqhEe
X8esh/mmIMZIpeWsU+9dor1j33aUUyPG3Jr2c60NxECItJLFBEubkW6uKs5ck7tj
EhVfnpTyX5NFCtcJLAd2wNa/1v6qj+O2Nx4uh809c1vtZT+pbDWpOWbN7sa4u4Mh
ykQIRMfuBvbx4w1behsd1kbmGBs0XWZ8wH9gT8oANFlCfIzg+xbBE1RM/TzNeRPr
Xgdk6+evTInJQJlTfp3/iUufsrFuDmvmsn0tmOAfg+AnoLtCdKgoDwGjDouleh6I
UPIAtWDWLmbIuQSohU7VIvSulIffdk2GI3cKnFYetactHL4F/N14Dtj4jssuNx4v
AV6g7C/xNSjjr1vjLw3l+X8daWQJjhlcu5R+Z5HOBQw/9LsIxRJatomBllVvxZz5
f5uUrIuFz47yn/95VfzrTtXqEzJc4yMbKdaIQccKG4X5YCM2ZmzsVh05MSx9ciRA
/td4dFInG89E5FbyUdbV1N0RiocrY8w0Zdzgys4xjPc4SZsuawS6A4J/lqthAVwX
/MCx0Xym6vw9bCxuXwrLRL5PMRmzcR4nc1ZIR0hQjqJUB3hFR/69Kso8tqNnNs0E
a0uV7D4QjO8/eSKU0MZ6iEKTG7jEhMWLuE/MZ+BlA+bCYE2hjnvwMaS2yHFTGbu+
3h3R7rk3mCREkE1gUT6u07QgagmR2mF4QO3FGiFFE543hrE1THmeA1CHpwLhDMZm
Y/fT8BsNH8t044JOARxBEMbAAbuBRJe8r7giWCy7X+7hE395gokV4vrQw/jQlqqJ
JCzJOIfhvOHL2zqr9YQuuGfx4HrxFbEyADCIKOQ77BLneoF+QG9qSXGGhiq4kzNL
prSwNcM58BsOatkys6U/IT26iXm/qSx2rNSGYKrC+Npr0Exaf1WUFddBI1lEnApm
e9oRSAkNwwb8b9659l3Aubc2Nl2B7culIhXvDCSXNQIkVJMxpqFeM1tUNaSIGy8y
lE2m767CgWN229ZGS4lKcMzm/h6ohYHKU+tqOm9TNgNTLf28WcllYw0Qxd5W5jdD
hJu/BH0/q3YbTultAg+z/qjzNEBgORJPQis7TPXaRmLMsn7BQtx5kZjSzg9qG47V
pooURMWvXAbyPwGKWrGEC5CWyR9PQ/r2bbBoj+MplbXiPC5uBnYzFBpwV52GWbG6
y3iEnyMZIQzC/cEUrC4RtvZnzyvBu84ZWa/7CZ9sgRaW2l/5FbYCUbfalBw4K+y0
T4wVQERydcyE94D9NL3j3gtgn8R7mJ7UBzMGE7cbELNGz7DuclfM0wX7S7kB/jGF
mXZf7+CD7+3j0n34zNpCVkRqcWGq72C7iqcn0kEcqqWRVjIPQ4EO5jAWK+VzVOq3
jG8Il9kQ8Af6cmcD262LiHgqwRKo7IVbOhia5E30y3Nx8kRffeUiSOnnqj4h8R6T
Fn3/o0EtEvWz9iCltaOKsJMHoDy9nWW5kHQJMGlmjF0PKHnT3FeOR1ZVEAUfYDcF
dlo0ZyXewTXkNgU9MORAhw==

`pragma protect end_protected
