��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���d�v����0�i�=\��A��?��� (��1_B�f�	�Ѻ+|n��y��Q4�]�aY�����*2�y%����>��������K������ �
�D��z�z��C�y�B����
_�U��hkF<�~x�ܕ�c�5�W���+u�k`�P�%b�L�nk��ӟ;v�a3bO��e�4Ҝ�FĒ�:�?\\t�Vޒ����Ƙ��|+�v�ϕ��َ� �]��IAx	6}��vF�k��ϋAi��9-`��P��3�����5:v�r3�.xR��L��kF��Ȳ�30���J�i�f�|�V6h��= ������s���?�����1��h�eo\�=�	Q�,s��F�?�� *����Ek��v����u�3�:[ۤ\�&���'�|���is��S�+.T44��d��瀫�`�<���ni�E�	ĻV|�2�㑒Q��B�?�(�����J�܆��;�e0���N�Eyk{�%�b���-�/C�<^���7���#8E��Q�������z��f~���R�����Մb
�r���?Uo2�J�� �lga5MCyF��#C�����HVX��=d:���Ô�@3��݀��oF�MĨܜ�Q#�\��j&,$�%�Q�Վ�*"�WT�P���<�'��_`��;�hPr%�pA�
ƴ�l �VL���wa�|�0�lܾ|����3�5�
+���!_�;�3�~��P@ܮ�)J����$K�Y���rҰ$�ڦy�-s�}qN�*yT.#Jl\�]��m��0*��Տ��<�-�:C0��5�;�ޕ���*yi��e�_�YlH�\P��甼1��է�����1s�d<��g7�sMSeP��w&���*�%��_������vv��Ri4�֣�~<�=���oi�1�!o%QȜ�?4B��SFQ�[�d��p�Vz�D�|���T	6<����,%�'כ�
Ư�}���)2!���s �Y	L��&R�����..t�H�B���~[�x/��:�a�~)�®�mB�ļRn>S6m��d��~�\#J�z�wx���1�W��w�aCE�g�0r�I�#B7�1�ݥ��?����܌=o9��eNw�ʕ����p�'��IY#��P���;�)���n���g	�R��:,�^o����-/c�e��R_�j(�`��R� uLdpa��(�$�$�FX�풎�ªhF�c�f�>���/���`��,���+����	�z�{���'>t� �W�z������mb��{�@�즅Dy�&�[����w����Ro�F|tߓ\>,���ꍌ�?Y�;?�|2]�+��a��I"?ق�u��֌���}9��Se�9���F���!@��O�J!���V�G)�p����0M|��Z�!�>���q�d�om�U7�=����������{Ǿ�$���b'x%�zBY@�x!٪�1H�.�Ǖ��s��iT�K��$��r���~3�~�x�W�F��_f��{�SK�r(�� R7��;SC멯��\9��c��e/h�,��Z	L@�]O���R�@d�f�O��Lm
�k�N�:� 3��]��(I��dNHrN@Q��@�ǡ��T5���Zi�@3�A@)ѹ�4�δn�Db&�TH���F��0e`�0�n�k��f��q!��;��iQ��;���V�0U�/@�R%&`���{���%��
���@�$�r���+O��`K�z�;�!�[Y\~|[�Æ�0Re�ɱGo2�H<c��O�e�`�G��,�_IF����}�}��atx�\�O���K��*1�Р5A�(T]ͳ}`���χ���"{PV�U\��`Ze�⋑푡�h@��.f��Á��^�#S���ɞloLNN�T�t�Is��G>\p(���f*	�9�s�;�B���WZ��65C��c��E�êLtB��\��A�����Ěe�E�hE���3�I�����yG��ز���)å����^�.�ފ✴â����n>?}�%5����Dz�< l��.��m4�)ς�w� ��,�u1��\M,�V����`Bht�߃n�M�b�g�	��{���Ozn��6�3¦'�?��m;�Oq�`G2�NQ�wE�F�r`��I�*.#t50
�/`�I��tA�8�!c�)5��� vI� ��)��p��k��ddS+���	W
<��u�Kzȅ導�$My�af�z���� gm'fWr������ �9����7w��&6��D8�� g���(��*��f�³��;ɢ�|�W	 ����"�$Օ]�jX��'n���h ����W��q�+P�`n��F�\}��LD4i��LMAgj|��r�1AD���$*�A�3�!�!�����J#��u���㐗p�Yh��݀�Fse��t�]l3��UV ���䓻'�a;O݌��n���,H Tr�r�!Y>�!�9%��
��]�:�7ar�$�tSqX���O��`���!��,�~����)�^8�K��0�L���!��d��K2F���٪;�M��ш��;�Qg�q��i�z��V�"x���q]�̷��7F#����iwk��1��8ۗ^��z	�K���]^�{����"�]w�p������f��F��ˀ���%%TI���2�5@�B)�#+��E�큊Y�z�hj�E�{#� ,����h�1��E ��$�_�oP �b*�~�hL�_|D�#��G�Wv2���t/o�y6�%Ѣ�"�?l�p1�32T`�E�-z8g��sǀ��fƙ�0�t���A� S9�m�� ���p(:oS{�E��ib����`��<ĆA�l�ufiƤFD$KE���@Z�����;>4��m�{��@F)�vx�f&|ؓ����$�Mq�	��{qkͅe���'��M�(]K����ܥaQ�艦K�%Pj�Kc6 ���-��`�%.��ip��pf�c���o�n�wҋ��kVRF��	;*c�) ��í��O.�q5�_��"r��&��8$�8�ѽ���������j�:��A�=��А=�Z��P�z��+k�Ҍ���D��	{7�V��@��饥�/zIh�k������b�%� �8,(�Yf�W�(�:��`bkY�Q�k�mk����+҈�w`��&y�'ς;A�����Ň.��W$�:4����#��4tE$���r�: *,�\�26�AZ��\r�Cx��E���n���wVբ���n�ս��� ���f��Q�S]Vp��f����MQ��=ј̸K��φͧlZ�2g7y<7�v7l��Ɓ�3?�����N���<��w���<�8�RY����c=�M����������Z�6��Ǣ����L���V,�L�v�����I(�O*8���nW9ݠ.@��b����\)�#��Y�T�٬	Q#��3�{$��$?���Z؃L����q�:�,���	�x�l���OƏ�e�'��Y�-F�h
�]�%KKC]������T�3~��X��Wl���g�XF�� ��r��}t�o|�+HRa��/�P��W��^�o�e�P���{y����ł���Al�m���3Pŏ�|q�RQ���Dx�=v���0
�+ƿ���\ɴR����oB�I��n:L�jz�'�>�����D�Y�m	F���4'�Bk](n��cH�?~��	 -E0���&�C-��� �'�J�>̛��n���I�r��{�����͵*��[.�s�)AC�����L���p�0W�UTJ���u����%��gq	O�7�}�7��\�8��ۗ����e�FN�-�8"��(��؎t`���3��;�,���X��gct-���J�O��x�ޔ����y�k@^��&
�:e5,n�>��H�ƽ�T�r��b���P�J�L��j7G��cC�Z$Y\n�O�3��*�+	����Z��5�o��e6��铻�{�}�Q�/Y�f���i�%���i�M�jvғ�/�eP_�ƃC�( @N��y��ӆ+��w]A%7$\'��%m�BJ,�$�D�ð�tW��������j��์����ր�FC����%��s,��Ԙ��WzJᾖP�2��<'wS�G�Ȳ�گ��������і��`��8m�x� ��*���Rܓ:�vh\�F�t%�/�#|�)��
�W�Z�k�L����@5�P'!0�;�	��N���F ��L�q�[�-8��O�O�X)W�a/)��f�|�!햧��&B��%y�c��A�X��פ�ůt<y��s�5c7N[�_e���:,E���d����}�8�� �,��ʋ�]�:���5���8kۡ��C��\I�������J�i��\�������i����Q]�Def��d�2}���!��?���L ���PU�Ł4	S���[P,���mv��ư�Ki�HvĂ��2҆Q%��*xM{ˀ.��C*���3�!��H��uZ�@9�W�:{�}1���JN�+���E!���l9�^�	bp�R�,D�s��g�%�0����!�G������(�S�]�V�� ����:*�J҄�f}�sS��$�B�
�������4���0k^d@�=K����갊���JE/.��C���{W��$��\��{�o,�#�Ե�$���Ӑ��o��5��UFʺF� ��U,��ܤ�T��}^��+3n|M�/ k���խ���y�����V�=J]�F�Dud�r����{Pt��R�<o��u�?Te\�U�oӲ@'[���[O(�@.��a7�*�s���Ғ��)�b�B:�[Td�ڕmĮ�����#�3-�e��2�ҕ`���s�a ?��``�Ę�5 ә���T��O����r�9���rU��t�+������y���$��u88�} cp�g��t�]�2��*�E�b�?�m%�Y��مX5�9(m~�"�pߣsU��m���Z!����D(·�(�Z�7�xg~�X���>G�p��}�S��-�ٝb��%��*^����0��� ����M�T��Z��icA�A��S2��)Frk�`��W�;43Ē��F���Ms3�`NZ�_z[J�< �Z��ũ�B����(<�|i@f\�VT#@Y�مaG��F�a W6��g�V¶X�q�Ts����k�5y�
C�_�3Qј��&l��GN-k����St��,�p�j֚����o�X�l�o����1����'O�/�!Mv�2��8�����J���v/\�NDVB3�Q�2�A))�m
 n�aW�.[V�=
:3�����D5 ~�|%+�yI��7Y}�/ ��Vt'��Շ��g$r"ğ&R�[�4 u+�+-�S�7D�1X��u�5ɗOS�3�@��	8�`OW��r��ӓ���O�A[��e�����z���p�2��uSʥ�4C�&S70^ΑTk?+�8�&��u'��a�oGn���3i��e�u$�:o`��4oB2s���V���)����?�f�F�@7�d����KT�0d���#r���y��Q���Ƕ��a7��l�X����Y�=��?���I	�DPM�i���~�u��s#!!�c
�}-�H1����Q���2�<��S�$�m��C� o�����*�D:�X7w�K��?_V�5P�k.�	�[��M�$+w�L�C~�_�C.)y_¡^kŅ���Ćy�ܩl�h��/����y'?EmnH[aq2�r���Wړ�d�}W+-���A�
T5f��lìvHekap�����M"���D�����h`>
�O(�-�4�_d� ȅ嘹���Z2
9M^|V~
��o �c��>n�	�����c�#r�Mhg��T3���&�M�Kx���ƣMd�Ͱ.�I�}�P4�l{�$���Y�mண���T�P변�0��ο�I;�'�����Ŝjܛ��t�?��:Dz�ob3=:��y�����mJ�\Ď�K�,�O�g�佛�b����&����4�s^T�W r��tʾҝ��i�M���.*��T(y����Oܴ��%Q�_e��3k� �'��؈�����M|W&��!���s��b��F��a3����S�E{$�)��Xm��G�Z˯�`�kۮ=���ӓ�47��m{&��R�����"GI��S�j��ȇ{�]F��m�AP�e���Q��u��c��"�P?+����g�Ӭ��O{��8�4���2��Ţ��4�Cv�iU2+�#oN�����OxHg��>KT�h����:R�s�t�2�j?;�Ly��`��U�)�c"���O&�аg���\!΅L��Z#��*̸��t��&_3��,�5u%�M6� �ˇ�1T��	�<���O�a�X@8ہk(ד�U�W2{��m0�""��Yv�J�4�)�����p��*3蒪� ���4���] �n��-ו8�\z-Z��U���m�fwN��
�Z�v�*`��s�ᕀ�t���y��A�_3�E8��|2;ؓ��<r���c�+��G����I�t�4�@�S�c3�'h�2�Z9��}����`�	�!ϋiN�k*�mw�|�EWU�)��s���,��C�
6}�D0��0P!x����R��a2��l%���Mx�e��6ZrZ�&l��7b���d��r��8r���|���*��o&�2sd��.cc.�L҉�p鰐
v��b��,��"��E�h��������ŗ�f�[��ЕEY��M�7�G�^ìĒ��$J�ao�����1.�@5v�����:	m)�y )'�E<�R!�&*R%�ªE�^�#rX�|VOW�&BW�w��L#)��M}�`�=�����A>�.z4�Y
K
e)���_ꥎ��=�هY$~:@��'OunjQW�>K�z�>�&�Ff�@�l-v��?�E0��8�B�ׄ��ۺ����~t(^}����А,𥟝Њ_�&�����q4��W��a�������|$��	`�l�fv����uA6Uu�[������l�l��_��E�*��|�t&�O�] �)DL�*���)�룵R���"��*Bq#2u8�A����X���v-g|t�����Q`�������+���r��=�X�k�׺�)�bP�Ufx*�垅9���9�\X���w�o!_N�b�D�iu�Y�i"��L��,�A)?G����&HsW�a"VJ8sx���rH춙N^Qo�����ͨ�X��xt���a��Mɉ��4x9y%�ftX�==���n��VF��]�7���`KpGUb�-��ߌ��oN�ٺԇʘ�i�B)j��y��5�Y�����9�߲�;ey�#l�����;t��E�0 ���1��Q�0��1�`�+3ơӸ��~�f�b8��L���^�m,�!�II�v���+��X@�%��>������Ʋk�3�`$�F*rX�~���[ZioN/�8B��S:�q�g��S���m�Xĥ��	.+�U)#;������/�u�;O���H�V�`e�m�����y�@Y>o��uL��0\��G�GŁ%��n�Х��ꑝBrW-���W�I���?�P=	�U��4�&@�wŁ�aj����9�@p:=�e��L��uE?<�0�6-�&�<�����M���o�.�2�x�|��_��o&���o� Ɓ`��O��C|Uvs�Fqv������W�^&_ Un*��m�J���/B»��(��8��7$�#q��������E�H���d���t��|�D���y�:d���u�8&.�1��l�� k~��L�ُpX^7i���u&�p�v�Z:a:a���L�!��:0��!e}E�)c�0^����y�
�zE���T�惧����&EF��ug�C1�멥��V,vXV��6"��3󥨑��em�{�ǹ�93;'�2��>a�u'����ާ���&�vji:j�«2�ei&I���vɵ��!��k�� ����̚,���ƭ_�㩅�,���([M��]���9BEX��3>�wQ���	%X>��౟9-����ժ���� �1z���
��8^�Pv�-����X�%������Ў4�K ���B;C+y���ZK�(o$��Ip	�~y�Y�������WЁ��g�5�ȟ�Sޱ�n�8˯h+7R�޻__�I1Cl�aS���s ށ��ïٯM���0L2�TH�H׽GQ ���w��o��&�Z>p���]��K��B��'�W�U�.�d�����s�i�jX ������:�n�y:�q]|N���Pu;�.=��&�\K�^t��o�p̛ӝ=2�Q��(�tD�P�Y
�FUP�w T9�����|��d��VIቋa��������	@����3�u�����:Q�Oо�����UW�܆	1�<o�@;���J쾐�հ�c�$��y��+�����C���`�J9J���FؤC��v�F�D/��L`v�x��L@�ҷ�]u2�H����E�ą�J�:�Q;fQ�L+dh�+}�l!�C�5�')\o���+�e�_N��a��ٽ�����S�ط2z�)�?1=��8����P�q�s�H�(e��=�3h>��b���!`���53jYoܚ���!�-��f�{ '�M��G���p�����*��-
{�`?����J��݈@~9M�$y�ox)79������v`Vn�!O�1M�Z��S����/x8c�;S�g5U����a?�n0{�kb���w=�l~�qs�Z� �zyR��	����fZ;����'F���~��ZC'�G�b��i����'����h�\� �\�U�6F�f��:�3h!d}2�3w�6s��9zg�1m�CF��W�D.M��cD;����>ZH<[&�yæP�X0b���3g$�B�� �WzH.�OP�S�9�%�SQ!f���L��+\]%g��>�5S����Ά�Y�KoKY���o�dY�b�Ge�aO��F%cI��>t������v��^Ii-V�����#�Y��2��v�t_�b圼�n.2�*�t�_��RI�W>�G��w�k�I����T���$������B�k񆟶���m���M�7#{�}���!����t�3-u	xQw[X�T�&]ie��~*q��]>voc�����Q5̢�i6��x�	�z�d�Wl��!���%�LL��|��v�Gl�y�f��3ǒ�gZ�8�,ᛑ$B�Y�O�?�o�Ŋ��l�Y�S�F\3o�>�/+z�C�gv�>��/�XGae��/$i8����F�=��_e�5q�ޔ'�{�B�`)FNC�jY���ɯ�(�ᶸ���o>�>.�m���Q��R�v���������K��eU_"̞�4
2�9��UAt�&��\��/U>>0����9u�i����ƖNOܧ���a	n'��P�g
j��H��\?@O�*�H�����)��������;��:?���"�9����W.Я�႕-��E��_�d��;7,� T���Tbъ[Vw�?8� ˹��<-���
+��}[�Ҷ��q$h�=�{��k*��F��~����-o1��Z�p����02e�r�b�~5���Q�� �'���"Dl���'�jkOQ��	j;r��`�)-�d0�@�
C�̚@q.�bɾ��	��x������K.�MWE`qa$����\|�e�+' L/�c���<�l�'ϓ�Ҁ;�N:tw���(6N��=`	�l�.	H���
/ފ
�7	ꒄZ�^��J亏_僰����cosJZś2@�'˧��a��,��PDJ���/bj�i�K�#��]j����v�2h"�#͆�iG5�����2$kr��F�o��2��׿���U���*j�-pK>y�q�殢��;�͹l��<�Y:��MCM�I9��q��eC�8�?C��sJ� ��?G��<���w�߈����� F(@d�6��F^7P��,[��/Y�$�,�(��w�MH��M����Ͷy��6�>��'���S�%.Ow�8�^����
���`�����B4�JV1���Z)�J�C�,3VR��^�ֈ~��
��Y B2�:��ZƸ���^=���66:,�r5�{����R&������{~��6���\�Z�o�ͺX0q��S��v�1��!����s4x
#z���9�D�����_��+�15�J!�#f��c�U���c�ZΫ1Z�4��У��4��+�7���w�����!� �n���hX���e�(٤5f�Z+@��s�b��Z��o�y�{=��Di�̿oE����e��"R���H�:
[��#�VV�6h���"�<>�������*�|	7�|���i7�.���-A�:<�j_���&/ғ��c��*r��1�Y��b��;uO�	O�凌$t<fA5$-�Ϝ�_c8��������
�f�����=��ͳD��2�g݋��m7y�qbP������	ԏ_�[���@>sg������k՚����c0$����}(o�'�M��b�ܰ�[=�$�ܢ�[���ɬ������
�ӕ�7ԕ��?���)E-�J��`��sa��ì=c[�Β�K�dE��n��*]����i�I��,B}��@��T�ӺD2�^($v�$`�JO>�C��ot�eHRMe����i��mQ���k ����)�p�ѓb Z�7�8Ť���_s��(Iej��p�z�r�e���~�:<.�ަpJZ�W ���,�?����p ��v6R�_�):^��{e���׈�(�I�a�B�q�'�\�+�����-����j�_�֚=el9�Ի[���&� �|9����t3�Nr7�"����|E|�O*Vjc��ޤԧ4�=M*�Tk�\s|�y������24���C|�I����{ ��r�ݑ�Uw�GMEE�ȫ� *!$�~Ô]j�i��,X��x�ю���!tkF�T�_{a�O�89;k�������� nP(�f�zo�׀��wV����uZȐ;�j��VTӎV�r��[����J��R,Ϻ����