��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���d�v����0�i�=\��A��?��� (��1_B�f�	�Ѻ+|n��y��Q4�]�aY�����*2�y%����>��������K������ �
�D��z�z��C�y�B����
_�U��hkF<�~x�ܕ�c� 9o��|�~�+h�PjA`�z��#1LH�s6�"���Un'��jg�'g��xwaķ�E�ҩ��:�:K��� $�;a���9�IOVy�x~Q�XJ-5<^Zq�gr����l��"Y=%�_����Z��~�ڦݼ����݋�O���.Ÿ^rk� ����Ұ����໛�4]۵Y�e�݋��y�]�-
�j��y<6��3XKL�~�g#ǽ�
a;ш����R�����S׿I��Z !�˽Mv���ʽ�R�ܟ&ht�˹�
t�a�kC�89�� |�`1�1�3�s
��s\�ڢ�ju��H�{K�Fmh�Ykk+ĔSSk�h�mF��Z���=4o٣{̟�p`ԯ+�&�}=`�Т��ݘNf����ujI���8�hzN�,�*�?�=���Ê9dB���3��!�2{�����D�dǎ�Ib�d���pـ������<�S��^Z��\t�E���B�>l�el�qދ�����?ZT_Z�ҫ�6"�\FF'��!�qسd`��p���c���5.��/s�o �+�N*\�C��t��-
��I��Y�b���m|`��������$<���.]tS�a|K���Y��6��:�R]H`,���Вe�T�/��������g������*�ʪ\��>��׼���7�E멳ߧ�@_�ѦE��8�r�1�>A8s}I�q9���� 	)?�� ��*�f�\�"��/�v�F�圬��t��Lt��E)��̶�Q�`��L�g��t=�(������Q��:)�_�mh�������G�џ<mM=��'R��!��kII8����`8��uz"�6��3��� �DA(�g_�����9¾(������Q�VIY�k���蝣��`�ܝ�_Qlİ�l�W����>6p7S�=i.ڰ�r���y;���ٕ�WF .��
�?���lF� ��ҭ�1�RdS��,���z��)c���<f�����Þ���H}�Y/�7��?K���g�||��37Tz�ő�����x�lT�W��9+�_���  �]���1���{�r��'|����=���pnk�Yn5@��M�\�A��tD
\���6(^d��@�pW��Ry�I-~�� pl4ih��."D�p��y]���P���������q�k�iV���ft�ɟQ�݃xRS��Ue�v=r���,��%YƂ�~8b��/�C!]����ޠGG�_I0��R�'��*�K|���;>�8�J��.���#���\_��%ZB�Y�'�����@�%���d�e�1�W��/�l��˟���k�b߱�C0���᠔l��I�,��F�΄$�"�2'�LH���Q�A\�����۵�L͏��$�f������I�ڨ�R�E3��Aoブ��<f��f���t��Zɟ��H���Ih���r�r_0�Yqps���T(��÷�u�/�2��[][���	?�Q�$��ء�$���x�(�����s:�|}W�b������� ������v]������126�N�rX*��ϓ.������sR�~d�y��߀ٳ�?���W*���VMc����kC 8܃6ZA.�����;޳{&J gh��ރ������Ï����N5P�Ŀw^�;?�3QAb�8���K��7i�m�5�e���M�C�j(�)HF��	$�J�	���c�� ��;�H�%h��lYX��W^������7S�l(�Nݪ��Z)L���v�p��3��y݇\�����+���\�����`�Y`�[u�$�	�S�=ٌ�9z���{,�m��|v��f�Bˇ^��&������5)���[���:�O�M���@�g�v�9��4���BC-K�0��h:iC��o��Qu��,*{K��':�1b�"�r��A~�ƙƳ�2s<�S�����?T��y�������ә߄��_ �=��ⅵ�С��y�hz�J|���:��k��c�-�%�yfň�p��� ���������W~���� �q�^�a��?2���Șg�6�_�տ# _
-A�;�� �V��PE�/�#M�i����s�,G)�O��l��/%�S�ڗ^�9�+HO��������2���ZʗP�T�����?��ܽ�� ��lB�07gpQ�	�#�����R��N$�������#���*q��VC�j]�C[�ʁ�NRNyk��Z*���ݾuAj��P#�<&�B.�75da����r���D5���"<ue��U�H1+�c�٠����4d��!z�:k#�`ظ�L}�-�z��.�ܜг6�_fH����� ���{�&/��<.�*!Χ�i'�W�m�^`��{:�U^��KF�`������h�r�:4�`\��+�B��?F5I�x����~�>���ғ��,=�f[�8`�)�&��I�$�r�ʀ�k�׸�yW62�-〦��ú�I�
t�O�svy �L�}K�b�S� ��$�%4 �� H�	ر�\[�3�}B�T�鏃 �Dwюr��c6����R��+j�v���'�����C��wuԤw�$A}�I�ª�MXl�^��$8S����e���&4K��D����ǁ���1��ͪxH]��HG���WZ�ww�ͻ{5�a �@�YL�]�����ǹ܏'.0A�lC�<�v9-;W!����ӝV��6�F?��D�SDeM!L���}.^x_��ڇ��f�ìC==��v�oZ;��Z4K����ѷK�.��iugA�M|�(!5��'w�,T^��Z��w��F �@�a#
^ӑ����;��n�<����x�tG � �X��(<��j��6�$�Q���jy���o�'�^e��|�i�*OScgr���=��	 D?�iE��^����I*�Y�fN�؉����GK�OGlP��"M׀�,��b�<�k�$�X5����#SCHg�2�	�"K�J�,r�d�Ha��  �����]{�4�U��{��mhg����R�(2�Ik�Q�m���2��:W�τPOhO��d�%��^E�~/ZMm-Y�m`����_jR6���7K���N����>�/�����˓rP��`G�6$r�:�]�	��x�[!M��o�Vm�U�fUg&����m�~vbK�+��p	��=f9KU�;#���!U�u�� ���<�d&�>�C�6ks}����?��f��#e�0C�ol��`vӡ[sI�l��}�6.�����To{��MW�K);ȨL֜���Č���C���i���U�Np��	f�	{<����N��C-��66+�#��TK�o�Ñ
Ŭ�ҏEȸp>���&��l�;��e��	��ݔ��x6���W[�:3^��A�j��&MBJ C�M�cV�G��>�>�s�{��ֹ�a��"��t���9>Z�!�_����'w�� �`AH����+%'|���c��4��n����D>^r�{��j�?.��o��u�+��a�R�gg���<yVW�vd<�9m|����cZ��\K�x�[\>8�s:��,:�9 ��=T�'fs焟�p������	��Lp���2n��y�+=�_Oe�mDxE�=jp�d��$�.�I<#�g�9�����p'7V.�`W��my���.��<��m��%V��C\�l�*l<�S�ѵ���|ӭ��6�S���(=� �8n�<�N߽�(fx��!	���A��3�/a����|�ه?�dk�W����l���Yfw��;��|ry��O��{hq=�.�o�	(�<\�M�\`T��5�\\�$	�^R�K��:��Faa!���y՗oHa.��k����)������G��e�݅�N�p{�+��%�LoF���f�@�d ��y��.�v��B_��ͨn_�����TK�|�aI���
�L%�?�M�D!h�+ x����b�J��*
�*�����rD�����/� �=�|�lԅa/��rO�Ϣ��՞�sX&�E��SC��O��Z���k�	��+ )?���������� {�;�� ��� �J��6��SA,
�M�:)NU�@��؇!���`*��\}�j�6;���#��Qb��3.` �!L����NF�Y!���L��k%=��cI�LF��?b�=h��	�a���D�@�FQ�H��@��H�cv������m��y%�u�B�WO�U	�Buc9�T�X0/�'r�? ��Ua-�	������@�7|![Z0N\	�������Bi���	�rޱ̟�<O�\������Za�� '�[M\�2��L_����hyO�^�[�
-���_;��5ӫ&�P):�<�#mʢ���G�#mP��2��p�H�kD+cN�vO���x��K$ѩd�95J��˯�x��.�Y�)W��W"k�~�3����o�Ĥa�Z�hJЏn�l���Ase�f\?��}� �����������XGJ�`�d�Љlߙ{rY{q	�I�l�8���L����6E��f�k(s�
��-����#��Y��� ��,B-�"�{�\�z""��m��U'2��9��ƪ��*��w/T$���1���,�0	�5����I���>�P�Bs���!������4K���p�#*�T�r�4U5�t\֘u�<��YTĖ��R	 X �-$?���P`�M���5֓羨�
Lx1�W佤� E&�~�j�� �g�{���o�&&���t���&�/�陂|3W0aS�����hTT(�����j�o(�j���	�GTS��r��B����GQC�r�Q�8��W��*�H[��yD��Rq���>N�#�>ާ�Ȗ�ȝ��H\��¹HfYSd�ҭ�\�	h��e�����M�믞�D�Ra{�C���J&�1�67��%Tt�4�*T���\�k�W�5�q�M�z�sN$�vi��"��*K��pch��	4��"��2��Ɔ3�ȯ�
v̬m�0�!��q8r �G9����FR�o�A�(`r^��_?��w�c����q�֍��d��=�y0U(��@����WS���h� tp�:CF��A���o�1�?��;�s����x�iS7�];q9���n�S���Wg�A����f�S�g3����b�`�h�r����^�nX*oЦm�����O�@cG�9�H1x�Ɨ����k�Y��3ZO�g	;)�u���	��VMĐ��Ȉ�{֪v'��#���X���!ɻ��K������\�$�'-�թ�r� ��[CeOY��Ѵ�Q�ObtZCx�� ��Me!�[8�����nˢ�l<��½K7����8�X�2�����C��!�\W6����.�G����v�0N�_�{6���Aww2�]Md���dc���G�L��$z�nD �������`�P�?H�Ia�'�0*"%zU���ST+{�KlA��G�ɱ����������p��P�V�L:�DH�����8��u�N�'��I��(���+�r�=�N�cyr�=WR�V�W=�E�@�Zg�{�`�� �oE�9�o��秓�Ɲ��;�!��H'&�SS�ƣJ`t�"ߩ�
p B��E���$�d^ꍩ!ĢQ���q�+D
%�$�;�Ԉ��2����xd�N=V�ݗ�`<���Si��>Ն*�e�z	�M+��?��v���ɬ}_�T�~�a���^ �* LܤE���E�77V�����{�9�Kl4�<f!�&�}�n�[���{r��a��Ul�#�uK=�A�q�M����B�]$���bTH�c|�RP5_ݾm��YRx��_#��!2>�]�m�Y�=�Z+A��Ӻ^T�J$9:@D���QhZY��s�~�����&j�
x��*i�bP}0���O6����e/������d�e��g��O�t��$4����ؑ6VW�'z���{�NG+�Z�A����\&#rRw\��������E�eG��>D�r%�*���_��~�����G\x�Jǂ}9�rI�@����K-C�$�b�.]�k6t�s�ף�bL�d����C*�V;�/=\~k㏱��zIR�-z|v+g�])�}du��}r�}/����|����i�2±8���f���u�}��w�ݍ����!�����8:�*h��R7��:ϯ�G�a�O���%1j��\�\�oLGx##�	���y�\�=?�0a��Q)�ַ��-�>�$7y%�"0[ĵ�j+�:˜ʨ�3��9%����B�����D�9s%��<V����?,פE7�#�J���
���sNi�?-�>�w���Q���V�B��)r����"�j���?���S�L����ֽ,���X�@h�x6:0��z�7i�/}0XR W��".�X�H������'(�I�VQ[����*$���ְ�j�Մ,(�/�n���SUЕ���Ϗ�1���-�d���IӚ!��>N���˗��!g���$�s'Lu��c�<��u��ǹ�
�IN����˛��Ux��Ƿ���:3�h�Tp]U�PC�M��bL"څ�-bj6!���=c�Hb��'1�K
%���S���IS0���L�I��2����U�
f���h.�Gϸ�`�n�͵cgy^��-BXl��N��
��x��{M��<}F�t0p�<�(��2��AG'�j\V""ÔĢ��9���ڟ@�T�;Ԁ�5�s$7�	���^�D.&��M�kz7G���l0�$�hu��}_1X���ï����[�/��H�ۓ��`g�l4(kbm	��h�W�l��>F8C��|T�j���݀<tc1VsE�����v3��yΚET�>l�H�h�z!���&�s�����N��97D���*�v�5e
���.��z���F9z���أd�����^V��#�a��UL��=�tZ���,�R�c��aYc��͵A£���  k/�AK`�����D�q�s:0x'�J>���M�-�W-8���;�Zv�t��gڰ2n�����:p��YVI<��T�����ۈ��	��4��i���<?�E�*y�0���^�/T���{ l��?3{-�Y��`��t�et���&�UH��kq頳��v�?>�g��H�n�?Ј�M�I^E$����w��ί2�c���p���:%,�q�oAs�0;�r��,����2�� "�� `C'�Ap��O8)We�u�o���]w������>���w"�D?��
�N���"E�e�H�cm5��3�8i��}Z����+>�R���(P8�Yˀ��~�����L�iC�E9��3��K�[�=��y.�-�#-�H����KP�5@�i�y�����J��U0s���c��2K�ٿ�a*܅���,��N}������)]�3TE��|eu�o��"�n���'��c��4C�$�I-#$k �s���O��`��H��5�+��o6���S�P�T�wzҊZ]rx�������b39����p|(>��=|Lej�"*�G�Ȣ�5�$B�洼R:�9�� K��ê�_J��+)PU���3͞��VO��a[㻺1J��}4P?��x\����9!�5���qWn ]���X�F���n�|p����/�}�V��F{��Tt@g�n�����
����a;[��l�\xQf)*n�~WA6U�(��m�{t��d�����#q��ty��QCSI"�$?�^���������=2�9T�i%u�`�����8<���������cQfK�֪���r����55�,@d6B�:�����~��Ux|�g�{9z۸��z��88i���p3VwXFT��\�5����N dg�M`S�Ջ���>�y�pH�_[��$�%w0�t|��+�}�/�zc*ޯ�Ɂh1j���B����e���	KH��m��A�>�(m3��ۘ(�7<aڊM�d�ցo�N�K)���6��pg-��%������\h��|�VY����fhr��5��{z:�8{���I��hByS���Ζ�G+����<��w�ֆ��>�~�N�|����~/��QU���;>����}U�Ӽ�F��������X�Ύ�����w����h����o&u�;��$���m:���!�6%ϡ\kx+�f}����A��EW˕�ԣ�HK��׊��uo\:h�<>]�W��ʒ��8P
����$d��Ǭt;�Hm��Mc��^�t������h�U�T�Y��H�G�c�����!���8c�3�Z�ANΊ�*��,?�q6���aD�V�<%��1yy�䢷���O�^n/�J��3�LR+t%���G���R	xY����1�5 >�V���҅�y�   j ��}#S��5ѫ�����lu&���-�e��_u��Y0�Tu���s���aOS����R��R�;�7��"�-B�y��K�����C�Ҁ<��&��ul�QZ��� i�+�������Í�CE����\=���aGn���� r��I���* �״xzJ�BυL�y�G����O͓�B�)����\�bR����_+wŭ�%WM�ߔ����9�&��x�-�z]�%�����e����	Q���߿�sʚ��A"����x
�����2�{v�30�*�����y�-:�*�ǈ2�?K�)�P�.��ؚ�:MV�!Z0��.-{��J�tP5�ńE^-5 *aחi�ݝ�!�9�W*�Ѕ0��z%�H�������Άޚ`�w���v�r2�K}p�zlvZ?Y�ħ��n5D��H��>��h�Fb���ZBX������p��3w� v���ρz�B|�tO�\�v���J�k�BUAS�O\M�UC���&c
4`-��8��_�~��N�W5�6sC�m�-�}�ސ�����Ҟ8wţ֛����<�#k|l���Ͱ�DN�1뢃}9��8Z�*>=��l��	��̴i[ ]� �F%c)���nX>%�p���q�T��?���"���מ�w������PM��n��/,�fo���ҁjL�W�i֗��G��
2�$ �̠#ψ.�^��ju�uάE�>�]��"DO��XdY�HdT �߈����."��O��u�#o�=є��+}�G�J3���;''�y��^����X�%��Nr��n�ށ�9�+���½�;�3H�"7��3�q��g�~fX�cR;�V�y҆_%�P�_F��5�>2�����-����н���b����nq������|痑�Њ���H眣�D��3�)��	�[2Q�w�I���b����][O�^���UUxǾ�ޞT���2��xe��k"��`ǀ�Q���ֱ9�%U2;��J�xGS��`�� ���<@���T�d��
?4>�
��I��<{�ȱ�c�Y[�����ڡj��;1���*�Bc�c�����:�H�D��m{��&��\q�6��k!���0����pK��G��b�vɑ��l��[�����8B�~���X`l�t���@MN���#T�G0g�,N�c/m��R��(�7H�@ޕ�ǵ���~7P��b��s�����jB`����1)\��6��<��Ԭ�7O��W��31'��.��C�=��[ <�w�(3��x��yd��a��4��]���5$d��0I�~�������E&��Ef�%�����X3��8���U��_S��'�0=��W�� �}(��q��כ
���7+��X�İ��5mп���>��J�ݸSCnN*��Vz�D*oDNB��|\dL��Pv˔���A����ȋE��f�3�<ͻ }-D�vۢ�Խmo��7yen�9;�r>n��N������r�V#[�#�>��P�"�.�y�6�Q�fA�ռ@�gg�CŸ;T�		��?���%5O��nD�v�~�4.�c�%�,}���ٰf�̫�҆��E�J���xU���~4��;���ќ;Ν�8S��'B۵�,��S�!��Q��]ǎ�66�f��yUV�0e[̏�9��f%�>�>v���{�!m��O���x(�q�^#Q����G9��E�����e+ o��v�y��|5�9e7?��S�,S�<fM@o�쀙�u
F9R��6��7I0����|�q;O��>/���M��j��rܽ�Y.�+3���F�:�,�������#_ӓ���O����h�h�0�G�:����DX	e,J����:3���Z����l��`�ݐ#[#`�� �0���ث���u�MRr� ����6V%�J*l>�+���5�	�t�����K���.��g���s�~���bN9�؃�� ��jZ�.>��Տo��c������D�Ԅ}93���h' MS��MŢ;��S��#�}fV��Mշ�`�˹�R*��ҢL^�w�O�
��[*�T`���m�G~L?\ �M0�