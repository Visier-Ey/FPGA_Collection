-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "N-2017.12-SP2-4 -- Oct 23, 2018"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
sUvyJrPG3iWfQeo4oKvkWupzUJfXRgtJbyqeGg/tjCjlUspxPaquQIXixR3FMAeu
BCPIkHoPjR5MDzEhLUzIcKwYrZHi+2/S2Is+hsq9zIoiCgAXXR3C810vkQ7s8AQQ
TPQ3Baf/3EAkj3WHVe7mLzGlyXLW5cdp6+tnBgaQWfM=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 12096)
`protect data_block
51RpQqAUf7bwZwzfJZpPnkZrRVLWj6G9bapmi7q2eHfYLgP7+tlvNDMs+yH8A7lt
booyhp8Zc6a5cXXCAmjAritlt3+r2hCDLGXzlVxAoKAIlCGRy5sJxw4PApK2qL1d
BWBBwvgo1QyivKWAWBCDOZClHQnPHeicvRXoXL0/llMhRKO84zYijLiCa+BUkwji
9B7wqSs69nUm/6NM9hT1vT7b418kzPjRMvzuSpBOQQeNnmiV/zoQG2ON0NvcyGpl
AI0zazwVK0lqsWj9uLJ9YahcsvqCtKBheUw6rhGpedFEb6BJ19RvG8YW1C4v4Q5E
l5bAZmd2QAubieAHQlffpQIkThiyZRkq+FDhAEFNKNtvjiqRRIqNFASPN5SJPtcK
VZMm4SkAiGurE6pu4YCNnkNMaDfgxaQ0lOdzxB1p6TRUgfoqGetiP9LOW4oBvNhs
+ZFBIYA0CGfI600O5BYY9yGilepeSUj9Xk8PU2xCFGcN1+GG8ty1cH88mla6CKKl
X/HyzL9ICSrmN4y76MyHS3BUtLzQzzZ7/w1XmC0JEJFjxAh/y9Oo+aAtM/CSZ8Vs
MgvqH3benK7usvo9qka93aHPpO357zqYpZl93LRl+GLZii0uks8OHoCEAEYOmUBP
XjcKIdIGY8FJika0moT9ssDTKr7eJTSXO+Xl3ULoW4SBG+Ln1Z+f0Kmc/c6ENRfe
+IYGzzwOAdPJkGOInc7EetoqvWs4gHKQGZ5cSfuq+l2H0vrCoQllnQ5F6YtlelAa
lMBNUgctkY4rqfVW5Sv5Cf+ofoDQWyFr3ZIkVvejZ4iEjM1Mw+ss2mJpUzRuiE88
FfmCIbvY0gx8cSyyjg+GJ91xv14c+tAuaq23G1h14Ky8N1nvxd8HU2JXzsY7dn9t
EczhE/BS5p0Urb/n+fa90fZqa0VVARhk6CiUFmlxe7N/hgHvSYk8aSNzBxDGGwZN
pYuCvt8EAbepidnZdyAP4zBmXMhnyC3o4oF0PKPaMV4nZkfy6S0cLUIaQawttl8U
ckl8gSBiqWFHyS6WWCpkkpnRnSQ3V94/tcU/cXMOElk+cMvLtCJM0ZmPz1Tc9lrl
FYJP1FbKGbXn6csLbhilY+g/jqTga8N2g5rEv3vZU60ejA+7ByTUTa/Z9IVd0PzH
sPnbWxzphj3evOjcTYn1NExgf3ce9RQdSISMeE/5C8lMqR/NqPnONMHLQ0g8H8Td
IzaNz4AHEkzCpP8/gu4KknHJBx7glch+6WeVw7+sZh5kKjWRizCnNeDSJSYs3ZOK
cXkhowzQ7U7SFv6q7VqgZXRBteS+DD7pc1ZkxAnDXYjgoSTs3Ltbgdf433hkVuzh
HIebIYTFD0wDg6Jks2jdMtuIGtKi/EQ6raCT68vt8biWlcXRubyIcZSUpyRuHKD1
UzoS1ApV59zOlmAXfjcwDcZlLh2nLNT+8ZGSifBz5Trb6cwSGfXFuXkBJlrl90Wo
tDEZh2OZtxeNqHL2o502BlXLQtm80GOiqKJLWkOA7vkWVxFUhVkIA4T/adW/hoEy
L92tlqPCj5e7MTu/fSElbPE8tY97a8pP4xQyxPbNmM9NxRJJ//qeaDMuGWsY1Gui
/Tt/zQrDYR4AtWRdb7qHicQicZnHVYNkssbwDgDNAC24JYpOHuMnfANTIPVGmRWS
ivT5RewfyTrQwnFM30s6lpgGxzllN6ndEmPMk7hMA50WTn4RVPe1fL4DYCykucTD
fkgZDuGmdPKEfQ6fNmdj3v2FqTDfDR36hJ1ZiQXOVX8h6wg2ystj7zMSrvLoRcqz
HTV6YoKhWtQf0dcXaYreYX8hHiWnI9qubG6ydlY0+GbUoWiE9PL3kmq32mz/IrHZ
6jGL/k+RtNjxqlx3TuXBbEBqo7KPKBgQ/4TS2nw1B643AORLCy6DCBGNJ25CKKIl
+nExv+SMSZuzztAJk6hJ5eykoyXkKkjAynzdbzWR3pHZEdNcpdujRVqO9xbYjg3K
VuFzpuw5edsptAgAODq2Zegpy+p+0zH1i52kXinJ/0itV5PwGnlr878ETUj56S/Q
qMxSUTeYTdorVr3rmqb+29r/XhByuEoCmYDR/eU5E3nY1f77E/+s6cSwowiuUvFP
qbGl/hrr2NccDJLBtdiGRYI05IjmgnZbalPxpuoHmB+hBA9A7uO7CZm1kWIHmWIr
YAylCvv8rgDpuYB4UTtj3S73XPL6HEiBVAqGoi6F0UGvdpGfRC7d+/v7zVDf8yGt
aDF7vaJMR8sHOWz+Sa3pWImmO6uTz4rUdJG8kHC5BfNGAyl6BNwYhASSnOk2XD/g
MCh1jXVY01XI7iYzf3Iem7GypXAr1qX9al+jJX5RjPAcrTuxh7KLlXYJZ3g1JPef
ccfTP0hUSWcYryhn/ybSNHlGH0rGQAP422c9NJCSFC66akiFGcKe9nJmujXD/T4L
Sfk8IDOVt7v2PyjmurPh3TvdDIJ7PwU9eZtXJRdCNJ9KZkQhE+3TasvgJE4dY6b9
mKCmnkoQY9WeFid+aQ+V2/Z5g0HtcRidWrRKDp+n2riVgcd5lPp8iH2a8mUmWpXu
opQ6W/9p6EhNnvZmfcC0/QUVQyXY4SwDR3jni0np7S98qXYbJq5oSYW/UA2cDFhD
9Yf8aXF7G3daVn1GKZ9weOcJeWO8ivyXttw4kTZhP4gFo16/i9CIezYLvAjzoIsW
nd0aB8WeLfxNNSofK1CliGearxFnlpgJgHKkAgbLfGSuHr2JYgUKH7K8l6M2rNXG
jCmA3JlVrfZNcphWwmQQwIlMNRrc9ytuM/A04PYfdn74XFDUHMwCWTrxMPTaJK/j
BJTuWj0SBctCgIwagiW5+rlW140kqFzyudwS9P/d1ZkiqkhkvghZSNhb1NZazY6I
FIr1An19B/mwK9asX1CYFL8muap3g98OgL+/ntc9gPVhLE2cLjrky3NgLgCFAoYX
4Md1juzm40TMNHkt4Xz5fcn+dC7kETMUp//VxMRHosCvVKZH8vvWAh+5prCSGK56
C2JaI6ygFPycCosFJvqg8bGHeVJmaR3r4otX+eZf0rSCcDD6u56kQnOH3jeGm5+Q
+BKWkjz07538MV9BvXUP47dgsK+XI/J9Ft9YSHcfLqi00brQ3Nm0IBTAVXRIm/R+
dgUI9xF5Q9jdNHfueqz8iZBhveJPlWcjYR6H9Tt2stwY7jjNz9ijqSKSgsrFeX18
STAeylH9tMJfkIW4y6qZo16nKbtDFa5OyxG32kn2j4BZVXR4x322wwlsXSIPLsOA
gwzZ4+49eiJ4XGGz/mfw/tYDgaHqIXF0KblDT5YBwRUcVBxvCPxZ1gl8Jd/vMIbv
kv9ClTlSZrb9skDoPEjfvXB+/520iAMHw4QAKLHoIgk2Rg510RQOYYt69EAflqi6
DS4yu+46+VSTwTkoAG/DZtdAGnl98ahScWUvAuMbrAD4/MMKnwoW5Ovs/GBywpUL
4qY10hPeZaGd+vWo1vUOIcIjfqHYYxrpGke0gIXJ8HKOfF/GYWONdcLZT+NJjiaA
IojzEuAG7ftpJx3qtfAK3bVmbpfXIVb1hEXegGtQFsz/qPGFdrcaceBHWwv3TxDN
A5mnuD24jcn2y8AqzqRo89H4FbD6m0YOrjfE8z5+yMWUO/bfKgmLK4uVhf70+08V
wmmMK17fTKRC0L3ifd3bxQX4ekKAG6Svs/9HftcUDyTTzKmHPFBiBCph82fsBb8u
57PF9rMWgvs+jYkUuEbT/NjUc8dmi+S0anoTl+o8k95RHer8Q4poTk34dhuTdtuF
bLASZ2NNL+Gv/h/B9Rxdo5ehSykXl1cOTQikC1flvv1VrIJ5UGnhRjGaTJ6qokku
S2ZX4Tf3pXKqzHJhE7wDqoKUxw7YQpc+Fry04MxDwNdAOJKcNx1dR+x7Gv2R0y1z
O2y0bFgMOadjlbwx3aJ3yj3PienD7ndtYW9UAl73nayWsiarvOaxA6HuRZwr+Pr/
ZEvQvW9dLUcFShPPnSDtdepK1qSKR4xsh7ZjWPa01m/WLhz/P1+Ijbb7BAGD1tlH
0QxFqELe7yn8AUmLxZ53SMgEGwEGhjQgt+eeE6kvIsosNT4KQi9Zhj8zIb883G1j
HgSvGtBmUtyMrfyAJBQEW+NAdrXkkhhITMITmHdxOd3CyZ9IgJmiZSqfBRCNU5Z1
2Wc6e72nDSoTDFZQCq5KFAEcUpbqoVPaUb2J3hNX7LURfJeHz5DpiYH+7s/O9rgf
qTDUAuH4lw00Kw5uphcI7r0jpdkdKqW32Umxeyj4WxjWqb+RhG06obrUx4srrLZ8
xChLZXwKmJja54TpUtMQ7eytnGcGql00xU4c7vKA6HA6bJ9LIHQfuKowYi8wXGQf
IkXu/iQgsb8qJ4j55vsAzHB42Z8seu9fI27riklfm180fylimMJYHt05U9TxPFQN
Ms1yIj6b208plLsVshqT+eg9m6KfCKIwyqLtfA5UeaENDa2mbDEY/yUBNlyCD5Pk
r6bvIpSHTDIZPAGawmWdYLwvxcAk23fDYK//54gTaNzP7UUQ82ixdkzcSj0dfaU+
ULQKM4tk1Iadi1WeQzEuCbtYXODgI1duGbPrlSQlAu09ZT1Kx1YJC3kA0TFEDHas
/Km0xSewMCQ76N2u86idMNzMvYW/cnzZcADM0+wYWdzqF6YdiP8v2o98MtbQWXcQ
o7fO4tp4ZRvJUkOgOdOaZe6NWVFMJqSyAM2VBTvXuVwAi1uWd0gTvIuNoUJBZN8H
G5I37i7BVtdBzV1iKbCDi0RNmXh9DDe8qta21hoSVJXgdKxLOdVvLZa9wnKyb4R+
39MFFUR9igWN6fRjse8RDVkzLL11DCIvbd18ohyJ2lQ8GxtxoFGAb8DDL2KfjqyR
OX7pHY8Z/BX+qvSGoNQi89a31tGHbHTsbeRT4r/3B6W1me5iMSEvNOk9pDskTDiO
r1JDCb35kfOvJ5My4xqnEVk+Opv6/B2Up9jlBXcSptSUqQv7JeW+Fuwt148xYSGl
6LfhqDMfoiUYnhiYj257jKMz04xRTPvuI+Bg066vH5ysCPMyq5I6LKpQ2MtchwYf
jIZZnfjI683C5JFPq7KrrSABVTGTzWT8mNR3gePLok5MnvfWsfhW7d96K6PxlRgi
WhY3Y9qKfodW6UD3Ved814kJIlzA/JAloG+g6DgGQtS+NL5sm7Ek/kIS21ke8SzK
ZxnPRewxaNjtZ+NCJa7RPr08VtxhAJYa+YSRCEQQxhLOaA8p+3G3h9U6LSIeAwrQ
Uymw//u4IOObeUHQ0QYY5/IPQMIYJOSXe2QI6m/9VCY0kB7KVgko+iy5TvD883xC
mpOcuxje2usEuIi5cNOKarM4okyfcnGF2JAsS5qiEBG//VMrEP5LfxdBu+3fK6n2
JethPyyYvDM9pD1xUBpHdC5bK/mkFNjInxMdFxb/W9mF82E2dveV9CLZSTEcERkN
hVCfRvXeExbYCUpWdh220X6kOv0X1x03BNHZYrJaEQ7ydCh3ehjsdZ08zNk+xl41
KoDOiRh2SSCSxhDQzF0FIRmhhjEsNNdC1ovsVFX2NV+Ek3r1nOT1YuQV8Y6cWDK6
Cfdj9/ZO33YcFW/6upmPrgzGmajanxkH1p373MypQjI7ax/T1RJyPtcg0KBDKYJX
fhGQ89uYwI59ULY1cuNycCNBsYFeTlkVenZxx52vmF5Yc7DhzDIEIsRoNeO7+9Qs
PyuDOvBqnntEJRWT2Vo4JMHM+7WachHZZ6TX3hz2fwFo/cMvKixJjIQWJbDVNqyB
IJxtnfS8Fs8M+dgaUuUrtpXVmqva+N98mVzteOvEVJc8q2gEQ20kodBVBxJ3y/Sq
Voq6dabiF6efgyNnjJ1FmJ5NGVpU1WmWBBKp8sdsSkIsQYwV3myDLI+D7rsKJKhD
4Ud26R/xWc4FhTgn/yi3IY+DRYkwtiEsFw38t2LP+wVYTMkmBB0IhPKVP1bvBefr
C5pTk9ckuMKRPyIcnTUvd+9boO21GNqCYPohxdiB2E9qEcP6eZ/BSNey8vElM3Fy
uO/JQ8ctG3kHA3aR2j0a6iGUUX47U/s5PwsIFeb32Otk30gYpyzNKtvSCWCYpN94
Q1M2v2Z5Y1em0RCfBTiau8/gWYPLrZdvQBBnmE7TYQAPxEM9R3WW5lg5hihe5j0N
ND6hq8ijT9wuyLt4voAM5xAt2mU61YMWSwzhJ0AptSpceYDSvnZCc+VF9FSVaBQI
B4+ZpWtyJCt9z4oLfD1Wz0MHDKhW0Xib2mjiDQ7fZTGUq5H5z2dVlWC/CnQ3gAV1
EDcsPysBaz03mrUU8eoAMO4AzRZAayPZkU12gSQbZQp31JsKkbfFb60gnLFfZ1za
WhfQIIG8bDPeqCOELIuMtXsTKW6qXGY5ThLXxjE1SvRzahO2ZiGde59HaWpoLGpk
VKoJVq5FkNowN+vob2VrOBXEbMai9z9R25Q8szKzRQHWA6SRF/ZTvkofjHZrA6eM
6DDFf+b4EAn08YK/MlvTqmMFostTVIwCYpA0ADZYiKmITKsr+n1kcsXXY8gHmj85
Ta0+3YJKpHYuwKSytOjDjN8DMjedq3cNdi2DyHTPIPpG59ONsyWV2fGJvYpuRJxS
K1U2jWHxVsOGn99W0Vl6nM1icUogQ2p/HrNWi3sg/AoCdzXnext2HfZ2hHsCYp4D
BcdtEeWJ5rxTJOUD9XVIlQhynYKF8WgHSWW+qT7qIuY6vK/x93JMARV72oOdubzB
zHqM5JXFIPzjP2Vno6SOK+nDCANV3Yk5UJidih8kLMGF1OtqheuMnqKCMCLZpfsM
pFvMJH5DB44mYY1JUkKThnz4lNz4FQnJ33GYk2GHBtDkzl7LOZ2mGq3dS5qeo0yK
IQ2fS9InZKIMrEogKw71BDZ8MLwx66p2j+b86f+BssIJZP9TOQEdYnN5aWChqi7p
UcnyE0U+GKrQD4073mFLEV2I+GMmXGi1thaJZBRaECnT5T4WntS0kAtS7KXR1W9u
bDTIrKkls0kRLhl5u7B4jBozZVthdqu82TTJ7F/7UK0iYquQHj5MYGj+DbdMdfpY
khYzVkPM82MKLoZ12Ro4rTphfIgDNkk9Ovix5M/RZL0AZnB1g8UV9E93xZZZuHpV
8d9pHpChzR6Myqt10A4858mUjVz9fy2XL2sniHoDh9G64SboPgXF8yCiHWc5hUy0
lM68TTVOoJdU4hwVMWHdxbPQaomRTlxmmFgAm76CiK1f4dF2q5yXvIm9Hk9rClNf
P3PIfeT2ym+/62GUyLDMK+XHxcTsTXIMiPfau6OBnMrBA6FgjBrl2HuhLVvpLcZ6
oDJ1IkElBYIdpWh3ypq1UB3a4H8U6qLLoTSoCC5FzyMUPxI4tRHCCUUKFxdGDA0f
u7UnyXqC8Kr+g5e3znIeN3MSGe7runD1JnIHXh7D15wNBW4NBVCdBGqHFo0xGIQV
lUKAWo1b5/9/HIprJ0ZdT4OGEIAYuAXi8xnJp20NFk3QVoa6FKRBj4+Kfo6J6NUm
7QDncN9D3/k6qemQ8RIRuh0W1qQF+HT8HdRAcdHJdd6nJTFF4ddGatiBNtEtrolO
qNDCNLFYAJXBXOjb4WPkQV/FAsBJYhQCQhdtkAbBUVR/C64HPhtqZwnuortLWFL4
RhxatGYaWsTddX7fjEEqR5zm3IaCMr85IGjuQV/1zzpy5uJnGW55SC71iTyPjBsN
+mFezZaB+y5A3XShWi8T+gkF8TwfvSW24aw+WtVA5Ub7iFEW610j5N5/ECHWGh2C
oP6BefXxTBilltQbeQzXizj8HQsMupA0P/aykG8kkzqLnX7DttwYBWjvqWwPmQVM
ZlAK1diOLmgS06QSYvoDsox6/BtJ56FDCdzr5iJVRyYji+bRAo+8loskIs5QUKzX
poHTmJpoXTLK9dT/WRSPJnmvSKXQmAJB3OEesamoI+1h6KLoS1kpwFGa6kBtikTQ
qHO7cx94lvpTXnwOrJBcIlt6QowgEFdjcgjnhTwz5YuAtyl9F6zNcbOxFJqe3jP/
N+L2GdC57AniuC5hVGTTcl8CPwnvxV7HzyIvZoSYR2Q9/sZiqOtNlQSV6WDZ+8P1
31/fWhCP/Y/uB2KHcepRQUsyUUnq0BhYP76jNL9AP/+CSJ1Uj4LerF+NXfvY49o1
Es1j1GqMKDgm5PA3uxoVrwQyXK+ztgX/ABr8kSMbMXL8KL1zp98J7fOvS5xYKpkm
LhgfZcQXayNf856ZJKwrlL49hWVu86eZIf7lGuvH7RW3aPUIUJUkXlqI8R/sm5BC
/0zKQ3s8WR0p7Bolc7seE5nu85hGB5qjoGRw4Kle3HM3uRW01QCZRK5aWTzQ4jk3
9SmR+Jq8XGBQf5eIY4Nk0If7FeZYpPNrDEbeDhAgRLOPUFB4LFdEC/cn3wjvYaot
SUFeP7LxVCeFzxNcT8KkhY9H5TJPKva9PRdLjSj1LTAIkzkGRZmLLgZ8Ea61XALc
BrNlza+weJ0EarAT5x8814M7BQSiHUZBdPvGNxA9QM/2nZAujnhx0dgoZRue9GLo
Gi+1AM/Os9orplXtrCwdddiktwtShX5+YJNbNvNxtbRGiWNi+mCiDcDjMT9HAWKC
QWbwo+56vE4oGMrD+yhJUXKtiGVqlRjytJShqXPhvjexK+PHfHUfH+xSbF/3oRtv
MrXp/8xKvZQFMa9Iw9IBjAru8hWpCmJp4muFzuy2LGwF0Bpbb7lh1NRRVZg7KBmR
vQbFX1j4AdmKa8Qfke5R7vn8IN/kXIHa8qg6jSj3Mkxyn4zKkYs9IYqXydbHNxTZ
sFs7/vQBjPcuIQgyX8QgsB4xfQw/p7yY0I/1Q3lv66J6Q1kCux/kmKC5vAwmG5m7
Ss/MiDYWckYhgVecAcj5LQAs8rfbFfkIime+bHtv/XrhxzJYtOSU1xBgfL4jEA1h
Jal+r0WO/KEtJFxiTcCQdxbIr9rlTHjVDmtcDSr0ViNwugg8esKtlekKaLDeDJB2
aV/isgwcui3lIhNrnvr+Yw5rQ/57padwWAYbpEVz5HIBgsafGPdjvIwV4MEpmiXZ
siy0cZuElQ1o+SUrJLlObMy1Zl9fIZdRsBjdkpkwhuOXKutF7sl1fzJyIM1b4Uz+
nn4GtS0jNxutZTXeEbOwvoqhgs0483lSjCOQJCnzBnrZlyw0JJ/RU9VajL+Soia4
pzyYXe0mk6/WVv7lLpGIzHaWfI+q8vnP8bIR6hT4jMaFJALGFr71LDbpJhJ8IJ4C
I4d1swZPBi1cN1tO76FqNDpixJ06aMycrE0oH5Hv6TklWnQl0SmmLePL2FfxrY5h
1GZeUp/4wzszn8MlAvzATghGDCqIZ9S/PjJkxdvWp2oR/bGYUgi2SILtcv7sB+Tj
LopxRQfEbzrc5Rf5bJ6ZaqEqb9Zq/YJ64UHKLn4KUvLW7/amSc271sV8Y3OhfN/a
NxF3ShSD/ePYQSINAARSoUeb7A+0QywGw4HlUK8WSRcXZ+gnZiOiXKZjXxQUL7gz
Tb+XU4+HSth2GUftU3/LpgOeFzbJqPr3NIeFOfPm1kzhxCyjHV7nvKkk7n8MMmbq
1phd/QHZAkjuK8W2lIIANy3BVWPtxFZ8Q82ohOx2CQJOAzDnMA3XcqiFR5jbzy9q
0l8fVQlzbmIQsI0bUfd/oO033TmKAbWkEMaTTF9HN84CmAGzNF4m3eLK6v/Q6H1j
mhUoJ0lhgbcye1RrZNyIr4/DMIKRE38uoTSnxWNLrOIDgxpOOFlRGKeI7t6ervcc
cOu8bHLEhYHwm2NGIV1QVZH83Vz39VyO14erJib5vtwLd9e4Km3asjg/xxx0NTpY
nP6N3gpGYdTN4z6dDZnn1v6JSFVwB53OfiedFpJnHlOxVaHeQWog433S5GhXSxdX
kWHjMqG+BgxfNcUuOXOezkBUehZAPTHTomEa/D2p7xjMMj1XzIF6+bqT8rYBI9uv
RfLNComq5laaGo+MZfMOoOb4IH2LosfrCiN56jXcenmpPMip3Ag4WIT2fRM1CnDP
hN9PPWn1ipdsWWHyTPHzaKOQqoWEma96Ga+AECCG18v93Yf3YmL4Xoe0dDgONzdl
WMvK6hvZ1tCoPqMRFxWAyUeIeaGb4AcwWTSLkZLdn3uGtHdBg98M9lterySSlJjp
Dsmar4JR5YDPyL9areeG/Zr0CviH4np2FKgtkWPQ2Hr5/vB3kVQKp9diDRyYF2EV
HBHD8mfE3a9FNOmXq233E4i+eZKSMiPUImhbZUxOp0WozEyrRxUStKARmxQolI1d
9Skwv3s2iuEj1hLzozxWbBmaMcx1adSkfVFOSn8c9lIcK5TRrv8BvyIDf+Jh2C8b
NDYVoXcD98zX+ZP3njSSt58LWC3CsTk57P6ZML7VSA5H7B8jU62fKSQwcneEiHFK
Q6mG1T6qtVStqljtJPsFqOaRbuVyZNzbXt4lymGEVBpvbr9/IhKgm5L12mqkds97
irxyVYFxjpDMKVfqpMZKCnGx4nA7Yo5ZAhQTReLmnMDbCrrzodJ4zz+RTqO1HJEe
lGiWC0vPQdeZLEHcQTjwIpJFJj3XadI5iASLm6yfXxLbm6dJzKQHR32yXqVNm7Zv
Jv0Qfqnoy91pEC85wEbsrkkpCw68SZOkK2+cdf8lpXkW08CgBmHYhAEtWk2SKPPm
gzH9hzvKq2zZmmMVPCFfz52YgJnDuGXt0QbPo8HBs3VXoDCmZowLq4gRYqvRQniX
eTFjddZhNhsGROls8u1mdm5TXAchVDhtYfiJV/R/S8jH/zwDZX/VYLTgvYY8z4pX
Oskj65En5X0bx9D3wy3tQWEjDGOpfkpET/0fT8QI1hOzVmw5T8KAFgh0lHDL8bom
N+GssGlQXCE0AfnrSaHKvfIanfZayL69J8aFGUyGy2djr9EZamaIQ8wlAcLLdBS5
Y14nX5Puneoi/cgx1Bc9aOYBHRFJ5w8xzCVDRW3UC/A6KrKaf3qkdbkTnQ3FJ+8+
9Ll/V4uRsIX08Gz+83Tc8yM0KMrI3NDxZYM/M/1qFHdtT9fb9Yv6ri1CttqIYbuD
Nb1WdHYAhGCwRG1UN8iad+A1dpuOJWyaGd+zm+3644Hw1KuupeYJbZ6w0hSo7/nM
69c9vI8Qc4HbdyOPCvUZRbnU6M/fAC6e6fXh6Cq5McikiFHzaaLYMgxbVhIzkCq8
mwR0FynSffhJ1quwO+earsEAobhN9uXLGWPu60rw0Kg08xbhrKFOJCvOr7Pcf1Ge
UZ+ANic5iIq83iTqYZ46xEmGWjaZ3z1qLwhGWwjodazRktaE1LvXSpS6TkvUHb8l
3K+1ggRfWa5WNqfBHIflMTgt23wpjT1mFm5PzP0fcEIGlSz8CufC2dYmLP20vmNp
GwksSbZMn5IvSi4wMW7JVWXXP2E5OC01KCKycr84Jwqecn21UrZ19zZoMlBT6TVJ
ULeb0VXMVR3frETK9S7N16GJATfFdRKH/IonbxXCZmHcGzIbmOquPz2IwGTqABH/
mbnnf0tVtA73QoKMZQIkuAnTKdDxmvGu0KZKbxuCwRxjhbmzbQ2pDiVfneRRlGsj
Ss0do7Jlm17F/mjHkPiem43gtDg1oSg8lQrrYyAJD9OSmlVa02f67gXnGophfg7X
8RNS45sQYalTOKEbrOYOc2EiGUmkH4N//QcqdrfMi2lAuUSklMtYWWjxjT8ZOfxj
OhQY68w0i9nblm66ntqosayNiSSILORDuTEpqqBZiC+8nvca9WBxJ76Nklbhx+9J
UjWjgaru58/0a0qNn7yxT7NTAaGg34b8YquRanFeq3eATxH2y3yHLLhT1fmEhbzg
Rc508yNFAMur1iP3iU5I86nK7yLtp/rwRKcBIK9UaYgScAHaIUo0UDP+uKBZ9Qdi
bXWQbrQFEa6JKmpNmk6+f+AQRoV31m0jsF7V05ujfrLRrcS4f5iRJl2q0s8i6ME6
5B9/hTypZnB4xLfvE1KWtsP3N/43WwSZvBHoMCYl1hFU7T8WD8bEKaA8Ohc/COGU
urL2KvCKQ6rmceXGkP5s0TyjLa/zd47WAHA6O6fB+5DFmmzGleE++2idujAWoQGL
sk9+t+S33Tqx0fs9w6xJLdmZkitIG75tgMHXFQZ0uiEV6pQALcMoPGPrzaG/crLT
/Qlq0ndzQX4pjDwkBUTMml0sIomP9ZLQqlmLUuxjbpSQg6/adrhcxtcwqqBmfyc/
ZDvF1paR3k52K68TDp9U2Lwm/0uJT+yA9DKrSyMq/TXSXqCUzmkJ9cKsNfEAuSIH
mvWAcNPime8Yjj5h2r2tBplvLCKZ5VIfSv79bajQlrsSjIcfcABRAzbejVuKwBu2
A7X2sdFt1mo0jLpNTop/2JM1ZrnkpVZc3+VLuXhWjMyztPCiuZzCP3JGJMfKWNnK
t38U4+yuk5sp0jDcfnz7hLHky9Tf6CyOO84KGam4p3cEvlMuP5C02n7qzTdrf4ai
Muwv1cNsri7htUQcORSV3iaWjoJgPutrdo8BGeBQWoTqf0/YDtrl7/ASWtPTsIYe
lvqUwWiQa6pSAVNEVLMD6CBu9rbTBr9t6obOxyThEtlFekO2mJhuIELvRAmq7Bm3
/cE7O+zYtHTfHSjoiWFD8T8G623SBcKz3eNC3WDhYMZOe08DIT4L2bpNvzxxocmH
5vzZHDGmNHNmvdT88PmdbC1NpivyoxD0u9pb5VsY6YBA1nks+1WnsmmShc7MfqT7
61l3LU44dYjIANbeePCCx3cJIdP9ZHDQ05c0HfwYTpDY+lAN0PEX+Kb0osio48YT
AEMzZv+Ldb3AyYBLsLveQxeDa8c6iA9mAtBXCDiJdb57oTnWscEXtGvVdNcqXqUG
hf2CJJZLD+d/ZxuFLaByoEDIPpr25N6DyaQsr7A3o/VmzLO8tR70ziJpYNVDHIAi
bE8MNEiVtfpRSDlNwlu+lFw8pb4EDVSQPGk8ga0JSDHan+FIjiJ0AUMgLg2XB9Qo
y9VCcPtGz1211pDBTH1Gv7UNhJakiO8a+ZE3HXyVeNqNMxoH4x5xkiA3oXXSy0jw
PwfigStUmct6LiWpnjFLeDj+UtyoZl77JM5X/DZbei4JBXMdLX2p68SJfkImnq7w
fdafigGZNx5RbILGcA/vZ0dHWEiE/jC0VEYxD0+scTR07D/brTjfwy90zlObYO1n
lan43T8FkZMahR2KSz67rOE/V2ozxyaLnRSlba2g+NTNiOfsx0Lih/vyzAmYP8LK
q6emGvgeBtSSX1d+To2py3tUvyZqy4SzwManp4OxRUv1O7SrLnvMnWRggBevnbB1
gnt1ozAq8lgrLWKBONWLEL0kcGBnZAW+vr9iifNMUq9XydzSiZNfglGNYRl1/5Dg
5vAs2U/jJoRvWp6izniwM2jwTl99qAwc4Rp60ppdWdcXuJvaSwhRWGY6hHhqiVfa
j5j2A6Yqk8wxOtQbAGNTR2BiorYVfdgYfb5XVKI0y6L/f5viXYp91SbjvfVj0el4
OQXTby7SO2kUUvovAyRNtEW20pFh2EI2GGUdbS8i2XcvtWHdskX104VhnoyP3rNW
48ac4Pia9Fx3D3j2FsuOg6jMtGPh5ScoTqd7C5grVHcJGyBJhum6sFUZZp3AXYTL
n4BY8OnSezIpcp1PXSyYZ8MMVNDRV3Ng654j90oCynxyd2/9Pyc0mR4nzUJ6G8SH
hT+J/JpMajLgW5xbelcBuPy1589nk57G81LKySfPxbBCjpF+2Tklm8NkE2Dr5mMB
G384ncWbvt35aX8c1dtvu35OGEwcFN2I5cLk/NVkeWUOQJpMh/KmnFWNXHjtol4Y
5RRJhZJAsKcTa8uJ6kvMqYYQHi0ukiMt/QQfDReBNzbc9IeuF4O8kflkf+oaC/mC
ySh6ESStARyXN7b3iVoKmThFyt1im695xhpt+dTH0eMmanKdGGDO7kLgsAAYeewi
rxSS/yreNJsKqtbOktNTGFVTAIfhkd7iBWVs79ZYjy6fFk6UP+0nrmkD5gk0M9X0
sYNRRmMJTESGZq+qxSSmqqUZEQkt6lduKn6eqSdNivRnGXBej/ip1/WqSPHH5s/N
lr08zrLGAUs2dO6s6oVC85aCdCklxqpI0ZKj+D2XpDMVtXtGcPl3ALg1urf9Uf58
5wY8IGJ7fQPhUU9dHCByJqvX+Jz/K+32lXOvttRQedIj1Bf2dWCt0FwkHi2eo8/Y
5sOgQ90HZEZlFeHXPS5rYet8+rYhyZ9jfRqqxOoyQN51rundANJP2QCU6CaWhIqv
1wLKOheCrOEgpGipTswCmST6T16lkgdEiSS3DXhv+DMqezVSZoD6hp0s1of0H5Mu
Tkp7S5cLgWDc0jS2HjValNixk2vu0ov45eoHvARXeVSLT/SDUsr2+RxX2yOWP0ai
HrVqRpHVdDzCMLntC/9wXOBbHiE1YZgOFGjmquFi3lebNg7sfRkjo65YeL6WORYl
e/wyOPlpVPdv+SX5SOcxrznz1iq8u9UyqB6ebgqD1SGe9wQPb+7HR/yG7sxsapbh
5aolLllxQisx2gdEnZquOlg/JgM5Sf1hlNMpVNlYQUtkoppspM8biHiCpw5+15iz
daftzzV3tBzR/tXCn45YO/5jFIZRHJIRxWfojsr6+AaQyYcNMCn6qs5J7j8eduP5
LdREOR+3hOoMR+y/KgEsROpgfcUdru8q/JRit5yTxSuTTp75Dc+ij2SDsUVPGg/B
/Ih4c5C4Pb/S9wUkRq+vKcyPtpzDCkByu7qJFbV8DgVXgB3sR6iJJ/U4Jxsi3A2b
ZmdeCBD6aykZVM+g2KKyqx7Q5uvFIB3BJUtHXSIlU460HOgMSFa5b7zHp/7q/jfy
4tYHXG+8jc3AjHBbGTWf4tPgwhwE4mP/ktNTsDtzzPL+w7G9Yld5quZuglsXjecT
Eu2FDla/DRIBimCsSC1nf68L/WkF/Tzp1uC7kbtCmf9hPzkheWQgZWpmkTucSG9z
8SAJdo6F4jTY7LrwWjfxt41kUJs1mHQie8KfSuOySnMoIvpDZ1JRS+oyUJlM9NeC
CWr7hByOWQ4LGVLDgnNegnaMnPq4+CuB2RM5jvAEy/kBqcV/p8eFXQFN2vgYoEMK
14zFuo5Bv///aP6txr0udnvOZTxPo0Ro74HiTXeFwHGNcpXXslg7TLoRu4E88JVv
zVblV80VCPneGzVl0xhWLxELc5i1HbcRHaHz42WBYvZmhp+lKJoqJ9e2vC4S2wo7
DEGT6npjr2Nwj5fK+VEWQWHmjNqpdldPNEWBf2uL4jzFMk/V/zETE7ls5TusCeXP
mBtZXbjO7Yqqjbt8pqmCIUTh1lSNwXmvUIB5D6zOS6niuzyMIRHGq+IBttkLQd4F
/6+V1NIzLBHct40oSRM5s5HML115suRKqVC1WS4LtIEC5Z2Tht8MFi4FkDMj9hXA
h/YQfw2XIzfPDcKBxm/gGA7dQrbvvl5j/jCHExelbBIbBPlgVwpoUvFxVaUHIRv3
jUBHBCBLGxFs7lbTsdmY48Q32Y1yPieMbPqgCVpnQG2I3qCfAynQlWfIFhsDPLgN
oR0pZ7FVt7Pkn5A4Ai5WsD6nl7DeiMWAIpovh0V+e7hoSW81A3xITdAseJEMfDeB
0dB4e/63lVz+eU88HLH7gUyI692i4f+A6NksKCWLrTaZSrvwbzwhoBHj49nYxmvE
DmIi61nOynPLA3ekCo/NiscAjZL+Tdpp6B7C3My3x/8YC6t4k/LJCbjPkXdJOVIc
7e8zwAbF6cwKF5jaKaHvrpT73FYZPJyhSFCuQjU/+ph2MmLEmGubgr3FSUA0f2f0
T53GfIc5y1IWwObGrRBwecLxRvGw99A76vZbfjxmXRP75YeIeSooRTqyFHCHq1ol
Q+zFZ+EJaU1tBDm0EaN2k2hMaxGczS5OV2oiKwOLA1IaYyxQG5iqaJoJLr3PUgR7
llOyGqIE/nACtQbtlZxhMYoeZmOcL49L3ZLjz8Fw+MtWObPDekj8T5x5GMqD/nl4
/9/PBLRgsSadViJEF0/jTLxx8SW01p05/7MHuRBBZ4FGMkB8yw/5jJd4p5YX9Yvm
APzz2s+cTJB1Aktm0QfcgiAi3tLhh3nDWHTTdsjPqi9bJ8y9QMxTXBdpjSoUK9Nq
xB9sJSD8UpjgCzJWawY9sDeoKJVap/ic8D3hoQqoXR7Y6Mhrw138QrHQ5jpqKBSN
`protect end_protected
