-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
--pragma protect begin_protected
--pragma protect encrypt_agent="NCPROTECT"
--pragma protect encrypt_agent_info="Encrypted using API"
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
--pragma protect key_method=RSA
--pragma protect key_block
D52vWY4O7jZXEZxvFBOoByAP6vo+ku4RZLNDw16+BzNqdsOgOcRivk24UnqModPU
07D2Cuc2r9koTz5HTx+CVj8bDlfcvf5Y10/iuAD2ktlYcODUNU0EthNK+AWQ6TTh
2mLbalzMTG8vvwLDIOyC0I+jfpHsPigSW2rMHggJ5kCriCx/WOpAF9eOQ+yzjv7b
GPkdzXDqku1HT2ig8ATNziCEQfhUVtAcAoLS7z6wbaJf4nY1pOtHzZO6WcY9Q56T
SKRIPlgsVu2vt1v/n41H6bVhgpslOXq+80chvRA3YgYRq+YE0zCMYtsQ1D5hVuJS
ZhW2MeWofg042BH4dN/c5Q==
--pragma protect end_key_block
--pragma protect digest_block
ao+B0RIdis5la2XM28ijx7eQQ2A=
--pragma protect end_digest_block
--pragma protect data_block
QMP5l++3WHH1cMqpFPdUTjk8vAcMyPPM0JQmH48EgK+qM/FDaMdOLjzMadEdyUH4
wxlqjPJTB0e6lqLuzJj8m2/14xKkGoZp1Y/c/mYeswt4C+s3MoHHuA5Upz0XeMk7
jT27cvNw4KBwEvC/Baz1HLjbDIp2rHnxP8w5aUhyOyU9ZNioL5CQif2OjGdOcWcp
2dtA1t1jqb+fYW7SBnKKuUxhdZk2rmM66XpUjOqH5mt41jsNhZL2htzgo+NOYFon
7b7dPq40jXYKddVd8PlsKha/+seM/1tT/8KhhQlBgcu3abI9JGK+aDwkN5Ev/j2M
m8vFrx7LeEPmpB27b/d1bBEi77ms/KUvKJtaZzcUwIQOsq2etdAIhiC6+bBcbD+L
1AN8k0X9YAIlUmuW7MDcskmQUFQpuRhkaHmh17GV4mdGkJpe0sAGmcrSPTDW3YJc
oHymNLkmS0EH+BXMOByYDmDPuMmAMrg4upLfeI9acSfqpPpTWpk2yFLg7l8suAJ9
AyMq1eRnYTHl0HeUSG1VkAmHl4ceBQs4fcJksyPQGvosv5HSJkCost7EA3r4lUFM
JrpVPzV0FNJXHMflafuwagjBezW0Eanm1+UiRZJI1l5wXY3rF1UmPyc+FbRgyfrT
3WkSux1c9KuqXw09gAkFZ6GcdbxWA6AkggyrY2AtPZfTB25T2j0dxzdlLDh58Zna
UHSF3a3pWH3ciLIlqRvX269lm+4OneoPPjaeApxzAsmMBWiAz+Ht9rKVVnChTv0X
+krwneTPP5XCIpetWSBViGRRjqNeC0roBsXOs5pz6GllY5MTFQg/18jFYzpf2LLi
STsfrzBvn0kkMdbhpsqigh/pPmH+IRC2eHPJ8jelJkCJDIVQbAPDwoVNxe/NsK7j
GhAexhMoP6FNH1XGgFizB9pFDAJMK3YTW06XQVwXGJoTTrhN4cc6YJ3LpnG7TrPu
hCNT13VrdK4VOHB7SfeW1GJ9FZH43vfgYuIUI3RCNrcd+tplsv2v3kFnwnYL1bhh
p6ekl+9YIapExv7ar5GkmiS2BKhy8FSHiBg1VgcoaAJm/GUXMJAMPdUVAqyralLk
LMNv5JmU9iNQvSroisXuQkqb0CuPVLQbSRuEPZ6NiSFWW0ivZoyb9bIVHoMb7UTj
LWpbT9zkxORbNL8bCOBZu3nVrs58zthgZRy/gBwwLuAGG1j5dwnmicg4JyjD15xd
SwgbAcOcMgYPbx2L2vaS/XDm22xxjAzxSk1tBWxJylfG4g2J+am3MrRwuvGKvzDH
xY/V4K163uxQyBvx7BnoCnFlLQOUkCrrnwLEjGR4rPwRrGC5BShesfiS0lj/gq59
d8LWeQqIVX2oanFzzPQ1yvaH8rDP1W7bxUcnX4MK8honGbm/EkPzb0C45lFvkkzN
bhpYP/1jluaYxx80xPTM1q5/RV9FH139dPBHXViYd6ss0RvEkTpG6lMwiLYyGF9u
Z3QltnLq87ddDFjEXERpkTLYJG0lwyG7VXpvBJ1ISxVB6HG123HY5chkrNGMLhHu
WdNa4EToAsHExJAGXWDl0rNXalJ45reCQisUHfwJf4dXBIkMVXsl9QDjnSRQmQ6p
Rl2QYQPdD1mdSob0saHj+MBGxHg/edc1Wd6hetARgszMYuz9rcxmkbYUnKhP0eZa
1Va4qs4STHk5PKdJrrOuCjKLUwSdMx5LMILgiqU1L8KJG+MuZEETlIBUic9X32rk
YKdOREUWlWmkm4PrMoa0ypVdj/UnaZHoscjChSsQm23g27DdOdLT4LbDafD1rbB2
QjmJOhhPaMh/psNJg1k0Wt4mjQHmgW5KxmXVJ3oGst6WHYYJvk63Aq5QJuMw8zZJ
KfW8UHxuA9sHTuZZlCojdxcYdIozFNEQXc6cuu0vpzWE2ER1rzu/yz3usLA0F9Uv
Qo9UUmdqeztvbhkuwApbSS6TEpbJzQx0EJ/+syecOITN0TIfYlArbT9e1SbbDzMs
Gb530Z/yempQhbUqcJOOP8qSpJ5OkaUlrg/ttuqZ7bAvymIs6cZuhDpVm91pprk6
/RzbqsYG4fSqbnlIrP/uqBRIhPl7HtkIf0aj61Zy2ZYvrzpfHHmdScmZAcpMAMe+
pm4hVc2x+hVYVgakZBuEY16/SOilGHb0RjwJjyhmuRqr5PH033mkwqD4+mHi7SMl
inl+r7i+Xzj5TpyH4UQIVIBksnYrWUf8otGdlhmN7D4GGi4EFawarSIXbsuiK4fU
7fgYh48/hENI3KXlZaJX5HtdJJ5ZU/6IfzRo4YjC6IBfsm9disu4Wuelpmggaceg
Tn73VqP8bg8mJ8tO42ynwv/kmdRZ7423Ap5GRB7qXw5qJ7ArtzzdcqOWTNIegGNg
1SoiLVTQcrk08Jc/RyXuGavJYyfqI2ezzq0GeLQphNo2ZRSYbsyDW0QRlqIEUzXy
QRXX1xzuypbsDuoDrC3bp7nukKPI5mCl9+2LDeUYRHvPOhwrVxAMh+DC5/tghVf9
yr3OxilXrLgmXg7MIEnswxMZVGcdodLtmt2i4fDOp8y8OZUxD/7mwBvTx9CUfAQ3
aO2rKLZe4KDYXUPTLTOY8IdFQIqmPC6HlCkFc/Y/FYyXl3MjXBA1DOlNfTlEmx4T
yTC4IIGXNSmQkEgxnGVC9ejEKHStY/MoQma4KgzREEqL7/QIPiqqZnrjO2kXSvT+
bekz5KeXYxsRjmVdMpG7q0y9PVAPF1JrBkMVO0BF3TUaNf1NHntMzSg8J58scT8s
f+ZnH2Ny2zVmIVYEHBfed8hJLudZFUZEKU2Hz7xM/XrYycINUWWZDSbLhkHMUaYp
Ps2AittlPpLlgaM2D1TdAnlbYm04pwzIM08mnZp0KDCrCyo2mvx8F1QaDpu8GvXR
+NXRR9Nz+511wgaSge6wwXTk28GeHEVfiocjrat3LvqjI94lJIrHBFzeAedHhjzV
lgd18wg6/2PnTAOLCugFBxOUdqlbZuYsDHjbQi4sn35ukneLZp3gc2v8WefJGzVG
x6xflFRaxjYJY1BoEx/l38o11rRiPPH54f+BdnEbkXX3NCBw9w+cwJUpo1lu4Rdl
ic9M/ocOr99/5sRRjYhe75GU1IxBpWY6bbTMYk+cT0FKWtLMYeI8anX/pqyqsNVp
vvywB2iC0UdWSbI1zRPfHVIBrcUK4gVEATQwclCZPSDOoDi7cc5icoKQgSHLRgMs
azDPe/0jOkY0u2NBdHfnMWyOsuTz5g4F8YveVCD282mIJ6BxUigUbkhiHlX2rmny
3gd+IkNw0KI965uVNX3GvDrmCRlxhbKiMr2TBipO7eIiQbYzvi5d3hxjahSHr2EB
ipAVSmYm3bOQaSrTgaLjaPD7lJ2ojeBfducSbdcmBtJp/AkqESfwdZ6WAkglmea0
52FWxQUcGILa3eSlpO+pHdW1x7d472z/ktvQeoLA7Z6tbp6PT+n9OpBfeNWbEezX
p0yTn4sHRfG9arYWhuI4THL4Qv5Rj9+EOo2LEaU/wvxLUpQsP8Z4DUZ2BgWVn9NL
GBcvKZ5gD+yqoHLhABmBh5J+FPLFOx/fH04v2RtH+NaMlTu/NyyNP0Ko+gD7doLM
a5YgddeW6ejP334wR68lxozJMh3XqD+mHh3B1eB0JCxS7PTAkXr/4XJ/126goq1m
uKudeMA6/nZasSUI49xDBFeT1ts3xNUd3zxRc1aoaoE2iBOYs6+cHLMtaJ/rLANm
CPP1V8+Nn+uX7OEP8mEcTZ1cUjJGuQwqywxChi8cwo3yW14JcgHtdd/6nhjK1CdI
eFMdsYCW3bhXeZnxzHEcOCLYOQRKU0ZrXxOrfAVJgTiE+R15okZDCdE3hQrXgahv
7X3Ac2z6wfmHzkTiDnVr4cIhL5s2QZa8nUclMvjOi4Wb/q00O0j0Zdn27O63aErP
TYFFKcH7M+2Viahyx+sK2mJ2UmwuTsu2/C7ghvfFDlEryiyNBW/hdgi6O0PseNZd
UmaOVv4079iFs1k2HYtWi3EU4CTo5JEE9Nzws20v/xGAmInmRFDir4laO71NOSEt
Qic/hS8ovC91n8YbLX2I6e4/LAwERPMjEj5OliF1ZG0C8lnCuflagSm96V3te7qZ
PDH33Kw7qO17TLImA45EhRZDUuMuZ1MIFbhP5NKmcyHVfr8+bDIMJHm0KsRVwGe9
X8vvpxqz9Y/NwuA1kqVjpM7RMzokDwsDygeFgIni8av6sjzyQuyynMUOFhh56y/7
0XcEZvp2A6E6xDIU9Wh7NBYD4Mb/MYD32T90+Ed6PFL1Or2+xkLGB3S4MMscAGc4
l2yhDDm0oNYXhqTlIUIPAyvlQ/GS+4Xz4eRCWg8dPHBHobBSoTnU8xCFFX8YcRBf
5wtgLMhP+IJtgfopKvS/YhZwqNpbU3HJurUA/9G6E2jqqFxSGBNe7RdrzQhncpoM
b+XHSiv7vCO5R9pMtVUqLmtEwT65cXndgzJu7T5S4ZBzjPpIeL/ijUY73kiVssDU
hNuoOXGLwtNxQi/AGAxCRREa5hmvy5eLHGAbJgJzwzv/M5+hTkbf4HAVNn4DAsxO
jc9xdzIK12TKI2IU5XFNkF+31z0BzqBHkP4X27Fyp+RpAPJ4Z7KBC5r3gbDfLKnT
CJy05Na4e7GrnhFX3lwrP5RAYndjxVYda8aqIjig9CcnCDx9CuNej+dVvwnHQ+ki
sGnxPYxT/dO0UKX07rI/wm3nrmlpCnv3r83yp8tmzPl2CJYRBfWGVxOIXG7obnxD
Tmur+YM7EbJOGlrFgu7gF37WesCKC8eqJDr2VLYtF1FksvWDQZoN3r5qGBFIRI4c
7phN/UaGGhVtkGE3yy6aYgJvICxUJteEWTcTVqgOWuwC6sGR+WhxTjijYLC43Ekc
F15iQE2adnZThTibfyRkmaDkDyAkmMQZ1/FOmWtofZOmv8/341p2RX9vnUKWrCaS
0AXrXiIpzsr4ETCzWydYRC7t9WpH9mSAyrx8I+/dFxH+XGANyKdAQnOjgue8ndVg
KJgCE+sHlu6engPcI+cFY+pfriy3AOhQbhFerkF2ii7Lbo7Z6G5OGg1GCUqSiiHi
rJAT1H9YsphOmVpchpf/Nl33uPihSaqhUaCem31EgslDkc9jYtM82Pwgjk94nP5h
BbxeN5JXNVd46PYt9eiZx5R8z3kqGO/XlsxjBwcry9LPaBCbh/bT4Am8eLwHfRO4
uLidFPGfU5IqCpeBntctFkbGICUVr9if8351risUakHHf0J1zsjoJAe1Od6/iDy+
ad5Fqm1wJYeswqrcvrE6Uppjx1dE+4e6Cm7h+NV1XVC0Nonk+dAPlqgaNkyawr7X
yuedTLdGrVZr7kBIUhvofbxQpKpyWH2NlbvWuz/x+MwB52wUWUIPYnAoBcgEq2LQ
EDjsMMyGs9v+p/1K4TgSIV8FKhCbB+CONwSZ73Wcx4JBgdyWViE4QnAGt1Wi8rQT
3a499idCKl2niEKdmDsmxR2IEzgCczumAgYzPpyW0yZbsEgV8W0l2O+eLcImd+TB
iQpqiEiSvoQjUR/2FJ0jXkjEN9iWPnwPqNvqy72NI/S+L19t08q/68bD4WjfKfOG
WD5p0WSqMLPC14n5LOHOj0f01YklUHQ9yCxV8OptHaeTSbMd8Qu96FCg8Zi2Swt3
uzElvFrGLvsIxmj8GJqUtlbJyKWyKwVBV+IuskJ/azAUM+6AcyF4NmLnLT84vu6w
DmzdhOvSlb4GVpVifHgjtO5bO6WGc9yIjCE8TvQcg3QhuWdka4e2ZCZR8oNF92kX
O0uI8Qi0hIMBG9euOoN5IeSHG54r4qkso2gqc1eGf2wCNIwDLKx2DBg9CWrVsaOQ
xgOpCNvenLc7OBSU1WYxxJub7qDkbKn4ogWnpGmPT7EdhbJ+3aM08GAOBK6Z51QK
--pragma protect end_data_block
--pragma protect digest_block
b9N5eHvWmXf75BTjkHz4HSz8dKw=
--pragma protect end_digest_block
--pragma protect end_protected
