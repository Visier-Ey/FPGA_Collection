-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
TA2U8QKHoBSv5q3gbGzePsZql1Z/KuXfacYNnjxxhlnmZYjLUO8UJsYDKrxRpp/iEMob2Y/rO9/Q
CVBFBNKyVaOFpUixGOCfV05Eqb55DHJaPq8adVPySssuOW2tF5WX7Pffqn+bXxONxHvcYQXL2xbd
35HLRRczXSCnNyZBvYKi+lx9n9Vn7BfZDya2gVL8zepwnWXd8G04neDFSUCmTXQd5IaGX7Ap3ujg
y4MmEHlu2xZbuuYaUP/VYYInlmyr8WlIrds720qA1WBTKXaLBjtisGEFQrobPc2tPwsVOu04q50N
ulvF2W6J4puXe+vu+tUhXWBqKNEJbtkSqlAvTA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 111872)
`protect data_block
CG3l9XExiAYoWjz01ZrLC61YIhsDIlF2ND0r2p091M0vQmIIFGGjGvkGFL6LUi2aFojFdsIdn34z
VjOV1dY5QC9usKycayWbMoyylVAfxYrA6uPg4N/odMM6DYCsApBl3/NCkAoE5ctJOq3KuggSugMo
wztUXNoubG8IQwksrx6DKujkOsjxJtbNW7V3B92iiHpgoraLYGXs0JNR7RDYBEKQeK+xswrkRsqx
N4TgFXPS8hnqbOZIRkbQD7iZaA1+usnKwOVFDwQzLbnYXZ0dY3Av9M/qZGZ0SmjWRu9EgyAsLmNX
wg5Y6FSWT2BrwUVh//Tgf94v8FUROvQSUJNRZl2Xg1sYIp6j4Y4J0LaJZLurCKLsLr/sbmCbuTwP
ZZTKm/pSJQYDhBzDI23YapwtRpau3MacTkmaaPXpwuMafAFdRe74GrPLG7i6wb8t69UUu75FVaL4
7v53EjjCmQDO5u+oDMUhUJEviRSCAjo1MbkuA/EkTVTKNfzLPfMYLQQhlm9d9qKjxfg9WvouO/NT
woD6bdLDsvKvJbaeoMWSBcaGJ1CcVBvBJzLAcil/6rCe5nq1C+6JoQ1xdJ+Gj6FxkzYWzy8J4M7k
aHCHAJHzWRtTRWTLaara0ylRxItD9U0G0h4s2WBqO/FYJKEjBLhbu1EpZJjUgv1D71oyZPS3E7Mk
fVQIG7HoMOEFem3movPUtadelQM14KIT7c3wVH+tcncG1YfV4up6bLSSkSF98OL+wRCETg8sDSLw
Hj+3Q7Q6JfZqiobnLTK3rZ+lbHCiSrFQJgewo7XHdwv1uOLTs4mkxtVTW6aNZPY9r1uVOsN3qfK7
CqjjFuDKt3QktODbUorQM076wQJwZsntsPuyAnNXw8f2aQLm7gn4L44V7xyRzI6c8aLmxzs9VeWE
/i5nY46JTK1Jk4P16gHQYhWADEfRkN1r2OkcwKD/L62gb/KoivdSnHLxbBkeS9SPCo/3zn857dlS
tBmAju9f8jD5HkUEC0vfaWrTctuGgv1qCR9XeSOHhW19PncN0QJOMMAn80p73D6RfKOzs/qLTz2D
lfa/FSDAA9kIdu6iYiY+aY0yd72Ocb6kWpzRb40nf2G1gU40zrlTRiGmdkNHl2gRvSAbjwJagpUT
FoWHkcMgiCjkApyuJT9r86I1JWKtRMF70m1J7ugg7CrHuHrbEpEZyPyHj9eSgY2E6aNN0mzHAbkV
48e62ZmH+oT+hfYHyKpCqofwqionRBjCgZVCfK5u6jgAY0Hp7fMEM/Cjj+MWc0jE+v2tlO+bKkIy
CXYI+qBA5A7xk52TaVh/hZr9CWqxvYToqKT9JKEQNcDKSyQWptOYms9mZonbr1wCohmF0kZwRx04
/UbjNKTNon7h6Jz92Xo0XrtjZsHOjg5RnIZL90GUTfhv1Al9HeQo7fHX7xDLahoCNyKWjwmYHWMn
L6lwbUw8lOflhGL7MvLcOIVlT0x0lLY2r3BYVS5h3AynH1bZX+pG7oFAmKSxjX0AA7sZAQtx2RUU
v+sWoD7hYY4ij/pKq/2tuylPBXASENNniD529MbOLYWE+jkKH8G/as2cHpaEUpyIH5uEDncoSgFz
p6k2M0bPJuqXenPVKJwqe7oVrFlpGOEXmmZMYrmx0Gy52Eqryr505I30FX4vuagtfIZtgBaLx3kK
X8H/f1kPI8hsCKar+U2Zzj2C1Q5FxxkUQ12YDYudIrwETEeKi0V3oETM0q671uXkCdqtq8k/cF0G
KVA2RbSC4xjQQ7J8JqBJP3prE7GUp1Kzg6+mOpODDvZqacjgbcYB3ZEycitdLl9GXx2DfDJVMs2Y
5cXIbo1dV1Er2TuFphb9K7kAtzLCtRZAm96sQRFF6oII8ySVbRsWEdRJ8ejxh7V8J70yygXrkuG6
IQkeL2aQzqwk7mUyELxlVGQ+nsicwrQHhQqxSs0Y2iQRvzzNiLLEgDXy+E+YABiw0/78FM33z/C6
n6ctfTG/PcgiRdlrwV9YGXJ4UZ/r/3Tlvf1n0PMK9rmnAgdxG9v2iciIAc9hVgx+a3VilY/2bXGf
oJ4Lzus7RWUZX9drU7OzFFnUn96I8ySgFUv1ivB/KhyD1sPpRrPcPZ5r7Uhaug7MSYnJ8FiHuv70
yqkLw5ou+8/WCrsEZVQCvZz0bTytpeHx7SXhi7yzVicNg4cvBrWVWjvTd004dj3pqoREPOZ9NbTN
QWIM5o86oV8rJwGNGYbxDQ8Zu5Cw/Lh+i6Xxa5THnO1TScbYxCj5lfGfitFW2OIG7iZpzd+ltB8z
NX555RwIuA4gRMhs6bmhVdHD1NmbyXIiOm40GtJNQ4JI8KUwT0M7HZXGpdW1vh8DbRSXerpgXGKq
nyXyk9O1gRqryiwNO0Kzw/4g/enl+YWHXBg3f9hYjH5ldqhMZ+P4ulxlzX3BrdHvCVsKi09BJA5z
lfzg42gnCGGO0uK+ebylzJqi20e0hYD1i6wmXSRQ69IFREvIpc2nA17MCmeY15K7+cf4sKIY/zuf
8A1VwYDpqhCEcgNudcmKNQVFIzIcUIKA7jFotU2PnibCO+wTz37VZNMd8eGpMBzp/34buOJ9w/sD
J0npYjy4WPbWM3eUSNtS5RHF241Yg4f/XF4nqwWK9tFJKfrt6/1AkpggdHp1btJIAQYYhZqlH8nC
noAF8diTExgNiDaDF1y922iyd5UzxYOrGCxwE59mZVbCwF8+IRId1HZLQI5Adtv+J0QjKh14qkcP
WAnql9MAh71yKQACoMu54oRrUetJQQKr0bxHtub9Nr3cl4oP2HdAuBcbQJ5axqWhFu2yOsdwvfes
YCIedDWIeGQHvOMWW+oo3o+IlOekWjPnTH7x9hH3BLjq/v7WbGX6iDZu5jbgHhYF3mgf2QPeBxRX
/CuAwESXVF7x7973w5nyCBm46+dnbUawRuVf2YXnYNVI07vftN5OcBmXUF1KxHsqrz7RPMX4Q4Uz
Ubtl3ObFQROBD+W28r8tQZ825qYXDrtUc5Z6MuPtYObmP9trsx2lK9kEUhYEaO6VaqcLwvN0Vu4s
NmXuhu5Ghzuamw61SEIqqFO0V5RZO9lbSmpgodEXAhFWSLJk14zp23iTGGvO09C9NO09ALnBWuXz
pOSJPpcwgzCjYW7qgOX4zakq/8qmr9yr9hNKvjsUsTqTK+tKGi1IrJJFd4Bd9fGkjJNE4kTdY9ba
es0QH3uC7ynudld1u2vaWtss/1qt4qi8aKEwTyxwsPuq20UsWNhmu3jWZgK3VQ3shTrkG/SR2VH0
XMoin/KIsq0LAIcbIKABkiPMwPPSLs0yrA5o1aE5n0SjIWrSWIKSyy546wAjgpT2NpWI8UjWvqDo
z0FByBJoZUCbiplDl1vHM9GsM6BITcZS2fLV6jWa0Rvi0EZSYwhCr9u/1au3LVhryclfi2538EIm
zVwN0QE+OPG7EgbsadVef+GA/6Y1fkaNyZhYvth57q4bjZmq6XUgytU5UfWb5gFY+C+AIQ7Q1UCj
yHXD3fqQfX0vmpTGwjO5VCfY2BLAyJgtCumNBNdcg1Xp6xZ8orf0KdiYfJiPsBL3hEU3ZikWkjwX
CJlAM2gdHsTYscgPscWRggJiWuGN/rMPYQ4G98MS/VwwP2xoCySZkkrUcM8uBfQcBHZYDQgf5+zO
BZvq3AR7v4ABGBvnPz0H8QlWJ9300yP7Jt58NLJEHYjlQ2AYni6/CZ4cK8gwVDtX/pBgSJ/p0diR
kg/eTOXHJrUvc/tmWcyHIfIL4/wi6MsiiAOO/YJOrt8qpznCEdtvDx3wVUzmbEUf2EyDATrH5JXV
XO4sNkBrqpaHkJOUGVw8fIdzofj3E73BIVuSsSFdKGiQM79OLbBVF3lxiaPaR8cdKOaqAqdt0uK4
y5CNoua23CI4KIpzV2O5llDqQMTGETAsFMHP9TLipRsL4mfuOcZaEGZvF3bjJCJtlA1B+EJBWjLA
ayEb4tr/u5XSpSCGmlKqMC+HVHMFgTK0zwqZxYl5gXW1+VHLl1YGhizp6Zs7+TXGuNFu66o/KNPf
uMIAAjUNpVsoEKOXZ+Wn3qGoatcIUTuamGfcUZqeAFW8yW2la3kBvblUdGDocmz+nZxo3i3nv983
YGVjBO38V5o6kMn5K/gW3bSFvJrpWkTFYt6kMuv02iy2Yn20E9KwGgTIUuAi2jdjYB4prUjBe+wY
mbv7jcE1DyqryI5khnHVzN1CHH1b/5dcY6qSnHjj2G7o1WpFVQt9WUTgnrh5iHBYjAAu0fZnfKvG
81DH6dDPlqxyG5BxkBJV9iDVGQXfIJNrZrF/U/0zQT71XbvV1VjTW2E22kbIkm/taSyqLhsmIaL4
D5ZuDPQOIIY6QJOtjakRGBMNVNR4Dp1i0t0R+yXMEydJDNvy1cBnLjNA2mRv1iIDT1rApunaZrhN
qRbCc/jkBlF0uD1crTKKacRE3Z67e2L/PMO/MwXylRVYw9Ddw1Hpm38+w0xGZUyJA2DGdbJ8YUc8
ityTMdyNoxop+BO2smxe5vlMTggkBy306ouGl8Alb0CMsst0fe3V5yNMj4+J56bgf8B6vhhS5hrQ
IvaOOzYI0TY3oSD23ARVQz0YwC7T4dx5iYEogiry4FeI087AF2coalTUy8rzkG2LxteU8cAxM8Zw
4+j+VJsSXesFAH6gfFvA2b7NnXGhH0QnIh6X/J16uG1x3QN41QUOz3xN+DCRCYevW6c6hu85EKuU
Ud6BAwWOTv6ze1xRqykPTJNXOUwFsEpuSpeiflRqv4v2l5G8j+YeOOxkkwMjOC6lSs2s+kguzwdz
e8dSU0dfI3LKI2qaTF2dGHxpmRDuCIO4DrRrE3UWJQB3MWe3CligRAQzLBKSbJE8EV9y07lEJNO5
mqTh+Hm04SF2vu4lS1cx/nbLG3ZZLNO0fdTLbteBha8j+v0SEBWHvcEAQ/m8OEFL9Kg6V3neDBod
0hnvZX19e6y9/r64YUAWiEJlZ8LwoyHZqEQfZdoU42ActFGtK+TSTe1oWtNt13rg4Pu6IkpRtw86
NhO0yoiRFoS75L014Zp6MptYhp4jwLpvmxI4KBrwKCtSW95CWpc2Pg4MtWjj0bdkIAPfCuuDSf8k
XiOQloqSjzmYmxmCpWvuh7gdZnlnEgzKlEZN5t8/gQoe6sh6G9Dklqy34+HxSTqalk30LXWfTHlM
hPr26TxNOvqry31xygDny1x1ANmYXpNJQU2QS4wV1akogXB4pHDWiMnNxOIHgK8W8Yi6cSqYAl7r
8YU7JVv1lBLABpw6M5zauCKyI+gzh/uhxDtpn61vP64vYYKdiDnPBLBLytvzmSowjzC5ujo6QtNr
sP9N4kQefGOOn49BjW4KnTLFSoCW/Bx+FvGcOyU60K9aE5JmHk3Ldnzrqbhecmk7F+kGi4U8zTqD
1WnsBXmZZsknqh8r109JIqLmMOqqCbhgjhtfI0AsoYLpx1yAD3QkwJ31sbKCp3al29IgzmBynb7F
Qk+sAEogOWICnf7FKT5MJhHL2ibcWuCDWRicK/tQgNCfL0DeMLL4ji5ICgy00t4aj5KvcYOzHcg8
GZkQ1bl3ZWZ6Accb2A1/AFOSoIlc4NbPfIrg19CubHDF+MnPvz6uwNkCo7KKEEslbPFleJhXowjw
jIZu4ujNoSHqEVEWKNIAHegyxA0nrp6uIVSShw1ltb1bAlKk+eDZp6tuT9rBT4E0IRVQKw6eRqrE
g4d/u8nXMzSAHVD7/RM0WWGNMdnRcV3cNF8j0Y+It4p+1jxsesGTIszQcZtLP1VX4SM4vTNTVLtk
anP6pWRa61NAjE7CIg87i1emOm+RSlXSTPf6XM1pFLpa9W4wD9+LHyj5cOrT9d6hs2cY5yaqjLFq
H8s6ZHss3BqOo5G+a0KSQLGBH6g8qAshGfK3PyURXbXn4EtbH/bESg+cadGqPAn3bQtm7lR7jWl4
h/pxro+faDL6ooyTn92izNwT8wil+WvdzaAWGqjqoU7iWElfHBzbyMLjBkAoeFldWQzCBHX7vJsL
PfMGx4HXVltMHKZkuv+KQNulsMqssGsJ/fxQrmM3I+3fexriwUNxXhVzVE+94Ab6nzbGRb7w0DX8
Ok9F4CKrV6kz9B7uyM8L4hki6Q7dVz4vdJr1CHJUA9UMUyNyBlSTkbkZod9UL2eiCMUrD4e/0gUR
ZzFTRlSDtdrbUI/Q76kFsXvxn4HNngAjrii4tXUuSbB9LR+H2A1eWnR4JBotwtYcR7wxaT3sqka3
P63dR/ez84ayo/Aws594rbqWD8A+Nlq0jo9tZxlRxQy00tmnGHjSJNJbQu2wpet9Pm9UhJv0B67c
1oxb73zy9sNE8RDHZ0K+oceAcZy+OqVod1bJ9MIcUZurqvJYwth4EKmDsXuT14F1iVDNQR898wyT
5eRWY5DD9ruNfrkLNhiSzp9D4MC4ieGKNRYgZbrM3+szBW7vKEHAX7ZIn8cPRBi3WvW+mVKJJk98
b5jTtv7HeUJmPcc+f06Ngn3oTI0R2u41c3g7ohbd3+MzIT/2EQ4YhSeBarauEvLy7fHBk0UXpNXU
z2RMLkuwchqn+j4s2L6ouSGMvaKrozijS08AQHzAT/q0oeJR0X+eGACTz8DiT3zkX9afJut2wg26
fH0WpQL5J9pkbzMitRc0XKUDYit50i+teGYL48w3ucN+lkqNs58f3xWwDYzcdP9kvmG1nYqIalEx
uugk6m1E9ic5GnB9/BprzE0Eh9ngejyDLcp/DWtnyTvSRYDq+LOoCmqf52hQKWpw+YQ/iLqOEvsi
xgGzUMJZ5tDHxh9d8lULW844tJfgBlA4WCvD0bnsl104PEvn0ekPTlrb4+XTlRlgHy6UUH128hxc
iC2VteYjdSQaFM5OHjwuLCCefA86nIVuknXL3zI6zySIwlvh9W7owLEW4RrpH+OmFE9E0zmtOzml
iWhowO+n2nz0YirC7vHF7sBCfANNaBWS308HmH+iOWKFmMru4b0X/XhyCMbHzVd7sS+HuNPQrXXj
IfcG0ent3ZP+sLC75u08SsGjLv1/nufvcgNNU6lAZOn2hB3aKUdjTuuBsEOJP7G9orSxk9Ybvr3R
6oFbXRjNarZaEg4d/pEt+35+7w136LQ0O5Nxrez10dHdhssmeBd/4PidtG/GwSFrd59ghR6oCs2n
JV5Nhnx01hASzsHMezY7EaNaj86aRZ98Mkj/iXIrAyTQI33QwajLKUM5rj9oDquYy76rTYP2eSry
OosUhG7KgmJQU11XFtTNJKaHKTsk15TplJ6+T9v2Pk7cLKFnw8fQgyGN0MHpVrS98Dj/arsXt0Qh
ZDBqYkyKSlFI1gZKtuR4o2jsT6qlWtSzXwy7jK68vp5xWJrIh4Jb51CRhJHh2eYSdxFi9R+vOs5L
8AvQC5IS+PvnTqxgEu6zdk4lSt8mbn7xniPtR1ef8T3poARASautBhyM8fUE0mwg8aadgH0PS8Df
QyOE8RvhWotHvPLvMTNaNXjUVdGRodO2XzC4D1MSO7jwuid+vPxCxgRDDQC6IkC42MFhREfx8o/S
XYqbsJIT/6JmbfE07Ynxqu4iZgtUkrYG5WXQepWhkbyAL6wN/D797QUvUmbGJQ9hvHzKMpLxGrur
AfMj0VySdqIAN30WuyLtqM4D/OQVT7UjfONTiZFm7BlBZR8RzwPXf6hiNKxz6ffVoKX1EHdjuMcy
f8x1Nu+JX0jJhQW/t2/S5VKhK04RczS1suSMgbtHLC9Jd/kI4nqmUNHXBuRZjlDgBdBRW8IWW9ms
2mi1WW3dsYZT9PtjMdS8w2bfq72IYUUE7huC5mRvkIgdSViAfWE/jsQVEmgOGxfifG5R87fpXWbz
W3RExI0EJDVSxULNA/8OWQ9N79OLBs3g4MaVlFHCDshFO4JKYJm3Q2hgsdwNadH+LLEf9ug3ZXou
4DDLzQQMsBZVvQ08AD0di8FLuognBr8ise1znDxVOMBkjcFSq+ec3+d1DUP0rtJygvsLF5RfIpw0
SXKzfCmJhsanXkXr7nu1b3cZtYzBhHwOArMx8B81j+x8BRGzYF8HEWirUpRf1ega2nXIFpxrHLqy
mmrbnFcXD2DDRgQidYsjRLm+wbMYfkUMtFCTCdcdiIMjMztK0A+QKq6V1XANDe1G+U/wxPB3kWAF
2M+Wu6NdY9EgarCFx24h7Q4PIwKescyifx4aj45CmBYLGJB0+QUzf2mjBsOrk0crba+zPNgGj4lT
db+dX5MHDExrKgbodPxeEEEr5z8/5aO2Lv86XAqzidn7GYEZyU3b/MhVvd317N+T6KYxYzSKxLbA
a/EAGIRDBQt8Cj+oRmCFBlzX6aPyN9ltA88gcxENioYGE8Y7rPBMF9F/nEWb5aVeFshtmAE3SGzD
2/T0QLknB89DVNAbQiEJ811qwMFRWuTBWkhIwPbYDxhiEeFN7ScIDk//tvfmSwxC96mUEgRPpXAz
pZxxGxyex1fRo88uu2JVF+QaArIxVQDqzEwTWRsGGV+coW3xY0Iv3rq4RiPJMgDM56PGgUguPvHi
joT/GoHUdOVNeHOXIJv5Hp1TD26xyJp9jyLShlic25OnDRoUXTzEO7+Ii+ZRF/TKG8bGRR2QcnzA
ajkNz4JcgsVHVwGCghPUxxgQ7qNlYLGHqpD78jF2wJjTY2hyYpErUj2c8Q2J9dPPsMhJtQeRwTDo
XVEqUeJW63b+fPYZnjvPr19V7h1I4lqcdqXF0FpFYgjmRh8CbR4DYjCCr6Bnjdlkh8rn1XsWvs3+
nxm79skeMfBJP5fePeJMGkJLU4451o0sFK39EK9lM0lHlCYEMWtyOwoVRPZhq5iOqH27ceZBkvtp
OL9NqrbCa90wVXGr9QiV1GrPVxq1NRS8BID5AHDoQ7E1hrYwqBr7fYcF03T+KZ7bqRracfQSpV8b
shqFV5hgloq8gWcyauJbhcvGPMVnPqD6KsIQ8M6uOJ2kCfiR73Z7cGrvzmrUhguKU8pQ01EIk7NA
Bs4zeQIesG9zkpvd0iyVeHdoF8tX6kyd/MDJJ+4f4nMEntmUhUa6byXoWT2xstBPXcjYBU42moNl
WLjInzNkA46G/l5KA1wBfU9U9dmrdPOCWINVVLBim7KWBy+vTLtrqHHHRCKKDyvSySfxqpgKu36S
pKRI7MIbV7a1ha6P4HXma4os0YWobHcvoO+tKHQNaGpsyCUMa1syBAg/ldJUqLtt77IuBtA4RRRv
j/sitOITrz2hfNiE76OJt6CnyrBian3zBvdxwJ/vSXd+xB/q61Kb1cW0GPsJtG778k/4Ma9gIW7i
jN2qR7E1VHx9KldlTZpNBNR2B6+1N1bJPBJAjW2TXKFAbJzYZr12eRWtDxkvLCZ0VH0nCOQG+T9g
mbeUc27QkeVU/N3kzECgDoslnPVgzhBP9scn+/r/i3/e3pucC0TlJ009LfBG4A2boLBaEMwJCXhO
0HbmUARZhYMBK/j8HcE2Fevx5uuOAYkvUaL/GQ39yTEx4EfsR/YptolK9qceIf+tjxTdYrvz/xHo
PZfHVg5zqupKLcRunZ2ytYCX0RVgn1dSeUeGLAIBSUXyP2mAE5gOwFJ91dvwdc+MQSBw0d2QqY9R
zz0OLiXuo4FYfdMa9KaBXm9YQLckBGKFsqZbeWEIY9QynSMfnrxNsO2g2pQaPtSfb26DNVZrWMgs
sEgvEux9xQWixAK60XbFQ1hQ0KNuGBOEcQd9nfFUYsSM7VTlgfDFH775fEV4PDaoZqKcXe5qv7//
WwRAmCx3eGx2/vWfZi/wksUQj8zA1VbC1ZdKnkXPSLtoDuQeK2AQwxFEme7srYxV9EFnPVgbT/Ej
M0uNqvoWYJn6a+rtBTF/ckcnqmw+1p7TI45uzkYr6ShR+6sZUFt+Edcmj41WP0Tr9qL8p5i8haOi
Mts73UB2wIMAcTSCKJKu18ocavfF0/tZGy3/CkaeGOszg+GT3JUW5xVQ2B94syrY5J8W2MaRWWD/
5xJ97DieqPMPyb2fVpJOxwsDI1RC2Nv7vE3QSl5AY9GiVWw+0GlAx0rGYMeTbgr/9t4ZqlkshNUA
i5JXfzXbv01EdjQYaQTSQz0wXE0kLQhJ93vUL8Yci53WAfDaV64FJZxAocrR8qangbQ+piQ1guv0
M92pml2GEr++ClB2IUxDJTUUINwc+toffM4e56bBXK4nwlYCNI9lYqVI26HdtTo/dNjv+9ykrqp5
rEy3UoVAqKQnez927mLwHlygP2EujTntR80+WMVVj9tTybyxKJDRX+EK9iQye4za94jkYYTsZ7Pu
736ELDsQeyJjYMxhLnJFkVOMvKnnpBxUTD7GSpBEM4Wae4VpKyc0QkXF5lIHhEkrqovmvvmLoqbz
vK/T++634jyOMKv1WbwbY7EJG3BimjT/J1XZkyTTNp0GsPcPfG/vE9QQTde8f+Ylnzq2yVMx8ej1
0Jm3/lTtRqL1OaZrgM/Ccwm6a8ou/rti9RDwqZMFg+SiJT8b0XEFCC3zt10Iu+NZs1dWiW4qPpE9
sKF+uNJBdRG57KzfaBSlsLLFmSpas30StzLTFP/PHjKhBihvWHc86DYSOqDQDbZj9BadIyLDKSUS
iNfxYMzbizvsvOd0uNQqRPeIsRwf7gj0X/qwewbbAE/33ckMVUzPFuz56v5T7PlymLVwkmRcEyxQ
1InOR7pI7p7RpGoFhufllQGsewqRrJm1/YSRjuBiIBGzgDkgAI9nNg0nREPdYJn8er21TyhMbz7B
n4qzKmoNrUhBp78se2ySPShEtuGE3x87rFXlKIhW6Xw3So3ICgCpwSW8jtZQm+wm3CfgtWfc6vRV
ZzioHgfyIAGUTbjFxyH3cUeaixXbemRGDjFHeSeas4tTYAVUDcPKNd5rLnkvGPpWg2IJ7LW9IlYT
UjTAnn9dVenEhS7Xf/8uHiadk6jAiFx04SiyLkTt5hz1mOl9GjxkZ5tvb+rA1R6jQFy9KZ2MFsXd
Qc7vKF+CW0vH1za+bG36RjM1Edj9bOaPlivsEHEGskmojqLxslVt4PU/n0PDok9A6Wf/qlPxl4Pk
UnYXO1kwjhMD3w0QBrgnHKZKGdxkvjF9CLCteVeE5D5JaoILghJTO6n7IqAw4Uwq/R+24799xEby
yKgf0fbTQsnZ477t+yQWCqfA9dfdmeX6pUVbF3LTLPlzFGYt4Ow/RSozmNZAPMAAhZA/zpTt8p+0
DIhrq/ba7DmXxauz1P7uPc4hK2l4FWMzABrM24/g2+AeY/43L9g6LEi9sL6oWJvKd0fvKCa9u29K
mVIelfe5yIq4z4aGbL/Fu0juEuPtVi9mob/ysSMSw7zr3x4DKjVcxmX3AmjkzxUYoyDYQn+sL37U
aUaR9Oh29Jv2MaaYLB6TeOqNi0pTCAIwRGOjazIH+fWpi8F7tDJjNt3eN1p0IvNLwlHWV6bkUVow
yXjRW1xNrzsDuN4jS2d4OiKnQAnOzOZ4w6j1WB5w+I2akwTygNWMGc0lP2IlXEoi0rMpZfmOW5Ek
LILkSQ2IxYKVBqbSxBwiwvmsWVB3iFA4rM+gtG1jtY5jWm58XoFw6FViTxHbf0p0qIb2frYKpxxn
NhUkwmsRwwf2FiSjbT6T9aoZxnAodyLhw/FRcqKzvfHWyro114A5Xc/D7IzsqkkKvKdkKcN5fmyr
Z03Kr/9gWYGK32xffo9cBLqJt9Ce/mwt5V0RezmvceDkZHduwOdVjRG0qJFKP897UPScuXynb24v
WcfsFoLB1vgX7qAgH7KFd0MQMy7VleDXMFPbPd6IAPDxfZk3yeG2FlCGr1QFlS078EatixC8ZLmC
7yRASpHUbIZ7cO5sa9+shOGfkbxO7lfDhn7g+Q7tHSxwPZ9O9isrzWMRuj2PPkBIZl+ok4ALv6Ez
mDALc0/mPDxbnP3rnfWq4FAeACfqwMh4U/w+qP4y8ItF5ktNYrP0VA13UlLORhRQfwQBZGNL1CIx
b+YioN6HVZt5D5+8NwON+221AgAnrRegpYumkY0zU2jtsA0x6RoD9j0CFdiAPqI8jiCjlKW/MWba
8vEGT4bMpOizTzozfzMk2g1puW29nIgEjq1NfwjaM//L88LYxsAU7ch9TRnvLwV+9XI6eq/pT701
7OQArp2FMuZo23QxSh6jItKX2Tz6hxNhWLd77l6CsuYuw8QHm96kNf29zp0Ro3wlTMc5DBCxVLoQ
8RLaKdbRU4ByEARI5CDz8w5Wau50n3ZUxxSC8yXKE1BW9YjwXlkdj/FYcsBasL5aqUFTTMIPaPZw
4Ud4HIkd7+Qztco9EdhTD3dlqLhn0/ZOqJK4h9NXcnzH3iq1hEPXOm+zIGpLeSpOx2lcVxvUdEqW
pIubHIgXYTLqWYS0bFQmEi3/HHsJ0NHQPBgrQAG/PkyMCzLsbEsY+zXI7vruR/0BLHjH4N8UKjSW
OemrWcPeQ1NRNlnznSzcotAWA1GUHMC/6HoqpXTH0mpYoTZQqMiV33fZEUlQ9BdelhVilOFyKD5I
WpqLfYjgR5yGGO4Ofmo6ZOt5hVC54MQYOBfz7GyU5kWuZfxhs16QZvWK6+aBEhIbMBj7MGrve8Ds
+saETayMYkLLrReTrQK4NpxsHGgP6eoNLPpvB4F2CRAwXs9bIPUlOZde3CswXsUrYyWb9vZ4Y2mV
6OcLqP4l5RvRCLMlAEyfk8UKFAR1agYzm5cTCBaJ2WYEjAoIws+WWYp7VfvVSpAqh1PxffukxLIv
JwtVPE+HN2nTomLH61N6S/fq9nyzXHLyWVJ90iD7oX7vkbgODTfVI9d1wUxTNmOlHm1J2RyhzXDW
PJqTI/WE3rAZtyOgMQQ/PFp1KAUaLLeBY7cZo52JorXuvs3qSvhfxPcGiXHXC8LD976o7+zuigWH
aRB35KvS1SIbxfAyftAkbllHvdTWOhguK3yqwfXVCo35nIezoY0ekIKpnX22uJosOLDvZ3n/nF00
ryQSSrxk7eryQd/40myAXTB6C5fQL6WLcw5bLvm+VbN0dtX5/HePrGk212MdYe6AarGJCSLYBOYp
UVPDQAI1PcFRMlNa35WHg6BFhJCw7m+XXIbPeiVzvzBPooqHNzSUx4gwe9VqlAqHT4u6QbIgzU3v
NQ0Jc9J57T9Y61o7dIKlK1k5RcEZrbFlSJ65M+4jeJhkzziCAih3xkFCxq1oPsCNXp9KcaAw9Lsz
CHWUO5GAaZ1GPV5pzE9XkrFEzrNzsyYwKnKL+ub7rA6752GTP3/7m7MsjVdCyEdVxDCelCQRmvz9
rv5xA9vqqxyE/tyjXQ6O4J3TU1jEEPHrhJhchgkb3RVRxku/4Pt222inXtPl5XSm+IMpUBP7RKTI
yHnnxOIIOVIQiUGt3pVX3F5pVpjf1njDYdZNHls5vpg2hc8fVecwcHb1dHemoJSNEZFvh5+koLhU
zqjV1F4byVDwsujY+aPfxEWLEQw1Ou2wkCeXX5J1f8SrOuyup2RH1LH8ofcq5OLR7s/eMMt1hQ03
XXf10VN4DOZ4YfxVMSbYOuZzNVDM104u8ekfFLHQq48M1nuclKcNiDm+EgNdtxlAz7AsDKMKytz7
lRb1rJuHBg6a3R9NSsf5m7u8P6Sg/d3e7u2RgoHzllYbjfHBhBUMBv7rjJzss+Wa1zxePhyD1SDr
6JOHf0MC+y0+5Tad8BcZE7IlaAX9DJBm7Hm60cuJdvZgtn1rrRt5Tyx65pvptYsG1+9/B6qjzGOd
Y6U2aFf5fJqk9gEiId4/rbn4C1Gr2jOwOuF0YbQyHKcFAhPxItw15ualBhjjh58lZp6sCmysyuRE
lMMIwqf75Xyj45Tni83+vXgoqTLjrrUGSkkCD2LWKigWyRoQ0kHxNK13LAND7MgqKUfA1vEa4qD8
H0h8Y9aJFcYu8VWIFUdv78wcVLKGdVzvcygvcKJWJ7VuXXhX3tQGy05YPq8utB6ME2fxvZG3A/cV
/ZI4MciYmHFjyZhFarnIOh/kkq5IyxftClF3L2PHDwOGyYTapCWlY1NOuyCwOWrVYq4fH0CcIas5
B3o+P7J/Y/KqrdM2sdq3Z3BpIq0JF/srvuWGOmoj0o6HIjI/X+YM5uPYMwjRdlQTD64KccV1YCC5
C+8ULRo75Zf1PTjyWPC8onS21Y7QdlO458XLTADcMkxPDbV7/WvG716k85uO5ptOIcIrAlZS1+/P
DWLPTagS5+mnUeznLlO4OdZqRO48X+/fmJkeV/MdDUJMREdVRSqVsi1u9TOsWwRcVj6IiaVlzeEO
DlInakDID3/MuCX0fc6WHHjaneFVXGztckVpQA6akydBoRRe7QDMWhRiLZ8BSXYdJk8qJtJ11V1n
r3CjiatM23HLsBUUgfiZM78f6ioZWCDV6pAqMgrdHnAnxY3q3R/ZHhp6Ud4JAgLImfmePSda3aVh
iR7m9GtRKEap7q6Tfx3dz1EuGFFKELJEEssCHfgu1OvWINQmau3yjmFXSsvhy/fZ49qDoRhXtexR
mCW96piV3LmrLs70vaCXkpynSYTW/1KYa9BXdFYbZiTgMmZKaD45AklqKNFbUchbD2TRdHoJ7a+N
BdWgq0kGxoHFf/azHicV0WA7INDs5NjBDtcsX68dCFE2/Bal9j0GgkgN2adnQ/wTz7+pqAWaZpje
dxetfisU9T5TZCfGFHNe8fd40P4gnlufCEpYOi2JPG3F9VXiPjCLE7fneeGasEa9H20cYPhkReS1
K37DJMA9kWPQAjG2ysUuDBHpkUbcKIE359k8VZcuOZWoqUg5r8+8vDqKtLZ4v6Nxp+t1XBgXR7R5
GcdRAvkXjCfcr9jkJecKb/WSD34gzj9r5iS/EgBo3njqsH2MQxcLMqPjMN0c3q/CN0aZkp8FGN8U
DClJShMQw0N2A1xCTMzkYnqloXer/jJCG+lSXSLeu3btnXkrus3X1hZeSCBDx2U3G0gJNG7HdtFw
jeNgfrWGD84QK+6FtP0C6UQG0ZyrIc0TjqRec4e3SHTssuFLBGUkP066cYBOzSH16gLMWG41ONUV
QkmqjsCBasF4/hbuqj4auQAZWWa+WF1aLvV0y3L/7hbH0ReujICvhYIZo8zTda7vd5bYDsbqbmTK
wFWQ82OUuKcHSwRNjIbM1k+yJm2OyG7CIK82xyrKM0eCKTzlakR1hKhjRv0ug5EiIo1Q2vWmScUw
fi3WTH1juIZLP3bTwnrcLBRkVv2xYLk7/9R+bZLAuT0nNWAV/h3SEi6gqk/MRtZCz81KA7GuZ7S+
+uPWE26tmTrmnsZD3Pm55wv2oor/uXuffGOIZJnmDD3ectKPZNTyEN7GCoo0oBuKEfqFVu0zREO0
9VHZXXvxBxIYENltXCDGK4X1RSOitxwZjY5cSHRhN6fCpmBYA6TP3AYJLE6i7oU9vIdL/2juxV5T
nR6fh9qdWFtTwPcOp+mw4bDE1xluB2Jmf19/za5Z3oKfVinyrReRaUY6B3hL98nyWfId2+T9S0MQ
MBM/K6TE4bt/ZG9gppszsx6GVTZ2J6PVe3Xs0UcglxehDIhpKh8pGWIJcQTXC50GHi7KfFS5FJVF
gp8oh154+LY+n4/iIe8E0h+RRx4/PLYxJTdu9y49ToAPpaDtaVc73oYD0i29vh43Lx7MW+UuYT77
Cb5eWsWB3/5odufn1u/S76QSpjrH1vV5OgEBpFcMBxFQDL8Pcpr8HO72/YoTxpIOYmJWWH281O9i
2SuynGJMBKeb3osxQtAIPU/LLWy4wg3J5HGZusOxym1rS8rsDTMtj79wcUNXXgbt2/hPMbRdGo1E
QkqbZWNePZ3GWIb9691mUXP509Ykgv4L8G2gRFojvYkuLx5Pbq5g0W4AIt9dF0Mm2Xxie05d7dlS
du68xEz/6PdDHIPU+vbcbLIqKD6xMooumtt6iRyfZ0b3E9llXS+A46zJIEtBe8rrODAgO8CxpabD
6cekzOFNErliGcr9gB3WGtfz7Z46g1WxAEV5Kabq1o0bzkAUOR/Sj2dKe/x8zQUrv5pcb9YzUVhZ
vLDrQUL4j+M3uRKi15Mp5Ap7xIVc9PDt+7dQGQvSLTZ9YVKGji82eS37elCeqStaitmT7Hq3zDQK
d6+Ii1IMaWIoHkKoTGVrtsZOaC3IRHpgD4QQO921sjRw14ZLqVJFDiKp+S9HkG8HouRVohiuLByC
WUE/6NKSw7a5fOsjPZGv9eLglFZqVxZEw17kUrZwZVhNd0vNHcsqMmEOvtcbKUq5aedRhL7ijhLr
jj98mJmF/VFSUQKMO5ljD7ylHPwqqCpJW10/uS8DG1yZ7Nkfss1Oy+7bBD0o3iNcjwF3+25uKYfF
jkhJX/euKrOLvMZkD/XvUDtGh137xmpBVCcQZxGP7NK2W/4xdl9BF+sSr2GaRJ6/bxJiKBwMS1xP
9MpgUXawGiEA49O5AFT/f6UR+DKn8jqnK1Uf8hWUEuSPwZYk1xAo0HThg9ftLHBjDM6V9ivNkuAT
HyetztFYb2DE+N4c0ypgCAVmBKlvF0OnF83i+bhCExZ6L65d7oL0GPAWwDwsiT3wF/3ESPUTnJA0
XTrye8xdPeS5UEkxWp/WM3fRZZqsPZmsKCvFk5j3qpjzqUCdYgRnvXG8MtDCjaIxMaxIOYH6Us3y
rC8+0VbGJy0of9/5t0SaWgw4NI6TdgaVf9yrXnrBigzjFgW7T4jBuSQJs99MRlJIwrgj6xsHAlDE
qKel2R2SN0BfVfWeMufr8hri6WQzWbKcVfDAk/B6WJX/P5stooSP7aksUDGWWY581ZUx0WDXYT7p
6ycNyNG+oIHSNp5AqUHRQXnKG8iTbSLJKNk21xhUCs5wyZvi+uyoTnoMJWuvUnuNP+HIqXE5UPVD
SxENBa55u3zR0mBdBUGmhSG9EnVsfm1hWIE3sH7tSIALDQWcazdIJ3ncSVg0TQxuApJVXvYd01Z0
bh+bosAviKQA2X5rdw1aOvJ9kWU3SICo8OkAx7S84uLwNoBRg9wjXVvgoxcexIIL8SndlRaKM4A2
xzqTIbT8noHvnMxBgyIQJHoAVdscYtOMAPEBKhEU37ZJrG3yXXpXO2ekSWpJWR1mEfiXXPMP1KUU
WL+zt/xL98DZ2CjaEX9FPb6iV0kYEcFEevBlx+Cs5cugsd6VNUUqybRGJeRQ7DMKyYuwELIBD5GQ
fUDBbBazoHX+aol7yfcX1Fav4XbBjAVCJ/R/tf5d9AZOdOkU5/UDMe0geW6i75hehxPLF8amEL7P
kwcDj2JnZukTQKrTZPrnQJ0Qb/sMTwk1m/8mo3YHApMhX7hFpXi8aT/PwAfZNqE5QVFCJtEwbp9s
jXL6IGzsYLhPdQpa74uRuCR581TSdoPh3jLQDfUhYOin+vixSjWyM3VSVQvzgtItQyn/wJhSUxLy
kkZmVaGeyvlreIMKFJdi0QUakiqiooPfKdp0p946f1qJ+Pi5FfI638+x/MG1Fd+LNAhQ41B0zt36
deXTjRjg7elxSdyb58F7NeZHUgVFE5cfHK7FcktQK80TSQ+yc5u0to69ykOLH+rGBrIA3a9Dfhy0
T2OaakOS9xuwsG2it0NAkmLJFDI7Q4VcrYiFnoYLR1JP9CiQuYKoOLWpeGoXNrVuEi4L/IkLeID3
DxVKokjmAVWdFo/G8Yi7/QxBqWl6iyW5i+uoU2J7S8LIVdwGjy+XY5ryvfiqv3cKokVXYBKTLUcS
qtsxLlw++eVgAv3OZaZ7y9L2th94YH/b9Ynn2EJlh26W4FAPgmceBz5GADEdcBDO8GQ0pUcJIGSP
1z0vWqq/B7Yzdxh4n9ltvAghg0ANnsJCjnStIEMzeA3NTZ2hkWJA1tlgh5ULNTtqFw0uF/fC6sql
eV9ALv29K1C8Id0OfbFqSZZJeIoMZZZmibzcBCVizmA0lSW9DgauoZv/e14UBMSnsg9LaImpRi3Q
3OYj9caiJweNMI3HdXjcFUW9gRqqoYOuFjlV9ZhYZbq2u6pZIW3etjvTfO3spUg11Gzr9xpfIOVV
PdjwZDoJ6sTvJlKuJnkhUowTvsUQCxu2FoYkpr4jRD/nIJ3iKVdIU1RGgnfjnNMeaiaMbDMVeZmf
Dpl0cWM2mywLRJW1QVI80gTzhMpjCHpMYZSWIMSnVXHe2Subr7oXBik/wlt5gZx4XmzAwiJjSJGx
jbze3m1mssoLHZZuLqn4tY8uNIg4fXnTe1Z9ip5OMPq5keuezdXJnbFmZyvcrQgqHpefBdJ4mNf9
qHCWjUiMtsJr5i4Mod6rn7tc83OWAVHQPSfHc1Muz+7uwQGh5mV+s9ksBH79uvm/grM9LYMlsI68
kMOqDFdIMG8+aEJkAipLeVZSYMVU5NE4PwZnICkynmR2V+wnAt1RMGI/rPXg92vBdA39i3nsqpDO
TmzK1OySVWAFl4cxn/eIx37c6/R6iTHtISt6K4pq7OdIDdKAeY98gD3mfUDVxuf41JliyJInWflr
ZeYm7ex3tGSjKcfFrOav57NumFjTEoSQVBdzkHpzkMfBdDfsRrVnuxIWOw9FOkZ2nCbbn1IWLlxx
MDQcLoj9FaRBA4c/xmZuAJ+c468Ztmcr78S1+KKP4R9UTmGtj815yMacHGVjEYvFPmPn4FK4npwL
1gi13oT3SkGlpih8gus/73THK9DykzzPQREgq8IY+q9WRqlEroe8xQWeHflnMleBpiJYnASgJk4a
VaoXNqpkTe+A/3wPHnXX6xpY8k9tvtr2Sl8doaChfvB3ZCYuuOQb2xExDXFpJSAN4QMd2NA9VJEs
a4HVguEOJZEcBnUe+6bv/RawTSsFh/zWBZNV1feWXV5pbGOaIdSL8jxPWj+LskfXHUZUIvBp50dx
9frJzr5PFLF+/soKrPCa9Q2rtJ4/hUWHVz57HthPyy3OCNjkxDqd7RE1Msxt8mfIi70budrgJpx+
KFjzAY6Au7GRjb9rQBeYWrE+ozEzfUkccXllH6Be/L7IEf12QO8e6R88iIy+xQzjEds3MQeEGdsT
kOy5jpT3lEV+bo7yz4THhemgbtitqqLk5KkwS4V+ZPzwHtM6WpzhmBjO67XCuqKvSpUIUvrrN/jV
Fmp/i4bNZHcDoiV3RdtH8M9/Y8NZQIzRWPNGlc/32K+YwyvULxpecGt1Ma5LPeTGMf/1/D487iOo
fNkf1obI36e8282F/Ivr9k4yFbLrqQhWwe1oMXZG3PUvVRHubz+wAb5/ax5DIPuDIaiIjQbdRF0t
Y2/fJIP27tOOdnG0U+gD2QvPupYDAvT4twy5vJ6weFOyctQ/cVD0Azlf2HtuBk0jxKTepcN5Qkq7
qm3jAOqrWe0CDLEiI++lib1S/8j3HDLPNp9lFTf9PY1hS5wLSK+9y4ffN2n3m+LDGZRMtKlrqGqC
CaFpLZbLk5DV4x1sP3TJIivv49mYGTGLBWxxHgZVl7WSIHMrhoi2pkgR66bCrftMG849SHMv+0R7
UPkFgWCQ4AqE9DNbTphj5DMIDyxqg8IVaKrFldugUnq31pQ1F0ZgwtEOmG9MT4kQQyxvAAcs9KnX
8WbCba9YNgeYQfplNRZhs3ZF8ReV+Pb6z0TmPAhPy1tzcf1S7OxkSSC6VXQb2QTznbO/RQlpUKr4
fuUdWE+5HqUHXd6CN1DTr/LWoYiqd8uly3i+FOKfROWFroixblazJHeJWV8QiXpAYpzB7mgeL/6x
NAQ/CVyYcog7zu3ZsbiK/ArI8VK2kvyBqYyRpr24RZL1gfiFCw8d45eUZHY43Y4cWzCKm9AomPgc
3Fl3/ZmNOq2LaoHA/ChzRBTuU6U6eU0ISFd8ppqSLBqKvGfolVEwqQm38Ak5bHB1Q0LqD9f4qzqA
Ovvo7fPy/hEiIz88WlaEJY+t+42rzMYD12/Yn5Ecxoi7vXvEfOmf2iwMuFKI8t5xR9na9Bn0doJn
GKpNiUDHsduTz+N9yC25B6jFoSE5kVhceFbkGyzu+iicmvgPHNCDenmtZUFJnkXknMDoLvUGrKqL
JuRTf3yvLOwLDEmZZK3vmDj+Jt7O96ijsWkMHI6GYKpJD5j6KHYnDqbFlSt9+afHGW5w2YFxGV1J
V4LmoVXWLU/ojk/VBLAgPFA8rehB9yMCxX/B3o/1xNpaYfbA0TzcW/uu5662pZOx2/SYzvEqcCkr
KF2MDSFdRAkBkxNb0DXOiLGc0CV+TPaYsvp71jdFSfWj/LPEgiLZvIIijD1l25LjYkC8FEUOwZnQ
OHZyBLnvF2eRsaAswj7dNDeSSwUxNzi5IhnZGARyjXobQGRnyJR39nzzZxNNuR5uvxvfQ2/+Sls1
/Ut4Jr9hKajPTkAPx+HrhEWyKNcfvbgENRBqJ5iUG3fKUCgDkdj+l82WEObk6Je5hYoci+zGj/Wv
R+Kkq33bdBEXmqozPCt+tqqYRsOAkcAji6+iyeV1KFKSaJEvBoY1mfHWhthjwZ28SGx++qTEqeaM
NU5pHu28faLDzBVR6tln671IdUaSScRFIhLmMGRKcNwoD5sVzSkiF2vwba2zfIhgjpeKZNtYMQO5
4AjEeUeOW+leL7G3HqlrJARETO6c8+J196QiJOgK/S4t4EM5+m7VAP+wJkFLrFb9EYmH9WCvvmG4
A1YlOkBTzUMvLdlihiwP14/g+IQqkzXnh57duFSYy7J1thGHHxwqOv4gvAJiuItCX2Z3FeUqkyKh
SjOgQ39lrJy6j8DVbXxvMa57CPDUx27KoQb7ZMbg103I9pbhaqEntGHC+eeUCls/Jqbo0cLo59GN
5YKdivrI65pC8+LycGLlzRXEYA4SEoCMs17jzS3w8afp+OR/iRJvki2zeT+yWdnEmcg2bk0eHKlX
ZeWLZbboXLZh2FB8F2vnoC695coTye4q7TO0JU8LzYVImopdAlZpkQt2k0Dq9uTWVBaQNRp9nds2
kbnjb4rM3c8CxMR+gh9QsPAu8BIlb6JF3pNBY78kHqZrp+svz/NODlRiNwmJDZtsZqd2zvOfHq6H
luEVOBuKR/M0Aej3w9FQe4nBFV283QdXTaC894yuSWG+fUQjAlkKDU/webyN+vprFDUZ7Yc5mLKV
G6zw9s5T8k0MSkr7C6cHc3Uaoa0Ua8xDUxCrCZ86AA62JfyRn6ivMkMbrmNNNa0KwHLEBwNLk1/e
1DaBELxnZ1Pp3MMgzwXf+6bNItOFxHjGiT9gDfdaRu5NzOelJJ1w6jSUdmVHWz8Aix4Qp3OBZD4V
fLHKPT5GAe8zUr/MTSaVjaQg3EP16bkopan4QnxoU3fRSZWX10pwA0aysIls0Cyk1WOa9zrpy99o
ujZGeKnULcVXmDx0qvb0hyIR+jycF703EffgtqXsnHfQXze+Ec/ewDYPW6c0znA4+gOzH0FC4g+z
g+5hMxbakV5SQop7WQ44AWqSZBTxPt8IKcL7lzep+m2rqE35zFQxw6eAWFs0dTl3ABGfg3RjZdXB
yP8y/fbffCYNJAYXpMqCQN2fE9wrtWek6O2LCGZLVfIx+TCdafhqEGyrArzHeWX0sZIvTBWD4Gl0
qGqjENv26ddkMffJwmehUQsJAXhM9Z5gxsNDXsw5lmV1gZ+01+OLo4fWzRXx4//xHkNvZVXnlcWu
0vp9cMnU9EgEhonG8FRbrNQmxx9dE2tnoyEm4DzkrIGZ3WqUr6L4K8AjqcQsI860C46/t6cBlybp
DVlceusYzmKHxxTaKUjGY79/VXLXvvwKvjBAwV9AT9Zsh7hA4KyQiFLZxIHo/tDa19ADgN1jHCvm
6j+MQQV5HI+rye8pAVAninAxoHFWYCne6wnqJXe/L0LnjsP2G2EJQ07Btspr4XdrYKwz5LgijLdZ
21Hka1eW7qCYxTPnkiH44LJSQBxyc9c2w7AqZHdA6qYYHW0uWqiQ3tm2PqtFEaHC+2s56m1zYOjk
jri/ZjNQNDRWlBvvxbdp4I/Jnarsz63KEn3Uy5IDGzGxHOTho4B2FOvL+SPHimJgKFhC9iibds1o
PH8Rm4nX7ff78UvHgB3CemenQJ16kEtSqqhPc3kdxQJb25VNxiruEL0mUIWX0ZwufKS+frx+Hm1u
fGpj+XJyjaDdbHPk/XLDmIp7BOJiiIfV5FPpJQcf28U0/Rghwyr0yDbTbWBTh2rU77N+R23LqrZO
CQfVMlrPdAMAhh3P/jYqGvk9AnTpB4sWAq4XbrX2vCy1SwVY6hhScLS5Sjs0nGNzjmuDbemHqo6A
E1T8Crn/D8RhRinEqDlwBttUr9swPVOKRyGIAVzvlkL/kS9STNiM/84WNxssA3ApF2s20dxmZnmh
ld9SnqUwdNBO8nqtbsmgdY2keLdwqAc6/fTIQaerZnvMEz9uhIJPwtvxrrwzZUH1BfqGilHoBZpQ
xXFq7hfvYawwkSZpKGi2WlRTlidssRftmpscWVq17L7TnXPWAm7yCz31VC9y3jygXqBuvxmjEdOB
MmL/izjAyPM+OqauVjtRoki8WDq1OMhNn3fHqQO1mjJBHVnWRG3aqLEoaWbHXEV+P10vrIeU2PDF
ljmy+Ju0P3UsKQglPbirsz7UlPi8KIbCm0YnLHYkh0doMzO8MVd9psZWPO5Uglw5QZv0vm0CBWl7
PRzOq5AxNCz8ehCn0T5hJlHml3EMex7MYhNOeDrz4PQhCO6jMMRMRUTVMDcKuYDROD7v2qbeLrmq
GsKNrBwlxr/Ll28+dhAap9ew/t9wxEUTBuN5q0Ho+BtMKm0f3sI99zFHVbeRATo3CJcSiSz5liy6
UoY09PdC1j2V1kUDB1YAJVdnd32RX9DrPEWadV+q3M4kk9i5qBfISOsdZi0Tx+D4idTJPqasfoOi
bPI4dJ+NQe5+zExaFeIxxeD1iJZN97tEb/9ZwZ84OJd+g+LpyFNP0yzteW1G8wc1LL9Cijd7f+eL
EL/U6mCIWPLOfe8YgWhIswMbgqW9yyb8259rjwLPkto730/ySzbuVPsgjjxoAH8e5f9njzJbZAIy
dNkRKY1F2tBN5MvMwH4WJxpnsxwYxpnsmsg520AfKH7T2eQEOS8xqVT72R7Cj+G2kMLtwOy7kpei
vLI0bmqgtSp6S3v0cOG3O+zDLieGmfJ7Ft5SROCgvkudB4fYAh2qLj9WypPa+FYJGewtWffl/vom
YJ9vprSsFSnL/lD4fOyOKgFrA/kukSyCOfr9vLtriYCSarimN7n/w7wftGvjKeAVFMaIrix2avNm
AmLsQbV9jClaNjXX8ja7aLUPU01dkWgGVbdGiIkep7GZLgcpftvm8aMJWD+fwB9RiZV9pcOgPLQ+
m/Wpg5QBg/K0c9UFhKqa/P9BipI/qk2t+VG/OXsw65TbgWFVMx7OmU00QXnwcaykkxAI392YUvjr
7b3xaiEEusnG5Rquazx39JwullfWV+56SXHQ6cBYPlDL8oSoHhz2779s0vl4IN4LRCkpYkiMzK29
lbLgqxyyYEpaaT2G76CRhAZiRYCOq7kOIX8BOy/qy04an9qK3gmtW/AMTXhMcPJZ/hWUsCW/8cFr
YkpaIdWFU0+E0end/SYFZOFHbNKm5tLFB4ZKUnWwEab/koALWapYhisY9SOLAc1ND9hApuQHSjG+
C5CvRAVfARoN2omCnxcoXVcHFThhh2Nlv0HsqaiQ2975hkZ0+JzzBeTZSswjyvAp+Uo6ibyqdA8B
s3eBtMHr+P0IEVAejeDr7vCAJArJa8w5W/9JLFEMh/uwugVqAINKs0SL46Y9b5nnY6tPUBA2a9we
410Sic+ypoW0UWrx+A/+z9cRdr6TWzyEHESnk/HHn2Q+pGPODkv/xwy3yv4ZLHFWRCiOVteM0Sbu
W+fCbILeT7wG/AwWWtCfmgd1xHvW/rwa0KzLT82awextxg+/0nN7iPXwehes7PYONJToAmb4X+pG
gkkZXxZcAOMYXrQgfAW1h5u88p+w+iBhcY8DjusMl2Ms4Ec2c9VDGdFhJU9ZDNgco16ibNJBjRU3
eoCFtggcfkmrFJW+KMNGXFuIt5vkDXHTZMgsGrs4Y6i6Wt67mg2WvRlsmKyyWh79RYOLDTLGSz/z
Z3+9GqGeCfD14s9xxVLwMPyeA2WxkhNraDApVZFUmtZNxm9h95ZHeApl+JaAjeXrXNfs6wcNZtrJ
D0VuEmFdIwl0QUCEEMG+cWsmyCVUaAfit6A9cp5PuJRq6msHHsF2GQkPupGfdndjBYZ99yPUKksg
WZm6+obPSfIcqykRr3Uzhn3shNYGc32sN3qZT6BlUvQ3R/yW7Jh8oAbqNhqYhYS5jTfo49StRe7Z
k1R1jmO+JLwomjPDelP/7C58sJW5wLS4Udr3U8kGMe/Zaoy8m7lcR7myUQRegvFXAILoGdLasxlE
zmzh5NX0JUwVc8WtC/KElE3wZSOcVlMWtK+RarzLqNKx6w40TDDsQCtlsHlEWpX+dVQt4y9OTgRm
GmSk5p7PTSiLiGzXQ0e2GKFSCiurbahvOzFbMNFzFRPsM2kq8XsrpMRSftPHLNYtiaxijcHE3y5z
tJ84xe5jsBpLg5okIm+YkNrLF7mfdGMf+p22klyUgCWALgba+dZMVHAz60a8w4zh5r21eY7gpLaL
A8gxoIQ95XAW+uhehtgHwpOBi4ywmIoinGHBqm2G79OSWKHMFMCplJhJwTntvRkQjJQfAmNFPqh9
gGnNt76Xd3/EsQuilEaLNSBUskxSlIuAsV8xKWhlNaFlgx1dBC6URMBjWLD4LeuczvEDEiFPyP5h
4O+BJv+m0Izw9r9bR8Mqt5CTH5fBVkNdv/dVByt0C1WO7ogj4NOvD3JPGgEWo4/mK+8FPUO2A9PK
WOT6qg4tkgZ5YxmKra6PVmMUPrv1XTa/rvfn+IxEclY/Y0xW1FZfn3P4weIP4MaSMgrU1n1QEgF1
itJWOcDIvz2YppL+7pfzSl/dS5MbUc99EV+uR9Xf5m7VJQoJQVd5e0J1U35mVaJxpStyuVyP3bFK
mr9gi7W2a0nJOAH9hXeRmR12ubWuKLx7eyBcgO2DMkjscyhuwwTVkct6fES5GTGvWLR3sKYf3Erj
AFm6KGETdBxf8dbUDUG0EqUaTYyUO+9cbj5RHUd47BXmssW2HM5fNnbdoV2l67X6EX0LGyUL79sO
SztA7/2kqaOMwp2f/PVDpoS5Zk7cTUhHCIXs50xJJIxMn4gHSik6MUl5n6O+O/Ahf+sOpsH1+V4f
rjaJAYZbwBTzM4d4/kd+UrrmoKrTt3wqKInTbBhgqG6q+D46jTLfuLPzrGgHcyAGHapxc5LUxUJn
GIGsjFYVfOUxJWzXvR66VyJxIdgCIKQpaeyCJ5YKiqFSfaMGMHDWyx/dw6+kgx1lq7ZJvFE5AGaj
8N6KnRRmfDIQN7EoHy7uLa3m8WHG3hFh2dHN+OwEk0m/Gykg0N8RsTCBgQcR5rsKij4FgZtGrExD
B4CFKMHqugopeWShiqd5cmps8+P6I6u7HXQVr5YAn1pdeSpXD5FfiSONVNu6HgJgTgv6qzqVm0rm
L4gy+KsaDgDpAbYnL6PY0vFgk2PtMrrsppF1Yrc3/IwMxgdBcj0X8lI3FF55OF69k+JPqXBWMpF4
nUbGudMwRDo/fv2pUGfyvkZWYAw+B2ZNc3zAeRAP8A0stVCDqYbVOsB+VtNmeLDMimj6Ys4MUE8S
MFfbuvMkUFhuceAP8U7qHwsuCuqlGChcxO4IHE9p0Nwcej8TAYWdXVAHL1LECDuUAYePGrJ/y9XL
f+BPONGfwGOe1e0AK2KdFHg3MO7JIIg6UIwnPf2Fj3BhzeVqemY6NPRYTeCsXJso/s00x4eFdVlj
SH6oI7uEcaWwX8+JFQM/mbkoJJ6nqovk51llQOeKMtgbs9qnheiSnPj2moEGsjjAh9Nt3Gx1Yukm
1zwBUcN8FLkU5kKo+fpsTNHXEvyxMqxVvz36L4NgYsaAfJm1MKxT5xNOGEHnW/5sFUPOIu7GIj0l
/jUeB4AcW26yHx/XJpUy7IdtaNO1B9SFYeEN9D0Txfa3+PwFeTgyT/1HMfB68HJ1LxOvuUF1niCE
7X7X00CrVSMIM6nSH46nfBymlTnQsbCvM0zYqMRpo5QW+HbJKR3A85Z8YmXh3arEfV48sVxRILQQ
VIRT0/ak6CeV3Lc6304UlQ4hiSfSmXwuiARJ9o9HCKaXKxHH9QoZE7SHnLO6DMme6eUSrASmp8/Z
P84xP1mMI8YDMu4QEceS7YBj5PFuNfVL9vp1vmaxfCPFE12EPDfEGnHOFKlVP99gKU1/0Z0U5scJ
gc4myOPM+POY42CSzFpoQ+cJl0atHoPwIJfsc+bYIIuZjVKYFV8sF3Xnec6GdBGCCK9atWG7o7tH
zVsq2tfuy+RVkkCiL8QwufwkHCDzvmykWXOdkCNrAMPOkYq7RkCENr1tJVxtwgeKP2RqNCce2Hn8
NTeiLPd+wMGcX2EONQlL5A/+1NUb7F7GK2/YtxWEYLRq0JZD10q2PpaUBcME1Ra1fpJ1dWmNP2js
Bu7GT5NxezsBJuH4pFwav5ETRrDOqqAj4hgzGHNXtlX/+l79wVB9g1W4TDmpqRbiAUDibL771SEX
o2WlIp0uSzksINAc7RQABjOGJH9b5FK3WG/ayNItC4kGrCQpaiMZc9foHQpuZG6l8avzR2ap+LGb
VXfrnmhh2lwTXKanz9DmjOMkOZIJQcz/4pIgvIFsSXmghahsjnrFQ8N4uuQVvTyghhrQyS8z2QyZ
awSHJS6b8eRrhDW694GYie2GKLvHatss3+xzj9u+66/AFDxUuUF/Pw44vPzRe4/NcjTTNe5cEmxq
jyxnloW6J7sWTJ1o5mVSTceS1nPb1GIlscJP0F3gw9kWKl/P14MzEui+udgd8bcBQ8Vj4NRZdMMG
Fwg3rq4uDYyGWz8TM/YWQ9TWG8rWt23y+l3qItSiRiy0xGsxI7I4k7qBXum1k6zMCBcSUWKczi9T
i3mHCCxDN1t2yAmuJgnLmE2EMtcUHKMCFENZ0ZWJdEb+3Y6xOLP7vzLczUHLjx7ZEJEjL5oOEJX3
BGs8lrnpfjakNSzLsvePFW0im12Le6XNuUqNBAqVU77cRVz1xaBgCO64TaqUVU6n6CzNjBHJ4/1X
Ma/mVuGAZUad6iaCBXji3PUCaRouprYRPdTxl3mxiYF06riLkqvq3ZudYBfzdqQVUixpmtNxyyfx
G4NCSdQbgtJHzLehgw0rbQrqEY9luQJIxYDDx0k8lt+zQ1NZEeCFJfp1H7qYthCOMP/LKZdAf7Ew
1S/97FcCiV5C2dpzpVO1ULcEXG9tpYvng/yZOdvTFNI/vHVpHc5oaGuN16htlRCwH6unj62x4VrN
xKm+L7NpnQ7p0A/66atAzvs9zG7QjtsbNYD+hajFNjZDRxqSKp6WFtlfa2esiGXuckltuHkxgAQB
yQI6LdSfUbAmAwSoAsHe1KDw+EXVJh0dftLjNbwlr2wCSyiQoeiyUwoQJ9FdnPJ8uUhn96VI1ldZ
VioSlI3pdhqZdRmE9KDb2ezjodWRoYBlO1NK7uDZFzzSVg6PPEuVn5TLtUmuR6voP1rllPf1R1B+
UxhyHpkTgNHk8Mp1lLnMIZGKisfbVqVQBjIUCIlAncvYcgrbmTzeZHyZakAcHTQWTA0HEfcXKjqd
K4QdgVyQpSRM7GXuI1iYhR1AipuBAzK3m/SBN/zGROfgLKPJdAch54gHNdRZscj1cDKMCqrefcbl
mxGs4m00CYtCqTHBFWc/vb6iwqw9HMuhI1Q/thxOvy3DagcGuVswLj/63C/THPpOhXN/rhixiN71
3PzsaVVuTBSR4UdZZT21UtQUBjp3YY7aIjt53xUycVf8AVBfd7UoQqF91lRwxFu8TC1HleuFHdX4
HI5NJfBtaeMiW0w2BglpJoDiEaehOJ+479MJwbO/4GCxHNaCqwHYfMFdW3+FxJi3e+5olngPopJP
2xjSGNGVBLuNcaP5mbaXfD3ha+Ahs7FHVI62b6hHp8IssfXxFEhUkXta1LPuDcXnEhL1oogTN2ub
maGIhczQJyMgNr8GpaMduVUq9JaqjlFlon0x7xrPLzFCqVMbuEd6EjSrO/5HM16TAvqCHlTsjplX
6rUOsfDrlSnjmIkFGmUftOHnnSp9QxzPKxdgjzi1kyEIZQFHRhEI42mx+5gHnYGc+Se8pRU40rrJ
DX0NB+z38Exbn06QzGrGcmREdbifYAVg5abofdjR1tFtjTJQ3/sxr8Tw/HqFfPkcbqxe/j8+Vdhr
GI2/x5tf8+mQfCM6OzyYRnL9STtcOk5gWwsirh92mlXLk9wCtTacvPz0/zElHIR+ZqqgXYDoSc41
/znv1DstLHoDNY7KxFa+vtqkZbc1mLppWhVLo8C9eBBkK0TX0MDS8jp+dWvVFtoOgKBhi4GT3YcS
8XVlEMYP0yFIHuFr10dIR0GGfleEt6EXSd0tieKf4rRGudD3e/O4uGt6yoXWBdDerYf6dxuyI3QE
NmZEN9CywF8vK8bSNqxm/vYUbmeWI/78vpENrztGL0DccWZhNjHBW4kfGIAts5aPPFIWSMWubE0Y
9cYaS1eEU//csC7SGrb8GkPkKjzh9i5Aeyksej0Aqku6zlnMUs/n9Yddk28ZC6jdC56tiyO/QBP0
EY+CsbWLjeXg3ls//SNU4Yd9KWDx0vrt/2/vnXH1rZVuW8znUaEuOBozzmYPK+XXkBuDnmiUNHop
eLCOqOiD9ojGk0nnd/AfTf+oCeiwGntd6rPObsV5+vfSbJa6JSG4p235uXNgSN0JDBYCZ8T5/jt4
K6IOZGM1GgrZQuLlsHJt16ExFjv7Ms3NjzZjCdEMOeRD3qy8/sY5HW45ZabyPUp9CST5gh4aRdBv
ZOp14NkiXc34qO9S/0uXQVeOuXrQTYRRr+16HkSqTpy0Mu/K4NpYF4MEnVD/iCB31qmGd38JJjD0
Sm5wQ6el8c2E3HrISVwpZ4NVHvL+xIOw6o+/TLiMwurWvWjk1s3yMoGyL1CQN1f1d5ATTcY261x/
Ua5lMpp0800h5yXNkqHbVz+/orElm66ofC/6xY9453F3rH5UpdH0I4/0X0QhHwuNmT0FQ2E3cVtb
tR3zQYJSmGl3lG9uf5F1OCLpylPVabt1UvYEDTEGb30m5bEsTuawEeI+n/WuUVTQDyyFvkvEun5h
ZdvU8M9xAWHkuIJPGHgYjrEE8g4JsMT94YkLo+vjs3znyRovtqnvhYCoby+N7ipRjh/isXMuOgDh
wqRaEJqvUObEY0+LcdJ7Ve3tBHJVJgxI/X66Ja06xRdxVGpEZh6AdIg7mEp6RTwKGJsKUcijcsJl
XHKTXvqIPPxcbVucD5/8mPy2wuhyRewTr8gmpw1aclxiXK86j/jSOR8y03kNGIkIWbirLgk0bdUo
UaGqK13lS+azBO6PKKayQCkLYncWbpIX8hAzk7l4zxX8Xt4Cue7n29XmVGf4Z7MMPBoVngU7VWRD
PBXOoLf5zu25klL46s1Fp3nZPVvMRrPNk5Z0/xZSQnlK6MMnBIYZ81aYNT3rrNd1GP30tlSInXWE
k06HIVhYRuaZoUKORWvp55XtDUzNqpvWHuuumDY0jVk8gJOwIn2Mn9/8v/XJKmwX+evMt9e6sIfa
KJaqvY36STu3ADRec2qvztAouKw5D+6L6KEP4acUnr3iUr5EcGT2ermrFty2/AlnbBxuj58kGdX/
QD5Fzv4Ur0g9u7KuZD6PQyB2aLMGp1CqbqAwY0XUeA6QgkZ49CN20fOZNzzI1YOQfbriDYJp12wp
UpZUACu/OaxXq4LEyuXhAV5bE5YZ2JUTf8HLaGuFc8D5P1uPV8hT0nqMiB8qwbtbOCQUH9f6vwGB
awY/nGLPrLov2eyM5Fd6d/hbOhVdITTq9m90PZg8SplwJZoVYenWQqD4u4poOgTzkhHbph+L3ozT
EDS/YvWE1c1jzcyrHG9eZorOHxC1IoHzGQfPLKBPbFKYucjt+2c+D/cXs34IIq6FSYVbYlm9yqMv
pfCCHPpAriDuP72FArtZ8nrhDAAY0+xvp3OgGkcswgBWq1mzqsgY/KPCzesJPZG/3Bj3M/Seuric
Gmyv74+5tlFEMrSOKLcYc3DoHRFK0D4vdiDmX47jT9vlyvdAVxWajB0EMizUAXL+joxAJUs7SPgQ
nxZlwxWqVwbPfaKSBHEbXE/x3FPAW/YRvz/J6Q/DwWJYDuGilHsWglkGUif8zSEO5qMFye3oC7en
6LZs8NYVu43sGBjEoOH3piiPPd59J+cAiL8a9JsT660z6mhGCDx4OdmXf35vj2YAAZwVvtqNx/2D
5jCjqtskgtpPQtKOrSeW8JxfiKGmoeNRBfs76BEW5ncxZJ9VckR32Ou2FwCP9wRGJ3UtdhjH6Uu0
WrftgnnYoey1Lo/M2saejQVyG0ytBKw21oryLCM3IdjmFiJnmC/uC4XKXOjrzjM6DFi8zwhEssmN
pyVg/9fsLjrl5byPZqvra0n9lCnglJQMQakWs63PYWrJyHLWCefvetrmvNWwXyslQog88zJfPJet
xBL5L6ZNUtJLEJmWr3yjuHW62MCyH3b2FEAjEzwuzLRP6bUaKMByiR8ICCsysX2KvIfVHV8V/vYe
cf9W++Gbb+A1ahTO2CbWIEJiSicCc3p/bOBIMJkYdYOTulrF4F9Q95/N7eVFRMWycB8H9cYwwXr4
2AEqeSLAk/k+QvfzHP6sKmWJaz/UnF8yPVB+cY/q/SpZCmM2Ku0bhR7nCXW7IuwZwrstVta6Wawq
bUS8JRgvTvUOgEeEPGD1Sf8v1X8Y4cjO5p7jvYIaF6dXdOORTd9HLGISv+D4JZfhXRljdalpb0NZ
PczLzAEhIq8uDZfvubcSpcXBj3rIXAzbDCzKb60fmW9YyXrbbfYdCyGu3s8/17Ltv5vryMySpILq
+dUTgU0eHaKr+BfzEdf3k6ogl39NjtnYZHf+v1p+25a9DRsYf0TJFtid+hQjHePuqmWro3cRFpft
DBIZP4uY1gPJzczcapATwgaz0XlBAsXy/bqEEV793YO/iwANLKrpX0fcoxiRiKMZYA8pRxHgOZVC
4PLaf04uWDpPPJ1ntc1hdheJn7k0cT4dhTkAy/rrhyk5fNFfderOQYwrbqMHMykQcQoRXuN8vbqr
uMXVmZ1lgRv4xvr+jynSLb2GI2p33UuD+WtHCNAyso93mBszmd2KH5cPFsxiFBQ5p7PeoQGJZ1A9
x/rwLBs4gZlhzte0x+Ic1zbBrdQgbAbueGl64rZPQm+iIA+Ga3HxzuWjiYLEeFigrzNVFsCHphy7
cP+xgC2szVvRe4BsVlp/cGzmLlbFoq3Zkt9VMg9Bi3wsQVpsEkQ+DreyzFGYBUZAgn4q2BPMvFFg
cZ1MewwIscTGPr3v1phU5kIoGUIlcTbfQfsTuDA/FHiJD88wQleOdWkO7s1ISa5n+YKq2Ex/tUTr
1gCFjwmHLwUZZ8pEBwRo60NsfNDYhEr9E/Yivxc79IrS8ErwtJDmyrEDkZSAiPu5qVGmgPZj3kE0
rtaWnLa6fF6Jai/wsyWFwpFal8InfkPT35iAYB9D7DLJzp/IKAgYT0/1r57QzPTC+BdjiKmJ4wMT
MFO2MAvKzC+SIs9mL4TK3nOHBfiex9l0OdKCvzLWf68lsPruBQlzDahH/ctOAE9aZpzIOrq1w36U
+fkErriH05Qu8wDTmujBlowx4m/oAs36ynOeXcV4hfmxZKoC02hFNz4uD+LRA6Y8vHFkd9CBq/Dy
JLAZnyzKMqNX1x+hhX7uHaTCFyfwDjmtGGpT4gstAyIxgXo3A3vQS9GRNzA8E7JyoIKMBswD387R
SpUv08UXAo0HsQephe5Us5dLIrW+i8sXYWBo3qQqPfLuIJV8oY9B19b2uqk/cbvTrYscWoYjSIXs
YIKY3ESO3NHUizBdGGp+D3opR4qvAuHCKMSJPNat+lcP7OLAFDs7MUnDgUJGLYxJI9iEDpqjyKDw
eV/beJ4OMOBvbMsiaXGbi6OJrEr+6AzqkW1k60KOqD+PSwkITaL8LZ5ugMTUcCxisoUmpEqF6t3R
5g+LV+Qhe+MPheSEd06A9jsV4It5/JDf2GFhMsJFaITitUnBs7qBF4G8v6d+Ym7+3DhWnpH9ki+7
Cuc9k4hDk0tENV5HNI5LTyHo4bNjo8lsBa6Hf8BWgqIFlM0KEACynymYpHxJHoH+pogwimTcHLsc
s5S5+FDr5TeVyC12qDrVUd4gprnJ3n3XBmutsv7Ahw7kheY105is81lTw0CDLnG1ji/K86FNk/E0
odrdpqAC504z7Cyu4XWHvMIB4NRci/9iLNchJjvJBRRi464vuX8ryccoOhA5iJY+mG8cHTzLpauN
129nhO3X3JORH4iCuOSZhNbQb2D+zYplKHVjp7GmZzVdYQkXdH7bx0Ca52XEMIdGhBien4ZWm6Yh
cd3af/6wCxydYeny18VuvH9dCxobXWBA+9YR9R5hPmzB9WL4PCMWlcL/wcGd9m+Oup94hBuoDIJt
olknWMhDSlQ2Vvcnsylr1wW7snHtlHGxplByXg7I5xr9ajaS57QsanPS5wMQpzafsUigHb1mDZoK
xy3NPRAJRf1RJqt7kX6uuN1IFCd8FahsWgcK9U9Gc0H0ksmBOhajfXl0P0CBSsOfi1iEJ8WG+AIU
BSi5J6DfuQyjl3j+7QGF9s2BpI+341j+sQMoEUjj7+JqAu5e4Eoo3rbL82dAOJhq6tRxuzjm6LY8
nVm6JZwYThB7dHoY/hhnKa4VHQSW2ge/5mKN8wHZ52cQr20cEVka3CXhf+fwWm49CWvOkelRfLgX
GJdB47ySyi2kbvmj7atSfK6tfLTnCiQpCmIvJR3mfimheK+ymzm0cnN4ILw39GsDR89dUBwwt3+n
u6KlHbjxuak2OTo4Pmd8+Ec9JuNqwDcEHzEZU7t2RezwPgjLUeXNBGP9zcOpPNowWiGIUsUk8IUP
Qv4Lyr0UVAK/UFcPRxjcbeMXdMZILZqU71dMD6Nx7ljc+wUQUCHw9tlUpOmQlqBSA3d/w1I2AEi+
KZrLjMmr4RCv5cqRDXkdC44Z+b8dJrtt3UGbC385sYPI1/4mu8M7ojulR5xgbIhz9zBG8OuNlSbS
FVbIYeDIGfpAxrkhUZNoCeBg9046bgeypqTRGAesQdTwDryCKuGiE/ULOu/QPjgbxs/lkvhWLX5X
GenqJRwUyneRHskvXzrucb5y9PKacbZgswMQumB96NQyn2QpEZ08BXjfcbiJi5Q5uhul3XtDqZQn
LLL+Y4O1pMweAkuZcrmYIH2ulMHrBw4CnH8FaY87yD3zQPXHSbwAEpRAvE8+Rb//F09MFYG5vSh+
zvBdf/qgBSYxf5qU9R6oHBCnxWzXcYcLERK2v2URkfQiMIFTBLSW2Mta9rnd/yQbiOLtqretKjci
QKwvG58VPASF3JuI9egYe9UD8eUScQP4KOhi+2wFd0YqCTZnVSXnSurJuPfMqaIWdh6ArJAIU4kB
fUFwFHl1eKNNxe0IacUSFSQW9fFQLtZkjxUqNcT/F6jAxnEw/AiB0Cp4p1Af/uEqWNDtKNGJvEbj
YM5DfAB2ToW7huKzhMwz83oBZ0mVpGelCLdYqHYkQ5IaXSNZS4Q3OBkJwtddeBnP+ATql2jWz9hD
I1v7g8CUOIsg2jSWAZkcemb6skH83Hd8A3fnVTT5boSz6nN5ygjniEVsDdV2Vg1C2uOI+GhAw+sq
Gj2wD4DXPFB5JkBh/+5sTRU6z3dk2GJEwL6paxWRI9j/7bsmqYMtaC8zT7UuEEtMq+lE3yXn+F3Q
yXfM/bFR1x4JsjT2UGy04U3uojWMeMIGQOsLP90FjjpmJsvJgThqH3d+WbVy6+ZcaOsSBSTcNWZV
i2w4h+o8rYLE/JY0X64Ldykyu73zlqVsBGWNxDJn2gg0Xpnozb1tWbiiSiIN5JkrKRlNd2FS3w3l
a4nPCDsvMNny/ZpDrkTUKSjPqLXpKMrjFRIhgCMilPReq+n7njWgqXJIBr+IeWlphW+4k0rdVg3b
dQ14OAsgTZhWgO83/w9OKm+2EIzrl2S2VpD7EELsvijMv1zkTTsx8GUGJ/QBHe2izTXwN/ZMyiHe
+/aPs7a1zUq7F/ruWlFaV+gmJHAHzCoPxheKVO16Yffm8pQd2t3g1t7izbp8djd0lrVSXjJz05xY
Z8t3d43Pcm1/NcdUrEKnDNobRs9FJ8fAdAHb6hyqCb8ZDkf+P8JQvFyL2iXNo/vjDbUQxfAcZkN8
aSmAvZcn7of6YbJWY1ah/lcGxTPtFTXjpzsrzXHMN4P9/9WDccuFDOW+DHobDbfQZV4PNEgMX81T
XIBvFn9/4TVZU0W4xfMmUEriY9ju18Xg6En5dbVwCg+HsYmVzLwORGe571DyDsINxxaSJCNqTY7j
RT2FaHDCc43vZn8UmPEi0JYdoZ039TYERQK+U9P+BoyDy4pjEadR0FsYUugXY2LHIcYfa5jg5I7M
Bx/hccf1+92pETbacuEXJ3w1znI4iiU/wPrgCtwwapra7rDbod9wE//lGcILNLtOSfdrDNUJpI6A
41aWjpcKqrPqPl5CwbohJlFqp9CsNnCdzT9u6Ooy0QNSS4tomo3Qj8H1ax9Ta1d+kUlYLmDJWMP0
gRJyf9LaWO+XS1kwBs76ql74N6DZ4DeHXXPL+1gGzznnLQe3zZIJRnx6dSTFFUdUvflaju5JvoHt
0NzmBn3QTiav7R7J8kmzPEHu5Rpu/ek7+F40KisEBuP6W5svQvIFK3ABUibHi5bxxZ4J8dLviY+O
iMH/TnJISoLedVbRi7khNedPYdoK2eyBntX8WTZ0rvn/He3ryKKRh19BNImbmTBFRm6PASr6BWgV
MLNhTFkgBNOG589BKa4RhqosWdc5Mlu1A2dFJQBqKE/YtiI4gMGVWNeo+bzOOrjwlQt4aBHB8Oia
gQKcPJDW+LoYoCfNYq/dkjaubFpZfl+QevUNFhvRTKQQv4u+uzzel300q63OU6+WL1vAuXOIlnuT
bwp7HJJv9unHFLe76JczZVYp5MPankrgGQ0NNmO5A6asCBGOu7YnMu6fDGx8FpFkztC3QYTmeATe
ju1Rbdbvi64HCOykg0qsN+Sx+bR+fhgwTFfyrSjGalO30aDDQAuSCR0c0hd2P6citoT81UAvkqJz
YFoEJ/BR+tUurHMz1T98HQc1HmVocNQbTU2iTieSYMLmI0poVS71/x8Pn45Dhr2I+ca5TlWkiTFw
1Fhf1R+RA5jfS0aHQ+tWgdD6beRNaJjkDgdA2byLSGcg6Wfpczs8vMs5m4aDnrfPVv0OFnEQ3ocP
0+tNR3h6oOks+Vzs/5+e54SDDmvHdwZFyC1ogWGcO4BIEcoVW6APLIS91A7s7YiG95qbKKZXChN0
kH8MCXL4MH1lH67nvpI3i73m9fFYCkjxAY2q3yCINVU/iys0qZ+XqdXYHAS8/2IOaiQBr6GkbZ+I
7wJtgVfVye3995GEqhozDc3ZtJAeIv88d7OSaD8mWrW6tnQ7NmqCg7CGBz28hr4drhU4ao+aIU2x
W5ljjfedLlLJ8g4v/ccYBu0GK5oNKqtpTIaB8TP248o4Aa1EzCPRh/rfSQ6axWe0C7tCseorcr1F
Gna7TyjHXaE2jbK+KDUOjQgVkHTFqEJvbs2qoRxU2HG6iqFNc6R87nNsla6I3U+XqBT4XD69wWMa
MIXLJt62qxkCPhlMxsHf5kJLR79y3W7rrgp4iedgJNJbAhtvONSI9Ycc1CXAyEUfR60whVAkDW96
YTVKQ9k+4GMqhzT27sskivFktRNzN7VPWrDu76hCZoePIABkaOASp+5hTUk5hQB/xFFEqlSOAd81
eAssANS2O052F8kBRsSb0Xx15LjEJ5CuwTEGZrUefhOdNb1X0VCC3H4uV0j1uuNbPDxMsR/hkOZr
W985sL8/RhASq/2mmQoTlnX6lWsGu3EnnR4oYDLROyiFkwvZxs8gthAbaAPw/8pCkKtMO+7he3AQ
OCdZgmRP7IilaVKo+/gBvaNfRTM8fQc28JlAZujTqve5FBIVPyZE7bFlBskkt0O0ZTqX7YKu/V6p
cYXjOtL1QJhVOvIqRJaMwPeIbPfTYMkXADftaZmJPId/2nejnS4oWQ3JzbUaV69++rN3qo0eQeXa
iqFrs1+j4aiEZVGqkyDnds6uWTjEMUtepypBL2YeoVgtTgg9oxt0WDRPpHCO8HMWeTGrnWGkwRpP
O4FWhSc3w+MmFFhRuOYN/qfKE4va8dyPEixH1eV+WzZDFGabXoBxFmcApIs5dgaKCF34pGftopFp
34bPvikohY0QJfRm3s2tGqKMH+m6gVM36Q8vAs2VaaIYxWqnY9vxq8T+gGrt0gD8fk6EZp/WbgwE
W3PdnLH9N+iH9QtwU+xiHkQCZbTF4EeT0qGEJFHU1CDfVLSj5KK2k4PxDINdJB9dNa0b91/PobKn
Jq4fVUb1OHUVStzsfWjQuaHecp00TaJ/8EKayUEfE/Q4K0HKF6ONCJLa8qdotOOVt+0kG9SwfjMb
UlGQiit9bRHAzJmVJMCbsit1oaGsCXZghZcHSbsfNQFAQj80XjICFk78sGwo3WgftMJUhGPpd7i/
c32C0iqtIvTTfwVHLnOn8M7G6o2+gtZZwzL4IhecUQ9qVPAlHPxAiIaURMEbG1EbqmxkspdBJ0ZV
xFlxuegN9/hZ6ydKLxUCI6i4r3yen2/Oz4k22O1yxiu6wug72sXixnAX1kFYS0g3wjuVvAUADscq
fN33c0O1Y2RAlq7s5EfPMwD+yB6U6UdCdsOEQhCzaFOuW5I/mfgeryxWC8qNk8VqMcMfUE44p3BC
wmHEsTuFgrIQ6+iAHPNh2f3kNZ/W2cIDAFoYpXbo+KDxQMM0L/TeYQtC9oXztUQ3LXgC9vTKaTZ5
lag0mSAlLJLIp37+CLyeNA0gvG/b+EaoX8YGimeHDpxubz0vGAL/gyaPqD6NfyH8AQjutYDWPcfT
+Rnc9sEYVdA7E1tWkCuSpxbVGcSguxBvCQEA0R70g8QPM2FkO4757zdkaPMQJOGBG6nWuyzc8RmS
8TfpOAJswSxgWWQ5OkUPEr9eQd/q5nPHTMMn0kYsu0Rke6CVDkIKZJpJlsWIlRo9d/bntzF5Nis/
LFt2RBHf22mqQ8D22kiroX7yNJnXB83ZMKzIAMw9faImp4uXLIRcs7cYS3NonO2IIWFYf5jKAEKZ
xqYJUeTdHpGCEp9aFavVN6+rCvffcW5k2Ai/6iKro6syHg8OkJLPa5vYp3clLcQAQHYe1lW6UvJ4
zCMs/RbSZ3mZjSTrheNfV+0bHooSw9eO/u3IyKGSgZDpuPGGb63+BOyJ3kIniaUkr3te1dYI8P3w
0KhwXfGL/gM+ffvFHej/8usUDLUIwsZqGGb1zHmGyyS3UKaPOvG9KKLL347Uml/6k/q2moHXuYjK
8IZoecDiB4HPaiUvzkmsnSTOE+XdENNDVFqAimuMdOuhL0OkpWzgiiuUTlVx1d1dzJOEl6AzC0wj
0Hy56P18H45+E03R7kSoczK9CAfO920X8JmPTAJv4bl28hnXNjsVWU0FpglD9e268HCfVRuEwfY0
pZwK6Qupn4zMCBrKu5NlKM/06PCwqQx6jCwKRVhWRhWhYDca9s+23STOmUgfYVPFgKyHqB7dRN0H
LicbDdXoPaT2+8UJiGiZlpm+49a9/w1bejCdY7Zl8Ipz2mNLn1rQ9VehefOKwjxqvJYHlOZA/8p0
cJsUancMpZqXFkhwJBlCSx2A8Zc6Kbj15QSteQZqTzRWn/DuRa7FbkXc+e18gzftcmltWFNZIx4K
LarlgCSAg3IDY649gkjWm7YIK+eJ1QLzcDkSCENdN/cIkFzibB8EFuoyLt9NzHg6vLp9v5O3Ecyi
JEqsrQnSIHE/Ik4JeidTauFAJBJqN+YutPbTn9WRAHwlrIrdChD2UnPLq6Wkzu1IYNqgzS5C/FTf
9RFBc50ubUOAYDmnB075bIZbHAfM39O9TyiQ5bSj30VZnEIeQeT1pxvxFvSt9dlGB7k6dzz3LM8M
Cjbigd7fRdu8BGZSNdn+v/uuw/Qi2r+B9QHFRNuJ9cVEhyXxBtWcIcZwwswAYumj6ooaFWd7Mex/
mTLRo0MPuBd6s1r29XH3LgUN/3cLDQIPGzZwEgIummQ0XIm01VpBAZ04GlwmHzltVe4ow1nt6hCb
IzKtB5Zi0FozZTwMnVgeuGSoUkzCpXDQZmTl+SIJra19HQoyv4zzowvut9uxZ7kLOLBpA48X9BHo
Y5yR4Gu0j41nE176WleqJOx3nM7Bpo7gKCx2wr9V5pK03UO92Xqjfwy2AJ4tJ6rB/9Sr3yPlC0E6
Ia5fLs9H1nC/hwkg2Um8n/CfzYEa25bgmo79UOTpCtwsd7i2N++wpN6WHV3c4FperjwPuJAiFfuT
NpxGeVU5Ddm95WJw1gD1nGsDS3/mizgaXAA6nVqFwQqvjTRAj5l6wA+PGO50ijK2jaEGwMPycAtm
EHlRVvViWXa52LHVv9rHGro3B7vmoM3IP/ETcdsE4jmwSVJzYU1Y6Hwr3vQzU7wg+kJkZB11Ez71
zczN6yxdZonK8Cm84IAf3u+MeuiYQ0P8OtCmFyc36w1c4PJ3pWfb4IMY2FcBbYh24ciQXeuH1gjO
F9T54vowPCI4FPoQtxujFFhU/5xBmP77EyviCK1nhulhvVH532fq/Jk6VuZ/4PwDKGwp2FvYGRmN
FO7E1BJTqNnLLCZTDsit4yOgcYdk0Y6R+4mCMssaUORHvboYvNWiMltXbDA360LpyLSF4Fr4G7pz
ueam8b0FNQ14UOoFgC3JZx2t6qhct1z4XdExaEecTjbYFd5Ol+7mp4nyXohql/2qO4mvL7s+XMng
DX0AommdE/YGuknn1yEn8cp9rryUBL33w2epVIvuEGMEFqgJ2vc1CR3MCKV+lGJMlXtksVM58Uxj
KJSyVGCBYTd/GJbpz2UF7GrVUMuvOEaMSZNlCh7fBjmy2vnXaBtyex/jcs3xLLats43vrheO7KgD
RKEzwxfohZvJvQWjMiT5WLklTRyG+aHNVMtPIA8HEobSDSJobAWzjdiLqFRqSkQXl4sDDd4MyQW7
7wwV4JB0EWzWTjrMMaJGJPY4w3yKEI9J17a2cH5oQqthPF/FU88+hWlzfP8sSDI3AtmEoQiamRMw
5kh2so8m7KQ3uLZ2wSd/vfN5QZrJL3rhsaaUvpTjSZA+0WQTLObrJgN7xy0+ZDnuhFZ277B8WogY
CE+PrMOFyjgZQraSgetrnNvrqjCPd3dLMOGczmUFWP8WYSZ30w/XwpcZ+hf0iQCxneqRofqKOHjK
yyUWgY031+luxtvmOgjj8vNQtMI9pPmSGSjEtsHDSIeGmkI+zgYN7OOMm9bGgwNCifeHNi0/LkT3
3EB2gDcLvJE32eEVyXSRd7KmnVr9yaWfM+Jv0sUZajgg9t/fDov585naAempJKBl1zZJFCFWRTA9
YJc4yr2vHuOLAiAoWCt1teXiXMOluANNDwfPMGrcbk72YUAVoV8V3/aPFh3LwY6rYoPKYzuWwvpv
gUkdO7MeLTgIO183m2fneZ8zlIPQXTtkzUK5BNXYQPm/65nNEmijAQ4FtihwUKchbODhVl9Ql5Az
RmSTwOSXzoV1iM5lEQ3KEdhB8vOT07wHQ2E7kRcpfvs/4o9mhtK0bezWHoX0XZZTcaix7JY4gcF2
zhDI0NoY7+H0Lgg5vJc0g9efVis/tvEPijXhBtXn3lUQ/vKf4gy/rGFT61dkeMlCuAV6lduEfvY3
E6zRF/qsIvg4X1WBfBILiNp+2sJlLT13SS5hEWe9Q3zHN64yDd+2WUJVEjgv5Ky7X4+PrOTjQDs9
3SJjAeen0DP9SHlRK9CPonsOvwRzAhmZbVRK/9OmVCf7fXxPKTwDvcAPEXYvPEZwZqeuhDtG8jad
HCBKJuKJ+0XD2aWF/USVWrqgcXzhE+YzwBBuOymegZb0ZwQ8ItfYWUhHF0CPZvs5C7+Ue/jIeUme
puaBeGMQFcJjC0BJCAOylgrfww2CO+UxWLApl64+KmR8HNfmnsGjlW5x879MHuji3YPyJbZSTito
vkuggEC9D9XxfRZST86vssbe9oVOwRFJv6g92tv/bK3a0KKWwb8tokAvxKD6+VnI/GzvsCGvFeFI
XVScYmV7XapcSvDWV46FBL85e30fUIaEBRsqJdWSI2vHjyWLZrtYwZlBu4A7YCw8v14bGMWDqYij
oRYNbA5bcdBMdM9pZUxvfiNnVI1fzKaczgc8jUr3ydx3DYHvwHIFnI1t4ypaOauWPjFWvwwADvW4
P9o8RuavPS+0PkDOwKcJh+Um02QomH+OB5ies320/gYL51DnWjUngBgiFLW5BE7pDLQI8btLguez
4+qnVSGYuCiPVbQDg8yBgZTL+/Ks/EU3kFSZW4imKcTo/99uBuxx9ZT466j/lT/nap68sti3NneP
iXOx3VuBHRzFZnfbHn5V11SUEWEtcX1D9llCoQtEphuKWvG6RTHsQomjK61/WMwTDtSuY/AW9uC4
2/R/wiFIJ/CYG4fHWZ4Z+3YukJDfl4KKud++Jxqb40r/Eo4Zy4poHPBaLbKzui4hTmrBkJCQ2Xz1
f51MJl5S6dI471NS9Hrwqqgajg8KF0W87RP/3Xq9OhVD8DJ1eUc1v14ePjXFgkjm1vOoI38JxfFH
psx5AjrWiRy9gakYsiWPct8raDi9YAb/yV5BXLE0CCyX8/RYEX2j4XCJsnI4uLr7GNPc+gPDXORn
APbZVVHy0qCsvSnUP4dqWkFtiw+NWb0PMkPMqInq1IfzYo0/MPzMjNYD44IHvqD7sDHPXstTbgwI
+ZbdLVaeqQ+Ys1Ca+Gq5irfdk07aspC19rK4QQvfrk32jn55azCFmqucrHgCsQLa58qMvGxFGG/4
eUjAVrK4c/iBAxyRXN1gqj/zfSc0gZ5d28trxgEwwNUb2qYz5cKIm3aQjeLRkwM311B4n9J9Kgu8
FxdPSn3j4b8O9hKOtioP0iGnU9IQRiPrtswQWZgnrHEcV/PrpDCwyPoT4cgFbZTbe/nRjWkG2FPp
QjmUGg0LW3BM/VXXSBjVx75zViNIxhYJUzdROj+jNqWOo6vE8FhuwpUOCzWBkTEp32WIS9f4x8KZ
ZOxzBP/qoIK5vEGK6j10FVc8K61G9Ei/SdmL2dkdZ1bjedPT+9Z1y+T3xcKQaxnrdIyWdASm/B2K
h1GFVLYAAgjFyE60/KDMTGRH/+J+YG/Sz7dKz6DWwFKWOjUDgzEbiGFGrin+65P5pfU8NsvANJI4
XyolFPERpZV1u2xEbpxobT/vpjSehf6Uq2G3h7cjV6xP533JQLVjxkL7dt5CqdSGQY34YewQ1bZp
6dseOuSj92ZATDpmpe/H6ffyNWb8WdoBg7Zmywi9wEa1vj4rXGPKIubrSrgpmXHkaCzOdzxNId4r
8LAW+Ta/xm4XmQnBaf0yU9QqfXAwWWaM+ZE39eFxJSJwSA6m4lU55Ffc+TXQWIYVfQGu5VOdJ0x/
eXf5nF6g5A2oEpakp1FFnVl5oPWgCrbd9friRynRIdn8cJay/MU7cGKQyt5nYLG4NCg9N5TvESXr
TP6BxCb79q5qnkERO8jJ03iKB/VNJKywcRmBhcrRzRhjNwjpwm4BkwTd6dNIAk3t7cRIj4r7au7a
LETudA2eVkbL06EpkMK6xccUc9PDLN7yq9HDoWvzB+OYz1aOgKqlmWbbMBoEDOTJLSSXXJYhCyfL
Y3Bg6lssSom7QWNT1cpfnX0PJQnh98BYnKBVP1zjCYU1Z3eKyMe72gUI8waKmQqyVuKPkJO5ktqz
VKecSz7aDAik415Jx3Oswm87ea6qDjmqdPwzBF0smQRgaMC/IFQTXhdWbsOx/PmdJlNliuyq6qNh
CDgQmSzBeQRsIWE9IllhgNPpYLwNpGDHJ3I7SH2IEqaks8A+IVlAFzImiHZtTeW8rj35v0e5eWq2
lyyDzAjc0aDbTG4U9vGVuAByt3/xJIYDxFuQWJMfaJLgtfE/BuiFinoFAGX7xhJjqUIQUmOR0qy3
FRmSkZtkXy7cJZTMAlyl+s8bcDEu64RyvxtwlYTgVcJ+ZS98k8GsatKe1VeHpVjn4rWbVK3T8v4G
R7AsaLJwgaQv27a5W5QOmdPZocYI/IUDvW1QDci0k2no+0GVJ7KB9ysnBkThqN0Jsi9U/kDv0KCR
eceErai8/hUovgDi7jtp8zMqFq8v2pdyiOJ+XlQI+j7Zj+2NwR2CdUPvXG/z27yF5SvSyLpgcWcK
EjNhNYaTOmCHljZReWLKIdWYbw4SveUe/WvssPR7w5nmgx3qMUsNu5kGcX4OmMGN84Wbx9KdEwqh
WRAK4TmX33g5xlQQYtCWhBeKtekX7emlAqPoKFomTXhMFPuQ1u+jXqMfAzps4o5Mgy4fu2qgt/mM
ZHe12JoJd2IITnhL6erBAa3BEVuOYeBI+d296L4tfZxBDsSAoYeCECM/OB7YQd86ZukjTHQAOKwA
d+Qf/fcToHtI029Rcb0QeXVf/s7SAl9gKjAv8Us6D8lzTKcZHUUmbegd7+AiTCAhwzYQPqGl/0lp
fZJTclN/lmo98/YaI7JLZxALlH5uchfFPVjCII+lpBLcs2f1niLhK/pSBT5W1Miiq0S06TF+spEX
ibE5+EOM/Dgpz8glGGmOO4FgYP+A5FcmxSAcUOg2pDzO/krGkrZVORfVTL/jDAL9iHxJk/rCNH2S
tdMFyh7ZfDpARoG30Ii+C6CPYc7BWpsX6X41Y33MOCogsCBbBQnhTVisP1H7abDjPZWTBhnRPIEK
e2wJD0PFkgwMiMlOmg2k/Yi98Io0Sqcqv0Mj5rQxZy/xiP6+AG3JybltULR7mmznF/YcgNmmWtv9
Op/IpI7m7exAPTa/vOMUU7brbJ6Ty2D5PepFzbdF8SynAsc1PEGX68ckqCOYvew39GhnDDAk7p0C
VDkfWiHHwgE/0nXtmdHK/Iu+7oUJhn9JXlvsgpFMTSGinspukyXujorEpdCNmnyTZODlcm1FgQg9
udQfRFMQQynYlJl9IdGp94XPx5bQPL6YBkiZoJi4PrqhFVmlUwN9zgGLNUCeVD+XoY9smFikZtBU
lvuBgkPbE2ge+f3M3p/8Joe8w4BY2qXlsvMAa4WLpLfc2opdwKZOm9w13pYjaCJEDtKDN0SOa8Kx
NkrNKL/NvyatSjWBUhQbyr0Pv1aJ//97JehZIWs7WA1F4Uq++Qr6EdDccX6b0hmNa2kFvXtneeTt
yaNlOxrbDB/r3WUO96iF9ZA5jfgKMD/EfJgNGM2OdX7E0GWwpGgIKhagvNWGhGHUPeflCQHALkJk
nl/zWL6l6p0Tva0W/ztzOsGNIYs2PXF/qrPSns1hglGzwFCyq9sjZonnUVBLNxu86pKZ3uRQH0o/
sWeJKUVbMsx72ebEC6E/ZT0OY7ewmkIXImLCX3Q0tv1ipTHHgr23Zd53bJhJxR1hyDQ/sUsemrNF
JR382/8HyYcJq8NsrMOdXiH+XpFg3ehTgKumx7naBukMOmxlCaVCfAk+g8OZrmGxy+uYl/RtzWRc
eZjvidzWbGQi90XvYUq8PMK6OCZ91e8Qt+nBBeLIonBhwwEAHsEUap2hzrS3T4WuRkjcsaiztXvu
fRrf7gsjMHbzF/38cfkHDDVKbaHy5ls2ZX6BoW//nQtjCtEvO3zIG7TmFokZOT20Px150fHhBMxH
9Y3WA1qBJ3twRmd9vNFTQAAXM5sa8ZCNUcIVkWpMLoIIYzVu30LuURpBuTz6PPHl1OgJkfNN5mHj
bvl0H+QOqiB74UUrEa/tJ97J7qlvKb2cDvl3H9BBvs7iQ7G778iVJYhBMKGDEc3ULJgkFuVm/1Pm
+evoIGzMx6p93D1DM7tXmJ7h/pTOBoCjM1Y2E8AG9JweYucpRqAI5wwpKDxpC0oM/rY7aHl1Ixvb
VNFicDHLwsoEgicNYp/h5fpfdc8a3+LX8gW8nAmaYdgziFhfh4gk1Y8cTNqmr/z2aLyK2C6WFk1b
lvsns9VoqqFxhEvFH+gSuHYzU8na4dTB3wOFYaMoUAEucIhvGtS2OGZlhV0XvqEw65yP2yH19VqJ
MLwEv8cQRZghtk5lApShwHYl0WBDXgWgjX5hoavLdKJPlslzVeKGyfUTYty39bvS1WFY3G9GYNHI
jzc8VqGmbiw5+jjDw+LgWqLv1FNcG1g414ypASbJ/aY8IGH/VGrafoZRg3jvOoaZJHlVmMvjlaqe
3YRUvGjs1DlBzjK6UPk+rlqU51Vj39C5lsvF59f9E+VQsaPiMTMDThpaT0QCXuCdnAk4HBpPkDoc
kLNYN+yKtImKZwczwl9FiFHs19Zp6beeDmgTJ7oQQXqzjJDoPWojGdaoRo8M2ZjZFp9Y4iGdGL9m
yBAUXo6Y9SszqtbTXJo2A4GvpNhFRDwnaO3YpfivPvcjLWTE99LKTfwHbfCB7XtMFtE6UXvnhc0S
ET3IcOsrHrDljIfNRx/vZXSSyekRNipUA6OYhVjURc4AlZstUft3Rym3/3l19RJjviCstQ7i7hS/
fHq8eemf359MEgX9UvN88iU8f+9HbuWNQmL88lnlqed/qKqccx7sp4q2F3IZfeMYFQIBVjYU1+dR
CjdmwhJR7nJcbe0LjrQUSwhg2OXrDig8SWeOwO+/QeiIwXryONorWOogxILmQuDdkyVOO787cLQ8
KH9tcFGFpm+52lBh/C9HTsdcwxtGDZf6mhAsYbLiSxGtXUjQFrFlTey8J+MUzYd7r8HXTBPC5HTM
B0dCaNFQqSD2V0h3TTy3OqYTmd11DTFbAsIXwRR5yO79VHpfu/yfiN/A5RIE4JRj8C2RlbxYyhRZ
foqXXbebQLAxaT6ovUJhhnPuELR+qFPI/PpzMhUQ9f1AALD3H5WYfCKjFUYLWn0VfYBuJXyOQNDX
E9dYOV098lOtxnxwHgv5h/KYwbuGs3m6kOxDxE/tLUl25SvgaF21xk0hO609Qr9SH2wg3Om4uPZA
t6s/kdIp6cJsACZMFVuGWOgYk8P4gUJcdN0bXOgVyq5XXraMc2jtuFnKhQw8ubCdo2LsNMNjSyQ8
9zipjyDvNrVuPIUuebD49tu7ArKIJrAE+hjsr1kSWMdJQSxpbUeJzkfq/maoBC6F/TJmWYwR0yOr
55h7DC95c0NVNCQ74Vo9fiuUQS8Ot3zyU24Karryf8A9gEtDBC1cr9NnD122n/5R34geGupIApFF
AZau8tEQKoI2FxIsbGuH0QtK2A0P4DwN4CkTVYiB27+kiNBT1L4PwuHQmUtkAx4uhKuBhlnmcNjr
Q3oszHIm6enNfLD2FMHEKCI2jfbXqXam9VLLZYntRYwnWWHcZaTg0OX7JOfC0fy93L7mQTfaZfm5
1WeBg5LZzTS/dQdbY5mTuYM+pfMaf9ks2A3L/S7rNXG/YQ5Q6lYy0wcfOg3X3Y3O3ldfO0hVvDxU
i7/h+EluvYTcuS0cbasZW9ih+5NhosHDgd1nhiRb8p2fOCdbNMO1k78zww6yPbOJviuUVmhqrF3k
CQd/h6u6i8EdJWXnxSvkYzKFeGO84YdyJJnrq0xUiM0+sIBQh5zHZipWgXgxOW7ES/T6vmFo2vxr
BdN52mW2mEAHZW+rvZsXoydx8j+ZcR0UB78J+laimbvVKtJ0V08Ah1457T+5T6VTklpvcczTKZt3
xcY3YUwAvNGR4VpdeQtlSVYRDmwqSLdalAtfgaikn0B1uWJKD4MGpNdcjCnk0lCL9nfDGLobB5J1
BcAZXsbuq8yWMiTbX3zOjq5nYSt3yXBSunlwgZulLWrRpwSWGjbnto/6DcVsa/DTPVzEQg1nGc/N
XOTEkksnoLZxhHqapRnVVGHRrhzz5jukjgzeM2GdWsDU83oSVOy2HNe2LSKQA3fMqgucfbtF1/kY
RXWQeBKGI7UAc3SJ/Al8mPKDqwpx9SI9VIoOjNen5QFHN8pGjxvVDy0wAwG9JaHTKW3s3IHZipMU
dPOs+9HyH0M+1spbS101YNFeECMbcRqYbMM55fyqIBXr9JfMYlvKY90fTmqKXqjkkSbNjnW7LE93
VNHh2gZYzkII3xEv6mqVrNZn/sm8A+LbafbO2KH8hKVDWdGT3ZlHHyq0JYfdbblSTHcXT294zpAt
MOjftgdDKoSNBYpRDRltPmJtdxKn/zfU1pj1EDaVT1HYlDMn8uPuCVgErwNewtpGFoL3vkNN5Rgy
AMF4ukWna4c1DO2ZZ/vVHZvxOK5f/BINYQwEgN3vGjG85iurKfhpjGXrKoD+yzDsQOls86EugsxE
NImP+NTecsxybkgJjuFVJfEDgS5tyIYxidKFPSSd3grlMHSZscj3A5TdY8oFMRK6PkoPjlltxSz+
/DllGCYcngriWE35yvhif+BFqP36+uEnin9hm2ephzOu/4Z+2iX03Nf8vcGxfFvqUnpsuWlYa0Lt
MC4yMDOphC5cWufUMGmmqGX+1aGKzb9qYcOMXfJnIdqf1+jzY10XgomZzT0h1/xbCs7vvFNaxFm5
Bfgp4BEm4ZavsBbzd4mIbkRmQmPpwCMG4zpqVRFxuRcg6EdTm63KEjDCuNQb5/70SyOs1KNhOjjf
EUOirD9uZDI8Mnal4CF9BeeylTEO91rNLs7Fuvbvpdja0QBRJ3M3Xu5Hpt1ReOAmhYqt3rfN6YNv
TEEta3a1L0fME56zGRm3OuDMb5KTFb3MVBn+AI5mFqQx/JoS7jb61UgDTPgKl0lFMcAubGWPRH9a
vRMPJRUhFt4700dov5mGUge4/uC/Loz9tHFSwQzdBKCeIsGkdBgQU7KfHj3yJGOGUX4NFvk8Hesr
Yz+F0udzvOgxKZu/7yHR/sQ/kHzGV9oChlBj0vg7ibv7IElFOmrMihMn3uptM7HF7JO6E3C6pA2W
QgINrcGyhLZt8E9Y41SAhZjvWbzeKVGex/kKSwJlL0VANMjZRFdy5Eft9dye0kNXefz01mG+pO+l
NRif80I2FVuipXN14b/IyVi3+gn+CN4u3b48AvbGyUYUwBVwu+RC/I3s9473xwJTWnAIrVTpQ0bt
ErId/mC211/oxnN7jAOKhPr4uO/stidkF7Zoh75yhQqUW+T48oVb5lg85rnjlIEikoO8eSAH9iF6
hQGmRMruwuOUT7Y9xv3tHwXxnYmrviu8uoaSSiXPM0hBU/JBVIU28DyTiv34ppV8SMKrY4GnzExj
AK9zyJg+BIs7Sw31FkGaEV9BdCcE7jPG1qyW9WpMDAB78CUc4IEVYU8lo6PsYJVvGMqRmG2eueqk
IISo0tU2XNDIJ45+Ewulz42iH05y/6NfAtG97RNnpVWiATHeviZQih16gKY16h1hRR7g4uAYZD3f
CjVrbKL8rwfSwNgGNIZQ7SKX61lROeGjg3iCINxMdW0hz0Db0iHbcCwfkYSnKqc7wILGFESQ2hAn
ZbGvrv6A6AjErwry/iOotmzDSXPwn2w5aas0JG2WmV+AjlyDc1GbvW7TeuCkzrZNiNdqYT++xhCf
a5BJRcHNO3t1faZ13LT4DAnkiLtvYegPSndTuK3+NC+i+6nft10QAgg3Iy46Y67XxvVlY1D8EB4e
LfaiixTVyT3UthWT40TQNMhk/uuNPygq9RfY2UDEt3EyZgXozQvT7G1QWYuFVxSTvYFqVZ5qAe5q
jptBtx4idiFzT4/hPZaK6eDBZsesFoOFgq5PgnYzCxhdyb7dCGtX07rw+BpA7fpWue5W0Wb4npjl
wGmxSJIf+rlDISofCHkc9RV4UCs3Myu72zLaw6elS1HpTqG9AaaQ//1j9pmLh1r+ws9Zz6AvC35u
UVdhld0UddPY+R2Q/rOyq0N/P0jevqgnJg+TgSqDQYaejnSDk/Yur/yV50/+Q978ijuk+bMWIIjb
bZlWYWmt6pI6WXx/uhw+1/QN6Uql5w4LsHNv/UqneN5SBDMO5P89BHPfCG1Vhh4ulL0ZbnfsTcqT
kva6YVBV9+IwqJ4V+bWv35yPw+3jXqB2IOHBFkTq1CmpIGMkF1FGScoPnr9haP0MXnzE9WlE3qsi
5fSDzWApEuM3grhK8Seun16vsTg0TWfIyQ8oIMEXjc6eF77/TsDu4WW8OxOJJoYBSw2ppXOFFZbu
kfJjzoBG6NVGvVatZ22jK7QvZs2z6RmcVpcfBGu1aPe4aTMhujBeTNuXq+na3X3q65nORzlaHMFc
bCkmlPyPcR3O62yuNQLM/6WLZFtewwikDiHIipPP1OLI5fu+xw7DIDeOehk0jeuuUrht2Qo4DpJ3
418gajef0iwcbmYkya2nr4haQPiYMd8gVy3dPEurwEel8z+Mo1EGsoOYiejd2px4cG3hFgYor24a
3jdp66jE2eklUqvb54HEFpUZ9F3kLKE2oDrPb9toZeztq1IgxMU0FU9wwjDz7dFlkbz8C/jCQKEs
O/zEwLShcgPAOKas+74uX2lCBIG4gT3/Gv32JFOsbiwMeSBj9e/652CAAt6OA1zzHlCZ2yWj0XUR
wIG3KhBFXgAry9GvuJPTzjarQBFCz4lQRfAgCq9GZwrTc6h0QrJpum31/IbOCNjFGLb6CNVjyk17
lqkueGkMcrB2p3QKihlFcFHqlK9WhnwQjwtm0wj7EoUP5pTY5ZnTyPzrzG4C9/DW0W33pYuv4SdB
W9NxdTUnSk5w8jbQ3lsfLhHBuKzJIdpSAKDcnv++tCeb9KZrNlqDglSG7CpFpnvNIHmS1prs+VYy
o71AC1j2+wvXuVrI+duX9aYGPRMZM1v4GEIbAlR4G6V7SIP6yUjcBsO5lshYq8hy6hKL6CE62oXo
XUhqX4gjz0O5Fj3Mk5wUGwMIpiaF6gZgG137KeRa3fa4Sd7LXlRKpN+56+y+UQRs32fXRiwGLnx1
Qk/qhATrvEqA5gt5bU3vBAJsgmo/UvOvrKmlOnMV7n+z0lEyTTJZcxiHWhQvfqhdkDCLWxfkK/Uo
hr9q3hDmo0BBZ/cly6j8j53qQ8aYvalmNmOouyFC7WDjiieIND8sxV5yjI56Ew7JTsVA2UNsMa0x
8Gg+U78Fn8+4hVu2N3y+snhPnO7tY2lx6mnSEj6PLNba0upDLaxRiQ/yjvDxgIw6WyfrSiGliwix
mG+LImGruzhrjbYH5bH3OYG+1pnSJb2Nos85pxnViialQdZKD5l6+SynxGSQBOPf+WSQkmGT5Yqg
2GpTVCNbvp06khaz/sBYmj5X/OMYwndpfbuMvTZctjAYqPFUWdIL7k952a3cDsiE6hlRY4RXAVlF
GEv0jq3Wlpu1JyPuYcK1cSFnwxOODSRjqqysBhba1rAyfo7ixELhShw6pQ0lagmG6okbNz93Kl/h
qpais+lkS7Gh6PHgyudagg6dOjtPiYGFrYZYyT/2fqAwSJBlWo7NF7UMc7OjArrYGhWKcd8rf2du
bfQRaMyMX28XWruK51zCu/TLpS7ONY6j3NoGs1pHOl8CHg09kaJTae8UvaSyfOVNF6d8qd5TOTrL
RJnbF+oKK+BME6ux1OqsUgLOLF20LUwNpLBZ4C7ZeS+EkkUMZ8iJKA4mvXTImNQlGrutAFjKAP45
G+/no3DeO2AiZYuDwZwkwOq86bQIzLnb+hKvOEiY99X/hzJ2JFThmLZIt2NmwSVWyXmaC138IrDW
hQXUF9lBNCeZvNOfiNOgY7G5Op7APUpvhsyGp8TK1CfN5QDcSk2uP7ulGsoBbaUyxxYoIsC0WGuS
DJcs/rht/6l+L//QU9ULIzFXLN1sBFkPxjBvM9CXM4ND79j9nFpnp2Bz2+TaHOu31VbrdWmscq6N
UmmkDiJiOVZq2RvIArpp/48W5bQUgupPROYxQg6BXAaTd401mbDBv2DiPVylo6vHDZYaiWOKnZ6K
Txqx6eI2Umh9ovcD8/Mb1OVGmQfruz/5h059rXO2cOfEA/VASrN0vtaZ1yanZ69DbpsOJ1j0tJRT
+aQGvpZZ5PeGK0X0fjfqYzsf6vOld5yVCLDEuQTlOxRBHcKgoGB7+4B+NOsGrv2H4naJ9NIabMRf
J3cu6x0ZgcM4XMHADRISpPq+IJ7Y7q6bUWkLgkcRvIrynKj6OjB0xhFt/2MaFQ7F5uT3ir91HLPc
4ENaa1meHnofRgiQSDA5XI9G5msCxccfTMf4fnMZu8nybFlPKR6LfTJxFKXOnsWCb+1R4wngjxke
RnwAMKPI0pNmm/rh1ydmEeRFNjcJQ9NFzgjAMrceWn5nijwmAltlBbliWXhSlnnjKHVXCwoCiJPt
msBhkNTCpJwfBD7tOlkUQuvab6+Zpo5m0bb+0QYbAHK7b7+Xyzdp4VxUW/DFVJocCHhdDaTxHVYY
qnm1vCGYzkV4H1L5poTmqHWgpXK9yqyp2hPtZ1pPLPTuTP/F7TTKARgYhDL+ZSTRTICJrcKHuNYj
Cmr0qjlCryggCXDYHWmL/pbIeBh5XhR8RDz2XUHzVj1jrK/XnVoH6wl09Ug7cKIFF6FfU8dyHa0v
/cUJJVvYXOqrI/ggvOh7I4PGJovj9uoA6HzqtnG0gBZlZ1bgVE7MnyUZJn84bz/jdmOdvUd4rSCE
XxN77en+5xRdBDvNNfJXnLcvUHRbU83WbiprdZeNaRwvFRrMvGVyHZOVzzqOE7fr3elToEURAYaE
9QU/gRjbOsukqHVJX1RZ9fJ73g9/fLVY5Rkm3riT4xrVRqVMXeX4BLePGN4RcKAe+KK3wDtas1rH
EO6Nx/+RYb2Nob1KwvkDZCRJNEgfCsLT51Lo5I4BTd6rInd3sEwggS+7g4A8OsPBJA7BJrhC1en4
+0Kg53Xa1IyKf0n/fzAJVGC2vVE6S6oMqowG4J2UjT3WiWKYaPtCJPZn7u7BFjAS+Lp20QcXOonY
/i88xhBTxJZhP7Y7YZX7xHuzXHHtw+pcmNMpVhr6p5HgFm3wJBL5jb/QsQj0AGt8zdBUSpqsrSIr
MaUoSEmBKViKTnGDKalanBA9HYPXMDofuIsajDqnQsh+YatIxE/J04MHLego84lbKB4gkkvOb5BJ
Ov+WeLOmz9RBpV8+h7qfKD7Z9EYL5eSa5LIFUrv6C7Il7jaySMeq7Hctjkct08fDD4Mx2z4DpbLH
nFC6rjtG2e+v/YMKFD3+OLq/e6h0pRu/zA0HJBNBLiGcLZtY5VcsCzfRH/4VvBY9SyNpeEDU0uHa
+A9gfwjzjOKzuYd4auD5DpBOOHvMa5MiudHSiBE2P8RpV0FcsDQUSfhx0BWVVHk6EPH0xTvc446H
xrQ7wY+idui6LL0T/v5b2LvBoTudyZmmLtMnPNvzuI43lE7Nlm1ck2L8aFTY06ocsAhMQbijzxpo
nvjP2GQKsmChDfSdSCDRL7tAF6YqRpwipGuBIjbLOdFELR3TF5WRf4PKB6cYzHPEa9VwRIoSo47Z
jJJCdAL1QyK+94dspr6roK3uD/ZkJYUdh3kDgz1aOLCNxBK0LrV2RB8NLdB2LXMBonSPEG368B0B
KNOcqB8HIzuQQQ98CN86yzo+sDczC3fWDW4WRCLN1oELEXlDoiS1NH3o7BQlgiWlllQIZ3rsJWB7
lN1os+KWbVhGcDKqcnsw5OCZ/kR2RmJQODVz93grznIbEDK5zQkIiHXkH5fQPzZ6vV+JrD4f9TYw
imJ6Ct1b2KsN8qh8oWVuwTm8WNBeooKQsPmo4dE9i+ctjQDme4H8/PleEm+6xQ05ZgmYkacCQaFi
QqRuDI3kMzBXistgr4F2d9Xpq38C/PkORnBEoZ3G0eFoBDDpv+4LL7kBLObw4Tmlj0ORt9QebISt
HlmOOXiXlpu4HVFpv2SVZKKCJGmOcg+s2ohB/i3nmRwKIHcGf99+Q5kcduJVUwhhZcwWfzvEUOVa
4bPooueE4zb/eTjIEiTE7PyF0KJ4v/HT5V5eCD7Yy5njAJ/QRDQotGTSCWmbZCNVpdW9xqH44h8w
tQPg7t5GwFUfVfY1EIH5jA1PRnTXRGFLIlsft5ajRJiNBgc3HdWVOf83VK/hjRZ7ZX2lb0SbUT8h
EjJ8eyHC+43zvsFC8X2oyex2pO71ZUPZ59ZRQonHnMex3H2/gRrfB4NNxhZdGrs3kwYPAQA0X2LO
ARA8ktrN0xvBOEK605tbP6sgwI5d3vHb0m6t6yn8ppkSWbUJMxEBlYtM1D9wK0y4ML/R+VEVxO3B
xdbwxj40Pk9SbyCqNanakMDZ4+eatsjdGOC46KRbkRc7Pw2/DEc4UgAusfWo0SU82ldMmLo9aFk/
mt8rClXD7WDPVvUuvqo0xFC7WzQ4bcxZTwN2KrGhDnh1GNKo59jSKDVUJQTm+vH4u+ARcSESt/mD
8B20MD2RdD7jD5RlAPmbQTUFnGslBLEVSD4KE+3G9kjv65g9bDLKG0qfyWD+x8JBm+tRNMEIWOSo
4OlYDqMqn9keyRB8BpyARyBW9qgxoNZvJJTnlwD+3xYcxXEWsj4jBhfrsIEYmSpYm4qvBoNNjw2o
mUOUCtHXPgO/rj0scWD+QJmXMHUMEbyokJPmT1bUoJ/RtgicAHEJTtJeH5rGuYqlIutWn7Im52Ws
CXnLzqBo5jdAUInekEoDYZmeMMW00VZWeW0ct/9EInmIkthsmI6gMhFd4K8bOq3LjzA6el9c1p57
bJuAtsh0BeCaes6FO9ikEjneThI86IZkP/RGoUX5thP2yxWAvkgkjyveVIUt5ZKkLDIaQBBfUtSS
TKzT1DySNfhxg8zbVwvApKaWCADeByKZnPU4bVcSUYlZ1lQmVogiSkObrA5DsEZvf/6kPphacyM0
lnxpKvIZlfubPKhBlOuUhmyyk6og3DwvG30ct51B2xNrHOL7OpgvK6l1r2L7owLZG2D2K6RdASH0
hOEcghqxvLkI4K33xbG4MShtIH99u6tXfLtYtS+Mw8sdTs6IWTdArRUkaz9PuAPiUToeaCybhI7Z
JOib9zhcd0dyYqqo8qbWxMMvwpN5mlPwBti34ptBbPU77BN6r/ifx2Fbwhy5Btt1VMhXjZKmhVXk
LvJgHRAemJkH2yJWG4GoDcOPzNxNTsjG3jDez6ut2IxuQcP0qj6kz08PqXYb/OzzGkjm/FgBg4jq
Qz29q2zP1kaCV7PgZ9QUix4oSh0eYMz1SsQwn8GDv5Zwu/sOAHrgZivhwiJE3Xflni2U/NfrYDA0
bmekvqPtDPyFgdSdtecxxhj0ULg0oBQnYgbe8w6nwKdOxhzFDIdduG/E1H040SQCP7NL4nJfPECh
/RYJ4y2kMN7SkGqLsMkqofGkl/nYbz9vRTd2i5WcdGGYBUXS0LW6tv6DJcKJmaLRDqw5XjqrcgsE
TwpAOeM7IHbhP3n2KU6iZpLwsn+YIpJznCHJoXIrWZ+Spq5Ufz2PQNhbLY5w9/opU1pSAQqexyDg
SI5+4mpql2b/k+Fe1pIe60YhTRUOnCnRRdzv0C79A5kQXgdM0dub+xtD9NkwBPo68j5/B/daB1Ks
VhNtvk0oVD6rpmD67LR54wtZ0zR5IWUQqvtNwsWghnuxfVFEn1FTHYwSRGKtIMxdcvPf7gPPMLYC
6qgN1aD2sW2HPftlAiKfJrOweb5j0b6GnD8WAwWL6wFuJxxuqU01MN9EnWq8XW9Mf998qJXgb4H7
a7FysrGxrJ5TGe35sAS5wVIytExIADIEGSvRXdQEjg2ayCC3HXal5rknvFx3fiFjzKf9DjN2GDe0
r1T8zo684Ep/1u80qbEhoTGcqNoZb+EmclQMcbE0544daw5E/HZx3L+VJIpEC8hoK2S3lMPUOjaU
OKD+5NbzeRTp/u8AeFhF5Yh7WFEXPuSGThicFT1paFi8ViuaIKCIFmqZELKLKAtH7ns3AiH7lsrK
WQ9+oplWj/PGjJjoywa8OTXS9G4+gTl+Apt3ypMrBfHxvWN6Jl23CzNY8N6AagzO1jtewgMqgNSu
tksF4Z5kFc2ZUUjSPlT1HuUNL7lod1CL0E/PfAa4Jc5/zSfqa0NDG/pVSwrMVo4tj64Jn2hRgWLb
IaQnHvD/NJpLxpMMhVvcGii3tWfm8vlcb/7jczQviZaljNlHb7VuYK2Ma6RTR2A4zwKyaQtfDpCO
QxmppzUE0lLKkOxXXhbqroIbinmrqDH7JGSWyRkAVzjphhgMOTRbNxUkKryB6irPa8aaTRIRgcK5
+qIFkFGf3YUzDeG9qdGj/DLIjtIKIRJMHrytwo617X+4Tf+w8+vBo6ekIgNBWq/aONZU9ZwsDBQ8
14g/oAiKOriBWkU7ip0uzy7cVY0nUynuwj/6fK/t5GLjUZ68ZDLHK7Co+KzJL0nxF0xuUz4dq7c9
ZgsR8yGkjgtq8Hon+u+oO9PBYhZEFdywibrv6upTepfLLqjNP+lg+HCjvn9t91KJL/iYrkKMpD+5
RgnvW9Oq47nPNqrVPayVJGhf3VLpQXqjmuTdCHp9iigAdlOl+PBvPghRdg0z25wNAAS4IDxugeHv
LurFXio57Op7LjnAGTa4mDjQcUevejg7G+nxYYv0XCU6g2Pbbp/gXU8JEhec29iTIGmQkiOOSi0n
P2UeWKy4RROUK14dBSy7K4K13vQ9ds5fHn612NUVKgfnckJW65r4GvURCtV4K6v4DjD1tJkG7XOO
x+eKnYReVgRoaViy5xBd5AWGDKPCeJrEVXoWVmsq2ylGdFJAoScr+Bulsuy8xeSIOvKk+aUJNlFR
5Gh3AkfOw6Gez12ea6GaBBAB34DwC83H7Q02abkTAYoyGW5sI70jGQ/fk8z12kZ3KUtx2oxpSZ6O
mVOv0p98+peFk+Fz9da34DRpB1jWW0g4Xu1YXjgq8TG4jOC9nAWQ5zoOgmS/V1fi1CPOTykCR48a
Z46yyiqGJq9BkGtJO+77zPej1Un97cL7FkvR5lieYqn+a5WxOx7eHkSzfNzoEVey/feT0FGEcu5v
cngS78GAwFo3nlca67n4KpP2IDLPoaAQ9fxaiWiKKGlQ1ZPW4QCRQiqZFLcR8/1o/SDxbYuPWcBX
QGGvfrNK6qYsRvr7zEYLuwF3AOnHbe7BDnvo+x1ATvQgSxnnfdqLa9oU94bHAJqp1SE6BeZ6yYUb
mBQWcHH3n/YNCCgesyAIGMjMU11FSZ3NeU2DygEaZlJvtJ2AZZG88Kp0SGkFgAdyrXMT0eng3GAJ
9yraD95o7IjzIJHnFfYYo50nCqSarREbPLcZwN/CXLPW3A+yPSrivoXNR8JyKWefQUC1IIQHHBQ/
T3wnzLcqp5mucrZqxO69z4VeuQOTxQd6emgXz7qJ8BXC5Vy2ZC8CGJvMy/iOt0eJO8uQAovRiQfE
FAuYGGnrPSqxHmX0th/VTCcyAzI1UdNS1p51XUwJ/1ROQlE9KutQR/CWnQGy1dYKPfJmYxtLolmZ
Ibpvnl/EP6hYWY43GP5B5k1ipPZEF7FnD8pEYniffARKgJUuLtRSPtjHbSvsysYxQElrRr82ljKm
ow3WBKo8exCU5cvaTyhlXRP8vDKQR5TqLp7owATinvJLfH4zjBhPkHLuRKHlcE0+edcQTlCy4RaP
TeV5oSaqvWL/HhB4nbr0Kg7DT2mls0yzGx3pMAiLyiFZ/NUHJ9XPpjNUNbUKUQOWrfKtyG3FJaFy
aIDjpjjklEQ6Q7axS16xuVNgK1WK+3URyQHJOOo9hkSf5Z+eC2qoAqfGnjWS4skCHOH+lkStyL8e
C5zQK7kbrTcLRsWNfZPBY3JLXFWrHmippQRKILZk4/lgS4CFayIg75aGoVd/G7BvU/bViasACuMQ
993RCMzJZ4xa2dYPbBt5MavI7BOq92Kqd2BBKxT4n16LUujN6W4+7IJmB2MJR2wuNLS5utb5dZUc
GtWsECMwkHnlYrPIhpvBRi1nYIDTKI17NwLPEdqWAK+XM4lye0o8zyiDunOsz2ziczKPqTJSpe/X
5xcG2m4IU65yhanHpJq6zawoKAJhM36ZgqtVO70CSCxpyBYMjU77rXoXv6qA92pBJg5gm+OTN9jI
1sJGZpLMULwEyFS+DbBehNUKeeY3BdxOYVXW2PTmvN+kg7VJbFw/Y2eKnXCYGR59+ZLwyp1Atr/j
U1ouIyjWJTGztE7OYhwcySwUIveVHC85yCOnb2icg5Mzda8reIJsmmZXvU4lAABL7p3/2aZ675XX
/YhHio2zxWMc2f8a/vwUR/CfahywMbJ6gF//5lxktl5TMdZ3lR9nZxi1EKRdNFOsqZCkLJqCAxKJ
xjnji4NnSMA9hdFOvD3Z3Ej+4oSu69vwE2qCaGCFKoQma+pSuapRCjshcvjgaSRAHKSu91uFRVXr
KOh4JltEuDXev+1/SCzzRoiBZgvAPkollIWFxV8sYW+pHb2LPxajIeb6Z4TmICZ+7gll0iEx6l/W
ANwwH+HklBHjMS+e54bcPurBQfbTqZEFMhYAmPCYsh8hC3M9ThvM21xa9OIWqQWwhgjPugevE2/x
VucU94CICdlLF1BP0MjvXyAjYq9eEBG0nB1hsbLD2OZsOPFF5CDpA1QTf4/zVKbu1sID6JPXBeKZ
XdyZlzQjVehLUIsb2+cy4ktx26eYYaWK3JPHjyyD+oHkQRHKiShO/Y99Hg0zSPLxGQidXx+LkM7t
0WZqElLqS3wrUkf8ZJssiH3q3Vndk7yRbM0IilC1kLemVKMqcCWC74REj8RGdDxvRajjQgRFfb4G
yTqr8sZCQNuVtdbBzckKf9syFvIGg2Ezutg7aH6665UOrfNesHoSSK+SH/aYzBr9rE8hLCxAvVsO
3DU/7fV7paQmEYaAO6zofgOKp0RV2FF/aBuI3nlVUM2FVczNAYLYXWaBhZuY9/mDo5bN+MkXcRZi
kxVitMXuD3DbA/Fhb09PgO8CPfzKQ6v0eu9rbUPlJD2IjnCp/OSx3eMNhs4VxQFSa/Sf8N6MC67Y
SytUUKaBkmXwyZH5zio+4oyRGLZFU6vh0Jgk73erHlJWjqzhmLdhT8ntcWINJV5/3zAROhqqH2DZ
dRKdF/FbvHWwk6mltfkRJpcNN95LWplliKWW3mQgH4kzHH5KDiJ/LhanLlFVOtizjlsZVIzgXBWf
caiBVJGg7vz/Zo5+GoQo3/nsddz0k+R9h5mDkbGS3r8q5IgLlmJxuuGsiwLRatbyRwES/QLXxPhW
zWvZ+lrsb5X7PUh/M4a1k1ETLvres1TVbr1er5XeC0gA/qUOQAIRj1Dl2yRLK9pGOWXBtzEmbYNe
OciVfZ2uePkpOtLGsFSEovZo/6QVeS+UEhl7C/Vwu0KSyGW00S1sZp0RRXOK3eXy4L4otGigJ5W0
0M2+sUaVqIXNk9hVr31mYPho7n8Fc/R/2+d4ay8YXpd+Yc1Gedc/hw6J04EWUZS76LYC3+Jc33rh
ptlnxnYqPUBF8r6ll8OzEeClySClflfcuX3vdvxkry8eOqqul4PlfBHctSdnY6m1yvZJkvNXOMg2
TjUp3ByFIo7c28TjNWAxKFGmH+y/cXD/RzBmpygXdN234RNNtXgp+Coo+kYiUZPvso3FsjaLrQ36
3tyU/7RmebD436JoLUHjHIdlcATORczR+t3VW4GdcoxRA0rNsogEj1sMlEkH/wR7GcqmYI1vnNza
rz1OXV7DXBwyQo8EQfxsmhIW8jXSVMACb1mgVWQ3iu45D9yTUNiRj7H+wXa+6Mm2V+8w/dmtGWxm
RYClVWcAf3DPjlveY8gxRbegc4O2Mpufe0SFBiaLj/h/e2d8RtMvB95H9CRNWjlqH8TgGwrF8cFm
IyHJ91ghlV+07f9iSSCCGFIAxWQrxoWWFnzaHVOruVCRst2XbLllZ/T534SEszHNuqFGR3Lsn9yh
GLGDDlSQQH1Jq2Izah+NIbDhTGH9F9nt9uH8K5khZQ7zti3fobdeN1j2MfpVYEFL+0larvz/2qem
B5bTWASmchAoqvtq1ERATdsO6URTgrsrsCn3FzEc/8AeGhb+1spA5Djt95NdhMfBFPgIMKBnoDEE
nqjf5pdF94KoudRbY2Ow4nmCi/OMvlmzORK7Gh1+1FYVIF3F9jLljCO0r+Oosj47xqt7uJqMM+Tw
/ObCxvu1ezLMDtFeWYRDBWSBbBoTmZjhQJDZcIeKxPJDBTVze014+qr8eXBeDnVRMunWhzjfahOn
dRqyk9OnCBwz/Umju0YCtfZpid7t4yDvYBDjuLmrOhhF6+VHN48RRVFdAtWWpYJ+7eIGJhXaGi0b
u5F6rfiHOpSWSjOGQvGEtERJ4A/1Tu7KCICPpBelg5RK8myITq1oMLgiXPe4Cpc3OHxbWWDbBZDC
d4TwYa5pXrJgxFvQWsiUS4PpYJAhdynSj+BIB4J2ZzP5W8ySsNwmQ2l3YeeknSY28aCSPc6pOMUY
WgVgj6cmZvFWSf1MGV5IOY9K4y31li1SAPmvyYUFqRmISeQqoTuTmL7G0kjW2pqqE7TdiEwywpVN
1FuGjmJxIg5AJ4N0z4n6U6zmILYipTUaYhyCxUkBm+6WKIPSecq7IFjHHVa95Tvtsv1akIfBA9g2
AP5YuM65L6Wn4tSWPik9NsOsGPURDHkx5A5BF8FsruF/SJ7exCOFzzcdxqswdYD/AvHrPgbFqLZS
q7w62L80O6dol6EulTSEa2MrByChxsXgpienEXxZOKRZfMd4Ni/6Cl0Jxql9lcjizqyfGmuO/DCV
SbzmT79gH2vancHRwk3hSTMqSU57ahvnxdPP2/tENdhAKL4PF5MHLUHgZVMYj0EbKCOy+6c/Msib
q9mVoAcoW8N62wUZEoK89jQEysIoF8r+A/zOGlMar4O4VzgWV37ho88D+wfpyXbV10SVGEwLPTm2
ZVO3yEjAt49pCQONWKhmhJOLyIKobVYvVgqZ4SyaTD0aoIhxMR8O0Bvxjia+GduM1jDFAH1Td8UF
HXKaHx+e9/OD/3feWRoG0Y6db/6xkxOguCUOso0ZuBFavIx/pi4/v23Xo77DYdFOhKfAwBYPHKfc
JKuTwWKJm0LkXH1X4yfbIrIqK5V5+w2Naq9UzGOqlLuABh6++tTco2t44+LkiNFd2GsNKO0kPm4e
k49HP8yY05ZJ0gtDXsbKnf+MdnvxgYr509xPPjrBgnm6N3VI/z0lXXZt3raeRyaBHfvCGlmsOOAe
bBSl+902UiSmSitkWy+GYdRsr7FLv8o7ZysXAwj6BAnYvzHo7DvVn3JTp5e5zo7D05tK7rs7WiUn
Gke2ozIoah4tr2LlLwPvx7jlhlyiOf1CEdtLBbyQdrFKR71UOOESTzHANo2njfpkZkDDB1+g8rco
fNNUvuvaUdVH1hPcjai+8oUlReom/+QTozja0TjAgecZym5COg1FKyiJjc/SyScYFPLM/I0/8DQT
HT+JTL0/JeWi0huhIGlvALiEFwpRO48QNjijMbgjrq3BDNFD6FeVED7GEkfuN6iO8/BWBMN6Ibvq
fL9rlbLkBiEme9fkfRsTUDqBGmk0gDzTMRG1TcK18+BnnQs8GRRacSvhcFiYqb8e5wMhZ0bdv8al
hech9so1IrStyUUGsOjD7dYianCoj9kgjwalTl0wE2PLb3d0h5tyCi+DIWSJCewy12XyVhbXNphw
xc7SDyvLGecsylxzYlzbjZwSlIi4tYOp1BwVghmk1lWMZgX+4cK+u4CeMewElCVWwaZlP4rKcJFL
G+PsC9qojizPEK0Mi9N9Wwhq36/dMXfuWnWF+K5VNV/DxtBV0RaCfk8DUFHwA3tnn53SsigirkYC
SimPw79JPlpECLnx5P6lThkxOGWDnMyZMQb7GBPmSCKwiEjtb/rfCnr310adLV8H5PEnUUbXgosv
LpdnBccwzFixUfe63RxnEAJsx7jQYTK4CngrQgkVb3KV/AWeO9ouNQBHkSL2uK6/+c5aDGUcQKbG
FE9IRveqYat85M4d4rWRphKGPvUKiufuaMQvbke/7v/w9H3P2eAG4KgWfHbWRolYEawLp/6OifdV
NU31VLd6EXTWs18Ujr9NI9gQrPHkiNL4Uh/F/U4RrYXu2ceOzzn2M6sTEM8VjK+Z3NHLLfmPRbtF
nN8NUOV2dRAzqKdOrHQfnsDizXgMRuN9ofU/HR+LVQtU2wi3Qug1Ex/2cVoDvmOufbPtr1NT6M1D
1ixqa0QmE+BdlONFgP9c+XSsspci8LYCJibE4btGr9E+Kn1j2/ED2I7yYxovcbAhwx7emqUxGV5u
JYW6xZ8Kvy6i02XWIe1fwMVqNP5Owtd4GONuwybHRbg+iHIAbkloRS3CQygMtkI0AkdLllDEXANE
CFZKr+HPbfoyzdgYa0f5vR5h3+Vw5E4eR5zEeUoArtYpGwmzBoZ3SfoAsWwioAvWZt50hoIJtf2U
nfvMooPbywV7fPcAhaJEjConCKKxtONB2DqELDVd6tzSgqfLboQftk/qJDfd5pWcRHBNJIaE6Jno
idwSWlJf83UFfZDRWrQemPE5AlIL9DfLO1PhLJzk5J1ZZBgpoINc14dvh21xIpv0MsO6ffCdulZ7
B28+PlzLH5PyFDShIiNxN630dOXTPvGjbarbqP5LkWPR+37eUyFdf9DFiVahmnH6+E3kqqjijWP1
BJEMShqoxUbsB3tndRD0G4vSyw2cDO6y8YcWAlZY1n6GwfmDD+0fgEduZewHSwPmL5jc2qE+Evcs
94him+v85AIXHmE7EovThgwc13kFZk0q/Qr9rRWVFZh/ZfzsbIbmTNOMEzWSGwkVZxBCESv3hXR2
oR760DZQ3uN7Gp5HRfhOwEqBhg22MQRnfYPlw4xZ6qHuBcSizGHRlcsdt+b3jMVfzGzU5sKJuFnh
tIqsvWtgzs2N/cjsasMsoxztJEjQXhBENiDmpOX8/tVrZ2VI+JDM+kcn4lyDklPTacesiPd0ON7a
UDEsIIMwB/AfYi+V0SHlDpfZQrSnbzbL7Eu7fAvUSzHHPkyyAUUUNV+99rn9S2zGKCemvQFEaY53
FuC3rO8npRJpRD6tOocdlomNun/e6idAOqpSbMrk28fvvPw8BBe9o1J61coMzkOtHpNGyFYLv+3u
SycW27af25nwJ9ShQ6n/hGPveYsSX1TrZxDycLyFvPjQ8qLqfZkk3Vo4g42doppRscKeCWsc9OR4
apQEiS/hXlQOq0o0YCG1+7BxDVuE8ewG1fBQ1T2/J55aQyNq8dblukgt0eJoqy/82E0eIUjil18g
thzuHZnNWZpLgWC0T7054qWMihmlqoSvTw5L20sBJpX4sCEG6BoCUUPHpk4YOhcQgvMr82PctDa2
MGE3GV4S5/TT33sUbt0Sr6zDgjnD5r8wm6thpE+snlCDyenWIAcIahyN0JITSmoNoMzoKqx7h8Hf
nWr+0akhBc/zzK/uwHev1qKYT1/ojaxd1ira/HpakmkHc+7yEuvi+DLE9/LnlMd+sIgoletFFxl3
dwG+5WYpaYskkHoqD2Yy9gtv8gkcgUaomHvLkhnDTMhfPhLzzCo550d+vHhr7L+stGi7PBH0pEM6
keYMrLZMzsKwHzw7zRmsSrnmtqaJN7hVzsD9J8LmHBdJhOBXULELarJwR+VtFDNeK8KPnAEdDSn+
v4kxwfiqa1W+wnBMf2+EzV4q443N3ivQ9m8jGl72rQ8IIFxTrJ7h07EB6yufvyMYXn5SWT4qLvg7
jSRDBYYfW/QO11Ez5Iu4z9FZtNbhamWLg9kp8HQCh6WyBp+BMDScx4CmeVN8qPEOkZSUbWRXhXMe
Mgmgva0e5sXA6/lLiiFS6y3SSdkCt4Po1gXqTRKOtBMPzlsOh9JQHwoJNGigC0f+fmHimZt9D2ZS
0U6j3QgW3sPwIryz76o7eqtcTl/iKvdCqNVUTGCMVsktOiMHVWIJ0v1YkpwkAEdmHUGKv1GJ5AFM
AkczIjmqhUbS5+xppLFimreBFULBQ3wi4QSfQ3LDRGlehuLF1YpIQH1VDmSkOCxHv7DDmvJo4EKa
utbZdUgZjxxzfsvx2kP8x5Ejt3IP8GqvtYsqH9fZqgfXI40opeTZGk9zDABujTG/sHDDId68kEPD
C6+gjj/9VaxSVHiLCuMKRS8E7Dj2lwHjzogmIcKuv71VZ5U3eZMPryrxhkLKGal9M/x8h149wNZO
NXpoVaJvbxOr9M1ULH0fsRBEcSLflngZvZ6Fx0pzV0cwz6y90lBrtQKImiKI5VNVWP+Se5JkpzNE
z9UEQAmdwLQscI0uXS+3VQRyLxpUgeBALfM0IAc8wsZXBPmZFC9thT9BI5nsMrAzc0h+Gne0AV6e
AhzAPVCvgXR8era+secaQLDh/YMUFBsUiNozy3E+stAJYkyY2kYgDuseDkGx0R14x1zydB6CtvQh
j+I2Efmbm8omgvM7ooze1lsaaxdKdb5W0vJbfoDsVbvlNnZOHgrDqWz3rAOxQqwHmpE9ck646+Ub
ukOWMTNcxTml2m5VqGbpaV77qj0Ot+7vZu3Rcg9XMD1EtUfGbOVPs9jzGJ/3h4HTX2uR2vAl+ph2
L1D1YzS3xNIQx/Ar2ZLOwKz5fwNJRFmqKbcMvVWVbe3vaXsOqCrTCsPmLYCIU7B8iyyNvk4gRMPh
Pirzna1gTqxk2Ok1cZbVxvxX2xgAzQgcCezg/Utf8GUSHadAhLlcdOfi0T6Z7id7Szld5wLoTZnG
C8UjV1IYnyLIiO8XJGnmDjecOe138i/yAhkkatlPTRv2V3by40rdRWhPvQ1FIwwN29nKmpmRRwQ5
DyTkk+5NyHoUZifRrgIHXSzGcEr7EccJEHva8aB7hVav2ltUiNGlKsuKuZCYHxQCkCKV3w7D3+rh
gJ+gjsvDW3MMGhZC+Z8GMVq0Drj8blG4F+1eBVPJzca5gkfdEbBtMHMO124GvT9rDqlb45nsiwSI
b3fZsqc9Rxg/JiSbHS9VkuqMeYNYzxTijuxl6uxEgF0PexE3AP93SpF3VIDB8rV+zklvAh11e9Rv
AStymtuWHAUEoM1LLwVM6TTULPmusv7eTiiwXbESZvh53gFeSwUZikRa8xctGoKr3Ko7YGRbzgNS
1qk7Nx5ANSKseMfQ7bSqsCHGvHycHalweZaWQ7/5peeQNDaw+xpKxP5soKUjAktE9csoLg3ER1M+
gJkYbrKaw6PFizV/K4mnE147vR50SqQvG2XQ6r1/OcsWKqyVWF8sxsbbGVX+wUf9HZNvqN2y9K+9
EHJ7F3Krh+aVYiwfwSPI1xOKxXS2mKeJ9blyf2bKm6mmLvyt019wsLNpcMHssRyZpKL8QP1kk8Bm
UCSn7GqLfaIwDxqrQuqLOAn7oIhTsOWVOwM01290yHk2uNx+utIeNE0MIy3sLMw97r7qSJExvIzu
AL9fP2caKGz7qXmB1QdE8YPm+cVeL3oX4JbT+srNqrGsaQ49PM0q9RXPMJxjZRSwVB2Rc8gBFuoF
Qg1E3kjr/thC4zRVA8Rv8XbLSt8la4UTsf8IFCUf4mlcBVkcp/2uTRbRKvhuGJBtQFfetrpTBbbG
IfdCPo4tbJC3NjWa/0wMk3gUgtS8eC4G5tEuO/tXaB6oFlbgvNZrUd4crcu2NSE+tNleQQTCVze0
yiJfsYkjfRez8JmyBDqkGfviIVsv5BdNbqUyoytDecclndfVh7JLSYZpekYAlxEybR/PQVNxHXyZ
dMuooky+xBRFZcgVI/DaLNfamtbXM6hLUTz7KMYBPg/OQf9nJIJUk46TjwLxPbvDa/o5XiHcZICV
+X8IavmcHEcapl35ER/jYdoZcrQesBgNtFE3vqDLRVxUwnZdZ/V+oDqeY2Qa6Ry1vz5Jg55o2Til
BVeO6+5brQtc2rOVRyaA7bEplnrbxcxYm1cNCyh5N1HrCtTkh2HoD80VFJbdR+DjPUGpiI325zBU
wG+7kbfOVOx1gU9MPOV4wL93onPm0EQ2eeJPlkUKSnSAZWQpZepnRIYldDBs9/v2sXyqP31yS37o
Hz7K37fTRH9Rs7CPlfiVJI678Rb5CMlGgZEBqUgAHbYpr38GQ+VPjCGWSjn8dYMyraZ9p/yRUpjz
JWhg9lj+EJvwWWZiONdCu8f12aS6Rf5NISez/Q2mDDFro8LxR2STHfQXKYKL0Uu37hf9kFpJ2349
mvU5fmTAtzvoBDCUTZ0B8UTWhBEJWMGYDdn2awZSgVgY6PY/Xtt3exfZQT1Aj9uBOdUv3SMcL0IP
u5dB90ItCoLm45NiHaU0/4aRK/y+iUqY6N7cf0KirbW1Qtz9YdbIZI4dMbSrjt+qJ4QFLTG/I7VC
KFtJwdSYPVcLBEqTW3IMQONzBEZwjrtZr9Es1VYSAq14kskUggkhlK3gbHwHZtRKYBFNe3cDiw+q
iyiWO2TpVQMHrQ3duU/sZsNOpd/icwp8TEYvu8/8phX2D9NiyqB0YYQX99RyAalW9eQMdbwnw1OA
XyzGKGeylO9Cq9XRLiTDXJMD9mQOI3pYtZ5HNrPUZHxS4auWDXk38tGNe6D1pAf1Ixg1v5TV8eUQ
MwbBwjF3wU2mER949f12fqfRJUmAsKzJbASiEyS3F2CinllP9dpGrN1hO+5GcbVRg5kFvHIq3qEP
pYQI0qX1yYkVKfdDfh4+nHOPz4D2wZoWxKdUTbgOYvadrNLobnUwEHqn22/DzvnDExuhyCNQwchF
vo+Xr/2KwMF+USjondvTMibqY2UtQFJpl3fCmTbFcKlvIbg7ch9are1HuS0FJM5HsXFnol9AgGde
t5GNe/r2q+cKrMupMSFYIeqvfURTFVEYxC5RqgUAHIAsKJiwVQUdGiBxIFbgT/LrxTEMap1mxrFs
6UGYyjJPPpnC/rqlKNva4ur684du907VTgO6EGWD9ZHAJcsQ5daHPet9/yAa/0jft1a+OE+Y0Yo1
7wIiAzVjqxvN7AgFG0FhNS4Nf34pFutaox8gMC5hLyppJm3Ag+RQhBonyBRC/p68LW3VxvHQq5FW
ONv1+vCt+9Bk7W54EeA9MycSScSGMvSD/BNq7ntBcO6mLbfjje0MqAUAYjpFhUROGazHJXAxMOXv
hNkdonFJeh1I93zRKb8jctC4aLmKlKA585ylYBacZ7vCF4xSoKk3qkymZm0Sql+MOzLWJe6kQbIn
iT5+VL9vBy7Gz67Lyo4xcq9u8OjgNKcoE7mZZjtMRV2AiNg2cZI5XaT8fkNXLliad3XPKP+AXo7o
iRxPfB7GKnmLBy1MzB8/Z59pesiXqU2BfodZLasrfdWbgSRJ/LCMsJtBxyfNaAGZwEXTp4fbvdDZ
s+RLrEbhCa3j/K2L3L3jIRWdq+fFVd7Q8yOWtlT2Y7O48TthTJrw8Tzz4uDQFTBWb6cYpzhItUi3
pYJX1OfSqoqRsxhDaEJ7kc8rLCqFAycnXczQ9+XDQtOEkn0Be0s1UG6w7lD34ezxy9bCCseXgm8C
n6bqDAvsGK1pBIcLoc48F9mH+ilqo8qwdM0V3k3/QwTda4EYcaWatOqcKsvYo1qFQj0dvQoANIQY
3fHSiA5WuOaqFHRHhzgwbuaTAO1Wlp7BppiT3Vz/B+5ibyb2yan4iFJDLXnmOgyjdm7W3g3tXg8/
EaZNEg2tuyRh0V/Ha/vfcbSDB8je1s/zpd5OsK1Fgh8nwLk6o4NgrW8lxMGULml1NGMmHXWTckER
4t7ebhsi6BFNhsPAJ5f/JaA66GTDqLZSfKNLhpVC0f/KrlSFatrFVhCGfhMTk3JT+scNiQgMsNPw
3Kfl8IYjZ3iqNBWaRzmSNaKlkxtBoHB8V+TJD+zRmhSvGJbWtsUHkVfTkvZbaM8PQd0n3Up76ejk
vcz/z/VRAjA6UBH1EwBW3sn70GaojYdDvxjOu6NMtrQqek/YHjztx1zteY0yr/snToTcq/Wk8koM
DpSMktEHYFj3vWCgZ/NKjP9chfBYVx6kTf1GXLr0MBAkpBNU7L6+yJVFrCSn6lY8veWiSXcylU/v
h1qQeCJw3VwfEG6yt5RLewEezVX7zW+oWerbl2wmqBiYCBr8ur4PGvihVo7a7xIqrYp6PH8kBfOi
fuNpsbi9eQRDNvFl+AfbDniP0xCtbWSUlAAPLHN8WGUHQBcByZnE5q53YUkA9Qs6Sp+H6x+x9K1A
8LP/RTBq3ktihoZUpTIMydIAHgoJzcfBcw7TfWpMjy0DHEGRHK3ZuszEt3EU1GDo4NXR4sfNEl4W
8so2kPZ6rKP4CsNwg6n447NSo7L9fVelgZgFQRfKA2Kvkgy7pRmMPAwMb8k20fmIZpAAe7fm8coa
AzlrCmc1QAIzRKZOhDnf+WHpuJANYnqv8HJr1vJ7rohZpuuSAcIfbiuiN/v8XR9gL80U5Jp09Awx
NEFuN1bAOUc91hrRI9+rHWYzCzZ/emwX/35KsvcEGorgkoY+m6Ceh94fjAmjw0oup4HIen92avCC
+++u6rIMHY/jxY0buUB5d84uB2KKKrsvcYF/6en736AGn4nj6ctg237PFXzxzfz0E2VGt4Iy0svg
b9k/rfCnJ2Y/aPgdGipG5ZPNi8jENZLp9jU1vyX9IIS0yNB2xDxw23xOrqyZtnns2nmJ831UzRET
h1YEcKMAUBlMxWzcIvT6DT3YXsU2c3CchdOnfSEbB2+3GpzVJIcMZp9iQLjVqvrLNGxsSKj+RmfW
y5jtMbVzxZUdsGXmI1NuLOwKraqED27lmt/capMfQlr5/xX3q4JeXwHi4xgOQ8Fy051qKpcz+3qS
GtVzmIUGJzStH+fxd+kbDruPwu7EYPpDP/SBx8/7V3gtqVL32gon0GcIAdpd5s9nMcjuO+SHewf0
b1vPrL9wBOohVnFHtFLUatSIi28fOd+WcQkMSUb63ADrK4uhO8ZmQPDmptavBVppKKF46EPctsos
H/cTSXac7uncm6K0bKD/rsq+xbrZfF4q7irIqk1bPpDZMFMrXvQ4MWErjIjOdUhdO7okcFJjt39R
KXUDNO+bHkibLkE7FpD3OBqBbm4tr5MQ90pSrDZ5rHl2wUMZv94yxA7lHA9sDy4nyjPrDCUTlRjT
v0WC3g1VVCtPOoqQrQ0qQzOZE2gP1hR37WVaJH826HGJ/T+A5SHKBhZimanv4N8nEZvvrLK2iAIJ
fTzZN+Bt0sA91Gj385iTbQTQvvD3zKrWNNq0M6xCFFjOkGWK+MvjuosxiBb17bhVmKyvtBQz25I8
Vayfn5+cRnSvo7LqPHNLIp4dxeYy1l3vwc4O08bbuOM1xn8ysWNshxJs6396Kgai9vu8kh5clGja
nZh5Napj2Vux5pEZInPyCT1c+EPb9O9AYL0nFGigaOdLRt2App6dwwTzRNVpg/dl4s344+qAmEe4
eS5W5gOWG0PfVgsX53MjiJtmu4KtpjPqsLc13t747d5V8TeYm+UZeTgYjiu6kuzMVjxmFmTuuBWY
leUT43X2H4bhawlocBkSUiVMiN9OYi0d69g5vdK3rSzBK86sES9SfmPHl+fQ/60b5g56Ouf1wksp
LyDXqC7U6qDvee4U6r5ho4KLVlSrW6GP6qUUKRCs6/j/84dsMXSXq5qx+auN9HJ2ST0y9zTkZTn8
pGll1T+qQxnHAPTaGcDqHlc3O4uVjTHK50DV4pj3Hfbilxuriy6Zn8xgz3SoMY+z5sXcSMEP0iaX
WNL25sqh3vw0ZIxgNOswAxttS6Z24SK6tS0VYH9ho0s08W47jvvhAIfV/m+CyoBDZZhj1DajW1Wg
cVkyWABPcFSWGmaclSKI7typ/PVEhutTTrNHUlZLrUagRZXBLxjSaBenMO941msd++AGlvWbF1xL
ODgfPw+cXjf74kPYJ7Til388uxhAAO8NNkgChHCk98tYjzC61nIGsZ5HkQQztkQOyNsYobEjQ6hM
gUkyGvf7kC6dcX3L5Z82LTSu05Uw3HEr1M8rTnrmRyXzFRKMBLOo/gjN76Jla5sFq122lx5Cr8G4
4Md9OIZorqLyICAKcyqVKdvMUWdlQBD2stDsR6+2psm0qTlejN6FbrHs3a39X0bMT3bimTUNYXOH
dJiCN4I5bbgDQg2K4E5bwkZKX7a+3xbEoHm9/YRRvnrxx6y68Pi7/Ij3W9dhWEw1bu4RD6m/ZbFT
st8sNaZCxB0EJfEHN6DoevS10XDq3RsFyDXky0ViLPaTTATAzMswNKj9V8pDuB2XR1lNilVzFz/4
No8OvEYGPEjorFAiPhgPPGMyposrPH2Vkno8xes0Pkrizz/ehXsJw7dJpQltTxhf1btdqlaqZgiH
Cetz9+nBR1G/JOXM9ecxedHBxXYZEhgoIZ0703I0xo4/eO9ykfPjF1VZ21UawyfyCdqhrcyjRcxr
RHU0S03YMnrEbmKqq3XbCA4xUxdODfpMlaEsdHYQwNgI2oEHdD+Xu1l8LLAIl8nd9DUI+ifda9vf
PVy6SfmxYWnQyWUgFDmwG6NQdxZu9pMJ4Z+pRA6E7MXM/X1U1X8hC96S3lb+OgciuyZosB0gxggq
wGfEGpWLWgEgrKgedESHw+I9efV9dp6lNDmk3O0NDaIF9W9YgLfOsBnTamyNyzI6eP55QGQF2IIl
zwmphsVsaDFa7xT2pQS7GeRtWOKlfl/lOMVOzROvlkN4ealV0EiJPxtUO/Xz8DOnVHx4Uc5luQk8
XYn8Juo9s+DmoK8z7RQJrLbJcwRDJja8VugdkouHkTv8A6zN0abSAbPuqaCy3wfb5wVZFJm5YQDd
KIWpxCew6rqY6XrCjX5fq/7qX5/CY9SupsUlAle88FBHLDOYEszo9aAaTXPY7O+oqsvTWEqhGG8p
9DhLcKUl4x+E2xpii/szCzbqwIxaJnrKFyqQVUiED/uWqv3waLoHyMEG1iMCXn0rcYTm9esNquGd
b43Uc9ymik9C+5lbf4xQ0bOaf/DgZ/llYgaXCG1eqluBg3v6sb80OfzyMRnRQS+tZoW0bgHlY7w3
GZcQpfGgoe0BbWhPoNQDQnuDAdNSFx2PD3w7iRay6fe1S9dbsv892a7imOayhNGJirsuGDjabL6u
eypVMxoW27f40/Uu0E6a7NSbb6+hH85ySDjEBIx0jyUAi34sf1fcZGcxCLjfjCPiUvzh1LTX+p5j
v5A3EgzDhvNnwa3/hCovW3DODAa7aE50A4TTbj5TBPZBbCShR0MiBAMTm/02odix7qtzoBr9M/q5
6iK4/+GJOzrC7U0uxxY6abeYVoJi3oT2rJgQqq/mIfFRgj5wxxlPaBHJLU+6sKKiCqqlKSFNAMy9
lpUU2qdAziQewllLNb43SqGJuZ4Dj6v/eUJwicPx2fczvOKp/8LUBunUfhU0eXkqResbBitgqTlH
Dqrua5q7Ldb02dZpME3/X6COR9nGbCxKMC8x1l1mIdOXuOLmi6zFBtEmdJsfCQO1pzhCcBtP7gLA
pH+RgwM+hOdK/BnoPRbQcsGNp/wTyPPV6a8YrCcjKQjkCNSM+lg9TPx24awfznk2VNPHxr9jG7dW
a/6feYAZ9wpkrJLgbUKzZPNtM/kFPUn9U8ECanhUar5u5m+Mu8TE65ILr3Lg2d/VFY76XPM7mEts
b2L55Ov0SJuf3/i8uHBxMFUHz/Ga70Bw+NzuqE/wJveaQGoPw8wslFCOWL7FhmGQtVyB0qyauPRg
vbzTt6ZwFaflCBPlxNbFdLZYaic76mru37bKzLzmxEyi04ZKXq+WIp8bxJfDVMOKB8dkNwm5zGXx
9PHuOalKX/5xsQT6MMQzdb2vnZFi4+8MXxpINVl1u7yZ24qDzJx5aFuYJtT7zr1aj++JHa0QwWcE
GZTu0QD++TEcrb9D4q8Q/P7ZXhiXSDiqbhKgYg77RbE8OwblZv1qgYTQNrJLnhANLdYKUnz9j/ui
6uTaS+ZJ927//3C7XhXg7PjOU3siN1a8Mt2MagHSXHBqocOydb9a3Ce3oRYp/gkPYKdN+PacrS10
82oEPScslV/Sh9RLaj0H3uKol+dzB+/G9uYZG3rxwF5FYozRnHdf9yG6Idz7/VCRGBGHe4RVPfw8
Lk1SOHUc1EMti+KWohm9LoX5ThONLgGurHsK1zmiy22mZ3hsEy6Tx52bRiTTl46jVVLHtqsobhCK
OA8deghTZ0oKk6+yRjRmLbsvX3or9wfdh1gdYurJ9qvB+Euh9JqPeRbLHrK2xRlcwqkAPFSNI9Qv
/halqc7Anm1uJeVsB0EY5v9pZnUYuA77dQyl95hnucZ1W/3MXBCH3hY3xrnrrqNO7EhAiTUN4hLQ
VipedC4TWcgT/svtDaNkh1ePzeiOyq0pzhk1jzJq9STrzsbJ/MoxVr8uiQjpnmnFWoEj8yIdE2Qy
jQaxNdOBE1BBGQo46qj4MIHklwVTbMdbRPDGXcuZdUZBy8fKr0UpLWYn5j/38+5U6LA0Bul1Jcx9
cs410DlPq8hZFNV0Vpu4CdPhJAlhaPUdIJsSq4i7pe9mc4SC32g62EGyhAvj5rTvuy6VxZ3+em2R
2vAVGsaGfwzB7cBgHED1V476BMVdK8lvohw2NpLT7PL6J8jvl45tTZ/WV2uvJWe6k1HIq4VOI/m1
K0qk/SjjskeHKKOloSqc3NIimgPBj1dvqpHSw/Uz6HoZ5zHE3c67sQW+EtEyyqX4pn0idxW4BkZ0
OZWN6VspI4LIq/S+2wPvqlIiqo6Mf8Y6UDxtm6M1onQzbpEykxMeOGOrT/XIIrSaKdFnJn2ATUyE
3Ywjy50s1+Ao0eHtWpxEvpEAtUE9G2cVEGa+vSSIh6hEDlk7wy2TE3nBqmPgg6v0V6nD6fbbyutQ
Y6bo6GPBQKKbQLWxzism6Vtgihz+CS3F6gmBdRvvJB9+wXuWagS4DgrboKVBSV7m9WVsLYW9n0MY
bGC1DjRUSuO8PJlPRKNA6nwYOFQ0j52skcOP/H2F68uRSS9EDK5YBsyCL1HccB0cyR2VeVcV8voZ
n1I43CL8tgHD3/f5mly4mdBUD7BrndBj1nTCYm2eu0/ge8NFEKDvnxSBzZd8mkA9sABm+l2ol4Ab
ZPDNn4Rm+i/PouKb0SMckdUhWdh2476I/6t/kGkvxLNVJYDOrOGyp/l5R7/EffEfTM+ZCCIl1vZm
DqijvtZU4n6rG63cvwMpR+qhjNvhihMeTqpZWqKFf1RG6WAge3ukbL3YOY29mzQte4qVEaYKecdr
oigixqZbWtQ1Twxs2ejnMqN213okahQcw4O/4IZYiTgjTCW2rdFWd2lAje6cJPoyGBqSXPRcD2dR
bGpCMbPOZsIkOcAeU2G8eTlVmYyFKJsS6kWwUrH78wJr513iTStUAzvFRCLSOeIg9HxPzItiEjgL
el6Ak3yd43ezVGbfW0/kF/G62zfrnmlHmNU4T8uvyiOtJeo0SKCxjt3VzpmDBMO6gOBKptD6QPG2
URrc+J5n75qcZN4/6dRzXhO8RGHdHSi4n830itRLz3EIVhucpAHMuFhmvNzxsgPt+oUpD6J41f6i
GfQR5vEHQx+4LCDJe9LS4R+vjYDkkPl0583Ih44Ln7hvH4GSqM1R96cVNC+KliZMluo2J2sZGRUa
IdqifhZJdjQX8uExMQJVqdNjfsD5A05hIPZG6W0T/0vojmjqHE+t7YwS+r4Sztr7YcSvKnYLFFaW
vzQBMdqAu5zkkq4tZZGCQFXBatNeyptRh/J3rJ2ABWUAyINfNftiKpL01VGkCMw4nX9HvweeMXwd
KrwGxv9+ZY6/q49iVkqiKZv+CR5xXZrgc1Dyi5Szmdu1I0kToneuZBzljbbeXBdXVFOq8z8EPJGT
L7mdRka//4egm8YkeAPUdXF8LqYPjgkEzy4ByefX2E6tqulU3AJ6ZTwA3rjsb7qbF1nDIbyS0yUN
Dm74kFakeuqSqyde46oybJTujq3wfqHfAeyi34t2Oe33n+e0C3vfCgQr33AnL0nqb4Z+Txt1v2hd
KZMJ2q7hs/gk6P3D9ZZ+dhSw98NR5PGQufiuspBJjq9leqW6q8ewFiaOY3B0dnva3LooqnHX4LfW
iqSSD138ZVvj28MDsacWYc3rKYUn7sRqupnZU5BCedbUH2BH8OogiET1zjgDNNpCCkWipyCfLyud
Hy83YdEaPYHF5onix0yPbXX8UKimbdGyruAyd9BOMYRQ12Q7psPk6Xn/eCtN0XM6YE+J2cPR59nB
odzjo1B4p4w8zlFtjZbYhFqky599jaO/8G9jW0Msla3lnmCm7vf8KuWvs0eHrqwX8v3jlOvzGTWq
G9B06I5rag+6Vuoo51AEEYxMe9E3P2qBenFqr67ax6WUl6Is9KENLsufdHIbnSSwzbHnpZMvUYz1
0F/I1sWA0FJCuxBmRLDOMI+41uNz6573S7VOs6/SBqb1DyoaET+LVgR6+kHwPicRlILOv6ALbc3z
fO+VMlYR/MPgiZ5t36zT6UIVXEiycSZnyt3PIXv2lsDzMm8Pk3XLlw6J1BFccG+EesXcnX0FHh8k
49dP2eMeKbJ2A4SAgB+cikCZoa+Nbsou7zLoO/vbYOXjLx82uhmUZ1/cxKuhDXKvTp6uIF35HxFL
RzD+JYey0Z1+eCHHYOonQlSopl9SHgkjr6yI/odCQ26HLwLyHRfTn5mDvJJRU3n8qB+b4Agw/hd9
fCF52pOayBKQg33Eyx8BrkQ036H9BRjObhLTc3wn63wegyG4TB6ogJEpiQv7vCIWSlaNrGQQ/Y+F
sB+Hnk7pXcTghWDlD3Dgh8SJGVOdSuI5FUwckRNYqjr92/2nhQTN70euqcasI3ProjEMecD5a4R9
aVt2Rph/eY6f/Ik/jD5bUICZmd/UUyypPYeVuwZZ+sHogh3Fe4W14Ab6Ur4nXOA3woye4q878e2E
glT3sU+K3/+peQcQZ8LDQ+wvuhEcxHZSGNpySxLdBL6/WP0nwcRAzvSTS7ANBxYQ5ASIC/CB23u9
mKDc+OU/pGdReSsxgcW7rGXu4OWj79vAyDYfjgONf0kzajzXpVM4lVBqnRjCsa7shWxJpPLDC7iZ
fTxI0mpsQ0Z8uBQiIrdz8CY9l6Loz8DU2E8oFCH04hUUpnTXvJ2vb1UMLKhjpF09Z20oTve7AgwR
LUKy2YSlNJ5Kpdm1KW1s3tHqmeyYIDJhBv7vLn37GidWcYbNNPKNZfReSkahc79SKu9tKv91YUxZ
2QqHYLix2LezCJ4HB0OWGf00cGd/LnSFO+kI/d2wsj5fcO4phgckTiSTpl968T8TrwOAe3EQisFi
KpFWcp0ZvlnjIEOdSOlFX8yjTyAtNA09dUH0/aQTZHwpvFNVoM/gFJoHQ+7TCxXe7fqe9IJBgU42
6BvpHdb+4tvplIRdI3Q595qQam0SwkKtYI4uEPyPg7B+Qd8W8rMMxd5HuYq97bQKHmAymM2wooMt
uWnXYgGZoC8Y/mYMah5cBpqR3wDTn5xryBPDkWjym2v3AHZ0VB8rLF1cm+rDhAjyK3QncRmcHboW
d7TYM2NILwxg2RvoHMtEmy4SfY3HOXgNaxA/rb2G2/GktPOT+4uthPEZYLrfdeQ5CTQUshat14mA
oj5lGK+WN+9o6eSg/dE3DEPFUAc1TDwdtQ0Kjx3szVzEHlvsD/9sTJLQI5AB2jdwJSyMhrfJLa1/
wDAIKlB1VhoW0Y0iRrWirmlHnsvPzCo4KuB9+jInL2QnomW2Gp9Tqttiw2BXQkl+ctx3VhSKd5J9
Rk66G1E6dRERWjXzVNAn1VFiB1XXDhKjpQ8uydx23CI/7SLsrwMRNbe4XnC+mrMdT0GQlWGoKBSM
fr3xO5yKuoZWnwXGW6RRqh0L+ugM7NkP7bLIoni+owS5Q1Yjsk3wi4h1QHZPF4sUMsi/BfirHXvc
VUNgUFQo0bDE/uUhaI+g2RrqPI5FesDTMH3vh56T8vT77V2ZAo15+kHQJOgNUtnh+tSyEt7kiu2/
qO1osQAM0McEGgCBUJI8PZEYmtdLd6EaCic47IMolAGP7TvZoETe2IaXG5YDxIcDGGcG+2GqaZ7q
0WvFiaR+mrCrkvlZE7gJlwf3TzbindklgT4rIew3O7qyHL0uGtnoQCZxKIsqIhTVuPCsYY41qgu4
fCjqiu0uS5NR2zpOkGcrVN48eh2igDpXjY848Mgm+ngiIS7/MBATuOKrKS3mwSBFuWmzd6L1HvAA
eARoslB8LBVeM+lsInZAmMazSqSfXuVNTwKZ1Qn2QFovDABET5ZeiQv9tJc+GnnwNx7U65vBTrcZ
Gys2dc0F3LAeAc1S/lsbc74aDmT3aymDCJBloddMXw6bkOrxZRJsVsmCpA9PAHVrqUYnFVCbWixs
Dkxmu5qy07K/O/GbDQWelx7vjwPER8KkWLqpTebHriYpStu646wJWyZTLnAIa4L+1tr/qoSVwSRZ
vm8WBLPgX3GQYfP7U7JeG24CICncnd2PnX802ejHnUbESBLZKCpe0Cni7tMGfsaDe+1+K6Wx4W/4
fBbOGriTuK86ATsP6DL7ngKb6S9inZtOOMT63RKlW4V8yVJNerOsv4mpqGb7p6oTg7W0uDwOrxjY
7E/U7Sb4yzOs6+gprMH6QfYj+2tKH5OAidAHWCHe6FxorAGZJG4JEKk5MSsi6zBlfPY/xbQOVOhv
iDbYPrbWR1ffbF7i93bzwLs3G3HPoBwmfshy3zvf0xMYiCAC2r3Yjua5f9T8wKYFw48h2dJWgBHE
vBJ+TKOnRFHqH8wZgs2TP7/WoQ/gqlsJCjXmHxuDdfB7/JTMyZ60IYuq9ez1Ef44uVYeWuftjzFE
2NQjQbAuCDsr01Z7HUzNjd8O9rTZ+CnkkBhKmvRuk0tg9LguAhMIwLo4CEU3Oyyqy/ZhHT5gabdK
q21gm1BqD5cCB6m+lpkVfAbV5n9pMd1sr1nNdvHh28lMTN/jgEcIDTpAjQRDk3qNUfHpLy59BdTv
Pfx32TPDZ3gaZroc8Ygzlp1FeIo18I4OPU0C0gus3OX+8ecW8Qc3H+PFf+Lk60tlJ1zB4V+y/Wqt
zMZFqWvZy11dYBYEbd1Hkucz+utY28AK7eFMdBuAgcSqGVTQ8xN6wFfmtG52y7NcAydii7AbWdh9
ui6urTFeTXmuVszA0DZo8m4X/1L1gA7qeLtkb65OlBBk0/kuVGh+rOpr/jG4kMS94ZdChbO1Yhs9
qmcI4dr5zPoBvnYc+x2P+ZlteyzM/V/gt3dD0vv3qgN6mQdkI9Vs28ph8LMnHIY9hYf32MA2ojxU
XpKQFnGQul62qRHKQhHqOdHaVa6XNisChm95+Vf8Sf9xveKWtFwtCM6Y0qwjGJeZ+K/5mI7SCHRB
E4ZTj+YqMqY1B/vNM5UfU0fDLjRoqHu0f/lumTp7GP0cvu7zCJt2JCBvZmMOg7VTeid4otUU+/1S
c3xnJdRslCQhfY91TES9sp+twTPEs/tDWUbYRbjKW3r6J/WGcaQCVlPfMKrf+l4hp/OAUATZderD
4PVawbwd+R/Rxfa01fv5x2nHKJhJA+1QpV1PKHeO4Cwi2KrM4Q58moA1SfuO/FGkVNhTHI8RoFqM
mB2TBeL99zrUd1q0IA/FiFn5HcQ86nbXFbj2Zse/3dtx7xipZQD0bMDwwn4mqfYEKTLyekk3IYfI
5Ujz+5Mo2uz3ITfErWFU56u/nX3K3xPQJdf5V+zYk4VRhnbspCp5m2VJuTmo8qaHDxtAIJxaZogI
/LdEl2fqAeAQOSZx+Qc130RpUkqp1l5VWtWhuHTbqTolC96BeY1GWev5y+sDXhDUtUWzSsInRMKg
w0sIpGLkPus2wqVCl1jsv6M9b2zWTL4J5uJgEkPBbEc4yXsJmApgmHgtS5LBWFdW8woeSecSSkO2
Q/r7V9xOV6kHsWkIGgCEYvAfWXAM9TU4A3fhZgjC7lNrs89JEmd0OyMc+puwaBBgmRuxrxQ0rQqA
ldpX3d8BU6qr8RmOujTft2uPlS+4Ekqaz18AOP+g/jJC5l4t0XjDXOVO121L0RL2LiQtPGGcAWkK
P0jiEW/n64+Chl38nAuUj2FapvIuT5sr4PdQ5l/KfdHtdBVia5CUqlcGCnwvaRwD4XLfQxlbQQl0
0M//jdcDboGbnI09521DCj33ks8WrB6ETRXRuXYMDdjPT8offxYoXPGVtNHVkZ67yG/ZcmlNgb/t
ZSDZsO379mo90cPlR43lLEBta9PTkC3MMPzZBRXlAlU3V45gsOjG6YFHrLk8ecXJehJr4fqXvC+r
XrV4awsY+lB7YVxlCohVsxXQi8duAveqNI62jJWR4Mljv4SpJJfqhl1O9cS9qwc2UcN9+ZU7i3Hw
CxOgISoG0ImcJBIC2jlq+EuGCJIwW5kBSfP83RuJGcb02cstiMY0h79k937yueP2smBfWPDJt83X
LdSKAoI9fzVszKQYgsQqpubeSFCi5SsMRTC3qv9djBLXWKQVlxTvyAMWmAoyccGLcTylbY128X6V
f4wvA8AYx3IeZsAQR/KxDhWj8mkCWYxSHNfES+q1bObFSbAK8wSHA5K9bxtRmAUr6y/5/a1GI6Ed
Qjc+MfpJTaYuSsz7ThJHVcmjSSeMq0P2X/xnSLd0oZKKW/TUc0U7hKJHX/xem4Th6wxAR5psCBzW
Wt8VyzxqTJq2OvhgPtU5JYK/FIOKVc9RQJrzdHvLY2WihAL0XVvJFuwUHbBd5Ir5Ex2VJbjh/+Go
OAIvhxTm/xik6lPfBKVcxlTI/1hX6uBC5pITzzR7XPPG6JOQFbSozganQcnsjIGEQSh5SzHojgj2
zqSLl9PwaDcGJGz5aWnNBUp6Mg4HiaN5U5jyX57dy2p2prCqc5wqCjc245JL6CTd1Q/xuvrIpR2g
4e+FmJhsuNuCj8o0tiP4w9T5V6d4Sas1S2Y1R49FNMSqKIJ8uswFAu68sMH5nyPRu2zDJKmNCHQw
oa+wanJfvF6Xj8XjnMvrPl5WQ/tdTeYqs2nxhhoOuw94l1BEqfr4c4XO/XtY5KXA5XiqLX8b86Mi
26UGFuM13LrfFQNTiQE+f1OHEpWPSTbdLNAmNhmhekbGXw4HZMuq4Law3lXAAsKCcjqVrbTt8WaM
riUPD7/dH7y8hEx9b/Pkmp/JV0IKUpWqpqgd0Luqo+fLjbzqo6lCKANw8S0ytGXvB8n4Aizpj7ao
iYaph4YCu3HdRiqx6o5oEJ9Vuix0IQkodK33fzFOW7pHz7uuhYBDSBieiCDB1NkyvZ6vId2cixJJ
3pGQw67vAnjwRT6CJjdyNxgq6MBkG1pkc41la/jy9P0wBhUpeOtY9PVqmBMsLBzzKnsUDCtNjhrm
k71dHfu9NvsCp74Nw1jUOWZB8Z5IoT95VGAI8AWYZOEruR+crsrhfLzP0Bd2gUB5wk9RPbvaPTTO
vMwvWAITr/O3cj6FEwP3nGt4x359T1jT0qYMtyCUkY5i8boWHbBSmV8vV3FemxreDkhB9Hzp86Ap
O+T4aTd5fLCIC7PV6iXdD0BOOT62GIi7u0UjbkDGY1emsAf71DQbIkOBuQee5ls/J33CRaAWeEyf
xQ+ePQ1p+zv+mR6XGATWhgfwHrcUmytB5IZ9XL8uQ4EXum8rxrs4i4WstpBDzJWl1njY47MJV/I6
wjdhxPXEWIcCmtc2Q63p8hwbP9M/h42EdVLAvDTad84+vt3P3gbX3dw87NhRrJuLgXoa6N3ze2k6
JauKVEkHNQ/IC6+WFf5ktMPr8+Bd7FmhY97VKY5Lb1TRLNwdvzHljt3t6IpFr3JlT7tO/d71Es1R
MkmxqtdvVUoCTDGIVF/2J2oarqfAeRY4Oo5BV4ViEyWnUvCCAGw3f84MxVof/XriZokkIHxAk3qZ
Nh7dMlCKAwGzBgxchPC3F38+pLQop9tMWwLZum82KSr7q3JnC4fiKuk4oSSYFOVBjRg7wsgSwNPD
kJu1opSG/11y0hQlyV94HcZwm1Bl6EeuBUF2gM7DAT0eAWlYbixJAayWtfVt5lZTtP15w/4N0Q4M
/ZR4EzWxpXkkCqP4jYYGpO4LA5RDbL04qkxGEj4iHTPWNNqUCOney83bUPD6sBxHXq/sJMleGWkt
Zv2lUTzYsjc4/dfFRCLxuvtrYgVUk9gI/Gqo+Wi3R0LxXA67TPHEYldM3geeVVZyhsjjB0cCHcnM
ne2k8Kt5wMnSuyXC2l3CRtwhiIxi+3t8kgCI9Ylya3BsBqM5u3adEMp3a0uLphwtEoYIZBnumzub
FXbp03F3rd6oXCVwcZ5QDGw42v71t9lpayEVMufXlk6r7u3XtkbTmnd9AJNaTyjIWpTJS2sqOWd0
7BD58wY4ZREjTfhX0MxtX7QAMkjosUZoyg2tFylFv2gpH8CH+wZSE2sIvJTQTn6v6lE08nP2YLbL
VpRNFsNHOh2U3jHG6iQse01guN6omcYwwTDn5FwcYe+F0Ti9igJeSes/vwyBJUcJQvOxZlmd1Q2g
6/jfs5S14ay7KEDq44/fbRklWlIrIjiy4nLCK5WEBEL0JS3t9TDOyFJqmqUd9b4UctQWl7+XEAHc
NQDLIM8D6sIHaYDjRq95lONICGgEs0PrrKgRaQDKisnfZTkEwSeBI5FTHwPyqCgZs7nz3K11X4B0
hpVvRbAxbGkydzlQSr05ocGeQNdoaMy9Ltajt+aY4hiqpr1gyjwjqAhukKLGTr73yKaLDTA4Vf37
tsC75QhVtoM2/lXCXASX0J3J7yTpkgiAtFIn60WTlX7jsuR8Ss97LLoMYWtUTJ5qJFajl/tpSQ8R
0ycGR4o1vwhmaFpbSHD/S/3MAb2e3GVrHWC0+LHLTO67XYmSKam0qpGola63WS2AdExS5lyppzAE
oBa5rtt/tdSu3SUXbHhv3NXgPmwur6pqfEbm/LzN80e7Pxoq6cRa1Kst2Z9oLXogx4qFzVLM7YTZ
2C+n0sbRr7FlnISDtuk4zH2zOEJfW3h+2i2vz2POldsUbvVXmPhJ3ezXTNtT9gRNm/u7EeGEuwQP
YGfubVMBZeY4KrNehmLg7JdBCUNSl+QTcV7YD2Yi0kP+G9e4u1fyjui99kn/RGRVyxLCYR9JQSTF
01/8jcgAdhaHAluifxW9yTReL3ihPIJQfGkfBFqj7CMZkBW0e+NDNtd1Yx/cIENB4y4xLISi7uoN
9qI61riq9HCxN8N1f8oAt8nLEweXINnlcfgTGx/3tRwzoERxvHF3a8vw/Kvb3uE8mdcSxHWu3BxP
1v2h+vAhoVRS/iFuLti+owz+8hlVNykOBYYRTkL9Bot4WSRcebrxNPERdnfK1L/Vc69QMlHrYMHa
ObRx8fJIHLvQLeztIJlLT+pqx1PiM4tTR9bJz2N/Op4uB+9nPHvFUhTwPcEmQy9vBiu5RX3pwDbu
fA4xr8kDR84W1O/Ev2avEdlaW4BVghOXxaVNvCYHG5NxkyPrEPNk1KjacysFJgnPzTSc5S6N2fY2
RPlociy6TvDLApJVs5fpsg99Y72NVLeV9Jcyja4Xh4xaVJN7hhzJF5t7Z8WRvbYEjSZURASxZlmU
sPMELGHMg/IEMynq1viYInILh/en0R/n9Oqdd0luhja5R2gtuZvw4CiRqCuNChlDh8gNqr2gbjNm
yVCRosmluz/tElEWrq/XsBneZGAopNxIEDA1ScU/Wt7JuyIVM8EFnvvCfuvCGrKrdnjUakt2amh/
6yVs5Ong1wdEpf27pBKkLGhvtEL7b7Dn0yLstKOk9DEYwkroLLHoXJ2tP0tB8ZJgGvihGwJDXZOy
GpnIjFLF3SiWCOC8JsuTJz6b0fyjPq2cq2LJKGU5o14wEU/dHG2jdtszctkIngF9UZl5sZsUc3vL
OAlHJBCMYJsVzlw4Jh+GJXWwkJ6k5FPhGxaxlM8sT6iMlFgReZxeDfMm4S8F5CSswhK6gZBRcEoX
EK+EjHhVdE1JB+IEJw7oQsrelcwArQtBdGC9BSwL1ZPtTJhjqEhn94fO6HklOJKp6P+v2UwDWvEk
c5obWcM46PQ5BlZmJZviECB/5XAf2sp3bHMjbgsITiDyuXH9r2bCYxH2Y6gvZFhlvcEiavjzRW3I
2Bp+8gk3gXvMrD0iUVU7MSW0K5SJKJ9zrALdNGwtRot2o4OBSoLwNqD+noU5452q+PASnQRpSSGy
0HsUsqm35tBBnKIAazS+5pKnoPnpYVliXBkVFp/UtP1pkatW8yW/+lpReFdkB+X2eRLZrWywhN9X
/IOf6xZgBufJiSUKoGVRdlsArEXauplEbUCBymL8LE1gS/y8mc9H0jD4wUsK9Fp2LuLBhnsK0/8C
XL2Iuaz20+D+yvqqCp/zld5ay6m80hbSjyVuXqNcTOyRvN+AiEnA/DR0NIVPUOg/lvm8BrRoUB2d
fvYZWG2uaqjBlWl+ax9Gy74PYbbYfYHV2lASjKj2R4h91Y57fQjcyKYw4K7kn4g9tn/bBHlxDs7R
Ck2RcuLAOKVsUyuTwY4sh450QW+rJV8/51NL2tlynOc07XtXtU7oYioKDew5nD1SdK1UCWNnmeKG
YZtYiplhtNHojH8eS+41Rf9wZ6PzrzUKSMY3EP0EMmtgmGPGriPSimJp/NFWP/MLKnDngGzGs6OB
Z0Dc/WfnavFWecs54VPNYuYZHm6WbG4iC6alZhcn8xMILnl7OuwDkyedfnzzNoDkGAYPE5oEAnDJ
LbzzJjIbUX5TiQAgNlu7VQl4ic2crIDspo+y1HsRizVgtlT3JBruKZLorXmS+HKHXQ+5Aq+eQ0y4
A554CBoT0uLMfzsTg2ov/9JsrfL0KCTRf9cxOOcsPtfMWWuEHeSVrnm9tUp5yqsGs2V138iKx/0R
z67tlZSWXcwIR/OyirPyKcRTRRKIBSyyoVue16oWtGWBmtkxD8p54cDwxk0vY30nBA8gsOvmvgfx
SoEjBA0vPMvB2+G8DN8OoIShvmPhCeHIm7Os69FY4GmvnzNoNSaITA1NS6IqqXxCOIv5rTLaJE4A
wMqk1x3A5rKaPmiFOoQwX9lDY+pP/Idvf8En2oqbtkPlOIbeQQaTZTSXLczTXaHw0GF4Uc28sfNt
jl9Bf5Vr6Te/mImoVxJ2G4tpnjUiZ3w3YDDlaWfRx5yKJocYcC0u2Nor6zZ9OMW2WPPhbAtCgkkx
hE8UEaXfaCI74w47xuYqrPiJ4dBXelpGnTitnECu2yTVBC4s0EFW/z0JEufPyIHkz1FZ5rYgjFbn
qNQQHNNuVehsQdjMODC5BS5wR+/vwzDZq3IQeJwA5DYwcqv6q2cNNgWzCfiPEawXgXv34uIVEAVi
5KCMoAqebPU4kOEsx84RZX5CSpmRwI5X0xy6JqnT9iuiKElQ5lZrZ5BjScBKUdErI0S4fmIT2eAI
lIbKXzS7b+jyyNa3aN0lghxU6jU0wTI6YOCF/5Mk2WBkdes4YcrNF23eekFeDzOi0UbLnZvUF3Tz
3LU+46r6cmSN9aaYaFER9EAz5hADNt6sgq9nVtuj63cpFYD1Rt31+udBvaFv5SWsfEf1NTA4R2GJ
+0Ig9PxcEMrXnisXKr5eM/6Mt/XyV6N0IFG6nlnUUZiUKi8WdZOl9mmGkGugA/V1eCHULfZcVk8A
CJPqw6+QIxRYp9H+U0+ky3WjvYAsKX/IcT6IDjDtUdlfXJ+wx7f2lx0p609nD8WLozAC6nb4UWbi
yitytD1e0LkPs6PHzSsO7t2+Rc25nU0Bt14IBInHtI57muVtt63A9TMQcXKAsKpzBNvDU4+i/uab
DxfRUUgwruYqlhJNsvoiyAEgXSTh1tPU7qvHN4XJApxrZ0J2+KFQK0ipnA4aiCvRUKkzyAx4iibx
4OaL3RIIluGXw5h93CUpfOtD/G90ypDsAuDcQMG5FiCyZwTOF2Ih24926Bckd1RHqhllScwBJHNQ
SVSLU0Dqx3I5WXGe227XFgX8qeM5XgLJjox6R8i4b3ipjMuBIy5z2OHDSF1p3vWIAYuQLiiMOROn
j7oauz1/PCRpeeQUaQLsQtjFMuRhJvOI8T96HHsQCmDa7yowz9h1pUewT1VcaNcU5E29weXD+ED9
d+NFYDS14pV+eZobXOdJMk05xE4HWx00cpy/CJbMOECED4NiBj2m92RCHw7gzUeEaZm3Yfh00amm
Z2mghWgxaardMGkWiO0WiZX+K3UiF+jWrh/rfIQjw/A5s/1O9eypwoIyfd06asHxw6m4SkNcifiX
JiWvnP4JXesioQsYBI5FVSQ0ulorfrU4Ji0wbeMysUDhRRYiZ2DxOWYvL3ia7R8UDD1M76xN7EXu
B9fFG9OnjByfMqjs+AiWe6/e7kKewZT9D3REze6CGNqfxXVSIvhlCZpXH43u67/K7QBhSmlps+YH
6sQLWlYSURZAPBw36wh2tNmIuylZ/197ccww5AJNb5cnkM5uBR4n7ZnFkzLDdBa49Jw8GTgTcQ6x
8OvvNJ/0LWLTyC9tEf/Ih5zAtrNgMLo4JkgUAukkud+9cvzESkaqPs8jXUY2yQl8fXE2mhOuGhA1
vaaiIVqS5EBr6YsSqXf/4sBJJXOsXKGhh0LL/kOJpG/zNnn1DVj4UJsa3ATcOEd9ZqSXGBlxuBze
0HBNdBI0oIMB4S8eUmHDKNOwrp6alVSGxYGWyCkxOwUzfDxwJIbrijL/oYwrDqAhRUPC/B1eZmqJ
e0TyfQeQrW1YEu+7qJmO9cWPKoPtJe3K2C1R71zfGwIcMBiNLB/Gih+lYZhpLBY3uPZ7YL5cYFjj
fHiehioenRFvCJV+niYfky+u8YaAVOk9Va3TC9wXMCma40wGVRJ0KDumsCxf2qA8WHJ3cCWlewaV
gkyYWyBdgUs81tRyI6A6ue6I4Z0l8+N3Kcn7BtA6FzcfWmogMbxbSD8k1tgdEQtLoi/EZM9+WMk+
uMrTUN4SI+cgRwCRoePgMMMkyXc3Yjsanvjd0hb8MFGKwVcL9peeaqGOFvUbu1Gj0R88k3i01WyB
Plg8B0JgQLK3yb2XOAU8bNV+vB1pwrgAAqg5hR5Bw35M1/XVyVQ41adTfOljmI+3+AJQO27nRh+N
z3+Rn8fWfiWldS24nsA3IwvllesclsYpfOf0Ef40zybePiooXpluXiRluWsG1S58Z9ZjbkqvHy6l
6rPR3it9dHZqkVJ72NSjv3OOtnQz5VGtLqb9BLvtGlczFxc4L5SG6OupmQaNJ90Upi8vYH96Q0E0
Oyq7974lmygn4Vy7XflTua3LPRbME8CJrFOVn6bIPtNAu1khIm0Yf5O437OWifKECptFZkpQiL2n
0QhZ5kU8dydIndpZECzjRhQn+FMvuoJm9ud7cNUNwBGAPHS8bP5DaQks23RqflE5UENZI4CWSujw
GyRfHrZcz1kIozmqTiFNxOFghqYf9gzOqzZh7439kdR5j4AghedoKsb9r6/o+8wwsZJXrr7p2Ywx
EJ2uClyOR60KeBMZCENP8QVBNyHXrlFxyfv9KBFum60M2i3R+myN59tijDBd+gmIdOz1uXuqbYut
/fItdpsUlrE69CX4c7FiClN1eSiYWhF/L/OvFUtm239SD0RwjjsPLxbKhLFwVbGFsZSsxdVN7HS0
HGPKKfLxjYjYdbUms0wlKixh24K3Y6GdY00lZBmuYnbpbUX3EpB2oOpbivGr3QITDGVnTdjMPBBK
789EZyntdQFN3FHrpNDcFli/rqvdFnPvsG3m6NRoX5aHZIKsckSWth+BVmOvNg1whYgGz4y5ogKB
2XG70uzhsxH/6tATfCbl4t44VeZlOU0PN50h7OXSEe1m3Qfqk8J9WHm0Kl5mg+bL0FtadoaORNWA
ipHNtZGYBeuLT/4qQD7aPnnW4OiGlnmX7NiA/sMt/eWyd++qiAPDLdUj6Ou20kTRUlmYusBPwMJ/
3ye0GsDBR5nuhOq3ABWsHDexTsRQS/K0WTIGmPlqQnoRrv4N/b1D7PvYu8dR9yZJaNfbXNCsI7Y/
tmGwEa/SZzbX7/cTUhFSUjeoFl+d4twLkfXykGVVMhKajuVWybrK0CEFu7FcE3skf1pZEwf4VpFb
7fyJo+oL4CsLea4Shemq7yu70gsdc3aLErOpvuT7lFzJDEuxyYPGzKUDqi4w7o/rmtwUVAJZWVhS
R9o/EOlgUiclpOGvpfcjNnYhsrnC0Vm3RAqdDQwqEC/vJwLSjLnB/vuZS3SDWKVFR1dJRbkn7pyW
Gcy3Tg179n8cei0IsbNRTldzIFYSROGdgDYhSnWtSKfYZ60hHGFGtv07RSL9bhf8TjarjyfNWIme
2vFeRZTHIMY+JpTBgouTsvfiy0E0ULOoZCem4V/tfuJsKSr0rbFricUPsaIMCV79NiWILSbK+UBq
04uEu4BjYC0Vz18fyaE6I1w2pUiszTEN+PLyBSrzF/HtVLFSwoz+54UsM8trtUmKALGBOJeaDXom
jDVKK8b0DMJw06IneT+GCSN9DvezeWaB/IDTHzqkeX89gKq/fa0MB6blDyYjdJn+T8AXeZHiEQWm
kNPC0PrnHqWVa1RKH6wTDfLCzbOsP9VPTNF7/a0wHD8hJ8+9RFpJRgNR+C+tDGA+egpfcGN6YScV
8jVKL+rkqBjRJ4/3DqeOtzj10TsZvzyigAYnMpTPpqygnyCAwdm4aKpCOZjMPokoT8e2bWyyIXW9
wQ1hlOmSXCOASGroP/AtUm+/tq09uNX+mLMC18daoSjL1WKhYKgGqN+IacNyLZqpkc+N7zyI42Pd
ZC+bV/hJHTz81FG+i8U02CHQu28qEZUpioheyS/5da0uvxqjtpU0UHdlPGuEWaZQUNhh9AtGKuJg
EppWdcS+WLPIc9NQ1kq77bR4Xdv1F391gSQMEazVoFswSK9gKS1C7x1HMP0ClWISU7UDCombGpLP
hyEGQAvyZa1vorqJyWYq1a8WYpq8Z6zcIt+OtYPaSO2ymsITfkKKO4GTd4nFfGPlqLVuXYYvJ6xD
Av7L3w3GAaRS7syNA2TlOI3rm9bT0bi9C/1oURDJOIih42YX7DjTAIqjYKrjmw7x8dPZYvVUOtaa
72FJKtghdkYbhkniFXDR3TE0GlDXQT+iQTdKFmuN1sEkScHypFmyfD6CWyjCYek5TLMHwIKEMCKr
gmSmhBl/7p2LwZcs47KlahxblSXjb9ObwgR4/8753iwJiPcgmAwhlmK8R9XEMUZHLJf8r1pwu5Np
EiD9Uaro/Xw2+jZ/VSZ2AZ3/NN9Lfcxp8ilxK/8ZG4KoU8Ae0qWnuO77arWu6IhPvo65wr6B0ptN
K2FgMTNYdJps4Mn6CFyMxDE021DBuNoFIijtNTLoKFlUp/06kOy/GVxNT2uhrXxZbm2PtZNf9SmP
UQCmtUhHs+bZ6mZuhpC20DJVXE8l9CIil+/V8eWUKAS69EeKOTbbzKQUF3mlE3zC7nI+YiWMYA76
Tl82qJfjSUU9ENCG610q0ItPGdveZ3xsYmZOIVBiT8hGtrtnlkikZlM4rTloVS0+hHmh/7Bqbi70
GA2n+bAeBOEbEKfnWtQ6F8Nm3tscZop2zxRjCu+SPbXjjmG9gdR0j9hilVwfEr+od4xYXQOHa1md
mpMSaZD8kr6kMWeMBgmGbV4UZQk/Eze0J3jezZsgUV7t+4gqBabMZilOnHlOrGE14oKN9TjXQjOu
ghl4g/CBS1IbUoef0qK5Qka0sUcUHROKVYUdK78BBl3XfDYLaRGUdCPKh9CVrzqmEBQjsxDo4HPb
qb9c0+B5RQBUMuY1rWT3YUlsDbZBPpwm6rTYcX9/T8lWLX7FAZxtsOTzJv4R6aMQYFLOru92/v/v
hF+cU8/gGsu4x4Ih/b1BFT/I6IkeYYPow16uQc/iG4zovidN0KKOE9hnrYW3Jpyk+cogzs6tV+j0
yuuzhOoJjxi42is4QsB5URuvddvtbDFp2K9pHymuViJgjHsYE2rF4ZXzXTXsIC4yhsccK8OSp3F1
oe8SF/HWnDSYRHPvtWMGVWVBSUT8l2o74X6+zqHi9Zs26NW6knzBiDgj8SKkl2Vm5999y+a5GdBS
IBguMbqVClOiXZU0rbFdE7txLL1GqAKbkqY7wU7MiL2J4H60dBKGdGzVJxysKCK3+btpKTD+8+cM
2vVQxrY+gRvG48b4zZgcBwkeRuURaOjPdjZnySaZy3B4ZR+KEPFOSLh17tAYNhXyARtbxwF8DZir
OudzTs8/I3fENAfLeUxsrhWbtZ+xxHSm/CT25s63+76ir012PFusnXLotu4XEnCoQnnYGJUODu3i
whvy3u9F7OzD+x18/X/p2ab3MJ4lQ/dw3RZN6ehVtpva9kk0iF2Xxt+lZjAv9innM+tC3r62ACwj
W0L8eRtP4BIZVfOE3R4m8GH4d1SHHSaGBo5IFqPo1XcV/nyo47IuCW7vlMSku9lAcUZ7dkWHJFzH
IOU1+dHoFzaJoBsIiKRkJ5Njq9tG23PUpW2UqAxRI8WejdRZNHIt2lyG5zuvPfxEUCltOOxyIPv2
5OGsDZe2B9DwI/ZkLe9t6/Rri5sFoUTDGyGhSC1lCWq7k/PFUmjWx28jlsU1XJgogOl0ukeL8Oay
CweUfhW6R62iN3xTeARUmJmCQmiu/gIBfzyBodtoiiJ3g15OAJhrnP5Xr//IlsimsHOX+s001yzA
iJodBMioEuM9Be8l2sWoHqZRobU1QSEY/d+iYButgWnmnTlsfiBkhIPcrwAOkbTVnZNeVdkYIV7v
3WWHT7y8NKKMmYhgV43/JayrE8NTZbVUhAm42FrYNPJjLr9Q0X2JYNyLC4LNQACijmOj7cUDQpAf
VQo3n2dlTT6hvmOVm1NSxOzzTJo6Ic7J3Sw+li5wTZU/xdIvMyms7p8uy6oM4s1q6T1y6aVV5t5+
RARtrm8Cnw7uMDwdC+RT/yYzRg1wjsJ/xF9K4bk3EPohPsUZvU5Kc44a3nA/6Ln3hxnAkzFoCy33
W9yX+ao24GEkWkNLpPSmGpc2tUWhjGulDeEXy/ubUBMIx2wQVIRPy2mX2s+JeUffQpW6pE7t7bYl
I9ERwe9ByCnQNTVY8HB06U5bgh+yMIPdJNIJayhlUcRzB1y5Y87XKLj15fg0if+ZtT7bDGNIyCW1
53h60rka0HZ9wEA33JzAsF+xvLgDh+X61lktADq9/1PTvQvp20+0UBHOPixvKTvLsKeIfE9UTxRZ
RaUBDdq837meU6KXpTPIGcyWuJyYy3L4OMcYiHc5M+rkFENY2GkdyeRbpCTtIMI6nTTmbzFHpz0w
jT2FFrb/YTXizd0s1Mqj/VoD42TGFkFw+P/HKTjU9AL2warZ3sp3JbOgKZOKHmM0ZIrtYkfSWUid
o9CKCGvb1eGqp5s48ULhk8Vq4+dHICHUzZAyQP00snU4u6LPaBD4Y5JKOF/8BzsapBmCVadI7f/A
DxVY4lfgY5eZGrmyB1507VWImlK5harV+f5eBkOwAqVFR7SJAh0kRsZqJeUnBitFU7u3us4V7ZQs
vFJmBHf37hx+9XbtLiIJp7dEcKsuybbwACkE0Lj75I7k+6e5NAM9hKihlNIjkse9+FE3DdZyshFv
iGhjLaxcCRGrCYQb0VaaRnPUMx1/NdPuiQu+OpXGmKpsQgX/5L03jBVsK0/fQRxAQMr7RqLXnN6S
Lh92sOldO6kzLiJGeBFNKgScMHTFgibe3Qv2johmmRokQEixE1K1CQLyuk0MoNa4JblYBFiU5hhe
UGBtcbFf3lumiXhPd5S2abQtz4OT/8+/qdM7nuLnVkdw4ES+IytCe7CkVQZAv446eovjD6cWBOuU
ABgvXq7HVADWal4/FzYyxpf2ulcjryuckp08JAeMZvzQ1+v8ZqRif0geEZ3eHBkobTnAoRfh4wHm
DvKP9/bQRs5Bj46mxXFW7N+jcyAyf1S/TLZbqAIhZ0zCOoHbhhBp6oGCM9ddcE0OvDLswViCDf0k
/n8zSB18eaPCveS/DeyWMKxs31mX2vJjef/aDLrs055FK1Lk/lsmM37of82ZNYleWV7OGqxbyIgy
fetdD9w99BGYaZ5ZBYldcG4UBcP1vRkCFWB+J7fq3qos1uOk4jnh9f2QO50BY5uuo/SRTj9goqrL
jwxoRR1VDZF44WCrp2hNRqQXnOjWNXTaqT4ASoxDuhA4G9wS3c64nfdIE14MAfiyZDxEtfeZLwJs
3mucLPx3vljLOD5q25tkDsE4dypAjxjLN8mXn7X0s3jxmr111WMD7mI0ETyXvH3UTfypRAXbZb3H
RAmV868V1rW18kNWSWz09ADZz3eZp15xvvgIRmCVBOT5+OahlInX0Pc2rSZt6zJA7AQ9VtlWlRzl
88xvOzWkI8oiHnKG1JmJxpdwIef7dbJIYEAavwH4psmJVFnMWTdx+DhKyYM1iNt5xU/MxMQIs2X7
J8v5J2CKBboA0AofMYaM/9XavH9K/d+7DxRpdZlldfFPESD5sJnSeu5rRuAYqzku0cwixywHomjm
SJ4csOEkgl7bYbz0nw1QFZ0PyNJafHA6MMu1GmY+YwCgtQGkMGAxW5O128rP1YacBZ+Q/ek054ix
y86BbQ6ygtbUMhf+h8SjAyCQbbi8+JrsYLk1bEi3eaOzV0L4Vxeh2ys8BxDYpqGdta9obvxSeb5A
d3BGEJ0AxoBZo5WvsCSrwtbk7Ah71ekuWGB8cFP5Mxu8Ld/6L5xq+7TaTfYLZQbkg63uh8Kcv8kf
9ZTWxnghoGCNkATuyX1ih8odc9k7pI4can4EqCrQ6ugxJcxk9Y/ARl6gGbKnsQTILHxSh+MCAQzc
uFB/7IzkYQ2owmby8A1IpHtSD1jLUG9iDKZ3kxBKYg7ciySlEg2dw2D3WZfhpS4kJWMspgCE8aY7
JtNSB/YVh8Sk7xaasaH9Dlen4QmJrneFds0kE6iCGZ4XVHW45C/2jauc6FdCS3l7OWNxc0agNRSq
5QYj1hir/ZigqiwZuR1VR2iiX2M5HjDIU6e9Dcg+mF4qTaj0X1cHh7rncxwn9HlWxROXW9vESAW8
0Tk276NJY0mQ2VKlLzVYt1zBAt4phby6aMDtkGGVuu23QJVFVUpcNl49qluBmAbhtNzQDBrUJqJr
temVknaCnft83lPyYh1w+A86yJu85DqOeEVLJsBpRUpHdjgPOfb2sZR5cf6PR9ezWgutwqWpKoTe
9qAviaF2arxHynuYPpaNafqcxNIxdpE4N4HgLS4aOlNNrXTm5Iati5GpZso/pieBnTw4m+4olX2P
hGv36XZyHIjFvgZWj8bAeGf/mEsTFsv7er+55Jsy5w9mZ6vyi1wzL1+eTrz9umu3rGD7Cw7de1uQ
E/zobPBZyw6dRYt5d9RnHw8XoJ1sGaqaWWtGEOzfpDmLrhCFPSzWn1iyl7/Y49Q0+289O0sumP+O
CIvHEkZJc3ZXbG4QsJ2LAShnV8Sg1Pq/rVfzwagcf7NaUdqk7juKfOqFPma+F/o9RslyxCX0puvW
cvslFJudgZWHwsj3dA8ohkI6ikyjtTdeJb5F8HURkaJ7jvbtj9aUZ9B0hqd/KACzGf1RPS3+n0wF
fQEVqCvKd4wF+IFRT0gueDB9HiM8Q4ULurGFRvJSRnBC9ubR5hCV1tpCzD+SGm2BqtSgRcKYlaYW
x4G41ATbBGJHMkdn+Z/o5vkuVxQEd3INHpb00cebLjhpIUeUiVBueuUt5Ed07SW5a0u+DJ+rniLT
nJMqv2lSC4bQo0euGNgahQXrkwFicWF0mwoXVpB4dJklvj7lQcrtk6YV66SPT/q9K3J9oC//iw6I
2rVsSokrUPnYiTuhnT6/l8uTW2F/WmSWCSXH1w9ttfOkKsZ35ms/gH7Tt8ASyudqpwQB8eWdTFro
dxVFEJFmk8QLNJ0RSxqD9btYGQueTJ3E/D7J+HGM3bNkr7PxLJbJ19/Rwe/KEzDZLvbMiZiPhxT9
bIo8/SlfJB880xAAFLCKfVj5YueCRFjayC85hkwAZ5YOw4yuno/wCVxKgWngQhSF/IRgsxmxowZa
xiJFSexPEFzELDOTtFqSUgabdCVekxCWz4jIo+RicR5K8eFsLOtqgHNelDZdAZTdkepOe8FEy63X
isv1jOQ3g5vFUEvoS6zQRllO/1HssGnV+RSwmxTq8fDO/REe1xtAhdBeU75Ny5cLoNO+7QOBiLZE
xGQAGbvztIRox7p2qibhqC/sez48vuRBr4P0iyLC/kzpmSO/OGGmzuLhUR06Mj2Qq8CkdBc3ITNI
AkquxxRfxtwJVh/ouU6A9NDx9tdxbIM82sNUlOu1//+MGOWIINuaTauxiOdlIsy4auVeLt9s3UGt
YTW2ehqZsN9YZ3PQxzHDBn70x3xucJ1RowLzWZXYujK+dP8p299x0oN+91Z2Iv4sVOExF7FPntA+
Ih3wWFoyn2o70cMF/UuZSGNUBDx8jO1ja36GN6jBkPaanyd1JGUcn0r54il0kyt5nAcroLz/nR2K
vC9iR2f2EFfCFcxG4baOBB8PcqAIw8Wu/tiRdLzPkRHTy8UTSOIafief0IYcf9uW+YrJDNF1CwOG
+JvYxxw+0IbmCYu1hcq6sQMtY2y3pG1PkzVtRnJ1lTFst0q3RE/IC4pYjdV/yDav7hjVCwNl4fjz
V0GbNEE+wbCDSh3i+DmwSIL0j1fTeBvuiBUQkk57mtVW95vTxnb8b2kdhcmEeihsYK7/M/NwPim5
1Mb3//t9kcg7/7WCfCjY1j2d9RiMNIA7svWEBcntgwnb8s+58xyJOw+f63MpfOtMMZsylO3NPb5m
kan3OfeOP8EmuRhlp/VvN6yw+Nkqav+Pfjy1ffxDhfEqmUSUele+9NcVjEvUuHjmkjjKyePf3z86
NnDsg1EiUKKL0+v9oV7/Hv5PbISvYWq8YesNMBXL/5cdfpDaV+K694sp/pxK2z05iC2I6yHK0evv
T/9K9Pg9fpbtS0Mcl7V3TSlz6hQMXJaCBnZqMgYvbzVT1B3zcOdZV1wa1VICYEXxaryx8GTsN4+l
gJaxw7Gy5pWbtPovlgpMeyqbTntKl4zdjxJYHEyAEkMh5tgxgImqJbPnk8Gzk9mGazS8nGzNYfWi
yskeMiB2iKvGILC/vRYgmNcLW5e/b1lMhESVyfZ0pgkZJOLVn2XIDfPWaYMS4cluiOOl71XVKy8d
caIFPHg9jmcwVPrvZo2fKXKYFWNRkFreSGULBL9fT7gcAsaM1bdXIUDqrdK9r1K/yJs9CegdqQku
OD5edBvyEFUwZUw2n6C3E3wFtdnwNYZbKK12QEUqYTx4tSKwKEfSrTEAKajVfrhHvO+fB0qQj4iG
1hWUOzwW8yZUS4vtnqOOhd9PMFfhvPTBu+qYbWVVfcONgJxHYw0tmmwlOs5Y75EOnQIA8B8lu4r/
VXhsz7sLLzGvnBpvMrBwuywdOE5EFMk5gBu78AR3upU1qkcwVvpWeyKVUeulfJ4eysEYyJGlRfCq
aoslLRiRFxabXThBI2sPAWEjipgh8wUc3wZPqcodrKbyRYXHSP2KSfoB98DwOXuOeEl78Mqvvp1v
WcomJ287ErKNh6KUMLSkIAbvQJ0PHgIuOZusjCaCcXqSGaPhisINRB6ej+7pT0fu1NvTsDnq8dqB
vnPMeM6z8kTBYrNyisnhx/OVfml3aQoKLOVYD7pdB8ZlvFchL2CynK9xsT+J6B+e+JvyK5QXyQIT
M76VHLbfylBE/12JkfxK33CfS3Gsmwl7BUfSIjHYzGb0gBJ10ZmfgJc6qdD3w8vMQbIxXqZXnazX
2zQ17USHRakylvuWGYGIMlAamyV1oXVwl2NPsol/dxHet5Ur7uxN8Us6PY6VK96GksqD32IUc8Nl
BEQ8nzQNcpx2+ReyI0GbHL80eJKulMyrKMcxrNXxAnHPdnjsj6wPPKNPQ7i/UW0ZFchHry7wTuo0
E5R008MLs5ThS8Jw2AXsv5rSpDhFL/FWcBxMlffiXPfDc76ZXP1gbOvtC3unXvPjs9vMKeDfkbko
OZWYyomTnFUgsdM4q/cJoBSOGYJpdC7vQRF1HxldxVwQanPzBvDo/vju7+qe15nGPEicGqPm69F9
pk5eptHPgOQufIyw05ZmVMrf8TRhMDH+zM1nUbr8ufV6jfVirlfloQlNXUWqQyFf4/ERgmNkS9HS
QgHbQpk8CpSFv7X7XflqpCcwZy2Chsomhi0ie/ZONlgngXlG/DMvYXMbMBbVsLF0GVj9zDTi220K
vdfk1N3/C75UOWmQMwdPg/kPfjgqkVBOqgNM/AVv+2ncW0S+HVn/ml/K59YN+Ojxy1b7Dr9yJRPz
mx5xrDcYjgYuRANUK6YRKRyY4lG3a7rZSYSrrMdtOJdlktVSMXIQr2JQFt7V87GCuSEuL2aYv4n3
uUjrlGVD0+VOcZZIx0YdkWYxcMpDDwMelfWRBLpVRZUtTZzhzd8h++PTTEhtC9T0T9c3X/7EoO3S
zTlWOfe2wPIhM8lPrkU1okFCAqJkcDqToob0BlG0Xy33n0Rw7xlLnvDrUTi0LnxMvDw+IiD0m8bI
6swwcM4zFYTcNusphNH2HdzR6F+tvcq1VMCpDhmP3hKD23/NEMPh2xTeuSBO9GoVgdeVI/XakHbg
Dx9hclqppM7XdvW/6Qx21/GMB/pilLckgiSOzpGzlctUxdy0xkAuulWoD6aNT4k3U7NVb8mpYxhu
XVF6SpVaV2xa8ZSw92Hi+0meBrDvWTBOLZonvXVFHvu9jDdsgTjga7f4+rowFfO6LCZmvp4x5FXb
NgrCaz59/xMB0a1oYudkqdtdpnjrIfkb+/zUZpsMukKV3J6chfzscyZMhSf+A6xC472/VdcAIcFH
H3XiELSz/IFRgbelY8x6BzFcPaYXBK9eiKZpi8DPvv0dLINt230YUv5Fk2Xxzc3NzHdvu1p14z+Y
4LAOZVvSTRWV6gu7b++fQUqXMlQhkBivgRKTbKhwXnojqG1bL9FS47i+FI3DJ2VqXxZQa8R2l9bA
5j53x25YcDW9/vdoE8552rUmRUPA7cgPEXJZuhgNbX8VUYrTUV108SSzHJgL6+R0NGs6pTn1vykc
EdChCA+Ro7T9q88pa10umNpR480+6JG/nR4+Nucw8mVtsxvr2gND5OrSzAwBd4gCXKRpUb02Ly7x
MLvhMTb+pouY5iEQKRJQFvZQtefpd+qEYeIjlHsUJeNt8Op+oAn3GfnwUeg5HOMZurmA8w/JVFXX
Pm5lt0Wr/KQB4UCEUPnh2wWzWVBCUcOvqyS6NzEcSpZ8ECxi00k0p8QcahbUMTwSOalnN96AcPSn
O6dR6NdCafSvtD3CKLx0TfMctolAC48UW7HCm++dBj8CkfuS4fYKIej/uy+VnVzAPlN4NXwXnqzR
pJt74prGOWesrWLN+G43RmoG/GooeKwhG/zNQDaeRV3v+KDlQL6pwFNozkprI84gB0H44AhwlFjH
aEglj37Gk9Deqr7acD8S9kprV5djlNKY+UwkykdH1ezhHugBOV9d687qh6zvM3d1Odlpo6IWUA6H
zRmwSHcWqMgeLptRjsRibWktbWu1g+W/9nZLmjVe7WY5Ma3nSRrAuCKU/YoLGxLFpnIVKwX9WGe4
A8j611+D0OMG70kkKcKFWmFRf0pwnV+65ui3i90Jvu3gBs7SRawsXNW0ZahQHnZ3EZn+9IQym8ab
DZtsiE11aq3wwVgWcSIJVskhPgLi+dcgmxzn2Z37N9T6WWYxLj2XeggjRG10eWCnlMo6VyGDvm17
DvYTWrPwFVXNdSIgL0aRbhIXz79eQzyzgEM4KqEgPbpUcTGDBm9Kmd7xzcrO0HbYoCb9M2JRrWYh
nCVT2OKFhjaDQ0oSxGsS5K+1tqebGBUM1orlJW/aQeXElfp/3ScYiUIvWcHNSUEwkJ8Q9om7GWwS
nkLYFfGee0WRcKSPX13ZONfUDiL7Qdn4oTRSMvlrFiOUVm7r/Ftxeq0h0GQfIrKCo+ahid4XsnWZ
TOT+4Y2dSnpdxc9MKbUuUzSvB5UhUDZjuz3+iIaIUIieSaSMLOT+fAXgcZUfImnssnI7qrIB/G03
v4WdCvg8o0bURS6iZOvUtN1+92CRQbXKwCb/z5LrcZJeScNl4hr6RfQOu+REqljete8GN0/+FkiK
ZjUiNlOnh+jYQszjKt8m1wzK4NSu6jatAH7Z/Rr2Wh/NUxjqYJwrxvZwHp6+TO4XEpKGd9hHsP53
Ry8+Zd6ovb/6o0biRWmFnROGK1aBxOMr1BCRzCtyasg+ciyIxe0RjUuXAcc12dRl3LT6YjHr8svf
WSSjhBR1oT9kD9gPe3QnriNoBFd4MMypgFWi6xucZbBj4/UXbC4mviVxAXB5waJaMYVtehxKFJOm
TUZ4o4dzq22ZAyIiocw7bqNSbrdOPZB9kcHa6o9nRhRAJ1AuLwAv69/r9tTtAO3/NV89Fup2IRnc
iuU+t1MoxADOnoob8qSLPBsZEeQRrqFHRlfFLQhRQ0itKaNvnco+ZPNcmwO+UiIMHNllFGh+fwrN
XMBxDlAY3X4BlrUjW0CNxqEilo6lxUYYNuZClwhVGOAlRukGwsAK8ijrKs7iuduhUu8a+HQaQdqg
pmPbxEVe4ZGkCaBZXpikH3UdJkLbKz+d2UfW9E1XYWmQTXG1wKJFFs9l1lIwqjUBWoF7zfLjOJfG
7gedm6nwhG9Ym3ouuFBVlPOWjIblnaXiX0Qw/auM8YeGbNOL2iTgvdGslH/QAjquOkky9RREGE4m
b5N9oO1/YF+WmBBwFWZcMy+95AG+tYwfGK9Vrus3YptaivwTm4STsU7XCMuwX+Sb7s9/K1rNI+mT
BnnmvniI/+4+REKqHL7hA498NPDqYD1OBl/3Fw5kAMNLxvSFM9y/e63y01WA8WlO4hf+RQahisty
MaRFpCen5A/gt+0CzpyRdftalKxmhciqv5mfswnXd/oH8LGVgD2q8Op6/c5pI5W/QFwMtyHcQMjT
WZEMCfO8eMwN0WrCLKm+lBvQwJ5TpVfUewlbcy7kILax9oWB879cj0RqaZIlaiXBIoEpWhaAuIq8
kvUuw8P3+Kj+yO72t5BRx31AKJCkTT6cBe9kiYyfsuc1rek+b0kH4dTiIrRhPfZvjerABQSzV+2f
SNci4rVFMyDHV6N7E7bkshMc7F5UckSqTXw4eJ0FsZFIzE2Pco5WvAQb79f4qFMPgIENPy2k5Wa5
tfQ8Up/vK+lMsgt/+52Lx815ur9gfXSkEo+3gG/j7BbPiIwgJVfEoRun8fr52lg3Lf5rfDXmnYCN
HJHp+2OQTcpzQztAxJ61v9RQ1YSlAiD91tROWTgnMMIzsq0RKY7fsEDN82YjUt/ZjbIr5Y/esBeM
XEap+YU8UzqnQBZCkTErMD/RmHpdLBB+1O+22edemYp2Ucb1vkBziB/H6WGhhK/DyqWjs5tWkrPD
KWAirEijrDhs/M6olGkiUa0ts8bRC8dJ0tmTHx4oFiUxdFPabw7g9YXiD2bYmHG+DUAIpVG+7+cN
1W8/8dRJ/KvhFu4TGAYme1L47vDB4PSE+kB92CK9HpvUciEYLPlhc5WmWsB59bv/D/qMFaoXTMic
elMFLYP+xEiFmTrNs3CPsQdLj1QxmdfPF2c+EOH8hxbmSqb5TLFmkvJ3naAai29ArQvaQs2QgiY9
/j9liITUGdccMpdUFBo0nMrOYVDZg+ZLODpg8kPqv/3d1PKz2XZEM8napmXU6oOYxMfUueugD8Tz
ru6i9TGjy/RPuHNM9IPrQm2CBzhV7pjts80P2ljcguAPAZea1lBPwU19gbBfmqQizxVji54J6N+8
by1ovbOqC/uAKhDzgevhRWhsn6zA72I5HEU4FZi5MHQLRnZLyNvadVrYMuDHC+wmWFHL+J2MKD3W
L7NpH7Y+ddEFBDy8UBlX1xvYFb1fodOxhXM5DJulqaLdRec4oKAUGNy2ZKLUlNcuwC3UJmRJPLwU
EmmbhnfH3Sa9ahdCq/RN0wZRIamoregL11lfbWdMe4Y9jkeNI0oiC/5B9jZD8fCOVubFFmssiaqW
qFBrgjSjJW78TWYoSyo+8wEW31sdWLCU9XqZBGZboD3Ge5oOpXTw6uZNYb9aNt60IZtrSDpZxQaw
XRipRdVhFIwrefgREvlm7YatI4+24THvoFEzrCCeRvP4LjkxoFTjttywsgAnA3qaIvVy93QnU24L
JWO+ozTfR3e3ckeENXq/LeARcMElRD503H66RZ4oR1Bt5tP+SeFLjq2jiyGSARXlMqpHrU1ef4mv
yU67UTaXH1gRY/j/RjSs0XuDpb5DhkHIGkYob6YtkLKUv3iMKDqNFWzArxmmIgS9E1f6cw90UJrj
iGk2sliymOTuYOYYBjhNOzk99UpNNp0vBAI4ki+blQ6XfoBLG46YKNBZPYCoiTKNm9rB4fiX1JWP
ErHmrNHF8j1EgS4DkBz7Xan1ubIkAiwAy8773AEF+75bu/q2I40YXUNCsP8Pckpjgg14SBxn3TP+
UAsfGgKh5ZTVsFZ+xQ5wfrByTitsZak5Mh+3uLvGHwnMyngvZAOFFA5xI07bWDufd0zxCEejLB/N
LEmJMD1SjYaM+XYFJp18pqHBroJigBiA7+w+BUmtlyewAQ3Ij+6LODvuTTXbCynEU4JxsZg24oVq
nRiR4YubbGZQP9hbl/0OafsH2uLSdbfGCcgOr9oShnZDk03RCRurNog5fc8tjEJLmQJ4N1t16WqA
Q4haWcNW0x42z7I06gDwU3nEcqJyR4PC7qgM0Z12vn0RhwvAlhCEdnRskJqy3ja0A479wCSsW4Z2
YtpGu8rsRhSQ1CBqAzB0PldrgDyZkFTCQPfM0Lscc3qHBtcYN2SCGaVJVOTW4ZpcPEkE5iehKJEf
aQ3GPj7cyFdOHA2LFjANFTSf6td1eirW1+rUYm+PzKCnJLG+dOBaCGOEuVXuy5Nwvt1V+Gt8rz2p
bhhC/YVlQIWdpxpZYnm/3TBuCTuVSd3mFxynlRtm0hZuXvQxer8whN8oipwt8z1YVfGR3tgc4ERW
tMXheJZhvk+nYEi33cQFqMXiyH/TvY9ypqFD1PG3h1DY2TkOzaIYW4/dCPTj4KXdVAsww5t2bMEp
qbdT9n6tR5dH96lHfc3TZnxunS5XvsjNR1eoqU6XI/yysZrT3OQfpSH9/vXbng+GntsgjbE0IIbF
Fm41GPvHpJIKFqzlXUsJaYyOan0B/KnnV9CjHRbhd8IwlgpC391bdjzO5BiBEi3j3ezJ4krb7XLS
byMjgwnPn0KqVFOm84K375BMslXVrkN+LTYK2YJSGxvMD8fNp3MQXszQg960qWeNsfAV49nBZr/T
+a9L+RMWKfRNGnk46bQrHKaA+DZpyHlxEFBc70a7jAyAbSBpzepDq0QZjXTssw+DWSE4TUEaNff0
uFqNBaJGzSqKGySbRNuefmjnx/EN8Pt83abAYGkypZLE0gTgr0/qjKTmZFIEdSo0DEBTEcPbw0zr
z9NTOSTi4jvabhd1JreIMYgNpWLspK44h5IOrU0r8u9JLAMd6yHuyY+K565BIAcgIyODKLCrPGY1
h9DXqE1dyx/oPPRcdYehZx2K/fYUyX87QqnTLIR5vdC8If4SwSE7KxXFPEeund/cZqlvRc85hgZT
FmK4KxKnmTNKGFGWh94ycUENHYzTi1LBFVc/+D2xWNKVqSwWmP32NOaOzxh1kxrR9mVA5eJNXsDj
HAl9c3FE7WIh3lUIK4o1utlJ0OuaPesEKlZXdPEEidA9rB7FjbUNIpdXb1t6xjtsy8suhzLNx9pp
yeLE8owEpacp9gtGAVbYjUaM208pjBeIs6GbBi4EL+yAw5NOiaP13gEX7UoH3uBgMocIpQM7kVzL
+RQHQBWJsrlHfmUalq/fPeuEdopRLUL48Iwoii1k5xAQfx4810+dfOVnvNLILwK3e6JSpW/3pgzu
UwGiCbK4SYNai4jT38Ae68f1j1HHbCT+l4ucNUgi18CdbO3JSBYUU457SDsY+mgX1G0qYATXf56S
8XL9EUXBhlCwAEm9QuQK8Jqmo1d5ylvD51e4PXt7KKnuTjLCRoWBt1SzNG9X+nXqb5qZirkj8PcJ
UltVXzV+OafFPw9wWWajeotuSNH4Parzg6H9/8Y6Nu6ZnxV4vG9eyfSCAuJx6Y8dHwO1F+fGHpex
etwjOaLPv4YNgKtyaBw3LRLD9cNJr6GnJfGcblkKQOADTch6E9EDH+NhCzRA90pGtY8ismZvKBqK
kTKbThAjTO2U6VzWdKHiJAfVpKNnGPwicdrIOgA8DccJFQJywvLm2sAREV7E3wR4JYiDBXwgbeil
dfH71LMb7lK2FbTa2KjHmq9xsYgSVWzbLmHKJQ/9Sut72N6LXFcM8t70xyAWvQ4k+98X09I9xWw0
q7u9hs7i2S7Ufw1eZ089r98+2NQ92e2GB2yed2vPs2lEcPheO/Twivf8KG8q+H6xCx0pN0cWrq0M
/y40foTqN0RuJwsZ3BlPjtvI7peAwm1xbBb6t2YEC4DnqhK5rYhOW47lwiL+D+bOMiSafjOAJLCU
S5msg6yOk/fChCnDOdHrv3HB+r/mpWBa4a856JuE41gFNadWxOawj5zyRE+vn2xrSDgmDRoHiTy9
ysH1YyAS4uMKRK1LcXTezsA0RHYGaPJNsj5oe54JRJouyL0Z6bkT7XM93PAwOzsfxdHMzCMrRy/Z
LnRFU1cTdgCgC2IrPnT+EoQfKTTHBWhdnAq6zAvGmbskJ6GnUTuECOs1328uOHmCWlffntSegbX1
b6HInv5nmitEQTPoFKaPeG79bZ21Nd+USgj/lO7QN8vBHbG331We4Zp1RIjbJY63wI6p1CRiRKjQ
2aM++XsHvar+n1S6m2dej9KYJhWsbwCT2U7j1wmXIyOrduF0iZfsmaY2UkDpk0KAcdHpYOYsz2X0
/9g425aUvVN+sMJwVbakvQNrBQniRO0e7gvFfipxFmhKDMZQ8AEYjJh+g5csbjQRVwcvbZ+cU5yN
f8gHUd6YuVR2iTZxuBv3SBUAyGXw9XYqKNyoz9I1IJPSjXPOClyO1Gczm9ptm0x2wvpAkcHDssEc
JFp8icriBTg7Xb6hi+1qDZo7AaBOjDJ1P87+CD+KJ65x89zPvZVm3pai5UjIGa+s6Iqm2yRjyMxt
XMWYBgOjGCJDN5HJCcAK42R07tgueYdV/nTrImkZlCi/V+VpuK9OWQxVts+9Jgn00K67+YRjSZFn
63+9whZ2V3nOOSShs9HiOzsKdseF6L/O85qL/jN4L2GA2V4HYA0IT+ZAxBhVBSTyCMybOFeggOmP
JS3vQYDnrYMY2FiA+dqfyXsnQcF5IHf7j5AV5Q71X3Y10uVes/Ap1qjezQcw02fPwrUh5vFdO1B5
XsYLPNkXWlGif61OKYPPm3HhN25M1YIKvlPjw40mTL+bA9LR6L+uI0rY9aeJpH6uXPiGKZ6RZT5x
9qQ/dMthwt3eryhsOdkJtFmsXS3qluz0iFNsy/GeW3Ip1+xlXpXmTKVpQLKApdP4HkdOELaM5Hj/
Hhb1gCzzs9kNTYDj/mxiIoHTH6ttlY/vGlHqZZige9sP7ZOO9QIpW7fYYA/TAHKff4fyP5xdLDEy
suH7d/EK3ctN34DOB419vD+BbWpb9KFNDNGHQ9fhYzHFsinXTRTZtZrkPgPpuTSgPzOV+HFj2NNP
v4Us+UA6V4slSQmYaZTENI3vo4E3g2Dh9pno9DNptqiz7WM0C5Xh2eu/gJoLIMfAlNtYpvcE1qUI
fykHTwPImSdmu/zwi620oT9ScplBK7TSaeBNq/w+EQY6ejNOr2KMKzmqG0dCaIImynpxZ6VnWTq5
mC+jKsSulcmCrULESzSJ0NmZmDVm0mzzMqByaLg8H6FKpqCdbZX99/sib5KgDxnzULOtM7z6RwV4
M4v4cbDt2BO0kP3gibBvQBOrcauj2oMJyGn/k56DOzflgRLG3bEE71sV7B7c9ZWFEPtZQ2U/OTJf
/WqE+4bbIDyQSQPZUAXUoiEzCmZb1XCP41YS68wQlin0G8ri9R536k1IgZIpCfXX+2UjOr9hCszn
kdREN6dSxthedWp/CcB4RZvvKvXbvSaxe8YG9NpYjGES8iSn7ZDCimV+3HQzR1ZKhBBkqqqm84Y+
OSe3NXD7XeGuPU7hT76x6yGGDUwW/4oeqTAW9ssGFtZxOh893NFC9kYoqUmYDViI2IP3NT6kbVvI
0egP7HJQ0u2TRdBq8RpIaKt5Jbbg2nsZUThjUS1BpVoguZoIce9SikSuVYM1i/3nXZGwCl/88i1e
ofkW2XITpE+nFrYwTHq0BFfemleqxFBrXrg7OLF94fWsPJ62PXvCLEsFUc1Gry5TgLWQUjjima3a
oC128GvQZEqKoCk3jVr81NmUF+yxkPe97/W0DljwPODPJ51paJ16ftHyLvt5x0Xu2evuE7UiIhZt
cpvEtD2QhasXSoxvIlPXcS3DGSCCszXapcheH9EPiIjusTu/OIxySn2gcEsHRiakoNwsWH7rMC6h
G3iqhzT34/emr/7VUylKy2FTrqiWdwGbHO0kAq1t47HlKiw9MhldFzFfpkgMNr8j3LQrJ+SMSzCo
p5H3FHySJ0IvsUmqFvVJ+Q4NVnqSk4Z8BhkmEH8m7juYh8X9vU0hDFg1lZRhQcpjl1keKekS0tne
D9vZwRYAvh9tHh/YSsXt4iOQJUfseGTjeVP5w2/yb3yaSZRXPilGB34iOXs7mKnQCeYi71nEqD9h
OsGx2uhh5wISd6k3x+BiriLoCUiYFbsBt40KJAOjaNguJAwmDb5aK4XeWfWSYgT0wiLbzX2oDMjY
QvUlMeR5JNdMmrM4VieoL5Yg4yPF4bDDsW5ZQ5w61jSNulEFADSwOma1gc2jsZ3hjlUmhlBgG3IN
Ox2w4d+G8OjpIeOsBw0LvRJjNcdPkylm72ReCb/zWdKQr2Tc4YUeTUpDnc5Jsli6Z9xNY4XSpWeo
xEvePBQRtFOpN8Mi/q4n/KPSXc8Ac5SuvY3r4YTC78P3E4VcvjHCJ0zlfvfx81YWSilS0hNzaVZp
2LSuJ9lCaYX4T4ZWoegjHNmlzUZZXYtEg+aOP4rKJ4FsgtHRumcPTE6PcTkBaZdOeCCyTfLSynSR
jAZPtTRcFdbVaQVCvquyYXPo3ekOmgpAyOIPVRRg04UG761p8lYZUaZ3fLj6nDE4dOurlY7cuwe9
oHJchiDHloIavHJjSA1n479GRu0nYNV2NJMTI7+C9l1MebfEQBBTgRtXW0jfWkFKb+V6U9UwMzbH
o8M63uAIgI+3dkkFVkepXz42ybYPaSAFDxc+fWCE20FOW+I/4sb5rL84zy+UNERnUUdFTVlatppX
dVDeKeWRutXwyJLhR1ZjkxIrdBTQXaR0KPSs9mmqJnkgQ+4At4jvxvzcWE531FN4bQH24JwE/ZdC
Xr8WfMQIo4xWelWpfob8eskTj/LSCXUubx0P9TrFF3O6e+rmH7goBg0pk0TbFKQhCelh3PGcIANm
9ZPoJpigJb2G97iayM5Khi8o7qyxE6gBN8h2I3NbwJBbdZgj5x1zsbSS+PVR9bpvp0pxYR5ra5pL
adreAjTOX/LcaXN8T7D7kH8s7MwhzCnxqwq6ki1w4TVF6NCwulZyfMWmF0o1ihRr6uhsYxHHAYGn
goTr6XLgGUnc041r8+0dyowl6v6clhohP27neURItT5vFZDSJ8ueWmgV6unXBJoO08SY6jWtcOuE
OH9j1n+8TXEbncF4XYRjHKkn9clR8Cv27uwJ56PuyaQDY11mB0cFcrnruHA3vRzrQnQONDRFdyxd
PuHtJBvImKemgop+4ecsAf6iNuK5rfb2x69847Ihy7ZsVcCG03tV2qmt6G3hhdm6Vp5Ug3CROlp+
bvnDsL2PDHIECkN0Y/OlDkfbujt7NA8i6+Q9z3Gam/jL9zq/9KJFwJHVJPOD3NvlQq3HViAiOiNz
OTTV4wo0CLodRMtmMUOwLs+prg0IAIv4+J6Cyu1R9B8DrnfqriL6ky7bQBcicBZ7ve6ZsCno0xfR
veZQJxckbXeyZC+yM6/hTNo9IrukGW5A4z9juB64uOOsQ5EPRH/wq5QMH2qluTDkHUIG4IAEvtEu
SylNlQoVf81TJ/8RTrKb+GFqmCP7xQ2TKSOwEPBwz4g/IgW99UrA24fZHl65ZcpNM2wF75EtAiMd
uiiOPZJ6MR7Gw8moeNfZSW/sa63CH+h8MtxMGopRXdoj58d0NP0aVnNUYLSqCI2C4/vSiyewKpWm
vzQAYXHi/WPX9x9MhrAMayWNK93BgOjrgwACOCVoIkvDgnxAbioU7IUVoY+qGdzlHGL1u8b6tKsl
KhHCw78oTBiuYpQFf8dO2qNC7khODJVJVZqai2vTB4Dtuah6RRf23gw9WpJ7ltzeEzfIrBZC5t/T
9omWXq5ArYp0Zi3AtugiaDFi7sq7Ml8/nDQKXO16WWi/OUI9VXYKUmsLlV4XSHzRDJJEvZkrNTex
TJomQCR1HC+p6XqQUq73xzZUO2B3KZZtIIZ/ZnjZSFhj32hrjZIXmXjR+Px0UFm8RGhhnVqa2wbU
oXTwZtx+8c8R1MwDyvTRZ/SMgeBbFynze2hj5oEoBGeiFMmXMTAgohZQQGl/qS5FK/2exVT+gUiZ
crjvbyHCjjm4aBBvTitnkk6E905zNZ/jzH877WuBiC82nObnnclRvd1+aVGf0etcVB/ZsICoGEyT
DaTuG57Nde4M99sAcimVsV8VuRJ9mYs5p7moErVGvGyIEj2nTbeO4sJdv4g6l+dsB6H0TqwRkhR7
VMQ3lk2X2eTilerH1EuBi6nDDU0s+/wYwl6B7NKzRutAN8H3tsFkAa2lvbGXglMr2Kk3sTqeZ6gs
sUR1EMpOmfMmwzL4z2jAbzabD9HlrPIyKEVQb4bolzMrqSutdNtHXxybSfs3DVKAnkKv3inXYVpC
KMOhjdHunYr65umosuyV+N4KR0/5BPRldk9uYhnJqIRPwGdQ9dfZcz77vbZQm11TpD+XuJjH7v9H
RGSWc5rw8m7SLuwiMeCVs5WuBkkG6Rz7N50TLAogA/2ZShsQUVGuU446QaDeuyqqbinwyYoM+9rQ
ECtqwqnp3Zw3dXXVM1/CSFirDqQmZWGq+aOZbs46kTvUlDZ2vz9S9LJFyl0QFebTMZCHZhh/AnjK
JWiB7vP0H1cnPEK6o2lUrkDNBjeGKEAA5onAwSRJ1nTmCBgA9x1QIxP2n/ltgC+6Qblwl2mqoUHd
vmfb6ERIwQFTfhu4O+ibZQNHqN7L915AFbb+mRWkiC2P5oVHVS/E7kmQO5GPkoFgu8mrFpUl25h/
+CYEfJRuB42T+LKL8sYo6vJd5jxrI8lgPHXNAT02asESStGhMApIpCzPcF7zRRqzK8aSHRnVeqFk
HBAh74e8/jhH9F1Hk5ZDxJd26aQP9B7uymulfp5tHCeCjw/lh9d4621oqvoLMDmOS0B4ed6wjYGk
rGw4pIV5Eb553V22vtKNteVHotwTCINak5CNcsnuLjlicxu97H8b2fkPNHQKjwFI/VKEUOa8k7YD
4KT9lsokOUKY2UTOakUVR3Z2tgDpxu0GhVsGo98CAPACE46dM2orzA7ddhemTRWKhYeIc+BUnOfJ
vKEpv2dKkNhu6i1d57jIRVW4RgEerqjElqkBMmc6hODcKXHLmhBYFlxS2YmnhOTF0+wYS9+9Ck1R
yVdR1Z8Pdu5QAzZVEQpa9H7SBYjW4W/sfX8oxPoD+fMU7ilETOGz5K5xZtmj+ip6s+cbxTmWSgru
yv1Qxj9qy7o1GeDXwZ5KCu0nFpGf3wf8tsv/CmpUWgRHqzDnjngMvAJDe6ETcGEeRBt/NJon2y/g
jBKZomj2l/an2xIGORatbHezWGX2yx7MtSEKuqLou6yMvEwIzu5beysVz0XdG5D1QOw++xXngA30
XRdBt8TQnKC19q0z2xsXWVCPEEh5L7uCQ3W2A/V5JiMlnRrZhTPoQTG1zbauAus5SwCRMn6hN+sk
urYdMf2NNC+HmF9c4L/NsYuDlce0LEzSaMdffKwV1JdPXw063ZokQZsnoyN8Yl19g+c2OKwzGobC
ENYtEG3kQonj73g7D3GU0ZjuuBK13tkF8d8perkRmrC9GU/tnWoMBxr0aWqIb6iA2DqFpgOse1FJ
5ysMjjeqtU278gvvNJwtxE0QCBTk2NXVldCpKJ8ZlrGJOch2+Xl9/3gFupExvbuX7m9MhYPEdMzL
v4FdGRK7ndZ37uk6Mrm/Pr2O3xgaQHdTI8+rutNG0Q/VhpMydfWhPBVuZ5cvPK6MdNQGdkIZZiyu
62w9pGwdf+yw9XqDnKHLsXADWvm4y/nFODvh/qmbCf5E3oiEgq/eKgDkx6eqIVMTCeCmCrTKW+oi
/wk3FL05ku08W7EBr7NUpCIWg2dgSY+YlQj+hZqU6dw/3JIW2u4kNozAdhOI8ZrhlCeghkLssAqE
G4dRjJlhdAkVBT1Lweq8R0EsmuZo8lQEbWrsWkChH870BpBa3AeLWsSO9RlBnC+TgNE8N57qZMVm
rFNqHTJkj08OXqRbsIe+FvSsvBGSJM9aSKEPG5ejUeKZ60yIxQAZdVjvmNyCmGl70gXLBekPzG6l
lGBiDsIE/Qi2CsNV//DYGP1/01V4gZ/yhJmM/5fwQEY/GU0qq+1/HM2iug20hOwuYFv8xQOF3C22
6ElVCM5OPUtJ9ZNc+vpUlBaczjBHWhh6z1cniDBvE5U2MqyV4CCNPS5YOBcOD/6AwXsVRqRqFp2j
2ivvgHrZnLpruEou9U0wNF383s2M89LoPSsUgutZ48Gj1QxyEjaBW70qLjBUxj+bAwXwBKOomhjf
qfJdvZUsWO+ifClLK/oezxn0hkkAz+5MlqhBIcqhYwP8CqYM6mqhNnPmaWVwbaLPY8/94tU6IS6+
bCKEA26FVzRBP514aBUK4z/62eawhHdu8Qgps90dh6JTDu7P+4SjP8R5mFKaYht7Yh7LBL/9Reqi
8j7ZvI2z2tkeaKqXLGTIh4kBZONdG0/eMjKp5mRuK76Z7M8/VwtIf08CeuUYg0V1eJn4ukrGS+tO
KQ7E/S9eiU36N0Zt2ZE0vaq9zLKz71tOx4KaLxslDal6+EWpUyQIzuU2APtEqrvlRpbjRVK92QGn
Ba6B58NaAPxvsp3ep6PB3Z8KEgWSSKW+IUxe4MYK7kLLN8iEhRruqNMadw9IBFdYDdY0vFRb0oEq
zZ/JE9FOwILN89ffAwuCwMA+TYgHJiVKEPfbhW7ZhlID4/ykjpEsJ19HWEAHEMpfBroOhsYEFa1Y
d0nJhNAD6CQj0DDc8ROH5beK18SvcNUGBlcFT+hgB/pK9WyicXY7eN2Ye4Cb3xU7ch6y8eKiDxPv
2hfjQ3HwivBfw/x9bfeks/gS5EI6BDunGHhyR/drUNzK48jAWP7oMyRm9KVnqj/kuvx3YHKqMqyB
cCkD5wLdywapR2YS4F2MOiJPMSwG3ZUdx7vGaNaLHtfu85K3Kma/O4g9R4Ubf+WFmQvbaaryE9h0
oBh38GRpNaLmgsYIrHGDYS2ms2Y8WkabNfW0zfyrQQC8W2ZU90NO43kqNC5QjAQ2GDwtv7rLG7p/
9yfZmKkhp4YKzHnuRwGzpJXaWHi58HHMi73d1ijO43U04/sOUXFRp/k3pGcXaVcSxZSZ3qakeOnL
EkoFT5f0/TKvPKhy+llebFJvGv+XrBtCXgkeB663/S7miXWbDXHFA4qeUkHTychShBmkEOzYIJWZ
MaKss0XSRFDp6wydVzGbKi4gv/Nwe5YNqddtci7/xMqMqoHJKRzifhJr3B6c1QqUqv3btH2Nw1Rl
pk/k06g2N97kpA1zzW3sLRxvlR2qKQTDPn02fp1QPegv8VEJpAI+LzTt8lWPA1z9nJK10QwNkd66
pqge8UVJDHeMJ4jxAvHN+Tq6BnTh5aKvM+eSfwznqgD4FXDxV71pwALmJLwYUE3c56E4DDfGZqsS
Rf//4fzZYxu6KcXWAPeiRD3BLDyJvwEh/N2IOCFg/MEoTaPhax0TWhL25kvVX0hH+ehStd+L2RiP
Fn4HQRb2d8dkC1ZYNYtIRAlM0bZqwlOLQyCM5zIWeviXXWM3RTZ2g4H4GohxN6V39B0yNJo1SwEy
qghdVw2vZeCH+ez9NkusG7K653nbh3lcAqeC01nMEF2dIYbo0D/I89hYnSxAWnTAFaCoBGb4aPOm
7Xv31Z9DGDhl/FwY/Fr+PABuEgjX/i1fmpAQwLIs1kAkeKmUfQivukjdnfFiycGkhzOHuX5TfBO6
O3q/jpyFAPCspnR3sM41MoKD8l2h5xWHjwW4EvnzPBmgNHzJQpYRqOnXj9y+Oj2DZBFldkDrfiAG
nH64dsVuyNF9LtMMk9CgHV8J1s3esZWZhCrVKBp7pu5g4hflxvyIsTUqI2wXEQOYotoAPVUzk0xh
8I81Fr8RCivDkmJK5UY4+QaAfzTVPJDo74ETSWmkiwh9H2tgTRMoyBhD6T9PV6cR8aknxXysisjb
nyf/2cRo0HurfXmTOCLLeqYCWkYhS6kUtqY5SvG5j6s4bakUExAusPeS1bm1/mhDm9sGNz7Ukch3
2oGriEXgbgKAqX9coR2AbwmEFDnOafd2ZcHOA9JaE6k269zp0MmVZPF3lZIXa3kLYKl+jBsPd1Ni
DbD5GwlB7X3cnkCv0y3yPcMqoQgCGlB3aE7DgsMtMk5ybiKOp2yqcttXM/ZjPvuYrUGBA0ZU1SeX
bhIIlMppblO7FvfvNDk5EJ8AYn1Yw4HQX3n7JSRiEuFmjGraQeDgghmQtZ+a6q7lXF+VMR6or8KO
FNi8r9i9VDQvdEco0owYUMD90NEnLOD3dVZ3wzIybddPStu81LFi3Jy0Qp7iO07ZcSixQroBQ/zI
hOxkhN1t82X1FurYe3wRc92Q9GYMunTenvUipkdFb3uSn6F3YqaROJkW5ptW1F7SL5fQMwWjJA9g
IN6lSgCqD/eI9Tc6GkewWMb0KSULykncdipOq07G+g8tYH1t3RzQUBn0M6f1Xhp2u6pKDjLgQ4de
NXv182BdYvc52NOz/jnnoLzw10m9YQLAzOXKEwFoAp+yrNiAduKhT9S3wLne6/WGU/yqkJia7PQS
bMD8O8SLUs9btyYewhhJus+0WGwa913r3js9aWvXwO+88nF37Gwh4ChuMs+PPBZFHVoVNGbr12rR
AlF3eV8UWwKkDGpPd0elItqckYC5AvEUiFUtFbSx2Irx/2ZiXlSsgNxHqA6ZP4KOZ8PahEoIDe1h
KoG6IYjLY3UX7Gu9FR0pkBhN0S8b3qSbqnnKRN3u0WRSbaVZWqddObzue0FdCpzkbrWyLwG4Gtwv
zxvM3mf2N5w1RbuFfjTWUGzTdEHPNwm4PgvLANOBOrhIUBJN6I1evu/4L0hOMUH0uXvfKebxNUg+
LjPa/VM95AIg4gPL/mdjvpFTsPM+KP1CekuDhgS5mH95ZQRmBQqOGa2ZJrdn1xf4Ik6rQj1sE0ns
HMD4Wg+BjQVWDNeGlAWIa7+G2EcjIMyreKswiE7DO8Fug0bKlO8tK4hqeKXzjYKC8NXplD9TxdT4
UnpvSIQDDljVVu1yl+cUfcpTNJWxrQLooU+LKhSp8UpZcWRkxXrqDwORuFtX1Zw51E50B2dQbd86
50Dw/poiI/R1NvPiF+Jqk+LI8+u3p5wBOQH1dCGIPhrPgtBJxA7jD8zy3ZuSBMmogQEAlUjtHlZN
CuPx36BZKW9mlX/fOL7b3nCBZShi8fAQHtWGgMM7HYdOz9X5hjKFihcgV7eHSE2PGL/epDtQzrVO
HMarCCqZ/YNTIz4pzsbWb41tpu5C0Y6MH+btw8pbyeZaLU4iB/XgxVZzTRngdxctqymFZXw83/BS
lehC6n2jegteOJp7QZOy8VEv0w4nPsY5bpP4wc4tu3boRaoFhvn8Y5njLnMfY5G5InQTiqS/V1dv
Mq2em3NyR6K19IOR8YRvItiCrtmwDFnuJvY2nuBofakmni1U3TV3ujWxn2A4phWeG2ydEBkGHUwO
NOQshaqzuccYLIsc43GWAO/p19v9EnasNkqyFk1FUgOmbmx6yCtI1+7v7ax1o90JqNkWK5bc76Kv
Z02ITkMgds4LizRl2f7aYXqdVdl3sEGj2Gkg12rri539h3qCVB0vtOODSG1y5dBb3KCAmBlhqwCc
VABfbA5xKKFFwY2fdGT+5pW8FK6W8tQz3hA3zLo5HZI4SR3/IQH5bov+Kqoi3xXcQ77kPLNp2+Th
nUY769Q882DE33Fb6MRuYC0De6GuxJXlfR6lWDp1bqi9Izi7W5SH7EwD88eURC4j04KguXF1PPoZ
0+TyhHmA+/xpCs9TuO8fKQ36Pbe3qIkFVoyJx5a764WLwV4lXsbdLuNJKgJJ498XTEiCTl5T+4KO
ARb6oCMG0oTNjJYPAN+mSKq/3V8CjdNNcpi3iW+X8iXgQCF9tOnh8e4mOLLfEnj0dGKVm5NWoygD
6scSmzWORowjiFNdA7HjC3BaQSMoCXXEnRAasugmUNkpRoyBpUdp3FI31qi5DA5ruwtbGt3+vxTK
XnMCqyEnUhsF61DiOJn1sagxKMeMD/Nd99/ETA4SVVkkuRevIbHMGEr8i3lWXzDQKsIVfZAm5CCq
13E5wsxPsSpdonvuoroZ+L8Cr/W5bUihwwV75mZsoz1o4sdPROTF8sYNVTYRnfmtXqptInyxPakN
kUmbZVRyyW62SWbhAebNM0h7Wk9BAjDJGDDj1XyX66YS+6EUxmlo0xNokIwY7lStkrHJM6dFPkvs
WLka5UruAYiFPIdpviRx1ocq3ZrosNwhVHankSHfFiyorW+F63DKKrZsljVkR7OPs1NzF/6uEM38
+UvthLzmc6nczSk0a/sljzvrXDszsTg50qvfpukJRNCKAKFWYwbzFm9FPlnkZurpxbYoBgmHlKK4
9bZAhsOCAbCw9YW+SnAOtxUcjh6k5CXTeZILVYPhEQcpAt4FQEM5E2tlj2PlCepzfVh5XCfMQXtJ
45SAPLtef3H8u9xheQN513dqpdbEDu2eTFbsUnQgkwG3BxY2vHeWLkdZX5X3XkI1L16C0Aw15aHU
Mz8B/6cLboTKnZVjCj7rz1U8kPzZwE0QVfMsfEB4OaFiiFmtz9hA8vLhYs8DIUqHtDRjYUMrd90q
xhhdybrKMhzJBe3dV8TxXugk4SCK8zr9kCWifIafOwE00Ds511TMaX07ILsmvb7eD8r+97skmMIb
woft5GgrTJU8wUVYaxf6BrVrN0Yp+Aj80bebutBKSyJHmQsGhxVy2KPWvjO0pJhGhrpXFcfyHk2M
Re8/nLeGPSuZFObEQDENNhdjXlptuFHLecgXQnDHHcjvKAsCp9qeM3VZZZ5pr3K+50b6BO2XPKW5
sK40aVzwHSU1ay8njIGajUOA7pSebUbXhSDjevapjfNOSutRO994Wgvtu73r68dJnAtFeHbtTSKJ
tIauAbfjyqM2N1uprL4rUgfZml3G/E77Kv+G7UzL9xei0/ho4vSUUcXUyoWILM9gg/Y5Qd0ieylP
/WbCco7U6c2ooM6e3P0xDmDixuzcZyWqZnKWwBaiJWdjdgumzmpJ7i8eINdBatPpzlhuSULcqTIT
zzkWCEruIUDr9Fw2+plpAE47ApZtp32fpl52+XfbQUp2ajS8xOSNmzEqEIBBXtBSlPxsx0JhSoeD
U7+TZUd17omS+KGn7hPoQZ4qffSEdYmZjPLQEu0NPLDUfbtRbOe/ddKQCLkcXhoO81fIqHiq2+ez
s+YbWiYZooTg03WczqVr+6WPPifN2Vw9u9AGjSQW6V6SGDzZfLAEaEheOrYBDexbv86xOzqFTJX4
uGBSLxfcAL++m1FTD/U7/k5p2+KwZzqONyp3CtPZPffjWn6/ZL1ekwWKIhtupDggo7i9oYwgC7ZB
6BuFT/T7R/QY1SUCW2Amfzl9Id6Qh6mHNH7s/7JNXOyuBZadFmhamA2iU8dVZQKT74XCjHe5sulM
da5hPqZ0+T548RbDvh9feReNbuJJ8WTThVrAFQ2NY7f5KHQ/ELjlCHhyvkWJ2KNxjubRAZmUSwzV
YnyveFVmnvK8KUTLDEMIV7XhJZ3YPGpexe8mpYnAJqnHfE05ms9o0/rqKTJCvvOTw6LkyTQdkdBp
CrgyTCCCBVB9umNRDYGrVq30wuj5/nzrbNi8cqtTlwp5jYFh5qxTLOYskmOPvwjkL+3vzGk1Wh0R
iem+KL5gc8OrutqpB23W5ZHYAcaZbbCF13gQpcXuzwLq8Ru3N79UTfYSGrRBhxQP4fRAgc+5bihr
mQzWFRa9/pQlthOKfGXSl2y3yrugdbRvbvfubpLRgcItm3ykG4+oC3/31HxGiwW3EEPUtntZYk0j
c7zJuK3JRLtbHCY8L1mNPx/sz2N4Qg+ciG1r8yjgt+cqM1Ja9KLPA9Zv3AB+2/DYVzqJIaUbqRnV
GUBvTELV2b4mY6b4/w+bUofteEnCvqoLHJlZHnOG10nyJhI31BHBihJ4Q6jg3qz08rkLZrTA3qmU
/9sEmeGhfQ4UjsslBjl9ZntN/hXgmrbsAE9LK/Ayj7UraoiLxE9cqS+C2Bgbda/uceD5JaREh7TA
l7zmEmDrPBSPKx929IiyUvVE/DpFtuSJDcnd1nUWmEM43wJiPhmV3kCuWHi8YnMrmLdNUqKL8l6z
pMHwOSHKNKU3qUFvI1FMy9ujox76s+w6T0S2mLNJa815x7LUcf6zLMkCIsaVsYnl8OcYX5avr84Z
S/6cd9kq+0LI+ktUOXY8dquGCMQbHzzVOlwcRINdXyDrV/M0ggRNzYcP1thZK+3CGNqUoLOSuQh7
vuGgKkfrcifzMppZ1jYqdWTFQYGmDWaf4dyriSiNWOI0CBkcKnf6RL+spx/cKsE/OwxA/ohb72k6
J8jH12Zuec8rdOxgUmR5tmsB7jTgrtjP/1iv8jOQWLw/Ipcbxi9684ysl/wD2DDb3Xpe4OxtM20W
dE+y3lfNvc/b0Mbg8O3FCc5sUlWc4aqhquriXpjQNe8Mwv+C74MIH7qcrNUIzyaDLUOzrNgNeHIP
LOum5OseH4+792rfGUKltGJbk72c4E/9vhtCBif0pwvi3g631lg9kO2CqT+xNieySjqv73qS/Mbv
mWOm+uuQmPBQDHXqBPWJYtcrM7gT4g36EFwSmMKVMdkAQkPPJ9Vp60ijJCDEw4+PK2e8o+s8gFIq
axvQ/vmNHYGle3pOC7DwXCEXxYvqME99YxoIt5jaYL79vzZq1TO54EMp6g3bfbV3HZubehH0NPuS
mfFWH/CaqC6aWspvSzacIO8re+w/MG4IFsTKsX5T5y4W9MTNY9VNVErtyDOBq0S27T5P/wPLL4M7
rVE7KlV2PlWJiDBxZBM6fXqqKcRyBouHpE8yP1e3u0AN+/9E4EFVzEEre4PUP6iRlYXwe+EYGNWp
3ls30HAijre9blA3K22b8iUuRWA66HyQAWXEatusOMBXybik5vKcJ+75Xo1C841FdtUOcXTX3Q3R
dbvr7SdZbXLEgDb172DQfFVFEkz3nKbSz87pU2Wvh6UVI5mf7QLt5RNowihL/7I9iVj5UiO/J3eh
fMCB4mO+XEnK608tp9aevHDOJ0q/4rQS/idMhxFR6oXV1t2fvVQhxuu5D79WVDujOZt3UoNupSp/
86pvvFGbv1ATpejA65a1GIDl6XhdjozUAPWDVcSaKA9IljqvSoZ6DlMtaCqNfD2PhUzZ3e5t6G5T
6mfW3BSHORgTAePcmPhRssN94CdaJVUrFn15euZef7pGYBmWu72mT1NIo8kkpH2Hwri8xQDkHp16
Dwgl6ys+uJ4kRC2W+mX9EUfbDV6xwj7DjyC5z7Dnd6wYep9XowYIpr0WWXO9dvZcBf+dNzCWmKX2
RdyaGAMGQzwHvqTA4VUT5lwOWlwf2va6xxi6Tpp7ll7V3iUShTZCs61QqGeCPohZ3YqIemY0pup7
sKpbzMM7ScbeZACvuacjsnyJq16zffiI8EH8JHliCTDdQcs50N1M32kR3d7qzMLUDwShc0P7fTeN
y27/09ml/Ze6CnlAw1ZoOsI4gJ2ybLRCalfKPs/M6lv274jwn5Iid929hjSU8b/ZEl9yQMh/S1ry
fH+DXy7Zv4F/0TDzVrDrw0UKBvt0vcIU9jLm4wQgEGjbRS6cgx7kVCy346BvCswkM4pFzzoIS7Pv
pY3cFPhEKNxtWsnxXyZlamt5yxoQ9DwlZbEVBaxPhnvx6SHnJB4f0lrCzPuTh6YbhWjPEyQBNxtY
ftDgfmUCVGGkrEi6OeH5nkqQCjL6iNjo94gQCLxfq0k66ckCSDq6i4Vvyqt3D0FoSt9yFg7L9fS3
WyEqoMXfpwgWZ8H28W75ucejWPdw5ovK2h7+gxJN1SH+FbJsXDKghRDBlXFHhI2DP0O+meax6Acw
syG5jeJboZVp7Ft+b4nE7O5wBnjDF5oRzdDH2Q4/5gspxggYsI/4aWaRVF3cJtKqKpGS7IQxPlEn
n8edSya216h0rjwDMYN/+bL/t+JB+RcRt4TA0U44OKQ77bcc5i1LIrzd+tdZ1oIZ/QmaZyDJiCni
JxyZt+qQfNHltpNJerA4HWJG/j/2cWPSgK+hlrwLS32AiTFUqrKHE43jMtJsaFaaz/7j6eXmMh5D
/taR1dP9WMJcHpOtUuyXWdsD0s6fNhlTdzyhksKz1kFzfUOzQZICVIFdgTNulaxZ3ulx7mbBZ4nr
6ax8+JDNeSNUcdzZ9nSKqwzVHQI72F9hSNrzI0j/CCzyWJl2+tfZMK1mxGpe0tgcc6CZZpraEfgx
/5ip7XAxd+DHJZRz3q1/l72PVpQ/gFrbBk4mPQbE09Xh1g3gVGEqw/Lv7eEBNUC/s0RBrq3TQgVL
hOn+C919DCLqpamOcXinmdUOHg8s/eHeBwygQWkDFVBjT7mmohF4WDG5tDwCTgdLcsN37gdfDabq
BlPj6R6MCK0XIaueaPFMjpQdIOw9bcfTDTeFP8AQ2ElXrhrFv2zyMYq4PHepwjkBLtNqRKF5rtbW
D4Axvj4ysMSR0Zo9b0I89sU3F3PKVM4VpAi/bI7Zoqcm1IdgroKdKCRCC0ZRKt9EUGNhyZib86za
3XpDymi8Xk9Q2mf1cuhLTgRSSCTJhvZLc+1AyrRJxobg8H7SCn+Vg5EvfzBV/nIedpxOJ0Bua1Pe
/ksJBJOW2qTI5NEWRhqQb4IX44Xqmhv/JXxUq6ID6DeKpXewncS+cNY0VLdZas9lgOYulGcYCWWf
/i7IdMTHp3fpbTtjwAqdT1cyc+AOtTDq8h9KFa9SBsAzWaQpXHMPCJlao2r/GOK28QCXFfM3ZxSR
35zjVo8clBUGylGCQO0mhc9gbJO0+A18glY2ljUYFR3e+P+WZO/Wp8PFqtwoLFvvdkyPq7Z9/KJE
p65LT9n5zuUGXZLKUmTCLGvbdyFf+jA8Kz86dAFq3vwPs1N5t4W6of81A3J2qhIRxe0bC7YiqJiN
7heAKlhrjY9D/KryxXHggvK0aV92klcQY0ZXzdCj9aKhpEZTowJg4Il+4+pspUZSLhw2iCnqyBgC
De/vJELomHErVU8TwVqTrYlsmK0ai5i1qARj8MVQ37dmWfH1OFNnPCXuG+J4wR/StNJFout3dS8G
pwtN7Fpy03hBa/O7wPDu4JYJ+92QtTvWHBzogHyunhZJ8X4qBef//YydCtNDQCmGdg5fh9YNtUNA
X03iNkOlJ/pQVq4zZReSwL/sN2+yEYmIYxrecF5YzOQhSXSqd3ly15foORhst6Wdq7iUccvPK7fc
63rCt0MwzxG/RdsKrrKhKj8E39aGsM7hb5+F32H6RathegMS+UI1FKP60KYGJKSuWEjllgv6lV94
GrugYcz+YB6fCZwDa61tasF1eDumTuvCY3qW6BO6f7IAje1wNkjqp7YjVmzDVQXvOgicWRqYwFMJ
A1s91+MQ166MiqlHtSK9awAgSumZzLOFE27oLQ9FwKOG+fBcIgtZZ3kuczMDeiunz6isQOYPGPEf
KvGR4GhTNsVZ2PSIX0HS+ZnqRuMObUYyf31PBc7zIRA6i+s2PJfcdBE9mn0wTvTVU48ha4wNhA5J
FJEmqZyjx/AEyYK4P9aOVnVMW5wmGhV8DmC+o9vr2/gVWZROXflDzqnDBiE5kDmYW07WfRSVf/nM
oN4S7VAxLdNT30MpSX6CY1pl8eQcoivOHFsrNOCxig215I8mzCrmwi0c3BN9sTT9TbsDltzCFE6g
5KDusyke9kH/6e+ySXBtiEFNoW31dKptWeU4JYDJm4ZmvsXtfQweBhzfIJv1qpEep9gSvDdsVaWv
6D6n6bfYCTRZqmkRAPjHnbznoB/1ahU+WvM1pnAgWQ4kdlMMstIU4hD53lB+Ty+lUucu8KhYOpve
Qh5fPCEZ8kFnFII7RT8GafEnIH0Jy0EmDbQ+UncuuYT59ktA5M7A7iGz+0dLFbTb/ddN2mlGewey
UOOreecOQPmApUsvmq5rV+MFVinbS9e5H8Q5515Wo601uaPlyhaHeibmGET3J6kY8ds3GV6glNyr
JpZ3bYU6HlR0ed0tNQ4C6Cw6CEo/p4KlfAO/d8Bnqppk8y3mN+sD4WOusJpdZk4rEZ3E9DY4i35g
YyeRBZigrjhSDOiXmnNWOO0MfgA7HBSI3qSbK5veLhGiMT+QGdT3voUPW5oMzy77drW2U/gUWjib
G58DZK1tfOqltiWzWWRjbjmY5n7RA+xLDDUdiKE6t/8/1zFAQ6slJ2FpAhuuX0FV5RGt4XqJW7AE
lxl0OZXL2ahdRMYMSnc+Rf+Lojs0xCQFi98cmTM0IQw3PCIFJW0U8G8kFAwUmmBpcSWKzhqJfs6u
F7pJmvJN63QPbImgG3lmqnSff4BTms5ftfSEEYm4K5LZ0I+7ftLRiMFOKJmFhU0gTpUb58QicPm+
pUHSeWkPyj0lE5aibHezuW3xy1jEWMxEyjRR+hU3gHqI23Jh6vDdUe4egB0syzIzbAPf4K5ruQNt
Z5V0BjqvNif4EOTzWubrUCs5xH78Gvj3NBjnZ542pM4UovYLziRitkKLSTV0uhxRxtASWqS1TSE5
4MVvNqNka/47GFAA2+71u4pMt0SbMjjn6zRnTqmrt88EaQ7B1ODM0+/nYWAyBbUohawMafeKW36t
stkZGw9vutwwiW9vBxvv/9HEf0qqRJj+oXU//XJwMlzb48c8YecS9zIQIZoe2EpPF0g79ub6erV1
2t7URLGUnXfgcRNxkEtqVwL8FM9/To2z2UMHkl+rrIwk7ShvmeqR6nosiki6uV3A63+ndNabzCTo
IbLHIToEQWfJfLFN//HFeCEpKFFmljos+3e1eW2r4o6xBRNZLgNo2m18jAV1PyxRJuyjLgV64Fx7
13QKYznhORlDVOFHbxCx4SUjXQac0NECU5hudjQEpvDPof+LTdX5BtRTJvzM1pvZqSpE6CNAhLmm
ipu1Fgpg7AgBPh7CruDk3Vhx2StpsDLGpXnq2k2uML5GbTL1e1lufVUl21gQnNOKRyfRUcNKOHoO
yTMp3h+Mx2AqwR377geFSwd3Pk+btkusS7uI08nxHHPu3vGOA/LvZPiEf/7KZXQbjXUY/gTuLiXA
o3h8045TMSW8nzRPh1qQ03eFqHX0hd9idGF5uDiZpYP928gJK6VWvex3yNUVYWjTS9wP2g0Ty0NJ
KTyqW9IEilbx3ASNrTqfyqiUFX6CIVuAGXbdDLdF0FBgMH1lzlKspfyQyZGHrxgqrfaQE+0EqM8j
8eoR8acUVY/j+jJbyCOIt79GJaAIp8zPxceTw2y9Tis41BdrAw6/PRaLbn+2UblqTzS25whHOUh+
Hq1QZo3Ap5eaCeGz7bHUD1IARWcVK5B5U55tdRJYix0tAE5UHaBvGyWRLbkkB9kaDQlKbbVa5lo3
hSjQYgXksRcvW+iHhM9X25c/X5pRe76dXVfmWpcSsp41yIM5t2e1LmXfHiK7x0RCpqSdZQh4ABN0
E8qRHrv6/Cp/Ix13uWNVgeaT1djb2xH8egMe0z9RoB9qie1yV0OCV1jO8ujHwmwnq3+7QvBTsn9s
X5Rpgh8b4sQgRd+zTRBnkP50SBW3pZQliLV3GWGXib3Ie1HQG8FSOnI0M2VNnrfeV9fCJl/zfr24
dzvMtYTCpqwoyEcBMcLx3i2Yu//YHDJYio8VkDmWxq3D0RG9ruyDLVMgxMDFTOl2EqLJo5W6k1R7
bHo86TyUCdoA1nW5O41fVP8QcMXH/Vr19bnWUzTEYixHj4Pu+sJjwksLtoVtQlJ3tmrJKi4lpiW/
ZZ5PoiSFrMa6dKilm0AF5r7es6iQbPa8Z1w1SbRFyOVADj8+aob6Te6VJSwNSYKF10OLbWS94557
83RUiL14bI2ZuC/v+AeCLqXaYt1r4quLocZqZNYUzSOLESfE4yLYFxFyydyZwrZp5zdrq9RiZyQj
v2KdkXTeVlto+fCu2YHs2GLU/fBWVbn1JAdQxCW7vlsruP7wMafzvq0ocgIRXKe6vYB6zM0mcSFy
pWtiPd+JEf/b5oPdA1w2Tplq9Vz8/LsXzyCxzqvLZJdVn1qEJjJ8WfLWrLecmjBVVhXr9dk18qzL
3eUgcwTQy1WUCKtXf7zTDxEzYNOOqGhiI5yvfw1bOSJliXMAOZw0WvWYeLy5exxdf7+FRo/OBv92
DonISiXRHif6fDolecweydsOStCfQ/txQgvK3Tf76tQn4okGOVB6l1+KyeA4G+eK+fAE/MEym6if
Urq7twcinFU7Uqt4pR5DPDIupUiYUAmfrtWsYSAu1Bb3Z4qNauYjcP4uZ4pMrCwjw/lYCp1vPZnI
dxm1NedHuohlpTWPOC1I/ghwcVVKfawA0iHa6lk4WSOskxaP8NKl8mcR78haPwXFl2kJM+kOKiHD
MHHm8hxJPVxLcoXKeKmI9E3iMr0M66I/OOf1ow5dijGokmKupbzT1qjNK2uBhTL3KuhOl1OzNYLO
mv3vHnEO70z+rWhAd+yU0sb3ceOGcLM2M4D+US2dgRmkZ65XFgkqp3sne+5tGM6is72+s7+MWUga
fWu8ztc0F7DwZFVi7qCjL55frl8xvZBBQx4mpCKIK8orr4pmLBCi19vI1vurNSl/7IPShii09Bsr
kiI1lIpCGbGcm255sCcuBJZJCx+MbI5nVs3IE5ZgD/Pow74pi3C4aFrRVEFwA7tkKE+7ZGs+X4rJ
F26N4vtj/Psj14yT3d2YCBvxzO0N9HMgrGX38ysaL3iX51lWao42g8Ni7A9RIE3O8/WWgdGHefJN
X2c409ZH1xnmPyHUB8RocnE9xmZOSgxGAeySDd6kb7SKW3zWCspu+Jfb8WLVduo2u93O5zgYekmz
arl8unyeNWqby2nmkH1nggG8wPn0OXnKOWC85EWXqOY7y6mbkDVNLQDhmgJygbEv/V/dPyisE2Xl
xWqmO2JXED1jBH2hdSY5XTFkff2o+AcvxL3w3K3FAv8WRepMBpOyfCGKMRaBaP9nLoxSbuXkTLBz
jiLcGJw9nqfSXJa2XGeX26Y/IlpYYPiWReE4jzNXe3UGWRvg+w+G3JDoVTYrULHSmORNfAbd36R1
WeGaXGfVVR5MaCMLvS8cpFRbWG0DnnF5wmo84wwn6cfrV6LGM+4owvqRO0oPQm0ncwEGxVslplvE
piu3wFStDEdou1zo7Wkp5gKvM+3yxL8rkJ4880gyOa23xIZ2T4QeeoHC+ZjySdgJIS9EdFv4GSAI
CIZVTi6dhDVfxk4zxLlAggfhgOAnmvBcD+ZmMYzQwNCT/lNq+SVaN+pm9/Ag0pn39K0lcCuffsxj
pJxrSPiKRpiWWDxeNqfnwBhc1WDt0lCUz9lOu7l0dtop110K4EFH+M02unmalHaXDdqXSFWENBKU
0CPvP4uG3p1fHSuNON6plhElg817I0BztRecFFTHAQ3ehb3hTENqDDHHHgeMyZQaktpD5nqp1AoU
4SmvEUYUWOnc7F2RmwEK3qCVXvBaBEXQFFIfu5MzNe/+f8DAjzMSGHWeFwgIFPLBOYERr1V6lm29
Dd1B0JUZTHPumtOZNNMZ3zkuqgqFOdm7AkU8sj0zEAkaeXsW7rTKE+0p9ShytZrkz4yh3UIIoTFs
i0840qQ0qO3WRd2U/wJThfiKCPrkpfCjGfNktvxCv+apdFVYp2+9YPsQwG381GNni1RP/1QxJLfr
TeSzp5QNLMwarr3lXWE7tc2urxNFqXz5iPIv+VKWK6CO+SQpZ3uvut/hzZfs8n0Lzy73LKiFoEr8
sQVQS6KGu8H8y327rI9UVAAqwJnzT27NBO/BxKozd58ppizOxTeAe2rv51Yugcc3AAnFEYJBsYAK
aXKnE/N0/LNq9UFimNx2E4tQw2BmEaaZZSCLs3K7oXi2nggboBKaZl/SnzPg6HYH4gybLiU02u1u
S8qQ8lypGdXOwtXfQcN1CouN5I9+bY4HJ2yF3LcS76rQNPOsggQDLL5XqyfXYtLJRRD8Od2HH9fm
1xMlpnRw/SHzHFUbWrq9Mmkr5G3PqwUhTCel+o811aAvODyD3K6W7zcIvGQcDlMl8ErdHrhSLExk
DtAikf18oitAErD21wSkoNmrP8lXIhMD5Hq2wghWCuzPbf7PiLK2yflJ4OkFuoXOF0SSQ/EcniJS
uAFJByaCY8j5amY2W08JS5paIPSKlGuHjdUJIpNsiDFid7rFTOhbyk+okw7XSQUeDYt556hEapsK
jLKJddsDF1di9LZG7qdrmlad8l1Ewkz55mHEyeWLLeu7PdPCL85gjWwI3Br84NC4cXfSQoHPCitD
ilaufeXZR6UrJCHHsmF2w3ckm/XrzkCcvsYbcpdZcoEImjLCKoKqeb+gLNAsVAjqCbu6DOxumh/f
mbWPBBg0dmowfXlvtRUbSsYUzWB1TrkN7/snaQB+b+F+Z8f4G6054R8aGY+166dsiOeHHBvrQv9r
3HzCodlriBXtvzylLpC34NhrnyO6auvxzDvDDaFR/+/jGKjT2whJIWFz7Nqsz0Ut1aFVawzCVPlp
0XlFhT6KIUlPtyfcVI+lB5qzj4dnsVGxy1joendDxzMVQhPViRlxsOy8iqccRQV+yI+XvWT8xe/P
QsrZRJnw8LD8BODkKWCe12BLNHbk5nWzHfRzwE465kvDRjq/M6rbn96PwiA9LKug86gfY8JVzZQS
MsiXYqTt4ez3QnmtPUIcdubM7WdrbtLrkpDU3LPDLLdoAr2caQlnO2Txw0nZfdcQEkyg0UVkiUBD
wSLCHy0eFkZhWxnyTQVGswzQGuJnRKckrrq3MKyGr9pkEvF8mAqy2/jd2MIARYtTGvClzRYFLEUi
eaXTjEh1sGqEmmcj8JFXLnX2pq8cn+OHOauOfaUzamtd/0OcygXw004cqEMw4Zi5TGGvGPEwBPVd
4ob4laB2KQ1Qafeb4eEVb7Kuv9QnVULis5UCaaPAvrkdBe6xFgBZ/7l1bg2jjmkChOjn/vctqU69
cGjCHLkQ76zi5/6j0NYvizbMKBESZC9DxZkym0Kh3XdLghPE1t267UDVKv4a2MKpfuC4i4U3QBp5
kSzh0RIR3mx/+kayEk9MZqlok+JeSXNjdBWgJ0vOoz+WvvR+fzFibJVB4Vj18EamrkGZHzXSrtJQ
Et/mCbcJAKeiG6C5jqyPd3+fpJWHO5UFAWWHK6biY+uXyt62c8fBuzpM+sJ/YKyiDchEWiOorj/M
pO55r71DV0TqVGQDxXyrpO34V0UDWy6r9aovD6cMoPYAI1rj8xYtAzbyhwd/zOyTxhR8eQScjE5K
RPQyT+u0HDOpbJIROudKQ7ZV/HMaDdfgelKEuV5VEni9pqGTekuavgC742MzX4LGyqZWn9PZ+SOi
XoXeVByN1FOJ6rXwjx/86EmzCDH5uGjd0hDGe8UTL7W1sUIIantgQ+nbgGrz+bvjiQnayajFZzvI
/PG0D94sPO3pauM7/6dUuuLRPiMcw2D0n5hCgPXSOdlW8CeZS/jnK4hz9JrOws4mjn3LZ5+EvPpV
khU9z6CAhoHwknhbTHXvPc1tbWcSwwYp7+fANIjLpVa/5AnDRW4znRtHRPjS6aiLApfvyEhFUw0Q
HONX0Daxo8x+SA5qzi4EODL5FdHnTlsDFvp2xbWOd4bvfzPyCKV537GS22U6QknuhJ4MmJXZqjHI
G/aKIjmcIESAPc04/qBVWoguQdrc8JoaQUa+9GGTm9g41faoI9mSkYDZnwoeOxFnCdKAuIHreocK
Na/Oc2pKg/BWPrO7whSo6OhZ7omT64OTHF7fnSpDNWeeIKK4yaR6QULHFultElo7p+vrCGnLK8A0
dMxOX5GpYRCuWTVPsC1Tc3Lma4nV5ONWrJnBPA5lNssLvOFHa507xRU8QlaPF2vYB10I2cB/GJqp
W3dLj1c9tatYGTkscjhBLI2E2neukUc2KabHK5zgj9DYOZG1zAMwve0P+WtiFI+JqW+eM/cNoWuz
g+ibZt2NIBN5n+iNIrBKEHmFa6CWbTDUWaVUIcgGLImsmzWUUppUpmoZV1/tiWsuNKBYOLwoUI8m
0IR+hskt8MYesSQh/DOGHR6LTolQgmiFXl8nLBAB2Z01zlyjIAKCaDC5wtYFpDIOzJ6UvPgHADlc
ylMk/s777GJdS3nrImmecAqyBLX+JXDJkggz3NMFLHsF9SlK+ek0+GHZfA8dlVHpjtj9Z7ovaFNz
l71f6Mnf+8ScQd2TxWiS3+CsMs9aFl/nLdeAPkJ+wGjNWU0EPHeY9LfjkzmJt9v2akMoHCXY2L2N
XDEnYB2mrgfR2THMiZRTCTM2lI0nBCn7scRxfWuoJmXpj5+2B/Y4GiBfylQBBQcCuu014ND1vXak
ZcVGZhVLC3OgHAsxlC6ucrZRrYg2StyVkBaY64gTpPQyBk6JpcHNEpKsk7c1U2oV5XpGE+sbFy2q
DS3QTwXP0RJjgcH2kxNOO8tJHyDR5Jht7eUuzd0tgrT5Tj9+7COl7XbZcR0s5JfSHQHGpt9NtcID
2Mh3OB2QF5/6VknsE0U2Md0S92uN/JOOY6M6DCBFoLY7XnZFg5XFgHV+j6TKHBOvlt16M87WFQrC
0pw6n6CqBkAKF5iiIbQ2jh6vSqxbaSVLpW9/ODN3yzs2lQEvmHTUwuhGU6ymez/DavJbq6yvHZgf
QtF2kg0ncOSQbDs2mbBJuVouyXJeVhtbT1pjeiZ1khtERun5SKyAUIe7UQ5Z2d0e10lrsxiWgFFu
du0NgXSiGCC6dioVC9Bq0LvmtMq8eMmURxkrftTv8neP2HVjHKfgtziHZI2nxySoWWAArlRpIH+L
KFHPShzGiAlOuTZ36EesH/CjWIsFqSID8Rlmc7XLn6E3uSMJbQpa6BRUOYzTq5YwKSgjjQ0BSUFA
4Sf/zZAMfmNOcW/4+9k8P7g2F5kfQznv5xwx/EX9Yiznrx53XYEF8TmvvaX2jziHh4qalvYh/bxQ
qlrvMDWIiTgB67mB9tNwj0rYtFNHZAFz547dp5euqWFNz2BRTMH+CX6xxMlgJgE6/1WNT+KEAH3m
slmir5WU3lP0Ui2gDd/9M208lnRQTMYTiIhFcNvNX5Vnkj9px6l5UyhInMMAKte4l1LIfSBavSSk
lFmMlrlGw6gFpJieYHOoP8DU4HbKo0ROxU7z1OlCHTrY+9kIFbgzWZoa/52DFHzkRcYRZkTJyWvi
U0cdE6GSXx5VyyLK99YNDaeMACEEuNrSsqe6V2n+q8EgNiPBl2+fXznVkJ+oYPi8lINDQ9dCgn5Q
3d8ErfHUZBydZGxD5HMsLhP1YQwQKZoV7W9wTNKE/MowegDOKjmDVhAfLnZzAFZeVcqAnbh30j5K
wWCrC83JqWNIZWHPDpfi/n3ZWg+AAd/q2j1Y/JkDNSKaQ7eJCEy3QkAfV9ADLR5hznNGBopWKKtL
IUqi3b2qiLJ2r0SPXyNZE3/RjKw7t0w64aFxn4es1nILZiem5Rl8Lpg2n/G5pTnSCFzpfvTkppDc
3Zongv50xK7SU6cTHiPoZ/fLSrAcaNxlhUJD574HNkQm9kUhaBdew+WLvbOm/gz0tdqq+dkMKGeY
vfmYsKK3QmjUaqFJReW0WPzhtcVlVUugneGgCL3D4neRKIQ2xrr5QlGZd9R49ds85BRxJ4p2oO0K
6uN46MlkBNLIJC/HBGl0/B8YY5gQab2BuOsN9bGaO3tTfLBd3XUPwNGsTAODZG6NTCjGSB0VXsBD
j66fOxjKSKQLy1M7e3T9kxNv/pAHBV4xjoK3flPwK6w1qOH7SY/k4iFDAwbi8ON6BrVlLAwS4S0q
Ifg/EAZEN0mKqfaSEBq/cEx7qxxCAFrfRO9SrDnlpOBDZTXto2zMawQ+idroyPU0da6fGMI1oICb
/vYbo0sqtl0rn/PJG8t0Lbal2tVrIon6QOXLZgmqek0i4tJ93mvuiwos1mcNrcp+lGRZEwCRH2Lu
ZWgaBmMlWvGcEKIqsIdDeNFqqPFFxLtiTlNi1eq7enl0tDbflz0EvhhNyXqgRilV+D/MQuiFAeqz
g6wNQYveubeWABlsOi0U71NQm3+m0mi/sMiRc9I44PczSdaElO5Vrka6UhR6KZngNBtFt6zmdNYT
rd1zi4pvREyODndUK122/C9ukAuT+x886F/jR8Ta0f1z30fXvEzo28IJzpxbxlIR9K0zU5ySH1VF
YrV8i1ZnIPeqkC6QT2dBDL2XHJdhOZQ7tJETeeCh84wLgnIS20p6DGxC5ypDf4LmYfi0uC8XSj8H
vPBKf07+bvjLsRntUPXNnLQ3nxmMe2bEt8URnegdRf0S7tvXURlf+D9k5XDcmcbHTpabQ52wuBMi
PoOCwfZmHxfW0VUYav/02gaZf5LmguEBYp/Y5KxYBdOQUasxoQYb4BdbUw7DrjmzA5SSaog7TvzQ
iakRndW1jrvGd/1DI1FG/yW7icmiZRtgj/AGpnlcIASg1dTRsaKh8FjDUQbgyNPy8HplvAORPeeW
pPWZSrEV9BjKywtw4GAo9Z34hjXV5KMQsykEy6gkTTXw3wFZlJHRv80woPlXjysSNd0+QXyO0Lt/
2JhjbH6yvq/Gap0ch/r3aEPcBC1yk/Yd03GqU5Wr/PvrW1bmCzzH61OInlgzNgsIGj9YCk4Pabt7
lV0VRRv0wVCt/nB3uW+ahVxDSMNRHf2eAOOZ6uxGFVFFO/KSSFb4+tCiAtdv0ZDpxRgHKT8jQfnD
DQ7iSzxXJ4ONiDtxNCw9Nj7LccB3JDph2N6Blv8MVmx0eZEFWr9YJ6+BoOtYe5V0sKjbZPwpYwgx
TvxlDhOT+92FAqcyW9dPMPnWsllAAaFmWu8EM/ODGpQYPBaulWp5sh0FoRmaBtaL1BylWyrZZeyp
E8GZn1oXW1wKmWQpzXa26IC52VpG/NKlllfTXdzuBdXBLqzgTdQWZDShYeXeaG7W78SJQabfJ+5D
9HOPjZeK3sOPD5D/WG++etXF3TVG3ojc38CmTTotVvG1b4zIpRO7UxWKUJrpN4nMuYas1XS+FkHR
OP6wNej+w3vhz3R+TZXi3e9IfMlJWQ7Ak8BIs4VUKnoDNC0BTIpOuxMizKErZtYgfvZsu7qG93FL
jyLH0p0gWPIVVN3ZWcTUnNiQ5XM7aFltz9o9q/cGzl0hR4fiTBqQ7UkSdX79bCJfoQLc+tUtrG0l
p5ZpRlxvfY1cTZYh9h2fNEllnZ8spzk0e73wo+0zx6jLfN3hmiYKa7I11FQaqTbOcyc6MCY5VEHp
dO4gfwb0L+XeLxgoY6IYF1N3JODhouYC8R5ZlBd4NCAryExMiJdYzyWSuQ13NUgzboNo2+QBHfe1
S2i5cB3pwn9BTQda6KMP8DtrP9NdFtuMSikYYnQmU9BqY7gUBFtcmL0RE/zQ8fiyu1JgTOj38YdC
LfL3NiTs0SssGgMOWfbPmJgMPr42ufVeDbeddO3p6/RFFGRB55KIl97f3xgiEtPNNZw942jEkCJz
8lVJd89V+31srKwAB4v0hza4Nh0XuiSgAI5jyt61iIBo6s9yaV4ZW/Hja2lwY/p3/ad0hHqFtxPp
+C6IK9Hya9qyJYefw5UAm7raI4EdlpSDVa/b03zPl60PYwi0BT8b4tRoFtxqmkBMSZQzvQ6wW+n7
+y/49u7Ze1h+fTAAWGNd4oY7LOiSuMbKLqBQmEzPAHAuzehg5BOMpTWiqRHufmw2CpAZU0IxiqVg
BUYGm4zNpsFc+cTKOPV/QgwS4bJLZW7zHlrFHUPvwslu+9av3TsI0gsxxU+g2uE6itK20iql/B14
caXbJY+EHqHJivVgx6JTwYXLJyoVQkDlmb6f3d190m/pNG45uNxSq+3KshV+4dtnSpUUNPcA1OBe
gg/eC9Wkrykb2hyQEn7Q/XfehZ/hphiGaiz4Lye45ep0cMbTZZXIWJe4EvUSJ/exUrQ1r0m36zte
Ii4h6W6a2if54SxVR7Hq9EHnCutFBHBexqHsLHS7vaF3HPSAZpMpI6RGU9v+DPbWLkCQpjrNCWmn
wK/vVx8eMJQ1vehzNQpph/KDkyrx1zaI/Ky/2g/NxQIOGkWRb9geDw5rDqYpxtIJE5eToXMSXHuY
j+pJuAX/cme3P4kLQkbLkD/cj0/sIzOpCsCZW5vYtUzfex9uwbnHzSqazVdAWr5sub3VpiQ8DMd5
tvAL3AdO9aaK88VLg3Oo3j2clmfr5thCxb95hs6gtWqHpm9fbw2x4FJPOIZOQkzsSkIKcAXhUwmc
2Mg/zTsb8yeORhu6Ws/xe7d4QwYqmY0zYTzd4WRlIixseMk1pHpJZkoYJhot4n66KzWtYIGzy2VG
8vVK3122WaJjYgLTSrBq6n6fZlgpBLr0kAMgt6lhf/1dWTrxvaQI5BXt6RsVBmayezZTmnfY8+tX
4P+yM3n+TSPZPc+PYQFGvMQR0lN3C35Wn1k/NBtasQmRgvp6TxLNYmLK1yRGvRrbo1C+MNIJXEfK
UQmyDyzytCzGVPW2yBIqO2mvW06LwDlIEfVbnn666gWMv1QwXxEqtZaCIoaiIu5E4geJ2XMQPCM1
hcsfRgYr/3vVK/eyL8+86sMx57D1zQ8pG2q/ZfLxWZU8JcGqfNHfFw/RW763ayFscm8zAPVFOQbN
tTvjrO8oTjqTwfB7L6bUGxMe+1RyEb/tyQJtGu+M+S1q8IwD2jS8PabIo2GoR5m9glxVG8f1U4fi
5fAgKpWWuWnuxxUnsiuELn0/tJJjNweT/wl/kQqHZeiCV3qcZ37tCQpJjcYcPPsREFB+WjFr1zKP
zvv5dg13LssM/XI8yLfvo3fqtbZxUUNfvWGM5xPIzerO9klKyxN8oYh4c69hxBgnsxEYh34p1LJZ
hiH4cXTsXV4ZMK3E9r2QOYz1BfNC7UiQhBgzBH2tLRARLXYgqiMREE8E9dsanuwjXCb2pJYBfr8D
qDcO0KeVnO0GQVXixFmDhwNg8nYlA/kqdBO6sh2Kne7x8nUIRmN6sfGbk2/jE/nI3L4K31trbEe+
sv532StyUcvSBNrKCVfL5lSS+8/PFYfl1MBhzCpNF2mSDoZvOaVuVigAijJRXKE6ZNDiD6oe2Vm9
IdPkg7Xj+O3KeH06Qe7KAeAEdb96/JQzOmw2DC/UPxKGsLFzSpZnUan+EXchi+a82m+C9H8SGPsb
8dG/reomWOrUyPqRVfD37uRcxxeYDxTHzrxMCImtROUfrSt4DoUrHY7OIy9gnojMUg2WZUXU6+r/
qv7gtM+LrhcQPihIVd4VAo8OhvOa8qKsTr8/81c/jnoLfDObcajKK0R0te4f+Pxmw2NEyS/6+7ww
vex5C2TMdSEmekQhBvtbBpMgMry5VpI7VRsj7egPWIr9xY/v9fvrWmDjrYs6a0gcSweRaTzJ8Yzv
B/fhpsBTqmHrSBv9B/gf+/W7F4fXHbz+YPyXv+16SRJEODCUWwd65008lC2raD2IV+htZqZkrNPr
ys8ieArpfjoPhi3HcDeR3gE1DO+Km8xvvPRfgybluqZTz7HzB18Ad7zkloyC2+d9AXjwp4ftm9FI
HgYkojBhyD/0DZA45ARs4WpF5w9q64J6mAZv6jpZCT1+PVs4Fw3nJbLKbGdwnw2j6bb6U6jG6j99
8uZ4xQkBK8QmONiYUocBtqOGH80wROqDG46EoyR/JEeAS9H6PtoRr3grkU5lGInjGwfCfAzy1bYf
O2+R/MlcLBAjH7TR324CsmnpXozpy/eh3a8KtBDSy/gCH99p634OZLZ52wxMIdUCduDqnIHN9wZB
zgHjbLX4Tnq5mdb350rFyt39zdvXt8LGQbe6q1KYNpo9HFuov0H98oq6hG+NhUGezudIJO3Eqq7I
j8YHJfZEASoN+3QbA571a6eW7LEn04xnfqnxImUTF1AYLd8HcFTAzthg45VgHqZSzCBgOmZTgRMc
XNcrzNGQbXevmYwJhBKxe9C9pRI17j8HgCy7Wiwr+qbFGB68oZo08S2rM8aWzZjC2NZLkALPpnJQ
hRzbWv+RZZQoxkAkgVWoeX9zI5qnK70pelH4XAYp4Y5DdTw0SQ6hT/zSuXXXnn7Rw4Z+6SZ0XgiW
SWpr9CWrOhxh46FWjBOrBaqauiKtlcE4apfGQjsTRdecf3+cEYbKBzp20oMCbJNFGBkdiNq0V35R
uy4RfOgjgRsTO2XGz4w8Pe3FobYHoTDu3qBJzav6UZBHn1wKMjFmgZfiQUWd13CLfjaS8YjRGCGs
oe2CgaJyvoKUj94vhSUeOZW1h8BJS1ohqo3+3Iv00/yMBz9ZlGURU2l2vAFhQk2STWfrBSK2y8gA
USHMXpc+ZboAlXppq6mOfI77a0827YxHZ9ELfGB+MW3feyRwXEj/H0tZ2Q9THKpFRhiGVjKBSMHT
YVNbWruPJhZcysXQELv960WMq4MGFEB7m68elAGtPN7t38OdqyQdNoYBGDSgniKiqXlbRv6kyE/A
AL7xDThbNTERL/osxIgyMlZzt2i+FbgLTpXlvXMCOSuOOkF/6g3H3Ix403HTLxiORdHcw0+sYIGv
D3fVoGi71ysyANuFSyaq9wuAN1uQODlJ/+gtpG0mg1QcxjKY/ou7PJOSRYN15GwVMMf9y5wcpsSR
xQTEJ1rS/fU8HPcSlXoN8dMkilx9U9oyc1XfGpQ5pD1gAOIxRBBU8yYH0F3of5K2KN1BfYk4mnPQ
qxvi163XfjMcFY2HmXrhwwvLa+mQE8Piu3AViyxYW613Kgo5ZEnzsmLLyMk8seyq1+H50eI4yG7c
9L285/KfyvIZ6xWMEXXTtAVqFf3GVKgzdSSCletltxfpI3SojkkJnfPwAQ3R1P0Cz+y0OzzTYGE5
ZmSWt37cBraxaTKkjmtGdGT5EUkQxo0MDdzfpqNh1JzkZ++WSPhtjkodBKYUMwg/v1JQUmxBWZDN
8F9+iKCw5n/cL90ZKBTAC6aPBCK79hNBzc0PVPlahCf5HdCcZ9FYyBrZovxzMpk0pqBF+0GIEwYr
9GpKA2noyqvDkk7kCaO3qNSzcJkJwNceETMkMlCUx++ItcX7aefIBeFPxBxLKsVirgEvBDBEPXQb
4tephiCm8DMmfYT/i7ICY2GXxvDiK8A8N/bN/x3Kyl2BiCk1u6JS1J3EuSLcNqCjxrp3zx5jh2D8
uGDzqYDQNvuvv8yfCky8GFPDKe7/wCjNI9CTLqfdkbI6BT655A/iw4Hp7nN4PD9caSvfrVRGWtXE
pdq3szitdH3cj21DNA6mmqjhprKJF7yoQh/bgiuZVLayigqWbN67rKg01ILYCPDOoM3zGKUO9z8K
jwtdoL4DjX7+wvh3Mtvpdc6a7DnfpJdUEF9O0YBjJ+I2LpGdjhyHL82gIDfRiwczRDyXgXlcUFqS
pFoWd6rFabIjcdFKp16tErHGNmYn6GvOTLgE7nh4uHI3eRebkZRnapKnOUvMvIkOkypeWSxLCmZi
dlKJUSGD/Yh9+gti3DrSk971AWQS0kAVzJ+K8pYl+F96o8DniYALqJzuPMVKgB12bIJhwJxt8A87
QRTTk7YTUQYK94f0H8sIF6M4r2JqHEsbzctrKwkGM+BXMQ/pPn9WKrfnP7/HkmaidSMz99dqacXE
9AhfUModVq9YCX8kr05YhABB2laH6Qe+IuIQx0kduJ8pVdImj/ImwOtQVL22gIYR2BWB8FPQE6en
uUxh5l9c+/jPqEU1KD7F+Y9DQGRtzU3OF5nZSV22uvY0ubTbMVZmrFzyYTBXVI8uvQ1rlSwDfE8C
tv7qshGNrZtS3XMLbXiQ9zISSl0iZsHQnk8Y5r+STsQXnaPxMsMQ+UKLXN7X9Zi61QDhfZOVYJb5
CzcOurz3ubMjMgzaM66RlaRqGUzLsrzldU8Jjpj/Fas2k0fZd5lKUABrCRDMm6AJjBaSmDHpovbh
VnM/N0UKaEZl3nCthJotglDc0myKxCOgf7vFMYSY7ZjBAIpTvZjCwGslnQPk5aAx5ifY+XqlRIpX
YrXQK9Ergdd8MiZWX/evuHotsrbopdjhqDFxRieHpibCaMhvPffN3jwNjBIrM9qQgCVdMm0isJd1
hmKgCOuiL/tTvH06ISFdcMR9kjTXX0nkNTfUzbl5D7dI1p0/9eSyCBay4NHxNo2wt/6RG+bdA/4I
rmvVQ/cz8CclT22sJVty/yv5fODM6NbZY5hcAeeaDdIUj+phXIWOz/1dG7uOPvTzhVAMWFgErqed
TF7ZBnEG8ILbIfY8ayiDBwvDSh+MHKzOA2NRGegDkSJiOro3IU0uKt5XQ9bxqaWJT/viLPih8FnT
zXlxkiBoc6tbY2aymcaM1UMDr5t+cgTxDuqqy8goDVA+0UE0+Od7eZ6yjE63LiZXprzJGauh0vip
mWaASgDwhkteqCRs+eW74K56aTdQsK2h4citTpGzxtyQg+F4JybbITyL8zZSdzOnFnQR8ZTqXCYi
ZVNBcSKUxXFPaTfWLyagodC8xn8nb9/rz1hCB5QjfGelb7UdS6ymIZXsi/AUBL224kvTV9mBoiv4
DtC+kSFpEtSTwIoxFNnWIpUlCpuigCDjaR79YP6RhKrWXUKRpriD8+pBiiYmPQZ02znzLPsT4E48
hcuA8vgFptAt9fSeZB0IGMAvho29vw0pC4VK8deZ999Pdm/v/R+fELwldBxlKsEmUY2/ZzWbrhnI
o7ds+e29IdCqndqpp462Q6i8XrlFqbNwO86AeqO48bqScEKcoBiEvRS26MXi5iTS9j0wuvhjlmEN
E4WMrNoQtsp8cUB1FXeR9+QUPxd9Bx2gGXjy5w4nAMKd33+tfQrTJRxKCB0f1/mDy6Cc3XHhqcKR
nXU8Oep3p8/PHy7u32IOpt/tIArlxrk9CqypyoEbaTOp8kS5weGBwLslB9xnfn+VMGXVr0qkxIPR
bYL0HPDS2mFYL6KiZz7CF8hQKEFkWg1YNxTrFw4gbOJ3sG3q7zYuPGxF2EaVMDn15PiX/PVQhhPv
7NfIveVizDotKmPmNF4mpcUO4JI3Hw0cNYMUhL8Pm2mnUecbMIMQZuTGsBaHatGDebz/VOi21lQA
LeHZvVZwNZIgK3Yw1btt35pxG/JR+/bj35Um96BpjUfRaQRGFfuXT+9Oe363fbtWihV1mZhOBhe3
9b2trt/fS7AvczzipYxvNk0UwMXiZ5S5TbpFk/gXNRplxkxBUmNRHWlIznLCHtIEN6l+w//WcqrL
3WiVqiDHDKV8bhppj0Y69JCiLlVX+MVIDygzJ/SaCIH5FOVJyRJOkT9WSE28ibAqzOxPC9WjdoOR
Bw0BDjAej5D2E9v5MBfzIqSREajjn4QxesP/kFx/FzSjUOzq/JUzE1WpxeafLZ/6FfzavR0if8wh
hG1w5+EG+vwH0pJfocuWjBFhdla+fYcqknOvUXYn5EutvEjXjKXyS7i1Cr9pxnhBK1Qkq45NZEL1
LuIHBSoeCc0D5Chm4KT0TBR+ZvcFSme7oCZPG+LQAt314meIEoOgzPb/hEMGbKMnGL5viq6OTImi
EpnMyoCAG1sBrIIE62FzHY0WHcYWiBCP8KpSDkeII/Am0RPnfEE+OS1mYnEh/WOF9yOXLr1bY53B
LMIkj/UrzSwBTkwLPOrUkV8eSGmibYOKXYOXFNocw5SkS4uUqstNU2SXzKz77aq7wV0DiT5SmPjT
cWB8IoWtIb+rvMqZKmpJSrPOO8hOdv7fafONnIxyJWDfFDbBxndT2JRltVAaEu99luUoG4OdT021
S3CAom/lLRTW2HuWja9egpA75jIZrb/hjDbhzLvXaSRgI6doSlXLBI6LFX85Vt5dfsDqWTxeeVBv
vsiqw1WuJY991rzXtD/47tk4prNC9iAGTIwO3JLcyG22iUEsbidyNve+U8c029T8oNJ9lA5Yn24B
9OZEBWfhWk3KOmXSU4jfaJdkbgjzPc3uo5kumBcn/KVBi36giok6TAa+1+aqJKy3a9YVxjJWElp5
+uFzN+efEFUxWb+OFRon69pFX16ugquY8TR3jEj62wYW3RF180d7eaFl0MhHvZJ5/+xf90ftBYzs
J/7RTBRefwBWV13KfxLCntcw6EcUL1qX8bwlE4kI6n4C8//RLgpyYPo4vljMQ1NEN/8UxNlXl8KW
TXjP3sVUYUo7/30GhgDeuIjEv+VUwzyKGZxbrzYv1bGa0Uu3MHyjBdvjpnwpA2sw8FOiqyROFjxH
+OLsu+DIr/uGzlR3JaXGJkbcrpbJqbxVdUZazGwSl6jEAntp2RJp4rAhr872SzyImU5sGMbFOWcc
BWnIXIUjBWdivnZcqwuAH6l/Rhc6DxYs6ynXGVzk4exBWrM/6YYiPkVhLvBjrvzZ28+BZ6tDbHJa
SvqiAD8QX9WrwF2NmKPz+NNE5sW3tDiZNqaIsC8KZ07PE4XAx2PNpajO4jEBHH2iWV6W6A0dw6gK
khyf86C4T/bJKfjlxB3As5cF8lwCWjywMneE/whIcYIikEaHYCpQf2vrD7Pbm0qZbTUYfgOl7nyd
CqB929chrGIP98PhTblIWUuyZV2JIDu2SH/Z1DddBxw9HxQx5OydJFw5eBIeyZnVO0SqNDDCyIze
r5ydjtVqMDGRSFRo5cgrcdwF7bUITEv4QHzjP5+jQjjwTE0dSoaPaDN0XZzxs6WQ95JuiM98/cMy
ACfI8OUSoh33OfNZQcIpzLXK77t47V/lpBoc3/fmkDrLIDL/1xK4L7zOomSUNVz0fl1zPKH2yPUw
d+taWKvZ9r/v1OktIzPonO+JJGzEga05UjBDneiFvYl4eH5YhRAW1QnzOaj6Fa769yUzAH6Kyxm1
Y2JJR64+pWtEbtW8tBixq4CZIFaLbZHQRNMyLouTo1DEsHk+yFTsW9BF/c1KILpEZ7RLPrdB49cX
4ZTd8/6no1bbAKjN5mUiYpCcp8WUSGDPTTGpCPsvx7xMaY5wYKOK0N/t1Te5AkYCQ3Q4PEEefoLW
fnQ5ySTPVYNpCQvz0Qh4QyjiIvWx5in1YBAHIKrM1PNLZHKPSt1Pv7oMuSt4bNFEJph8BJotOZ2y
+a1fsWuO3ooe06dC02M9OQ+fEUlKpZQdEkpmPYtFZn0FIOnEsU6k2z51KqTKGfFKvCsjSa8fSXwT
I4BrWLI1yWsqRob+ceIYntLJQdh2GPYa+8cTRYTSQGNqGDaByW2xHN4KyUmMQ/F3ym7XmkVZiysq
RqGyh1veE/DSRVN4KlaQZD3vi/c6S+ZDojeEIsQYf0vLCGOJJMd/V4Th2vjop3odetnKrjJ+MLtN
rBQJLXxE+RsuxzxvfGQowiECUin48TC143NSFDkO1G45I6K9uYZAEWpmnJX7iWAPoiq+KjZ94EcA
kH7y4XFK33Bn9JrIdbf0qMuPDUnyiJSZJ2vQxsp2/zDp/0hdAbSClfGXzKn6riiVz8wcE52Tku0O
kr7WehIzCm/zUgRUPIUQjiNn1WFqcFIQUqt0rWgXBW9IXXvs1VH62qfPRRvDymBQEvTIBSV/nrmV
jF0dUCY6bt445rGLvUQjXrH5H8e3zsb3TvOP7BQq1VbAOeemkcRGPdgDiDgecZiBzRaI197pxvJM
zbywTvkOFO3DBnotCIvVndzgCnfxPx6HliPBl6TLLPF7HBBgj1Z0BZFc//urOUOPjkHiWRY3DyOL
YknhkqUXASBzMGl360mjPBSK5bKoT3ZTcFpLuY1APM5xSrp+IE8lPQH3lpedqOwn+RwmssiZeLXH
vgCdQiHbCIoySKJ4oPZNj2Dcb9hVu0dGAfTFwS3SOarWKg7mNVyTIsFuuCLfP/3uwWr0yuKsxswp
SAl2sJvgz0XOS4B95qBUzgExGWZ3Uf+S/N98nW7W5LoJMgn/4pFl3FIWhwCDbHnpW/uErjmHNurC
E2196TmloPOkpg9ro7xvmAcfj/ch+8mcxoOHlf5rl17/TeIVD3fpnT+0MyU6wbuB/UUEP8NaNMnn
S1I7ogmFgJoKAQYKroJIyEzeGfRpU9uZjh1JSwlCQKWj/J8dTHk8e7RiI5BKtYeosStFyxoRx6as
xljt2/TNg1A/Efj4iS1ZCjgHGI26PCPzGBTZuvDAxwwkRahvjNwd8fVMOdwfrijKS+b/5REGIDvK
dSyAYdPVYhp8V7++QfSYJJTVEvirWsHs2bpQRErLGLxpy6sDDAEkyCBEMYXirJ27bblh7l6IiAZR
we4BbG9pg7z87jKiPtlebIPBYIEVVUsCA+1DmjXAD+UxBahVcBbwsIUMA2cUYKHbHYkOpPcRfNwt
HULj8zE6P744oE79SM3Jbqe6dIOfYS+9sLcXlb4Zqs6NudMi9/LG23oM3Mk1nBTi26ihS5Wr5WKX
8nYb3qalEwGm/ze885tweuc4eL4E+4VIRDoltDmd5ZKIFiR/Ltu12qDNECCd9plMM35MD6JM98fT
d6o4GbsmcZNxxdPYQQjy7bwMVl41GaSdMXGgyYW17IJFJzYCO1Ih6R8EaAy/oSCAGwU/rFrK8zeB
F/hYZJpkZJTe3W1upkbckZWmqXSUeM5JKpR6ODvtP3pi6vg1M48Efw/A9ZX3i/jJFTiQdp/+Bos1
jXKYOSW0zM+qxEzbxjLP8JKsCelPIBTbh1GdvFGfSFhwCnVfJUk7vTMjNC3QI9X06sXuFrdp/vXw
wUOq5vqWAVQl2ctOQu/QgbQ8uPIq3GmhkQLqd4Pw8Ef1omgUmT25mnW0PAW7WaPY6prmkliBJ6vE
+cuUoHvD25NltOvLHw1c6nxT5sFgCPETI5Xc4PVUlKBpXZjXpqlnLYIQHrR3eQ4Ed12MvuvPGeVN
k3aAu9mamKXlXWR2NVDJHjSfG8b21MehiwP6UWzQCJA66/Q1cUbWDEBE/tD6wkAVGVjYsP3jxhjn
Mbnsvib8THZkUp1lKHtzqNuY+5d4HbmlkyBwMVL1ScnxqIKG/x/Rqc/oghFr1KNOx4hJ97x3MZPu
Rau6Du5YTVNjZW1CtW28Y8gWko4onlswLWX8tyestzQixpPZUioltYDrfj029T0RJlU/HLOW7yiH
HCU62qngvP2bs6WCz6xXlp9VuFDuQ3dpNyW/PrcHHDOoGwG6+MORqjTle7CGq5SCdSLCdot2QH52
u791aPTje6eGWR5bIkTS+pDbdf5ZicoOWojzPrafEX9fLfNeGVLg8h6+kckD60M8m5z+EpEexd+E
Z12AexD1KH0lwnUKps7eP5JUMR2CdOkRb/BkkIN/d7I1gXkZv5XIuXweZENvFH+OYATzqACYU1Ge
tfwRj7xXjidRAgv8YMFy+Kplfv+61E6HjMoeMu+oysfYcjNNIU7IOPEQZEfdoZyWKlaTEVwIIsr0
vWEFcctSWdhQ+C8n12eA5Q/l0F3sjuUtCu9Hy0aE48AyV4EFXSgkKilcr+6qettY5zmLJfrM8cWD
4jLMWETbGodOquq8AX1lt54f8kOjOqwRGak+6DEm8Z9JWO/Lo5PJ0Hy+7XaofaEdZcp/qr3oIaKD
9ZYVOuK4aauqVJ1TNmIvrDHzkv614FvKq3Ie/8NxKfDmi6bjF9mcGHGMk08v05WbYUchXoEz8MDc
WeYdQ7mgpzZnY3AKhndL/LR1V6FuhfQPXMJV/FxfJXjuPAJzbmT6+GwQoz+0/1XryvUkj2iGSt/Y
tdemh2YYOJvcCsFG5ZhXiHojjz72HRjahgvnZFi904X+2YxSkoxdU24qOG2JF+MaCUrJJLp7lvz5
0UbglmolBx5gwhkEGOP/lllVlviWDFZsQIQg43irCgASvj9/zufONoJ1EU/Tvoos8I40ovqrm3jm
uNFaxg1xoDBOwTik/MWlptVoEPAbphg/yVT9dEuHZcMwmRrto+1MptdNyVIhi4E5NOt+H+whJOsc
dw4yHMv49J2YxaIqteEQdl/6Acknpz5q+uGxalc8s5EaEtJ2PLO9sctFwBW8MlDH9SMX6LTBL8vr
oRFefdrVkBJcbZyqc0q31/JN805+EP2kJaWo3hFu16dHSMI0EPRE/VL95RfX1aev6dkvj5usCiip
BGbMsbrruIc9EYsRBpAafI6JLSfPr7oacYWRDzdzEhmdVXEbJsRQgaljWZZlKEe5+DcyAsU4+4Ez
GCKp0JGmZQj/y5SumCgjUXqzMSMF9rfe/sBnHHUWR3T3boNDcY1277dV4Iq5jPpbWLSTq75KtRrr
I5My1G8rgopw/L2SehZVEIKuJ/GqmztjIT4CaGRHWpneL6qOT26W7G3Aie9bXJ6RpgOr4bvUujz3
5LKqRl4PuGjpUhk3GOQGe0VEgqCjmo/iMZCdZnG4j/JEHHpcGXYV+OM0vl/vmb0AdR+0UOJpB+tQ
RIF7Q/CtUSxn1K9O5Bmqj4fzq0gx3F2ZYBnZ9VEXduSbOgLGG+vNFpOzWKyLsk5GF9XKlvuM+WtD
njQQm2X9jBAHM+6SY1ct5nFBAkvfRnvCpq2K+HD9H6kJu9nZpoJZ2Flh12ry9eWV4zNMj2mhZ24/
WL7Iw2G3tGsf44D7t/Hi1Y+zAf912E19utx9NdV/suwbEVk9fXIAdGQ0se8ur+15s+Ii2ihmNhdG
Xzz53RvRlRv8SXV6zbL9KzChoO9UmYzY4qbcSNjeDymXQ7XDWGWKs7k1++iBlwgFeHlAsuZhwHg1
2Wg7JuAodWGC2SyUlhLewvyIpq6SHDl6pC2Q/EAvUw5uwE2UH57+7dorJsrA9ZZZC+AHZpoC8YZZ
6JQ/7ZTvoX+ONpxhEyj9NEAcXI30bmIFfVS7OyBaSLbHJSbTQ5818x0ZYS64roi22+yOBZWmierG
F02ZUn1KPqT6b8QnCRp6eoqYTHVrnTclUKWbg3e9Aig7+eMyTZWDg+Eope207YmZqVc8sCpHI9s3
v1lglExcTJ22OZsL0AUXlYGXDRg4N8O4z7vqzV98lWGrSF8WBs/ubAJTJpzai6iofd8kRUMfIWaN
D9ZNwJ4QzpaCQizEmAt/Ph+HEpTuWIgl2d+y63vni7H7cj83UVOBs0wZPg9+M3BchhvZm9I9ziSf
mg2stQQzY6mjMwCcaBR1OHOT8r/bomvDWHfMRp21Y8MWRUSLEu9DoMX1o5qYsSSLfxIIpnlSAyTq
3FpS5zBytzXr/A4Imom19thPy1erA3ij+ibj53Q31m0+EinW62Nh6U/kSoaZfbDDCP+a9nwPUwLL
R+RxOgmLuTEjA2V1+181IbZnapGC1elz+C6pTsYKyelgIEYZfUd4DjER5NyrCUSvO6+UDTkJT2Ty
2D5JSQCWdKBSNkxradOS0ibdloJ9D6EnjOKj3SBDU/gwB2fwzMVPM4zAcGFhnyOAhBWX65dHqota
smonXdKdWHc40o3qXbPM333ZqyIVbKUnym3OSgPs7NcFp1xK0EGaR0ggz1aktLwcItdXZT2y5JFw
lnQH28KFPo7IEGRGXheF7uVrfWr4gjj+k4nkAaXex4Jk4knA+aOLh13JtccsAiHnv8N9PD2wTBY7
gyuyX3r/duecZ8ji0Hggusn5Zvz3YfqwyFHgp/R8FF+yjCQVTd9EBsMFNy+FizxUY3S+5BtzHpBN
B8V5hb9uQFWhTXsxtVBrLd+EyeNPA+qXHXVKhDLV9JmFRu6uGEI0rqeoOqdmeMNdJ+/S+XxRW9wY
/wB3YH0wmKDUAw6LlguakbGGOuC/fLSwWsfc2c/H9KTygZHtQvUMR2vHhEySo6BSFPtnTUOTkwlW
yE+g30ENNXZ/B+JpFEXL5A4lqWJFHfEn5GfHa4a+LxM4oUBC+Ikj+F6aO7l7XPs8Wy2UBqEXNPNe
qnZkrQQ1rvNpgSd1t5wpUPvMoBdVc0+HQd4NfLmfYoaP0VBUsGtqalW+Ldh94s9chojDsj9yd0Og
PCCOZXt7b+DRjgAIvZD/FrQmle31f8KLpEK8eyaaj947J25Ch0eZddU3GzzgB50tU8VuyqLx41p/
MrgqYrCJy+ldQBAdA2+IFjqK5FwiD38Khzem8b8q69hpW+EdZTaSXZzIs1RCOnNquznGuU7NqIZO
egzF7NffhexMb7ZOnnYoPpG17fHdq9uBG5+gfMz1HpTLAJwWLOdhCPQGWwBOrSZJ6XbJO0a05NIf
Qiz9Lt0zpunQMOVjH10VI0XP3SHtdo2DNl1R7XtKZZevXmQsdGZMo5BiifSE6DAPcm/Taiu1jlXX
xFKQKSWZyxA2rH3UL+w/ZAjYzuplLs2+9WC7z7DQfK+WmawKVsy3Tpx6y++slPE0Gyv7sZBktfLl
n6O/qTMuED7plLwx4g7ptepXoapScAJSfH4TGRl/SjmY2be1wMjsxCH1SDgaLpksi9Ju6oRrnDdN
fo31nHTYREDeko4OVTVU3zO9l4NaDEoR+hfVHmAObog3z44bAEvMAFAtpa4JCNOaLOv03dV0q8G6
cPN9xcoEfX5Iu57CoFCqKSYTjFqpMKd4XOaR5rtaIvio1H+FRpE0fgzyA7FEN6IcUYAmOq5gEa8t
weMxtetE5+PCjJI6Vpp7L/TofuSfIh688TXOt0JJpvdYAGC0F5nQSA61cntq+tzyRvlkStO9jN4D
wQlz8sfsLMEmnedW4Tp4LEr/Dd8crXuQ49kjUD9I4q9c5vImOPwQE0rHyWU1K8wX8dm8WuPSgWd5
EX+NGTOPkUCrjFIWraJ27NRPnWN/C+kNPxGJGx8nINmSYCHOGK6kzPPaKfVAW9CBZfmas7Yga01+
+zeWVDAYwmyAtRf9wdbkC7VvQPVtRQcpdAqrXlyg57QFzzk1JWGFbbmI2MDRo9cjgVidifR5GbaO
WqvBs2icziDkOf8vR6Szxdxm1/hc2HXYiRbzUjZZUk1/syyH6h70ZVDe2mNElZb7is50bEnHOifO
Qfd8ixSvwp/rewivzzgGcolbPnEGxwdTI2NBF8nl4MBhK187s/LVl6W3FKTdc5fLQgXvdZrlF2dt
WFXZE5fNyFmmyfS7U+nn9/THpNi0QKTmFs8InkDcYF1stt+F7KfVNKtvBk3rfx9nVQX5hvYP+uR9
iTqvricQWEauJVhusE1wPqvEgFCBH7ItL2png6s93Ph5Mf7OIrFKYNTA02+/aVA01HWhAbYP+7Bp
nSYjHI8wrDUQ4d//ay/M7GtezKAzD1n8tU197Eg0nTPJi8KdtMHk7iHExdaVLa8CkXpu8iUrmZw6
kBZEkSDOFWm5qQK7YA4R2tiFJq1FYZVKHe8aBKvSol0wUn/tsLu30uO8jNFstBoqF6u8H9sqj0n4
9/aeoZzqLE7wnFhlYIzScx30JlFwm1htI4aCHoedsnaeUWpXfBIuShlLOBoVuoN7OPe4swwfihiO
84Bz1jyehH0dubPs+G0lQPvMfyG1Cc8qO9Z8YyJ4AFdH+MO1OjRjilPIIC3y2l5Im2aAqQvZ2H7a
nCroGX/Sf/1KD0cDqRDqT8U4FpbgAm1bI5C/nz8ZI/iual/Rsbd5um4sMZ5M1ummu1hJ5a4bqYxA
FAArAo0yvxhop+8+F1UOQHxTTkN4BHHs+5cM7SiOCSg5qN3EbPPu5e55wBmgplZRS3mU2jHZ1BD3
iWX7oAOoVhNbfX3K0vQ4QDyuO94tvbKzczM6pBXt2akrJ7jPZzcEoIX2Ovx2QvIKsDXLDLnO/qR2
E4nX9EQPZ1rLbtvQfZvjl+tZXJl0FGmyflEbqiF8oWh0I95vbjn1C4LzgI5R3AMNQgGH6MzdI+EZ
Q3v+r+QGcb/4hYea9CmaMGqegqI8n4z+KMbVL+vMTx+gGIxZud2oYyYvlUNI0Wc1sm+rhsje4BaM
m91dbW0ajntMOWhS16CiDPuZHGshddtvftOwP/pbDTNwuW/frO6PI3TTjknTFcfecetdoIpcGgoZ
cLmNnHM2Rbyk8/lXP5J1Yya6jfXOvErCfJUyw6Li4q7opGomvhgVyZljWSutPgYEvu04PAEYLVPb
i3e/hLzAJOt3oIfvZxq7wmEZ92Bmu15unh888+94TGdgfY+HGb34Rt/aolQX1VVn6wK5JWqqMuLY
DtaoFyQFpCG1MBREHT7tMOOsUXWTTSzN58Qs/8QIygyZ7Ma8SwNHchxkcGc/s/68Iy+pWYeF4NWK
oKt0tjKYmtlCQ60J/2sP9NAxbHjmRoM+6d3k09JVq7CKM/m+XpnrOnQ1bVjHfOChAL7Z9Uz6k0vX
zxME5TCijt1CkBTY7hbuYzmdN4PYmYm2+J1hqgbMXEGR+Br/7uFtypOSrU2UvlKadeTNoBuynNfh
PDrekJ37z4s/7V9MX7XLu1WhBCDYAVl5CMgRq/Y45KcSuqvS0fBxkECgH8imcxL99ReuE5Pu3H9N
+AG4bffv3MttFnT9kJllPJw5sglBSDVfjDXXt/j+myqgL0hEqy4hRXCvmtsYETtEdDygne5nJIIj
EMx6KYEMvU2A2j3daCRUgDEvwZ/caTPd2BkB63rU69Qi0v3e0b64h25j9NxMf8LKFEKhOMx7pZCA
AJL9hsxFzIdbJrTwRYTqrecjkdBFR6vZaoFdKRJxLee3fMyI8hlAECZajiK9y/u/wl94w4xiSbcU
RpIn7xQbdvKBtQpdleE5sjuLdgkdfKvOFd4lWeUpQq5mXDK8LVqQgkxAfi8mYXPGXL8AkdjUrzN7
rTjH9ui3lDVZ7i9SQ514/tvYQWUSfhkgz5HkXoTbq4bUAj/cVoxwVEhnYhEel/gh7Waed8GJqIf4
2Ra3o6V/rIq5ABHcg4dvMp00KE128AiipSW9Jly9L9Mxzb4JpaXti2hFElf+B4jqQIxm0A4dJywQ
tF23RTXAAjZvLiIezYTuZk9GMMTEoFQ2NhBtPqcozuqfzrCvylGtU98qsV5TmID9Bnz9cfppY7tl
NpEXXNzbJl33zDu9wCQ3q5hawchReCTljwhT/HzLg4XI4iOf+rKZkuqEydGOSoy24VvvDH8oNxCG
A5HncVf1ywlbGG02W2IzoUtNBSg5yUKvrfApU9CrX7b/XYJaZQuEqh1DQF7bOxDlRGyJ8z0eBosi
prnQlHnZGB2hCBheyUpVjkmCQ5nnau/m2zYD4iDcWXTUrfc6WSrjvifX/4UoMBbS2m8u1zX0uVA5
EsFTMF/Ng05ZeishMEnTXSqa0sGLsoPZe1quhwR/N13z73cUXktvgDl2ssVg7yj+RgnbTvb2nqKe
dAlEbdhtYuS0zsr/sBPgYsAa9HMcNTzHd8akALQZB9PRy8t/PlHt9tSAiYv2C7IKNrAriBmPWmSz
olVERO6aOlSbNZN2DYcUu8k7Pp/YJz0Y5JlHM6n45y9iyVqczlKVOol+37mk8ABYoaFhjButWsA5
rzx1bZr7mHWvWJISCViYJraoizvL9stFynJpx8hs0QkrPt9DHUSUlZHQRH/nSo8EZUMuFWXfjUXv
M1Ue8z1lxPLzs1f5AlKtsxv42hnXxppkg7dB7KP4+UBn4yioSlWC9ow0MQ5XoV4nMVWcBuGULOzA
/0VUuMYtpgb5Dcfg48RCZeoPca7vu589uJczbViAd1DeySkOxyytLQjRvHOAJDFgRVtyOJ7H3wRc
bp7L7K+3DwJxZ38BrwrMpBkbIdmqjoYVMsYVEfhDO2Own/cLHRD3/tm5kYjNNnwA2BT85JwYQCFR
9dcp2WFAVFhJQxsngl46x1aEZuozV/9vnrtazMQ2nUuAmhoBePc+9U1gdisgIifQvixShi0GAXrI
e6o0GYRQl9lOapDnR4BFyHm+GhWyjZgOU7g8x9hq8JCSgB4qdpp00HQbcQKuOQwbZJAFEL59VtXO
RuPWv8UKnF3lOB0AlNju32iHFLThyYZClGPS3oT6ziTMoO11dM68VRzude7/v8c8N9j/fX0FthAo
8YNQ2a19aWZ3ShkKq6PEKXGRPDjEVMykvH0c5QMrwApa9/eFfz3QTRaMItbqok2fuXw57xe+24hw
uUtiPG9tL8HlyFOlqHB1xnlyAQ3cUwLB1Qt8OafmXHJjUYjmcWbTXFdd6xgM5w7XnKpMh30Ncbng
E89iDtCyVrYWVYmv1a3pVcgZjjASZXo/phloXfHeD0SMQUJy/O/z20W9ARsCNssou70fZjxMxdkL
z9c1FVBQuYlJgkMjXnLHU2E6Zfb9q6L/B+COMPIaB9hbrOLdwmANf4s6/9VaDC5UPsEA41g5OAVS
dxrSuBKwsrBK+BAs07AmzyjFBA8qIiABfcg0Z1lOK1E0ljszymdKmCfDjzBgQWPQP2js8MG5TyUp
24kd9O53BvtfMBGCV/jizaM37WnGFaPIXwf/xErP+3jdT4/bKqYcSIibFujmZxByzdgqJWMvEYfY
HHuxdvhGa6C5KaS7kDFuU3tT6jp7d+ZwBXKOIX0igJ+zynSlK0ea+nUP7CGLhAZZiixd8mV3hz0d
OwgPFqmHW0kW07293AdOnfTxvBn48sr/MqAC68co/CZVfcuJGmURy4iSf7MmnCNUcnE8uTjUi88Q
Iq20lw4wIU1fL/4ZLIP1Yv8/HIYWlcZO4liaIBUI3yHhzZ0dnqCnbiiFd5y07zdQLjVHDJseodu6
j2gl2fWWFUl/uC4+hno0L+F5U7idcTcOFQYuYXRQIf5l2DY1SOrjeLeGclwP+gGpjnlGgpp3oL+v
5j7ljZRmqyf3y365eO4SV0CchkIhW2X8xSQBYjOPpfIsfcHyxSNwkaqPav7GJByANlCTsLGly6Jq
NK3stii3J2DPT+qcJllVUr8IOHmw5gxsuttpSLLLNmDbTQ9FBoGCkAyZUg8tB7fymCFSj4nyPcqd
E2zCd9kqpyJ27KgBpzp1ZULslxl1tsAJpCKm2hgegZBtb3g+/PnDn1zOFlW+lqTKHOXbDtycybEd
rHpFBO+BvPxs6x1oBelg/8qBzaAOOtdx7lJl59wIWWZxkxSxkOcxI2DDNNZpFZ0ItPYSJiZGWfLh
6JmPnnQgybP6CV8qOZAtdt6+FL9SlLDqQrgFqvk9Qh8C1F8txx/lMGq5EQN+c8S1a8hKI0FrJBR/
czTXkcF1hq4/+Y35BJ44nEI9r27wUHi15G6TdAEarzsD8m1yPKuHl52euU7oDr7ewS/CkrmCIXj2
W4rQs5l6fL5rfIvBtG8WnSzuP/JgR/FBIrbN0bvdyv4W0dScRaL8L/lE0AJu4Y9Hz/PAM6abL019
XPzc7ptcj6PhzDt9kIcjcM2tYZtNCW5T5kxzb9QXm5SLSocB1jx/nGTO3y5629G/NXEBXPIR/mF8
vHlNivdlwRElS0sv6qfMBTTm2KbSlDDx1Hi9cu7SD7PdEthl1mtw94QutFtgg1NaOqZaGgfU1ovl
mbvTqLM/aMdWsdCrISdgx6sgMbUSFOyz7Kct4YtL/a/BWw49Dqd+NrCIgS4ojdHuLdmJ+GxaLDl/
Kmolp+iZfbYoJ2cVPAz1brNpCkFPi65GSDbb3SqJtJYT/Bq7S1PXO7TNUvtowHc3S0yrWpQRcOvx
ctQKU9L0HlBu8w4Gl7a/7fcCChsIW/u9NvKlNryJyi0gcxkelurQ8fAnaWqwkZG5cnvd9nMmHX1M
Pag+7DRtpRdtLZ/ltw1nvUh6i+1c6LdDzk9dUecG5EK58UU7Tsr2NdnexvjTAfWCND3tzIHU1fjQ
7mmpXIrnWfmU1zlOPYsdtgQE8t7HsVmFLwYpuX2L1Ik1Id6qfc0VJJ4cAcUPUn+iQOQfta5JQ4iw
2gKjxgDLYANabE0YcS6Ew42aF5WEeecgN2gvwiANSQ14hfvXX3vDCpbM2bCudq71utUIcbiL3SWK
RAhcMxjxFchLSOLoxL24uBQ2Ui+b+49cHrtQpgI2OQB3v3/JZ4J6wKzvNYRvD7fsbG8K+AjF5uqR
Jt7hDHDflOo1dqNbjkOefk7F+1ScUjZq6OgLzl6xkwjAt5WrMkf4pDnkPcmKNkMoWyQvGI1AtndO
SfEPREoWSBWJDZnjkb8h/ypOHiuOcuc4zV33L9xPHumkMa0yrwElWJZTdoe0FfimM3O6jsPrsQ/w
72x/pMLpj7SAqICMzJPQHUdbRA+o2kMrqA0lgMh6cO7z29A4JtZWY76p7hV05q2UZci3x60QbS5C
zhEC21wBYlemKDE2aRoh1p6bd+doZ/oVhLjlSfkfrxA3mpaTIsNhFVvU6uACInJS23ldYQpf7oZY
pnThNRilUcPOoWQz6LcuZWPexTcBiCaa8gIrcEH5lgutCKpFGZdTYGY8V8hUry0hgZdMNoKNv4Bn
oz/LtaHEaLtyS2Q6qUFgm26KbD2d2znA+gdY6YvsPl6MmnlZHDT6R6e6DHyLBQpNQhm+yudSOPRm
OekbM+mTMO3epiEMUzMLfnBYZJZMUSnoQWrRAFr5Wj7fBsLPNtcxClcgv1yM+bmMkD2RoOX3+2zL
12v1ggX+iT3iPjcX3MdYnOzzXsqbC72QW7RvtvWIGeX/yFumUgQd3qe6bXI+GOZBkfKHimsjP3FC
dO9qjSlNAt//GrFamZRQqqRE/6pMrXECa+8hl1zQ+3NJt6resFVN8KDDE3vgdXpz7kUWwGz/NHlM
YvhKlGqLdUhkIuaMbWL5XoSyo48cK0AerVse2cRzblgVqU95ktDMChmfwlmag0ecZqBhRJgr95OL
DRpdDdB4Rqa6SEsW3FLTitELMv7J60fB9HrCz4YXskjWPHZGuQMkSpolzwSx32IOLTqXU9wDP0Ip
Wq4hE8NyTepDepxlMA05ipMjxNP0uh0Q32DL2dQtBWpr9eq9AdGCiIGf+5BgShs7Hgb11YRR6jgt
VT2cNiC6T3X9KrxupnYdNF0wR8XwdPA7x23DqbdJx8njjG1ncuwLodEIxDmtDHH4V3iRviq0yiNq
c37UTwwFAHIlA5t6GgRcDNMiSF6x2Nhy9s8OI9yoq+ciHV331skg3gOxfxufdvdLO6vhRtEtgw/3
P1HMccmkf9xm+Ys1syy6au0hLTu4Ti8JmfSQPKw3ZxP0I9Dmdmr8bFzQRJTmVjuFMPQYaFCvlpoO
E0kbLranDBd5X9Fs0ZqYnqw8UXNdec3hOJxN+faJrB9P45FIZ6eqt080GZBzI3FS3mx8nWpdcHMD
RJdnQYYipbL0iTXcl/wnQnv8UCXUK0vuDATDdd8YNDFXtuhVGoAT3/pzuZ8JkpXt/56ZWseuJxP4
GhT0uK+qfmdV1hL4mVSqXmaImyvqnsj8vl429hZtK3pgznMXOyMTMWgIkT/MFeREePB6Rmt8V9h4
gdiHS4DLcE71NfQnqneN+7pFZc3VPqqiLOyC4peyw4Iiu7ABWNpOTb6cGHAJKOv36EnLodITdssk
5w3XpvYSF5DJUmIll4bAa81WH8hhP0D3FAd0BMncCx9PKX8WQ37wUgCIlfB7W27wPU9S4dMaEaxM
/sAI4SgOE5gigmjH8x2YROzPOYZTLG80MGWH2v3vCLUDxcvTqJJGV9H2t9VqSrMGMJnOTKWtgoq/
33MsW1pYs4AloMu/yr75BH/Z51vDqWOn+o76SyOmIs38d8ds+N5CRhKwTMWmVn9A5bcsrUl3kump
L5E1eruaR9G7say6NOlXBy/2wLEEh3NCw6aTWQJLaY1ZXFRwxFT81eHQ4PZxrRQNvwq/npXtpOui
6LLPKfPJYlUVS9wvLZlmJh19Rx/8EdELsN26tz6av/+46guX9RzrrpAqJg1ueINrMGkMnn+SKc8f
9X/GreCkbFFB+Ajp69uE6k3FMLwFpFASz+mQXh8y5fqmfyYKi5BEzAdstKJSiuOOWkzxhtsKhAQx
6Y7mYx8DNPEodU2C5ASrbYHYYrw9XaGL6lKF2iVqyjgYdrQ4YFBOImwQj04fkC/ndWL2mWUFL14n
ghAbN/nESXZV1arFadOmE011Fj/OJc/aKTph9f0WDxAbAgualyjL6iOX30PHIgt4mb9S7rLuA1Na
8jgzHoGD+VFRqtaQFYThBoySo/7mTODldveA+Kt1b9yfm0TT1drP7swUY8vW1H1yWgFoETW9LpVS
0D+SQgjBVwcXwz4sQ65j8TJpZwIr3tn+s/p8HzawjxF2dcZq44/G4pht+u+IbuKBD2UmcvSFWsHk
ap/2xGiYr/xxk9hU0/L+0Jroq4LGVsqygd/mdfbnHw1gxWjRCWaAwZWbInBgNL7IdJjkYyv1oY1r
PzG3SyincMz3yrt803m0TwBeylQS8MDScWmeYIpt0ORkRIgimI8xck+R6q5kOSNvdk4l/x1Biy/R
Lm/ubHBRkzYEbSP+zZtueNvRXeCFfsUlxUaLj7EcoIPfyIXdkv4/76fGzO51KG1m4ZgaiT75bTgg
gMVoQX7lZ9wwFmQQlXF1L3dTI/02gj/BxTHY32sBnP3ZZcQIapMtXirlhAcr/e2o6bDZYOTD1JwD
aRulgze/gVdZfTpqjQwNWeoiKL1JnZlyu6WpjC3tmUWDdW/DX4CbmJuinzbNtjnRCbVbkxpmTUTR
pnGsq+vFyj1A5snKKEo1e2Ha0K0JOr77MDTfHweLZFiNyZAMMe5V1fTrcX/hM2N1x7vwEGxiXkNH
iu9FR9aDmoU2RBTXURyOEyJ6qcRRUUe33ArPoJDMvwJWfD+QxFom4nkMULClX3s3dM80FkB5yP8T
lhP4hQ1OlG1wLyox+mcBZJIl5A5F77SNR+xKX5hpfgmWJy0F3f0oBCLJ4eGVtpFnLb519wlEkqY5
lm60MrhJ4rpi+YxVkVBtQsmKJVunp6j9eAXy/S/lB5ffpxXVV3jc8aUH2meVlmEPG5Kl7JaJ5usH
5dukbIBW1r5KUxOaA3xT2lhHdOMChHX9bcyk2ODbVrZy3YQT7893ZeRHzXiG0qVgXDylXQy7S3XH
oiitpIjFDWzaKyPYdO0XwJVtVEYCfoaUkMfvcL+/tHnxx+Bsg2sjuLHMGsvOMOmNSnQT33N5zXGZ
mN9kKO0djOSJmWYXi2uUkMk9CTF5Xpv/6xtXkrhvpRDf2yoj3YBTwk41EpFfEHdGoIh2KbdqYdEJ
aIyE2W73MwvP9Ma7QFuIuwyJHl9m5ku2JlbjtahJMLDfPlqjNU96usU/HSJuICDfbDhcsqNKNyv3
uMopLxSyeUgWG7Wb4n28pBZd68YQxSgcixxAx+AkffrHT3CR6wPxXQMFfNwtcvZ/sQH+sMdVN8hi
//5D5wIDrRlWhfNgfenqlEVoPLngq8L06lQiaNOoGlCa/m317RTh3vT5oNIaBxYc8rC/3GOcBjk4
p7l1283awNYf/1IsW/kAG/RPMJ3RrmDo/4tsLTeAzau01Zph4G/6uo0OoVY9E858CIxIhKbFShSD
DXu6EFPYDC1rB/T1Rg9wmzXvkt+7oaqYQuaZSo22GzlRFMwzu0Raolt6qFYItbKH+YjgLU2PRJRb
HrFI1KV5xciVXWzkEYUFKqLYcRsFHlSDF9rBVCYiCpdb1MiJeT8UWxkCZnZa4aNjpycZRTOOBlfw
6Y4NDbyFDi3FO7YWa7OuFR61nY1NGGDOuzX3ArYL0ebiRP09CShvPC5yO9lwuDfVI4SeRILIxwRE
4ZQ1KQDATBOBF60uRJPSJrT0gGYd8mY2Iix7Jvxr3bBSvY0H8qmJKAx4xURLgcmzv9GCAKZEHru8
7u9tqY8yCeM1eNH/UUuiaSShDcmvN6hPgCyTSyxSUOkla/cCPe2n4oi/fpYhcnowRJ6fnS9HM+U9
GBFzr7Eer7xE9YUwiC8DPyxUUWgc4bFNxqrXCGsGBFdsuOcZOj2lMQAYHk8xYt9296G8H4ZuFJFX
GC67eKL421fUY2d2qEXjpa5E35gHClJ8EOK5/Embq1DXB6S74+0CVwjF02gkx2gOcD0IDUu3HY2j
CT1T8Vr/Rl931UKYt44KJnMbr9Wd8bFWJhFUvQXWwLlfNWbdYQEhiCey/w+uvYb3+1oEpqiCITFV
k/S3qhJK89Qi+4OUDc0bNDmGqL9rA0hs+YDsdJy4cZSSX9+hS0cvyYzTR/+kfsPL1VrMpuvKoMqp
Ksp2AFYjaFDG9eaJuOe61paFdhJidWGYGPJpqhXhPIIHKMVFHJobz5xLlMK1osMgjy/3CJv5qs6e
DI+EIA7exN57Ahmwf/UHDJKlMHajSFfYTC+42nn5H908jKAbUrY+obRLnECG+eJbB2w8iBEnjmQW
0TcxLcoAF4Ml3OxC9HtYgD+C8eAxPZGfzwf6lGNxLavAJsGxzS8lV3BTINHsw+vJ00qAZvm9JIo6
AEERliBV5YPHCZ2gALSy9AN5GVIoMk76kmXTnG20YQCWoulRP8L6CvYot9Kikacn31cZhS9jFiVw
Xc3IBvrsh0K4TtqtRDH522HBpjg1GiZLUl3iOxPgxzGJBrunFW6xC4DA7D/w7eak9GOlV8pCfdBh
YYLtmQu+LpVk4XRQSDW1z5DQeAAA3Zb8k3CUbrA/u9PUcHNexbse4DQVnONxsNq6agZ6vgpOkbru
jxQx0MT/o3m+x1kbLWGLbl3W7c68vXTupIzNBlummdMbUilCKFSuThPktHlVqwXXGeT3Fuy0SQ6Y
V5cRytGsFoiUEVIy1Ik+a1Ad9XxpNExva0vMi4MGy/B2q4K+Oig9yOW3OO4E1zn1BIEIuErv/mZB
+1P7NPGscKcopGCfUU+rU6wNFJIzcJGbhgN7TPPmj3ytrdADkbm/3ShiM7KFV3ogCapTK1W1GjrT
GkYr/ary/sE4HmewyBO55i0PkrjdVc5YJHKz72tJkl3qQJO/LgqnEg7vES/dcbP5x3m0a53kj0TG
xh2sCGzAcyWOa/PwsIFGqal7oWT5+mxsNo21TeZGs+cX2hhN8wuQFsB5Ce0j5eFwMqGET0iFFps1
6D1BRzSDi87DdNkOmnwz2hi87GeDirqWr/II0eWN39dNdKTY0dEqNBTBH5eDlfCAnXCzCU8FGvLH
8iE5vkDvU8mhdwQwEjH0AW7zWt8zjSRmacE0pJE1vR6f6HaZHJ+Ehg1C9WQSYiyAGC4K50CYSP2+
neaaFFZmK3N1UXTir3Oe1pHTCWCEe1lRO2WVCA7p3IdnM8wq48FG5fUasUI3isk8pLKZ90Ip+p+R
f4HSZbhDDbSHOkF3iQr2d/gXjlS2bRxVKKNv+6leEECFrvt2WDnntfcdX0b96vg+HuhTr7vH7atx
EHdYHy8wnI7wADfLwZQQEvLONm2tcOtXynNTj0nkTjYDz6/JsMH2SlCZq70pOlowxwJ330f4lANo
HemJZtZlLMFm2Tl4wokcsZW3pK4ZBYu7+vISs+pTdog2JeiFx1kUblTxaSYDfONLEbxo+ZvNLsxe
6DN2mKU2EtHQw3nC+RVuwwFI7/QwWNOC++7qbuAuuS0V/YKFaamuGNU32v/+9sjeNyrnFjcOcZF1
hA5HxvDNb1+yEYYuAYNHvHhZPW2dht63T7P1Kdzwnrpd1OR158bc/6F3BWn/eKxpl+4xGQv7pS6W
AU6oK+yCgUhDJGarwko50zxgcL6lThRU6gSvCDPnm+n2j+2lLcnFsi71mBp94ogsvKaP8mg37QTP
v/4/heYOpI6/bHQrScA222LnPWF0++EFPGVULhSZGEkDHCw/BPT4UAP9o6ksiOeGyxxDLwG8ONSV
kY2syU2BZu2aXD223GVZPTErLL64G3qgKf2n4kV8QO0O7MjYtOEJuEcRKt1OFRxXxwcz/Vqe4Vwn
oj94Um2Gx9fznA2rIPZZm4DD52jv+253WUOuc+ubh3VMmtkAkic3wR58KTuH26kHw4PpWI/lmRdI
gTy7Vh0PnnTC5QARu46zlRY440h77SF85iDWlLt6Ywy6VR779fg2rXvpC+mZAI0G7FW3UJAGlBb7
8UKsatyVK6DdD+clVxrUvtvJ7RmCV0y1BEdZHPhymffaM4v/MLAdBu0W5CJOddFi9MlIBGxZpL2F
dj6A5gKEf2yg7dD3MfEI4JmutKf0avFrg3WVTOfwMSsrrDQUx4QDsUsd6exrUnDZG5Hgq7FQlUlo
9FDkgmMfwckxp/oq7dQlyLuh3NrWYU0Ic29GkbEN5rFHog8ivLb8mq0quV/c5VeoEte674cAYlvs
L1n/GnGZL4kqLg0iYcxYBSURlAARi99XZHNO/Qjp4M2qpIUJbUOxE7bRXAoL0UTn6ldEbcrIEDo1
hiaGpoZnJFJ3+tg7i7Kc8TJcSvHbvchK+i6ScxlL5KOH+H/04P+mDNnYidt4i1cQXxd/mrfs8lPG
lIdfI0PLoMgVtsnyI0atraahtqFw9T00nx1L0E+l4vmzmOYv0IcuX1p9smmkz9VcWBtk+6dtn9t4
LZ7Gr+0FCmworw2GLA8k5r9v6ijqRFIHUEmFTyitRgq5smTErF4LWktu8DQvC2BLl4lrzb5VeKFl
gZGkTE3mjWBvFfYHqVYuvof2/6FCIeiIRa5U7Y+CCV34tBKG/3yE4k1BxxFq+Tfl8t4KOv2gAI0w
m4+W65qWbgVggA2Hx/lNM5A62/X3FInIhRxrc7f0562oy/BVh4XNTdkZ7HIdxdS+ynjias7jpqIX
k/jxpt99viW6MdRxZK3ehSulhq78xSXUGCkz2RP5sXnlV5X/fm2c7ZB+ScyHLNB6gFIGRn9dN5Xt
fTK5xY/J6WLE6Rz5pph4CrgUS4LeR9cZ2oFlmDtxkogeVpEg4DD3baBz9JPDWQFrCCmiTHt14e//
sfFfLp/AsW9oJbk7fEcmLLzi4dkqlqOGHCvrAProuVe06WabXSIMIAK5ydgU2IubE1aSxihriw+1
sKuvOD/6DIEMiGzOLUhmZsLCZo25MGsxzUCCKNpSPebckTJndVuZ9Ca0AP9m0fTD+H7kam/cATXJ
SP0Q6MVqPAGMu5q1+4WKJmvhI505fbRzpn2nzaciQE/2AkhFikeVQI4adBIvZ/kzETyz/CVQQ/+h
J6VRPI45h7SR1DfqURqxLYLDTCvPsmvD+i+H2M53Mz2iHLxLxhSms6g+lhwL04AEZXoVD3Gi8GzK
P+/20rXvhpuARJmpTxMd4iTOcvn8TrCK7XiefI0+zEjT0xUYVzsN6n5CtKYJQ+B9LzVWWcTNZp0L
yssEqF9+3fbO6+k7Z1ejXoUPDecd1s0NBi4diTOFw3Y7YKiFXCh7RDC7it20BsBN98cRKL0sY2Ij
IPWj4OYL4TBaT/FT3RDISJ2rZBivgD/LKuEtvAZv/oxmVt2cc4ORhoat6PA2w9PQ4RvcjaZN9Miu
+bF5c+VVa206OWkj9kl/zmk5EO9XpPwWFaKA6HdMEQ2K5+M7Mh4=
`protect end_protected
