-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "N-2017.12-SP2-4 -- Oct 23, 2018"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
osxJcXeZnVVnGNdGmUJbRduNxyqeV6mlWVI4ImrJnOgvncP389wM3dU42zTaOFJf
URqz/Qy2/D3Bm7MPoBJxBZF+2M/ravE6ehJjLKYWBrcYm/UlLE0HbJ8qNFLI4p/y
erzL/mKi/5yutCjAAqkI0aas+Q8+RknclEqfJuWrkV0=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 23392)
`protect data_block
3yDzeormxWWVsDOWJkkneFh3MGi8nBEU4TzQPX9ArIykU1+vysaLL1ph8YCPkOQ6
zxEImq6YspnP5mYi5I8n4L75FVhleyA26zjNz55z2QrdeBlOXQrNzb6o7y8d01UC
nJcLNtPs2lvUbXFCYjC3CfvMX8V1rlh3I514rFOStxlkF4ZWEHcJmmMYPBvelyix
gOoPFiQ5DlVfm0ApS5B+WZM+IKWvdEAWioN8QSYwNIAxz/C+SiO2/wovclmMo8IP
QinRYFWHWTfTuV9trKiVGhTPhg6PE3ZsZ05gPCxcghh87wgzYOBxJhpD/+PM32HZ
ZNXI1SNikVp7Hhv1+mscPAtZ3LcmO51Y8umKB7FeoHSBb2NLGMJLDj1+TGLxn1Vr
ImZ4yqTbVer6J2feRjouGjBEQuc0n9j7lc5DTk4SsCWi6sKGWc/x/iQ5MWPylYYl
3I2Ykd4e2nA8zVvUQSNqUz++CFFoFgyQOm/RQGI1ibiXjsS2vIVE3Z3lxW5QuabO
DFgZ2p9hOdaTAsm2KBqo5rXJ3G5cBPoVvKt+o04Lf7LVgdBAdlID51Y4Y8KZszfZ
F6xWZI6OLtF2g/5I8r0nhhvQVXK8GuyK8Yn90Z6KVTodxPs0qdmKkd4VGxmhRL/E
EV/tnEeBthM1UwgUG01uKFPN28EhayH68DEoQ3dMQMjpvPr3g06bytHSHbYxjasv
Gobb0Zvgab8fyhbVd1uo8WsWj75Pe0WidBYs9D0OSjnN+XDfpw+edV8lbBNaH2Av
BrnThn34B7MVIppex3MsvUPsyphKHQvbXZRIh9gCkB1fspl6WEptos6raHMpv0NB
za0xEhHn1lKbfJ+advEpvXR1yqB4KgRwfnIVdUy/aVvxL2Xwln1qn3KeCxaATxpH
3lt6PGhaUBfUbzJHLjJm1Ql5g031Wm1weB9GslF7I26eka3YTFmlTvG7gtkXwGfN
M4GO0KTVQwiZl7YjwnSpAEC7EmKfE2ssbSJFpbyYV6p0ShcMPYtNifHFkV+hOCCq
jFtvkbSSyDZjStvViaFUpVbgLl3+20/6ew2fObfo0d7QdB34lpvbpepuaRL2fTXb
EqbJN+L1LJi7afSB9RMUdvdelhkqB0UhfXkcZGiHULbf8CUA101VNBEuE9S13rAI
b5ajcuOIYE7CJmRuVqEk41GwK3eti7z25ptPozgdnI1VfXJettZ37TPh5UMU4ZyI
KV1GSl8SNtbKCtAXQbQsMMRqFVkbDSFOsGTPonDbywQZ+TvBBSbV5UpKiOHZ+3Y6
2chDE6X8g05aCK1DKa+zRD6JqngjxtWGCj11KoSYrWplIMjD0mjPcdpP19pFnabt
wYvc0ZIoX5I1AMkTcA9BPcVzAa8pcWvqEKrEoXws8H88/ncpk8rYkjwCz+hX4lBv
JHfyVjAxwLh/gdo5w3ypWRK5CJAxhwqgOXIH6JWplmNqHNR6DPV/Mvo9Fq1uhHPC
OYxlNyqLUKwlIql3IBrOrZhMaa7ziERX208FC/a1+x9G+5Jn+cGo5kYvNaFJIKWY
qsijSapsaOO5CAfcorhcjW39E+iWN+oM2me6K4mRWB2Q78/Xcc3gRbErV4sjl2Xy
g9iHvCcPK67HFQpzeuyi+BSGA4FffR/WzzVqxNNps0LHbget48HfJHrahT3Pa8lN
PFbz8v3CEZ84G1HfiYej3emHZbneXKh2vzPcLdCv76cwPOew/C6stzn96OkjEORw
bVeFHjHnEK3nrvZuod143uWAkgcaEE0avZZab+HgLwA2sFd5y8oQBR6L93cQB/o2
kEWF3wR0fx6NHlmE+eBw+oY5hXrSvG3HRlUidj0ZwhhezSOY6NMleL3v4kHCXF2L
JtpCzQqWVyj+WIkCoqnF+D/qZE/zer8AmoJGVlJ1DaDWihLHWGCDDZI3esGMFK17
vjn1szhOJ8BkWAVBpjhKPl3koCZaG+Nc2IvlEIcIfGC5tl7aX2RmwLz+tZtUslal
f7O03GHcZr+kesElMiLE5N7uBTaQ0FIFVokOdZxT1NJ5dHD0NiaZwY8EydsSIfER
xIma1nbs/VvqoAm2zo9pdiW4jtlD+MOYIQw30QSdXtlsSu4tq00Hd4g4Eki8Of15
dcvZIJNjMtdv2PR2wwJUEZrniY/HhqMi0HdpDW84PZt8IeR45g8Ku0a9rsOQF92q
ZQTkhmrTDasX7OObrR1YIsBWyeZSYADYCdexhxQLAnOaAVZQoU2ejEsMwNrcpQYT
hH/FQ/O/0Oi4307TGhTxw+hHmhzLdt5fGxPRBharP/kMz160AJAp/xkhFOxw5d+u
4W0w2YBuT9J6nju95oE3ucjn3kNmGuTtgtWRU2ceU8HHpXhB4gxwq0s5bVv6GeLt
Uw/OSLpGnsKUM8yCmCiWY0BzYufDMv01KhoXl7NvE0DNumGXBqdfTgt08VdHBeG/
sGg4Ort2zIlshEhFyvcJX4KZh3KKYAMH4LVNeKYys6gkfjYwu1Rzr92oVAkBCjAq
W+R+UtNiRNS3hFpZ571YT+K9gOiiOpO9R9JTQwdRpAr094hIr9POa4suz9uO3gT1
AP3q7dcoF+jI6rPfIJXCfkyE3/qH7l8iPd++DCXZiDlSjK3DPFvNBnF+xUIamI35
SXAI4qBdDaVGMIMmy/V53nnrWqK2s8PMXRemjbnn/eopX73yQTTaLgpY03RZC2NX
GqTSP+rfYhb4dU8Zx2gXVTkNynGiqim0gbH17cVpEk0WqqGudgADDCRBbrAz2qS4
rv6W9THbjOgO/Bez2gSia0JIe1+iuKdJXLVFV1DnRCbbloxYSZWsHR5Nh6bbnRJf
ItY59KcAAt91siwLyI8cihuRVHdNssqe55XfJjs7vdcTsy6tnobXjp8vnE3rhZqB
nyyaDKKIsY4xx14YUYl9VDYTADuXojWKzX+mcaJwKUt4T5ugqjHHlLyJfn/qPoEC
E9DQyCyKnUhc9rvP0UlXCLrlcMqEjThGHbOhRQZxacIxaIhheTQXmHTkAAQNrJiT
Zm7bl2zhbR/wIzVWvxsctbUK8YpmRxhGb8o2m2pJys29CDW28DIMunLEHQb4Z5Ti
/0xP6O/t/1sLOWFYPDaFxYSUYdlsghVIo8X274P0Nj+noSaMngos+JLWm1So7JV3
NX/VfBG6dhntHD95ABaEm+5V+00wlKWeDHTG2qRvGi/Bsmrvmc1JcjJJ4L4Ob3bc
WPKTDFOievtngdGTcrDkvElcfgMwmd5Rhtqhezdb/GgbVZkvBKa7wFRWDzBp6T9+
z9MUJZApaUfPMW+mcNH58Ddgo6PS3+sz+CeUXSehnf7t5x8oR9XUYs2sBeN8UstX
MEBYWvTCSHidyQiary+HKlhwBckNHCf6A80JAgMI82roB92GNwUsVmdDkMaJmWVI
tylG2KFnEkIJNGyb51nu+Ktdg2KvBdr1xwzDvdWC6aqaKHZNcB+rPHtg5h4LOG/I
5Q9oERisZXYEnkjwYPubIQ3aWy+ui4b0v6a1FIUG/pVOCOZ5fYdtA5E0sJRPNMu/
Ys5UeEE8JG8+qhSpJCd/9KyFMl+0FE2Pc7m7zRsCv7BkDvLS5/NtdJuUGBDG6StV
38JbsjeEbDsvu+gCE5kpSGxM8d7XjTBulyvAhqt2PsLI9xZcBclMOQFZyV6wmmRU
Gw1WVbX5NEHREpMbqeC2xqRZJlsRx08alOV+HR++pZfAfhp8atkpHwCigPrRGSB3
Xb4I8SF2Vf5I4Q0r40MM2jhtJxTUHPfZGeE0kCDZD9+jKYYhhZIAEvcBgR8AGYHG
Upr2lOm08EP+vfPcxxOTY26Pb9xNIsHXBXpU7FxYJPj72pzPvyW1CXV9gKS6rm8s
FxbLSwJqz5jeqrpanwef04VYC0D56sO5ufdNciLmoBGIWOaka6/alWR2zZvpus8H
ZEm6ouY7FwCMK7OSg5xCh6eUBahsudRidPFkDyvSrG3F3qtqtrg7Zkb90QqbCxFG
1z2u0BXyBI4M1vXG+NtXj7ugNWwUEqwbBupdC75UxTv5zVe8jvSw26P8Xp+8aExB
PTZEILYq0VT7j6/7zwS4deBhg/cubNdKpDCGeDpnq6ksOjEIjU2L0Vj6tHfxToNW
pHHWgI4yyn+wTlio8UqvLCQvXLYSZ6a91q2AtqZTaZF5zxQycdKTDaIeh5CZ+yjz
04Og99OD4BJyJEd8PnZy5AdylUaK+3enA+ebdzY868rsWpFzLDQ56CCwWFvMJNhp
3j+YYGNsL0yl8NMacY7STT5+bmh8K15OsIQa4Q/F0p0Eml0Y1hVu7TSPsWWLERnh
I5nzj33wV9X2M5C0F8a/Y9HlR/jyClcBfsElauZDHWuUuZtdjiKkobs7vCtUVr+n
9uDcZRifIo3kgQCjl4A+2Wn/AL+2s+oSFskpWc/U2Bxut3Y0mwvPydLobvjMGtke
rX/+xFBdArbfV8yR+usFcZtApoQnrNGyeZWNcv3Ye1WfHF8r7kiKwGMAEh24aXdP
4/vNs/p30xSogHsy6lZl+HSTa6SNKtmvPc7EKsXnj51SgpwyI2CY09qmjPczD2kH
bFKdJ/44XbIw1MSp6LfW9chdJtw1Fa/l7SGpmdClOkzyz8e9Jvq7NPC2Gy27Bugp
xBPr6DoI2O8E7cc9r0SS79RELtTIQj15Q8k+m1q3WKO1GMat6tyBL37vLJRM5L8z
GWAueWg2HxzcqnH6HeKITPlDyJqIBZ/Qdb/Fm6MYdK7WMHqqOxowRQ0i0LiXym8L
Ny+yMcJ84mK9STZ8sjK+uz8F5NO42Ww0YFkq3fD2IvsiV9PcLaAj16CIQgKVKkBH
V7S87wjimeerWX+o7I6+fSOml1zJ7S/StbN0wo5Lm5lLP1CYtMOvKpzFCEGkPHJg
5u0rCDzynOO3XT+3qYFLDmCtvCibAwgcRJZBcgRCzd+Q6dMQUBzYsGT9rFQ/92IM
uYxDEbEJznONUS0LcNFxo3HjfJ0UXcjz5La9pxFfaWv6YtCCYyKHrDZidb44QrtN
yV1M3Yqek73ZuoOXtCiNTWmtQOkhSPUHhV0W5OTXJiM1pwGdwIjCtDt1sw9DUJhe
kAgRnVtKnpmRvIeZEXEWQ6SWU7klTpXcBCJdMeLyZa/jsZ28aO+bM+JY0j7MurJv
FjZXKgo0M0AbqfDVYfE/xSSR/x8Yy2q/7/KueuM8UvYEYkTwgo/vY9HYb+mvZlhx
F9D1+43cNfuJC+IPLdB0Acl3L5Le0lMoNFdZY7Kn7CMO0C3K3bgThzsC87fS9LzE
Q6QhWcQ++9enTyC4BbxGNW44snONhAsjLpV1Q8BcJhmi6P0V+WIZ7eQzUG6SDUWT
njFRm4CYB0y2Vrro59DLFKl/MISUHSK05jbysqUJb0Jyn5tRnLp400BqC7cgrO3o
luoaUCMpsE2/RmR+FGYMX6Tv8QS9T5Ufxw2clXLaprj5uLWJy2oMOUIkn0o46gb7
uVc7QdwdfgojLnevD3vhflwLDuRKwgTL6GdOA3+u3zaw/GFRb86NdhYMyRTmzY3N
eozy0YlWWFt/7MCTRM6GsNWciaJQV44HvTGFQLr+WI0ouXpEHG59HxdsMdqAiXAl
rbyTB3JSsnuJy53pwhXxoKIUa4rUOM4muCpzO6uf/h9n4LY/DLT8AkdYVmu+K3xA
wqM0vPm1sXx1UBvmqGoBPK5eQjFf04/ROK0XF4MXk7giNwhQuEz0ckTwbtEL7oge
Xl/qca2FzFlXU4zp95R8TTzp4Nd5jFCZjZ6n+FI0pvggMMpw3lRp33AsNUzpOeGL
tUxzCOe4MErs6xYeaMwB9/imr5KOyC8FrOuZP7zO5GVjaUKnmfmBKTlY09Vm73mX
3ZfZ9TyD4xpmg9j8i1JzsbE9OzlhCVFCIv5Eh5Gp3TzT5/GhTyXvMscvOy++Q8tg
WIcRw0f898oMVOeNyjsQef9iS5Gax1CcIJU5qCmvc2qpPis5UOfVl0Bs9YNwuAnD
t5L1zpi9cxriM7AwKp4ZMofdrJ1MB+JMqMWwgNFn3M1Rwsre+44lQK/Fcu1aQSfV
/2Gz7KqYX53h6KzAqVUn/NXulQJBBtoPz4APxQ9Tdv4AylEKFjSHlPZuHFhmFo3s
Cdc7aN0p+lYQu3Rj4YhIJEGEelwYs8qXXAZvvYHkVTluH3QQpHKnBVA2oAa5VCqY
gqnyXR9o6UqS2OVNAK/LX0YQXL2DtSCiUwx8cYUnrMrFeJtUvk0NMCwwxSjWG21j
/rPI4Qey81koc/XasGzUI9+u/M6Wp8refHMXStITe88/0sq8rMjUrQIyQz+jJj+A
VPCVwbYicfqd0KjcLRw4ZVKX8W+0m2mXi8cKdSIk22kxrqHyCImeQ2vJhHs2/xiA
zHx6GEUo6GCFgzBZpmSDzE3b2DHxE1affvH/Rbza6UJ1haYHGTWX4vyFQBXhojJs
qzoLulacWGs+goZ6pKPrMO6qC9uEcgRE7sO7CVQPaVmKNX+KRdIpLid0L47xcmNo
6byPX1tga1R+IGz9pHZbH5pLdCey1U/0D7V7bEQwZ3Y5qG128EcO9m9GTsFMhL7u
p0mbVJYzi3nk/HfEh5RKkdDsxlWrVIuUJKcddOg7Qc73DZroD82wk9pjarn45k5o
SJsDfT2+AlWY0LxW9QmdVNEA/gl3VEJq2bdddtVJCkTnAyDtWit/xXpHjQ4SKeQc
SWorgSXaFWK5OnkUvv6RuOpDGKMqyVGKtQ74n+CzdhCjAmea4JNUzoQhTNdpawn9
xKrbojR/2RkMaghZufBrQ6ov/X20Ie2gtyGCE1N97z6E+UE0hfm9JHeIKvzhMW1R
h0LAAVrLPMNUSpAPZkLX6E18IHoe+PTpXJzQEpOUF0lSPFu8KTPxItYuTu9aL1So
CUxLhbgTy36pJFyo8fFow0DU5zl/hnYI57ABfe6AHXsyNCEKenTzzxmEtT75URmD
O7qdSawdy9bGOpaf0mT+Cw+5wfz94qbvmcGaDLgdOyUD6H5ROArVWK+sJt9x3rh9
O01EnW3B547pp3+Vl2H2UECBbEBPx4NL9Jnz/WHjOxkesWwb8iLptbsQ9+dN4J8Q
y++MIP3Hf+4K9+EwTaOFb4Rqc9ZaPpxOhe5x+RlMLi9uSQZYi/0WVNg7Ads97h5V
flYeT0ScTgn4n2Aw9zQO4azTI5hsxXAiNkhemy8HpXXL5/YMwJM2ukcGch4cFtXa
npHZv4ZE8lj/ZYLVBhmB995t9zScSurFMiSSYD4OYu94K2Cau49yhWpe2lUlLhRa
DyIOZAvjgonTuuyL6pmZhw9Pp5S5/kfMAReDRd1vl31rLko0i2gRKqYhp0rQ0aRq
UoTmmh0RHkMKTgdCdbquaiEaHj2bK/6oRbhKah8XaeRVI1/FqxTRx3nrTVbWuaFC
RFZQnUVEns3+IrZOXSwFj82scpOcuf190L6aSu0w1VNTrw4O7WMyxD3usUFxcnOr
jUFywh15ArA65yq22pnWEGhRuL4FxFGswuqjvhQJNk14iXb0Q4eRSS8YvyJh5lqX
pUXUSaAh9gQBKrrjItVGO3nq18qeR4GiHDLS/G6Yfzzk+pbDxF+ojfWOIzomHUlS
hRZlg178d7X7Xy3WBZjdk1w73krQsUfPx0mZnsXk7ceG3/LUZmx6rPQFl80Sogtn
tf2zvdn2XKcHWL5axnNyQaFzIEGLO4GW4ZMIlBmRUYzy6fvf/6trD5ttOZafWCUr
Fofv5yfttHolRU/KRf/Xgix2nqxBdcnhZozU4Hxlj1PrnYwWUr9ccdIwfouc4yp5
KAoXRNOQplc6Qt8QSt1b94fQISiKQlmdgD/Sfwg48cukdeT/D3NafX4TNsHF2Yx5
AFn8X+UPbCO67dgeJZxjddX1H6xdjmHaY7MqAbhwL7+P2HUS9zW683VKFX48Q4xq
4WpslrJ/5BL9WBvrrzsXwHs2BcuKmblj3Ll5N71Gjc0mFYIyJNVM8wksW0TNpBhC
j5hgzHJMLtb0qGUNs5OYn8qNj5Hq0Z4VJFCrpJX8zAKT/O8k9YBIm1n5n/pN8G76
YUicuDNITp+kCiXA319xY15wLKei8NoC7bV/t5HfYvDVWKKIVarSyBDxTA8+4nEn
tQGDwLdpJazs8dqQg4DcnIyLIzRrbO9JIk//zrw0nHXQAyN0mN1ZqsReMZmqF6Cd
sQdmJjhadhw765HmmuebeH/4a3U5R8dP+KL0JL/T4UtYHSg10tE+Y6Vg+49zKI7i
ppgdBf1drSbcXWgMcuJdobp9FAvEYhYBZB8xNott2v/KkcJmoe1sPcXo+kNHZ5PW
gRsuH/vN/npb51eB0ntDmAAYfRaGHDkbkUTsWrhkSjdKouv7lZiPEl3ui7CZYF0/
h9SUg6R6n54P2pG7qhFToTXK6AMYs+xJg03BZH3+Q5m9v3XTirurP0pXfkN9NnYe
o47WQgSAaaFTpEransVaz1tWdhNSGaRCLbObhfuAYeq05OOfCBWlklNXURLTAW/v
b6OKlc35vo9t8qdZwZSRqHOlUz0ulKP1GFiND+2Scj/7OFvvSJ8AgoFJ0tMWlfDR
2DM4xXol4xZh3O03MK4T/yqr1mBnfgXD+U38Shvec/8xqmX7LadS9SCH6n331goy
W+cIn93QWx/tGm5Xlo5Iw8sDySrNL5hAH0R0l9WfkghpTiv9e8D+fSX0SYzJjwL2
oVIoinucTZtd/ti9sRpKPsTnJpSxWjdroq4j4gyInFWwJd0LAuP6tzJjAsWzQSVk
P5oLEMdxdn2pg0KXDcf9awcjWvLqbOmJvuo54oxu3DBlbmjhwD+2/Ec25t8NiQnk
fsZ4Muu+UXmDVgV+a/5/OgUbxUp09PWDZq1xJLc+gocdXb4kq58CNGwUoFPrbX45
3RLyw54leG48WLyvbUWxgtW1xP5aYFTX+YwtsLfDl5hK0Dx/ZOgXHkE6tnvVqnOu
Z0Z6Fh68w6A8WJ1ZykuxLr+Vlp2DPpnGogIvxOCIHU8v9PYQDkvqjKr111WRiXqV
NTQ9+GKLndtugM8RkWuroOVjTqlMirEih7go64lCPXRoMxAqUl/bQ41g2+DNURCU
GTFCL12YZDAYivv8fQdEBU7HnCUMthYZNQv0KReepqercuig/qkALdfpHEDn9voM
FDBWJF1I7KH08vpIh7rfmwRMmRem1nndsP9eAnsyj4BGyEoej2x6NH204yXmxyB8
5OUN1Me1vcdXv5ETr4m8koxQxkBMlfog1SzNwrsrTMGXrKb36oWq36fHVwEcku4w
vNc4E+uYT8sOe+c8wWZHA8IMU+1CYvbuQeJbcJoauM/yEfS1sOFZuk0dBUpTUnNw
sgJ4HmG//KVay/IwMvnax1U6XizoeKk5y2TqgE5bTORDRHoZ74saNV9dFW1Amwfq
We4DYQybMucG2EFljJqr5PtswS7QQeNJMCvWlD6ZMxFgKHeELREp6Ns+AGV+Uyki
YIr29KctJTfZwoiYwELnF4Wq+XE5bx4q8APJ4MAG+OrJ0Qkq+oK8YQMhvu8zQgYo
VlyWb18/L7kc/Pzvqg6vq/6f30suFFws+hzu0/vMPFQ3ICo/2AbRoV+zHZGB+gDZ
jRCMhNIzGGAdSYYifZxUVPI2NLBU4xBN7YttCwjrKIi/hNbeND3rAxEOHRxFVSW1
+LB5KjQthjuoAJcHSUocsK3XEo3KVBoHczS7++Q85joq7Bym6CfKcpNArUq1EpJK
Gv9RD572wnUi75nmFtzTHn6l7BnC98oOGHIUpDikv0qGelqNDzJBhgwYRvmRGh53
iQ+ESDwOKNE+Tl8cRoHjU0ecvlLXJV5Lrn51pkNTmxeC3E0/EO0V1i1T7+o4bFUR
CTJ6S0V+y/kSwJFp7uVqZ09OM0l7EHMu6y5cFP3+m58fouOZpPiias39zQ6QyKfO
ng9g8uPnMhBpTsKDTloncuG5amOKQI7P3ZTxW56HSLMEFpb8Q4ounEdX7jMayxNl
pe/NPyGVaNVK40+rkGOK+GuELQ6AERKW5K4Juo03Q9kok0TvjPn24NConkv6xuCA
/pQzC5CYWk8WJrMLFxUSp3ohMDWQ8EzpnDQm2rwjMWqVpF1Rj52siuFGdqAoSjnW
ApHWTSZunLFGTrHuhuSdVGDRPFcxVYcRLvkuGs4awzrtTGHANKYIZkufo8S2YvPa
0YTrJCOSR6gkMAPEpt/G+x6o35gjEbbsIwpnVSxZnSAhvaU9jI2Pt1iiwRrnV373
xs9DT4xrLeFBfEhOLopzVcfZw/AXFTR6nWWr97HwfuphO5izJFkgVKCKiJrxglOn
20v4fjuMWWSTuyNjODh7a/DCUSgtLxeZXYIYfQjoetjb+pjydDgQDX4QhOXgPfS8
3ScuNjBci5iP0XbNkQ1C3hQxIWfFvZf4wAkBnq7LXq1gQjUjC8Z/pyCy271ukmSZ
UiEyMVRIoHP5Q8/bMoPZWMrNLmx4/QZWOQ9OJwy+7bEJEBOdTSj4syr4p58wMMjL
rqKVMaoyPD+6ATIyGuQ2wXm2QvHEZkKU3kQ9doVUZY3Aq7l9ZNmwJvK4SzTw6Wl5
ISTaVijS4HqG9lNI70QN8Fdqzgm1ajUSpE41+bY6sHn1HEuLIJQXwBcF6knKOoqM
yssdXwjeK5+9tFar8UyfTc+DZhB7ZLprS0wGkOP2BmXeavei1fYm34N19JLJBnm5
74soYS8BmONgx6a9ddCP8bAZyfQiEAudgH+SEQCrg8Rfw4rwc+Mfn7oO97CkdQmR
148CuaKZXPmih2sQ5mVe5XKFE1Go7EUYJ6Faexv344haRGCIDMCmpRS+iMXOBd7n
O0qB4V3X+Q8ypTz+qKONfSLKQuyXA0GYy8hng7PvjunZWb6emNUWyoLbsPXOoK55
O451+mrXE0jdE2GTPBelG5I6ZK8lJJ0yjyos/LF14FDLkjJXOz19CnMGy1fdfZ15
hBUaRdRVOo3c9b63R6uuQg3s3bA5m0MjNP3UW3efEChAtlVcdoiS6+q2QLDIXKB4
5QbWtQp1aJRPOk3OaYuKNvB2qyMKycs4bl603xHn2N+fRkNCDRUXzNDH5ckO4qao
SkvaUuKlHBx1fCabnG7YxhRv4nd5Dxtu7lq4KMcUKVS409VSnSuvAWxyZS2sf3RI
hVYz4vhUxK56rAIdc8V9CcZKH8c6pUJNkvq8GJEcV0lBsp2tEuZdzvBN+rR+dYvI
szaBvQ3MwCCJrwTVdcIyegb0VnEddiGsSvpiORSespJMM6okP+Lg5PsSEFdGGV4F
8p5njI3tPJniaFyV5DQIVNSbbxcitZFhKh+xlchp2SXIYej/4Sv9eZ3CHbQfHB4t
JY1rp6TA/FWOJMyOgWohiAAO0s/RCIRenFycmQUjyMAvKr2wY4CvuscooxsNmm8u
drhYQP5zDRy3lasgDy9kf4n/meqnjoZ+S4BNYWUk0hw6CTim9WgzuiaskYT5p8pZ
f8aGer40+QlsjXZPagFpmRFNWAG8aofg5pnG0jHsBlgLxF864yw4uE5nNEmjRcr3
02yM5Lph4scqa94R/hgaoSn3nYW214jStMakQucC0jTIIcUMLGHnxo0L8WSBM8Ia
475NsWOSyv8TRYyyNqD1tJgLpXx1ivo8urFnObD4GtZyzl2nhqB9BLxCYfaV673v
fbemLNaQ9plgl/4xvpF/p3T8BHIygtTCAZmI58gl4qQ7LDf1t5ZWf/V9caw6dZHu
NBuGUuVCtKMboUXfTdYex/9ht5wEljVNVFHmgWoBbmJRaminz1Wtln9xKkhyJq2O
I55wDgRw4/KAsv5mHA4UhHoaXKXaIQkbJ8yXbzBxob/0Ld+SRBMxr20n6wFclRJr
8G/lAc/dKjoLEZWhrizHjl+yxNT6vnmDK5KA4dB6GUt1KNBdrBH9S4rVAGR20+Wq
J2tfvMTbGncmwFhliQalR16HxtgGmi8XKn15Crk5Wsn2GQRyrqaIVDsSje5ScD7/
5cQ/KJhzJwIbexdTqj0lmeroQahj5bHsWsDjV8gQOKzPnkf+3tpgRi9/838cxcQ/
RjuvunjgydX9a+dOPS4fTnIKmdN03jyKRFS8QSt2fUn3zqhc13s7D3NuLdzlK7NR
f42SCCRtJ1MWNXMbnCA+4UvkHSSPNu/n8c2DP+KrwUo5pqetOD9CtfpLJhZ97Hfd
/gywuRcf0wKdHkUqvjXr5uMqKL8hUsiA5jilYz1psrmzrPJFAxGqBfz5BVVy8hUC
rJ9to1wzEhIFbTW82fVPOynFeAzWeBsbTAtd7tBGdF/wUKREY/IZ19LAk0IYDCxN
j8umcy19MIVcHxlFwxc2OpSIhSn84D8aIqM718oNJz+0rslZRK2/g7xOW4kTY6QI
HU/vISHJLfgkY62C6SPr5XVTICKTeJ7nDz4OACyS+g7cSckFKc2eSXa4YTE1KQOA
xWdQflE1hN7ZwYH/LHMqcEic3MV0cyHa4WUmZZSRznsm6NZV3V1TANUd9Sxd9GlY
oYQKt9KYwvhGcvRz3FCb5cE1AABEZ4lK3MTlRFpPBq1rVva1/uganpb/ESoekVfd
aq5X9QyGnwIE3LIq+w4LMuGq5G7quPhJEL73xOPFRB4MA9PV49kHvQINE3ylhXXL
jIodOcbgdSQkoGrCLywAM+IwrJkKcHR8dbUuEDmA1SGQVVGX11TKmcxhbeaKBmir
DATwx++OKmQFHrmBq9P4dvjNCbSDQlp5TTxtXRyMw7cIasx5wE35fxc1lfJACsQp
Jm3dMrSSn3PpH5JUzLjYM/AIIChwF6iET/6celsQMDJMEHnGg8MT4zi2XexEuwBW
E6odLNtrjNJwqD5SGT2ILZCGnVY1EavnhKpiGcPpOUI2dDuH2iEp7OENOE+fLiDB
jgSSupbku1oOcA+IyNMZMbctAaWu8FjV6CJKCsb0SUrMWUX/HQMTT6zj0RkjJUAw
meYzTZaU9msGRH6lXv1vNHfCO0acRx7ZxhgkbORuaDD+KpMJhzCccCG9bXRIJQC+
LCa2BBCo4XvRflH5Qusw10vUDyUDxXXbtTDqRmgYDjWRzeT6S8oljE/YLaAo7Rhn
QIgQ6ocaD/kHQ2v5/dt8el8BvWK58n+4gQ10/glzzjZLPH89dZTWQhY4fIGrxrpL
ZqBLjnHWsy8IoJgDnV7W2lHUdh/ieqy2S86ZL9DXYud7E0ZM/WlBIJUAHBi772QZ
vGw9c8ctfOszKkOSK3RMf7XlwBP9uT0iuY5HRduZ5kXpfbp1NCW6b9bA2Vg51s7q
shABCYYbgqGY+Sc7oH8U5WeFl4UM5+KBbGj8+C4jutn2JmfMESGfC6TVioDxXgUz
gbLAOCy6GsJwXOYNqlRnRsHYX/hBkkhjaWcX0BZUYsLSeQCvc7WmzYdrXGWN9zzq
7JlPRNfNbflh26McJ9+q+oG8XzsRsrFnGTGRRzWyZdeLeSXdqXhP05g9mdntxNLw
Lq7krHYv2iRTIBccmkHb18moT/CrBu0w50Ax2QAGWecH74AtmozQdGG7TBm4T8/f
iUYeW0DjLReaFczEvGd/BRl+LkB+1bkonA0qm/ECI5LPtWlXIb1LhqpyG9ef6w3k
E1PmiCZayW1UVnnNxFhS7+4BSbgDdpD13Vnrma/svq9bfKIZxxGI0ZNdZe6vUR1a
uqz1E/0RajwAds5q42V7Jy7232hrWV7Sn88Wiv+J6AwrE5LdQySXW2penkv0IZfC
cbnETg6AiAcIoF641yypySOGM9Y8sbRwIImQ0uzR6Ys+eiSBFJcus7Uu9rZCF4yk
pGE6XkDQ+GIZYLZZjlIrSqY4Se0cueTF36XX9LvWCJfg+d4q/+BY6WJ0VBEZsHTq
ZmuPdNtnWvCOrRhEowbYC7TChla2b8kp7J9i20Q5zTjjjhzDIAvAy4QqiknSi3hw
oFy+9IOgTZ5IPrKN3oIQjhNunaaF21T1QBaaKyHlslMUHFX9LoBeiN8PiRDGPmVg
LxYHOkycrVnmqKqvtJAeUDbUecX/Y01MsmaT1XAfVWVxLaWwDFoRKaufVjzEbenz
Qh8XJdA/md1qXu7wVs7pT68C+wozHei+uXsxKX9zkkiL6H9+sesrYe+J1PtUmaex
Ok/yVSBKaJ66uD+5poQ1J6XqaxdM7fjbLpwuqIlbj0QExrtORn46AhpFCO+Uxgym
5xwRRlni1766NGyUxJRdt7JVlRpE90JR3jKHw6b9zvhm1VNZ3JB/L4qCxhnETKuz
PAphanNXkzyL2lwZZB0KjZicMdisApYmN7MBWocpLIbq0/NFrG21zaMTDsAO1pgc
GWTz9+QJFJp9VmBhtzJ8PJjmwhNmXzuEVAWQxYFU3itnERrDROZDBnvLrLrwOsE1
nJ9Wg3Q4oYh7d4BBnP0/G209oohsvsMj4zvlsnGRctv0Ovp/cFT6KEFdVewqP0jJ
o4KSUiGl1hcXLxGWiBtVp95UuQE0yTqnh35pO2rEf+IUkx7sJtu/rkA9ceJJyKOv
JuxMrDco3R/dYj1VYzV17kpIVAy1N/WWBd8nKYca87yZ9cZTPo8XsQId8od/zich
CCg/ulTir4W19PMHOvMEzjoHj119LQ5oKKEJPcdLLT44dudq403VsBmTushF8JjZ
fIkpbXgHqLtjZZhSGNJ94RoYdcgpWMhHUFRXNnTCe+Ly5hgCSWl2wqC2r76ISz+k
YPLi4jhrB3sMDhn5vwFutFE3zKcH5vbbCSyJi1kMHvg4R5gieDjTJ7evMMG1QaMB
frHm6y316I5IAYWAvfCHAKgi6h0yTPsh1t6L+zGJmObTv0shf64hPmBN9YLBnXxk
Q0hi7rNB/VmLx9DscSTef8S6FztHm60jGZWY1ACD83K8M7DVKDVjzqsPLY/dksc5
NlUx6bpAyTPOcpU0Nem3a4n3uU0hDFl1jMh+y/gPGyd+vQHkbvIMi9WSjrP4nZw8
3vKnfpi/87cyMZXynHuCs+w6F4AttN+Rawlh1IozcQu8VnxkGKa5kuJFfPGRuP/l
JItF7+oHLSV3s8yLj0iZ9KXnjAjuZ2bq6K2PvX01SPoOetu1+omnzZ9p0wfkHaZO
dy8LszEGhLDUCdTGNGNadb+0b/nzTZvLPwYDPb0vgFdfPtmOb3vt6Xa5MDUsMxpC
82S4irEDts+4TtQbwqnhkCtLOM0S95c1dhC6PExxBiotOVUCy5Ny59UTXRBFdbOM
OPd9H5l3pNKAhHYR0ArBkt+aEr7R7W7d/qHjsruKmb0mc/ukPOeqoVTSfw/eNrcA
UgiN4aTldMnhih0bRjxV/GI3EZu2nV9YpEE5Zm07qrvvhz/OAIPvIAvT6QuWgAza
6N27beSKmuN1rWEHsCuHbE7MglZCzqefi4/dOaZoWpJikpmXH6lgy37Hhicu0WSH
dRfVO4fi23OuHW+6c0LR5eKrYM+huqmBaGiQZn0S8nPZdlJxCDJ1zrWuenqwbATR
PpT7OlzfFTtH2yWUSmC9ReP4DXQ/03smaKNjQOYXRIK9MM8LSbmE9e9kbpJ7qGGx
OLDyTgPYfv1FYj4dxNesWQkb1KhiMu3yNo0rK8HoILRCro+2ThZITBMm68nf4iXv
1K6pj2D0FJHdkJ8cNoFv33FLHfQ8upADEJxZJjmxC05Pze5OCQztyfT4SL4rP/nS
APdqffCYDnnfJ4bzerdaLWo3JPHMPtPqKjmiUM1Z9P/4/9xa21F8Tb/meyp7wXuB
HyZhNG2jPqjDkQia/Yww0O2DDSyJpaypdWe1LYcTqF+1eB1f5/0WeWI0VFbm9dH6
Q2oW3MbHM3h6XBjp8x1lwA3O+fdLYp/zjjhHbY3ftdFbh90IGWXymTMO8gI1Lqwi
oGbPnZWnYDzBmqGrEgol6q+lLNXFlGUwhrb3lX86DUQM/Z9+hk4lbM61PTzqFxPY
m86i38iRUdoBrUjBtriT6Vm/Dz8Juj06cwNQHEgII6qjUjIy1kXNzgZ+yePsjs6F
NBqRo650air04t/YgGcWPulaE6IuoRaremc5IhfcskNUDu0F2sPeQ7xiAJr85vFx
vadAFmKIsgUjVBej0Az7CL02mbeN0wOSniURg9jaBvVSauH9d0VtdOILWQwuErGp
xBRTkwOqAC3aLcg0GHMsypGZR9blB8JQe74Z3BQHXhv8trP9/h3YhNDJy+LziTtA
ovB6pKQWp5eKx24tyQyxtU+prjBOLnxd0lrfkxez5PLbOWqqAm4iWGyQDi3FdC1F
chupjjDNzMNB/8E31ZicZ0c7fJC/IuQnxAdlzJZFQW4tmC1D/SpYyQnQ4rDoekJN
CJibQll2tjXqAzhyTpKrk0QD7Ic7LakmIYtuQ2eGamiVTiOu5IG1lSYwG8uGazV5
BCMRblWEUoCfFNT7pk4xD2KvNuunN+QX9DvWMSEyCB5/E9/IVeWv0R2N38DPlwM5
k1GlHBAp2qcuFutQxg+YqKfkAHtIp9susI0n+CQuXuth0rjzvLw+PtL1XgJ/OlZ8
bSrO8J6G8fDe4DxeEs8BJHogZwYEktOHTfcVw17YdRzeCpbey4vQEXErEUtkzLcH
eFmK1G13i5TO3SGjI717W1AjqK4YcMWCfbZryxRB2tgo/BNnNzvsj0aK0zu7wWF+
/BoqnDj//0WILUsGVquD0uWssimV/ehOaMDHKZvZMTNChUczDZ0i6cCudKmcUyP6
bjaIwJmyJ00j7Xu37Q9pOd9muVXi2iKUhmsLC+EJFj68BFDoLpJuv0XhDPabT1jM
KGgnTbltzPcfVFN4RKJTxObnPSdnAcOBPZVWEjcTKXvn+mbNOZOMvCrSgorudfmg
bNMpA/Udti498i3k/AX/v+Rtsm9FrNx9obwSwYkUUODxQkXIaTPJx0ZTfDWIF/0b
euGbMRanJh2j2mA+aH8L/tbbdvk8BrdzRr9ArpWgYd55axqmfzFLzQ/FQ0mNpfhB
lWw+APZXqjkAWDGeDtN5GIR4eYLf3x2LNjFWoDOQVxM1QWK5wrmjN7YGMV2glHoZ
EUATIsvd42riwPYEsLDva0hI/Mv5Mu8O4LVfCQskKHAFzlCuYzdaVDGLARmdb8uZ
joGABzTqPmR/s8lhTA6NgryYf+YaXUHJ/nRn5HvKds8oMjJaSEfm6UPYxfrfUAXP
vEAwK6mHVVa75e8KrV3LbFRPetGrjJksoIl1OIftq9cdVVI8I42xRoQAGYIFEcwf
pCfw3jafkK/2e9WptYqdWwwi9Q3c3+0TvA0+n0Md9op5fCBgFl3/EHf1+UkE8J2/
si9WDkYzxhL4xIeVVWNXieRhYI4V6ofrPd7SQnLBs+StbgIWdmjJIIpcZ3UtSlCg
4brhbH31/l55JS8mvHs5G0t/rUHeplMsiVsU2emilHS53/ptMX30S3OA95CDZDJM
AN81wkhdgAycZ1Fh7HKuqkAoiKHvTciP7D3+B9QqyguQFZRHEh/Fh8iHy24/kjla
9l6xTEZTfRuVrdqBn36nklRLD5pgAvMkqAFbc++DRc5GcGC8o60P708zBPvO76AT
/QhLJ9zZh1hLE+3S99sewjvCnbFPlIACeTZOFq5PwqEexXfVhOeEjh5Uh64zM7HP
Zr9qvx1sjeO3KrRZ5MwlZIfMiIQ5AILPAfvGiuDOXF3yWcbQ35N8PFl63PZBL/n5
WGJwaHwsnuxmc3Pcmql+ZVyoStYmoZbz0vk0QrPJgSF2w3HZsoTCqTh0qWtsHJsa
4pkeQPYKm9wZHeSCsD2mC+zKfyXk4AsQVbuPNEttcVZoNyzNBu2NC/MxhTJxf/MB
2bQGWu7uMzmoLDB2hR+mz+au1mulfzo802eAKdG552ifysISdTStcCVyXGYFQr7d
99x4dnAcZx+JLkkbt3pXppZacZrLFUu9HzB4ChCHzOkK/tib+ymiFjFGYS7i5xeO
aHIZNUJX78Mecut0JFKSUEiKPb5MgGpvjHqSkXXk0dhWpr5pNYe3FnKWq54pY4UE
eW/95Rz4oMz106UaU+laThrRdCkT6lK3bOvYAg350mlq3lE/89nzlSOqlncHBP/q
9zE4t+8icyWPXLcSakloU/+XEVR81Z/w46l1f5ARJKkXGZXYJDw48kb1f7qrMNk/
f+aiRH4CoU+Hj68OLzUoipH8BAoQ/58JAekYh9IE6/zqO/z64cZ+HV1KYKJ1hiAL
r9FzBT4xuhyi7cx6qBG5tibxkzJDDyduKQrlyDjGVB3j66a5WFZX4FTninDbV0og
iY3wTKiI/wKH2wSNCmAeaE8BZoLxwZelnBxXeK4nf8AJHR2z4gmj6jakIUxsAR64
ZOrQFyIoF23b5VXCNCSeP9HHxaOoKwTO6Q30qEhI0kek5595bujq+87YPgdNCF/D
cbID2yT4wZWsRxgo2BeClSpxQHpQ6BgxzV8hPb04besj44JX92ZqHxzueeV5Pn0y
74lssmm1lR/fOaWjBGlxx5qatzVEIqHjSRP+5IdqJhb4+bB3lyJ3Tts/VYcHUmmC
YdnAW/Uzm/mOWKmOY28BOILlzNdkz3ZhFT4kQagQdg9K9hg8NorsDi1k7wNYYEFN
RhvLllbFT6gU3t1qZX6MzdVswS7Tybmi/BV6ums0+M9xy47oQ+EgIcpTZgSlHdj/
/giGAmrKv5XgeHPDFiwJT3iUKmk43/b+tMaPWbKcymeV2GQvSCYm0zlwQn/jbThC
cnNK7FyW+cKr0KA3AhWW+m/aO8nuptvFxILFj5Dq5ZGLpZ4UQaTYhpe4PAUjhAvG
9Jiywph74NkLIuCRzH3mzdf0U4BzD0TCx/dDTjYQmr8/pniH8qWD92TR4+bZMqpF
WmfxD6BwMXXA63traQXlBu7L01bi40GLUG1kPIuDCSED/UM0Pd1SYFNCRT+VHcQ7
pDU7qGe/UgYckDyfwCpK72n0Yo0ab1gZXsQ/v6AleaafXCSBcp/jv1IjXFX/zhdQ
wvXoJfO4CHlS7yvrfJSvPyGVr4Z24yOA3hCJN2J711T7Pz7nQRFYPUVhoO99CTzc
2XUTUfFFSR4FHKSo0GSA+GrXW3M7Vh+QBAXrPvF11BFJjgixtabunHMp7N1B63cG
YyCEUNyc1fIfet6ef9/AWO3ArKnyv5l2H08ZaqUnaQtQu0Ngo1weHLBefwryE6PO
QfkTN1Dp5aHmzWhofUx/s1tqWklrJf6e8MZD5HMppkqsknbc5aAjB9ykpk1UdDQf
S5LNodc3aM1cZu3P/xNFpAaZ3FjgLzXGOlupTaNZzmLqsu/pxmxySL9jMCCe2wiw
tsdnO7Wjpor2BpgO3gYZJEjoFi6Qei5TQUFuaim1ddDPkMkhtrbGhgcuBZmtLNg/
ndqCiq9x5/Es2uBeh9/c4ppF5QJ7y/UCvkb2+ApePIFVPhQYUL4Epj8ZrO2Q+sFt
lj5FYweQpR46vjbHLGPg7NGllzJcS6WgwpfCGmPQCusBbb3Bkv2GtC5m5JKyMZe/
WwKYTdubk/yL8S3N3IVpFAHu6v65rYatK10gDOQ4aXaecJkAWbuLgHovnQDPkAIl
CQa0v/Kwb7HlhqUQEh1B7/y6mC+yAHophGAyFxqT/gaCYo2++FW+IaZ2cTVkFAUx
lWGeOC174DoSvRWQNeTtAp2RWjNiz4+lS98ceDJv9Hp1Zghs6QwnUc4+ewesdqxA
GLzuureXpDBZPqzNPtvRhUcjjme9eL46/yarQLEdObXXN2PvAv5uM471KtN3kOx0
0JxssoP/8UyFl0YJUge3Bb/QNyUH5T83SgNZfL30VpQxkNYm+WSSwIsSvoqW4XiB
Y3fUatvvtGBXkk4cF7srbtXc1jgbglS0kkrpWOw6rC3wVRHF7L5s4lGxMvXEJohw
hjMuA2bQOP4duVGhW/K498Ie29Jzu0h5vKsFVlNDVf+7aRgRtQzKbZOF3gNvtT52
yAZ9jCgNeTkP3B7crraOsrpnscwECtcY6S4vE4f9ZuJEx2nshU73iCLwvteZ+Hji
zn1WYOtHXFuy0+AyxAjvZ0XycO6v7R6pAb2R5IwCbiKI/4Ruz3CZY6oIjjAvje6h
W7Cle9cQzt7LFlloRAZqxa9diJHvlF0AJC+7hC9VoPJqGa8PcpNOSLEjEPIuSGDg
9vjCzegFvwicKlXqbMZaQuXKgYXxvHfYTime/d7Jh8g78CCR4NZ+CcdzNy43LM1s
X6JsxhCdkYpY5X1H381U5u6dEBdgXpCDi/R6q0TlnQEMtZ7vBkJzeQPgnr9BsrfY
dvAuknFGvcIfs4/7W7P5Vm1ZtGuzXb+OR4EKj9vdrkQhy9WJ2JGRdwAmt6YRmZVw
+xE+Hw2fm6BQFrOO+0A4QI00Zt0u0+wZUk7VNvcObEpPkR1/nKCC7KBoQ5kvUtmk
UjZk0f7SJXdjaXnjT4QZ/M+1H0/x7X5kXZxzuQTTzt5aSZhbxVAP/DXeCvxN3ZZW
SRsTbfOh3s2R2EP4OeRz3Ja6Yfp97TVm/5gZpOFTJGXm9KePCmdDCk5wVcCh1LVV
UzO6+AH6LMdGGlf9QsKZ7ck+GuWHuCbnB4omQM9Jv6WFBchi+2aisZXNIdokgaNx
pJ15J9KKZ3hjD5Im2M1yVScSlZ1SSu+PWSG6pRUhoH5RX4Hn2li/pqhF70nfZqB6
Nn5oVl+SbWHyrIOap52tXY9+VJrdhd1bxorzAvkinQcxZEAbfBtLyYLFAZOE9ArM
b2FSKmQIjjAQLiSQFqUKl5vEMsCLzlkwVJAN2BHJUZHlQDaJzee934mmdQstVRX4
AkTPbF7ZRYD1ne3c79WbJuSaETstjjsQuc7IZw17XOckvXDQ9VTlE9S/i0auA+D9
yfTOS1iGAQ8Npi4027lNtge4K2WE66/c0LxnAnwOKDsQdiMAEOkJzwgXVTCEBDko
+UnnUy3u7ke17ZYjVoELB6G3sgoCVlVstMAy+iMmKkzxIGNJ965VRx2UQ5cDbUxj
OCybZA9aM2MxmSBtYOdkSb8ZZc8e8XGlKFyhQqNDY19asSAkXjUq3XSA6jC43b1O
IH/1Z70qxVGrFY2G6JkFfooU46QYMH/LXzBg/NhYf3TcTwbIkgI/JAa1SarwMI7x
1YaAsqNiA/fYCAW8u20Q4vlMkcJqLAyTbKf92F7WjtxmPXWUqboyt6Z7ElmhPg8p
McGFXXHg2YJ2e8v2PwGct88ydp2Tcm8RTQakMq3eSX4FXPnxAtrI0hXRfny+mRhh
s4UIjeZKwDfqJWaRwVW5YZPndyYs0clGCefuu4uBDuSi+wiSO4AeGt4+sfRIFyjh
8AUDXirw4EZMVgbOMPLT1h1m/alJWVz25cwevzaPZ6uG3C/IjuxuudAc9LuH5fN+
vE7wy9M21EbbxKN0XiNEOtIPulagevQOxIxkBxvZDnGHZuobIuf23m1BtGogjP7G
/dSkqHKOG6Hl9vzKUHOU1rjGaf7RkX0rjR6B4XfOzeAHsh4EAagqZ+vMob45vbLd
LGzksCQHDbX57l9ZgN4FOt/g9dfA3L00a3h6EuDTjN+aHjrT+lLhxPix1Ib6A5vy
ax8TtHzUfp0Y93m6nlopx6MaRTNg+W52po2Ml/cqleDDXv4Adia6vgcy7z8WglJn
BzsBZMFsBcZ1TJICLj3PL/uBqxF+yyy6PWlLmaVReCERpRPAjLVa+nVBfQk64VaD
BVhA26Eb2El+FD8J+2m0JrQPLGGtH50m13V5CzvhzGfmSyJJNBbIxoNY2nv2lb/F
Q9fV1rt+6qqhPKUn5dI1jQmnMlqFR56U9ADVQwjNtrFL7QbJLF178ewfJcFkGy7D
fsFyAhrKBCoezZBbHvOGgrxCg7pI4Si0mudvmJkrlS1CFGXmAbQkj+JETlJlLxCr
5+0dNtEcDD/zBzgul8zNb0noKJdvHQXZz8oVQ3UIp3IoILnXBq13rKM9MqsA/m/r
4bG/6vbsDfS8SgjK5GqbUlwrwai0aCoSt4qVWSr/LznGq824pO9VeSdFbxJfyvNQ
3XNGnOmlLUXiumh6U3HKxkXCeAjhGleGP/3v2wk2DK+JCddFsCZEhAGRvLDxNsun
sqnSMOIROnUHxSvHESF7wOWYUYZpV67X4eRwNp6tihHa5SW3Sa9qt1EjqLW1RYJK
UQBio0YA5vAHA40RlaYm5xwn52ES/m0a7wFNsd/ClX9XbZxvKU6zqrVNmeXsRyFP
67d23Wlr67O+swol3p0zec4otf6LC9khblhFqKxvEUqiZcC7VBCdFyROKdqsvm1U
6BYgUtXhy7kbeiatCKCrlSpXwrcukNGhpHZQ34pSQkIV+tiVva0lbp7QbIQJP9VE
vOqubxbXfTssQGp/1gbY5nxmRZBXfdPJaAjy6vJIjgcmfOpEjFhVrjDCA5DLYiwP
2b9p4vAP2kx/mgziAYUhiNRysEPI6Uy690Px40uJ8Y6g9djX6DJ9mB1RWkPfHOPD
WodBsw09LJ0Yvsj4VuJsLLqCiQyvIYsyOKraJjQ/2QAKW0xVU8Ic4vGQ0tBJIYOo
dnMBfxKAGH3WT7tU/1lknIWeKZEsL2WJzkZqFv84HzT1qzKpZyelfJojTzZoStV6
M9uF8zKJb1cHm4+xcpIqbG1+jYBayhUZJ+H9a//pLjilmZgkSPf3IRN6K0NYyr+i
Bym+0KHiygr1AlRhtzDUfQHoiDNUyG3dL65/yDzK5EPWlA9iZKoNRleZHFYFULEq
uOOS2cx5TeEyiUIHTd9Fds3chNv7xn10xbhblnMnyklXK953h9dyduIY7wIWoYd3
h4qlsEPS0NHU0ZUCGx6+c1VXkpAMWoQtfrCPIdDB5YQlxyENG875YsOG27l9PA65
9IZvQ0QfqfkHx/IrhBQYKHLj6rk7y6rh28DD8q7gZ3WkS5q+ql+QtXAVL+MA82A6
N3eHwniuL8/5ioJu8/F2fs+OkC/XUDW9YDOseLnYur1TpVV4R43IQvKIhBgaCCKq
5EkvXOyUkkkgF4q8gxx+YHmhQ/G0yp1bfzM4qr8zRz5obUEjF58x/qA9ZJhR7Z16
xF9BzRBY4g6VMPjOTEHdH6tRpGlJZQeMjXF4W7SFQPFA+iumvRJp53K4ot/awI88
UqC6shEBU0BfJRR5QD6uEJoADR+JGKVnmq7MavYPn/ZNLcDCy3XBVvk6c8DHhaDp
g7pRYuVVMgq3pvLbUxoPvUpMpB6FcsqxMHUngGKNK1vOv52lSgg1k7XHtUfzjxLW
KUa1dFUldpAwdpuu9dDHwkYUnWw+MZDXl9hqDlDW+fC1HZ3gfstIhn3/p7Vb4y86
YYSwP4Jy08A+fZtf5DLRoM2QqFdpcEyBiWJR5tV8SFBVQyDR55k7mP2o558Ymehf
d3yZP1sQWhkBk9FMVF4GhfXwwYreLyxh2LkeyuEEEPz6vCA6JptfgdiFxaTAB/QQ
jtr3sZhG/zbC7GgRDjPK0A2FDoNSeRG+F9IjoHOU/iMXZMDQDXEVmtu6oUMuHX+z
IiwZ59Uv3cF+/Y2UvqelNS/1OdFUyduBnldgU/XvmJ+Vj6eqHkYVa5uTjVc7diBu
5hBPppVYjBZsazIoC1Aaz8xcLKvTz3FcXuh3nHyksO9cVhpUCVi/9JhjzegfHkt5
KGVUPK5Au0609uV8sD3l49/m4OWgBr07X27G8OOgx5NdOsYl2Kt/dp1pwGqjvHF6
rv90/Bj9+/UyZtn/nVXR6jJPC3BKxuB1F3Vgwzv2vp4WjqHx2IOnMibC5ctMFxkd
DqgAEp6AqA2tMJJkGp8cUGgy2iQkTTvei2cW4rRftuz6FAQ/vK9EG8tgXv4gjU3F
Kk2UXqbIlNwZW4BMHG0ulgJXKJQaN9hRqp7lpYe7ZClXcuPstN93QIKtc8mFWwoJ
DlXbyBcdNIzIxoK/WS3P3luka+LWiEaPp8T4hlDCr82ToOwpBzPLyg+5Vkgtz3Q3
Y87CAlrSkB/r5VqiBP392UF9KKeybHCnw65NoX21KKCeT3ZKfe8O2VGqFG1g53Hh
dYiVUCbt82Lz2BtA/xdNysO1PPHBYeV339dCYm3nzk8a150gen3/Sw8Z+k8aYoPP
KOLQ2YqE3Qwsbu4XWDf7f5Dhd5zT4ax1Od5E5H/bhnDm0+0RlLk3vTKPHhD4rYQp
RMGO5IkS2CwdP3Aoq+KTle4uLCDiqiQzx7e3c3a3OiNZLL1MYzzL9RLxcnfIPbnJ
Ft3OcJ8f8MsCESxrpwFNQbxs2sABvfMCgpmEZEVU6yiOAULfLbaTYPvNi1f2cJwz
74ZxuKNldL4XOG6bEzbWNd/YEO0JDdeXx7FP/zOwJIpFqfSBtEZzXC2F+vW5Cgl8
qv8Yk4BAbNoUAqWC5Hj7cG1jE1FoptOuhA7Q+O0S9uIKLfWANrgySy19yv8c6U9R
fDureUtLLSSu0puoLYNlvNDtVhaQWn/hOrNoMsHdYItB6cD2iKBetFPWKdH+YgCd
KRn395pl+fAxZ9Zn0IeV6OSuHJI4KIyNwAo78HlWkehA7llaZJQYraq2g1G+tiKk
nIwfK9Z5ENSEmlNtxWSHJfgY6/ItRGI5UyDZ8/7wARRUokaSH4hBSg++ZGJwu8DP
bjQOkWpPJJ/OV6oWWFAczkMTJX3tNgpi3I1H0W9NfJWyN17EwYS1g+nJdqJ9Hxpo
8jCB0PR7r3GqW2Ll/3Vpm/3s5ZeAtLuWsHKrIGL8LfHQMQnPiIPZ1xzIyQqnpPt6
ineo5bO0QCeo0ktwGTLNVz12b1iOByU2EHiQTNbdvx6+SksQWpMFnFoV0D3ZATAO
884bGpL1VK67AosJMAn1seUUaVJZ9ltduwL72yfIOdALhYBx/boViudc88dJaLO7
DZeg381HdlJEMUlfFQg4FZfW7RkmyQIErib/6or7ZJbt0GvZ3bQw1Rh1BSxLvQHh
hqlHkyGwj6a6Dud8/QanjNbH4ZN7zr4amOQ9Oso75w5FSAihGI5O6k96HFCDZSYp
RLrMLfkmNL012nFXvTJy2S9RC5dzHHiXkvZjh9Ws1ylOzRqACiBwruQA6L4mQEFN
MAeDSMljTXKAfhPTux6qN9Bl3PwJjRyDlPvgJgyqANzBndlTO4CMMnHNlHUqaS2H
1TMBAWaXhx/QAwXSCv/woGTarycZWuRC2GSndOpzQj+mZjrZgLvQvw4Jf0heNPkr
3yacShEbxd5xDWHt0bwGCFxB5g3y4QjhanVrNNbWame1+uwooT305ygL4yB67LTn
eNC8smsVxpSKUxpSodLMS7625abann30anQtoZVNqT/5oXQ61v5QWcNQ6WrwGLUR
tLBWatbtNeGMEq+StZEGJqg5Alj0LJKDhyO+ogUvC3GOTPjh8xTAa05c8uY8108Q
q3Fhfd3IA0OXLA14dr72o6e81cRVtb744M6w2F1TFqqfWCV2YPre7WP3FHMdHbQX
9HZsePyRKXUCXAMOu50qXt64wYGDEE463Mxsktpp0sObecvtSF/FcyZnI/9wWptk
upohQOGelteHCGdtB9Ik5Onh+S2Mpojr4DgtQ6nX7f3ZZ9zEtVO3uquJYi7YzTS8
CNuZyhSsKCHdhJy8oefBEQf/av5HmawoiZXPTFMTfH6KNiTJb+APNiQcuGg7obpE
XHzvmc8xjgYV4hEyLP3DeBkFPB9VRtErGjoHBUtzZ7gPhrB/EcvHL7ti9gPFj0P3
2eIorj3wG/oKVPJ0QDMEq0QekzVWmfgUPd7WCmYhVfDM9fTinWuCrv6Rx5+WfF5L
MywVnpJGk8CimLnsncnZufKMckAPrpy9iIfLe0IOZu12+y0SmIWa/CIlMR7EHfOT
7w9mCk+L6pI1/pvWV18Y/mTt3P0fVTKY6brZ8faVyHWwkS+CC2JPjkDnWNyFbkkZ
6YlaCTvJBWe7+sQW6VVQd++x98hWP5Uxlc6fLTMCmcOt0tpnA6ZGogydP27G6EjV
R5QgBgSfn6A4ogVGAtOiDJe13CR7B/VJ9bIcqbubs7JY1y56bQt1gCA//zcY5Q6H
vlKKrbLwTyWeGrHh1CVR7857wXuhE0JK12RO6dJyrb3RdRJ95LBUqb9Laj7aEIh+
R1I0f5eZjxk/SKBu5f6+oSopqmLZEiwhocAofeAP9zj1Wd950Cfbf9RjKmHiobd/
/lYgl4QbmYQbBVy+VGECWSkb8YOLUKiZz/8BdgDIjsUdaBh4FIIcco/HhrftOLQT
Yot3YUfQO3AIOlA3JtE6FDk8Sb96mfFONRBIXsfIZiMh5PkrX1JGpmBs3fagKPm/
hhvIObTRruVxMyvR3FFYkhev/gAEAaUNB9FYmqlJAQQQHV0w8Ke1V7jGskbw2gyN
sBtCJyWFS/L7cu0vpK1069verCN0NFpIB4cKk0lKIBZH83b4tMpmyJ5e4dapwirr
hR0gIrTb582su9i29ampdSoNGSumMY5oIbTywBBVWc8pS24HJPI2Vg5Nh+O9bvIK
R8dVhe5U5P58qjOTAq3GQp1PUoiZEDvK5Mym75XnjqxZdtUUUaT3yCDdPrvTNBW0
JvFnLY1jmI2/ImgnNb+E7zVkjWa6ziFmwhL9AMwUcQzmGhrw9hL8yDdxwEMsKnOA
Flvk/Jolakb3N/nBcDz2YlEqU3qEitu0wUQcBcdyQ67YGjLGqJB58OEc79ZzYMjn
9tTOv5W1/xtJ2upgsfLNUnJ9dvoMT4LdFcJBrk4HvYyCmsJCsfhebQzdo7bi9CG7
3stpR7LFWDeWWHyrYxD5JfR7UeGi2PFE2LSxSofEhOy1cHVa0op+bQPs8uhsgp0o
s2YrTiA0cD+Ib0ieqYPBcDdoxbek9QbdtA3VUKzkH/3nS0pfXbV7ksQ94OFUgDc5
7KV5XcrwNUgqii6gf7unJOADzry5EtfZ8Bo8IQeGCaUgzGwmhw1zISC6aiUWpbwN
OwfZZZ6XHr5jTtjew1X6/WVQmRPOwkzcbSMb+iWoe0H3HRZT/Zrkxo38JqsaId2y
XniyIHdHN1HNpLUCkIdPxIOjFhv95EOqaapNakw7v7TjXj1OEgp0cBGiEDN1aqjJ
dmj2hZloko648ZSdMLyeAhrNw+M1BCgpHXifv2pbIgMTtWjXQ4WuAE2gRO1PQzjP
7KChYECJVDhU7w9mcq2O4sZqU9MqlLlnveNUxzM0vu0BWpSF7pM5fI8MITGFD1oy
61x2Ynykpc4SDFixiunVmkzeieIXXz5V+nL9HrWv2o0JldunqwTCjoiMnT2m8OC8
22bBYhSD8pqELn1FG1G7nLbMi484/Mc8SI/E7Nm3v5fgGYzHtjxTzKIH/c1xLQf5
4N5vj8IVn6fKuF3wky3PTbfn4Akg9muFZNkvV130DqggsKcLbxz9IXh3qNnmS23Y
ywc/EBrU+EuasHqZQNbj3QlQGxRbCual2nA+BJkC/462yINUBgwDhpzLv6HuyCv+
EmlxTcGmwaikVV/AzReUmOveMQhgAmU6Y9cNnJ2svbzJ3M6DDLjas/ZA0cNdrAWU
I/pVbKjISvAsHWlou+pFaeyYXEj3+mK6B/O0y5d0WetjyNxHymPUZl+hfW80laoi
8X7VzdsmhzDCsDk/RHgHsyj4j1oEcLZw9CdffkO+HAH3JN7d7I/bHwUFHmiBvRix
lhSwRZjlS4KppSGznvnw4Iahqm4C5DZzjt4j4rfqSllCh3mstoNIdsXqfGHa78GX
n9STD+ZNNHkVeDyg6aTTBaT8uqagbJ7tq2mHiZgmA5j+7iWiL2I2Tng9eKjS0yBr
r5QmwfpWR83cuNClcleolFO7SYEIALtehZaW+tnqVVQfQOxRSubtlY92E/cjoKsU
qhD9JykUUn1in35Xr1ayfwbiXNN6CI5/rlpxdtQL9c9GIyVJxGgHZZxMP2Zm1dLJ
NYNSwKnay2HTLJ5PsYlV4TE+nvPhS3f2GdD3X23IKFnZMDY9Yk4nuLW7cfcIwqtB
L2k6fQ5TyAtNPBqsycb0M57Ue5hJpk8PCb9DdfQ1RAWylLnLyTuPGaOIJWlUmCxC
NIpkJh7NyRSQFtIgATogIfEHP1b5+FM+imVmLlNP58mJMXol6jGBdcJC2cJFEDuj
4MR9OM9wH2nJ8pHbRlBj1iaHjes2aC7H3b/0+HZsMf/FwkAPTg5RE/thVFWXNnG+
/fXzknCvUr+Rmxpk0ngcbEkXY3mHLsX8nHITork+w0/VgIOkiAeW+gu+j8zZYxAU
lGZ+fCGe9oQZBwrIWRTyvykeT458aiNL0cXdmahqMVzOGdDEEU9MkavGhYd2vizl
1PZqFHQnHb+LAQlJUeZ7rwHU9UCIjx6uaDTApWNKDT0We1zyxPzpOqYvo1dVGWKn
3CpqikWPblHQc3eHfJK9DQqD6eeBcdZIUh7ODx5/cGO2iRxqfemB4qr51aWok9TV
85W14gyh/ve1N8DeNj2Z3qOBCVpjiGsLJq3dGiceNIkUIAAzvYylompWhenuVl5G
K/aBHqkq9r/bZFEBiHehjWRKt3Z0BsJE2J6Y3ZRktEag1HJFNAF+NVnhsA6URXS3
k+7mr+TfB4jOCjNSdEbwW9nY++1h83sMcsXkHN3LuqFfVQaUyapYcIsrq8qQ36mc
KRSJByQn6bITK2TGLjpJLJChEQpVT6l7+v/qssqiar1Q3z2bGRNi6z2J3KRZc/m0
w3h1lJI7wltTPw4I0QdIJQE1fNKik8hGlLuCeUNJe8gT8wMdHW3gz4QcDNLVBhE3
mtRPQFJK2EXATwUCzXrTSmMSHOSMnp+VCJ4WR8WjXbnPGj3ry2j12vzYPEoOB/TU
PopuU0iuQphFyEnRbME45nFM6oTm5KVJABkR6ZA/iJ+FCxzl/Eg1Km1Fyr1FSC8v
8pbEQgKxfkUuRcNuMlZyzZ7XKNs6WlgryrRQ1nZFfuZEgK0FH5dlNmZUs1wNz6Tx
re96w3tfa0zEMfF1KEUeZwmLVCyF5Cdkr/Vz1+m+s9dgT76f5W2PfBKfh0ORX3gI
GhdtEms/7elnpBGR5+Z6F6Xi+HbcZi9MFMmFqxnydbYw6+MdTsAYHSuIYYSFqBIz
74zNcKtNKt8S80SHygcwipyG/0W2Nlzc5jMKj2gxPcLgfyydvRILrX3zZV4Fo+os
j7XtmT0Mw5RCB2jYTz9Jbz2Q7pKm39C9APih7EbmNgOakOUiDcHOVPawGrQUQePh
YCZwf6f7EbmXySeGUKzIgobKDFsGI/PPw4qAUx8cKKMbz/adTZGVVyFpkbZJLzuI
3JjyaA92yVZTU5JHqr9weU6BBgR68fbnmLuxoKot03FpoWDBZ7Yu0a/dRcxmqsvM
0em4rn0cTPr+7qCJ32lV+TKfdVFZhaD8uNAc4PsVEVgMSLIhqzjxep/8Ch0KatRD
D4zLivl0e9EnzC5m4x+u0IsTY2Biy3Oqi1GiErmJP3bJAZACS7UjoMZN13WrubYj
FQACAvGlGGhQfU17FZAcTz7APS6sE50SJKhhGq8wpHpseDVqJiKWjnrUV6RYKsfw
x3PfrlYRIea+Eq0grO0EkV3wNTRny2v9UEwO4qD6AX3hhFeHFRrkg/wSzhKBhQH3
F8r3iOVcJVVgVYTSAXRueS+bXjfrmp97pjVrocLdj72orxC8ibIJobZZRS/MMn2j
Iw93nru5w32hfDn9M9iWN/Yza6XGM0U9FQMdlF+3LFE/himO81d1ZeEeBtXx0UaH
QtjkdFp5FKOMAd4g+7gFttCCsjMWRWbMjUHjf05FszV4Gczc+aJuQ638Q0B9wwyw
kUtll1erknsQjLMieG1hY5zZGOZ/dUQefoIVsIp+UYaqrYhfrLXKkWxlnedbSv05
ZA0GCwp/L/gBln3iyvdfn94NV5J3dXeXYL3dDgRpWhhXcU9NWUMfydBR2xJ74wDY
wFOjDZrtKASp8GH/fXEOZZdk2vSVkhdOhKLWDZnhTpYrskL89vuqFkX/v3/OcPzo
0T952IRCO6j9jY/iYoJU0BeNg6lopdeuKl1eDjf8MsGFoilUl8BWAZ5KIDhFZ/gP
7Vh8Ru4s/OZv4753gvoT4SfFhWCwsoQF9wcY6G1lgxi7ALbNH7NXOZfiOXXrnZXk
F2QU7UWabYlq8lBFE9Ear0Q7cZ0xWhm8HcpKpIGBU1zpT+LfpD9aQczE1KBgGfFX
ufeqlKQlbNVu6IlXSpHnGMA/TzXcabuBGCAjFdZI+57AgqnyVI9qz43xKxABJJ31
itdTN1rM7OvZWJyObi68yWLdbS5Gk1z+JgkHC6fsTNhKFtQNjC/DLnRmmLBTwALa
l/ivm0FV1LfOJQYknT6Ko+jKVd6j7xZJ7lJOPNlDxQ2mEEaq9QpN6wqvX5KbjTMT
gD90cgRKRkt/yEqGz91d18ODPxSDF3pvClcgLMyDevC3enVquaFMjminmGCCUwGu
YHisZKCIBh+kOyPkkjKGCGIa95jNIoT9KA5R6PyGTRoZ1H6DhN+cVympaN77pe6F
gnwYMCOvx3RqxLStXVQ97D/2wR08oB5CND+eemcAZuTxpYo8G8UkGpDxeUh4Gqq5
brtCvTpOr/bk68YXazW+Nl43vsyup5QmXKZ+/Vf+jrdw5b1yArhIgV8p8iU7iPEY
nCk4fUF5VSI6lGuKeBoAGuf3ZFqDbXQJhaGgvdI2aeuwNxFQ52oNub/BBUk3vPBy
iGvWYCnJ6XrBsRWhKtQ/PkXptzzpvqRId87vEBo2tlsWevJb1+NqqC53g+wapRwz
PmKZ0KPh8FbCzyNYeZ8cXjRdYzuIHCBi+UUyeOPMFPOj6HxuVkntmNgAM/DD1E7B
w+V3jxWeFZI5HA/vjW05twoisNrGtIhBWPvzhonDw/P44py1x8EkL2JmKcPxXrJi
tY11t4EHYIwjBKi5aLbopFYes6quJVxmNiWq40uIlGN8LPLnD6yPNVkCk0enbaM2
qAStbF7yVq1mM4hF1GTiek6rCkkbGwuSLqfXW4irAnJnT/FDBXCC+wFlPZA9IhnH
hCM1uKIQ4GSHon+e0qrsnv10+l6nnkJnmUVDqBUy1VOhTT4cfx8YVG3j6DxT5fFn
+7gE2KLU8h/o9807gX3oBAwyIYwQWzRVR1Qc1hredbKrvKieUovkN6siwUS7W7sG
bpn2mJcUrh/+vDJiEdzC/xbFk7RMzpy7g7qhw4deQjO1U3K5iTHN/79JJfPzrY7/
kvLuKJkE3fQdGW7OZSjHmC64FeU5+dnuOWLkvy1ZewuZMEaxaOrBHf3kv+qLrrIp
pLOYFcdQzshVTE7bChNJrOexdi78/2Uy99LUev+QAtvOV0UW5RFsnDUCA9AdyyNx
YCo6huSKd+8DgKMJ4Eer8sUB8+cBZ9yf2ssUfTm+odL6PWips51DdhSMSMfHRtH3
ceFCzTo95i4L4iY/yHnPvy4aCtYDTjAdFg4D7sPYCSU/xJyR5RnC7AorKZY9Oscw
OdGAwL4pxHGTonX2wwwFwA==
`protect end_protected
