-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
UY+hPmij6xH+ZFQWOArIpZ8LLf0nT0j9/L1WNuJxbYkFZ6koch+KvcGXRDkmfKz4nU72FlMZ0zjE
+ONZDsC0GljQF45YzAjt+5php39dvJazDS7ZN3fl7A1m9cOy+FLlPWSg7dP2094vGIw3ULmD6u4l
YFR78R3mmhyiVRqpA4J7vQaBz6uXNVE0svru8hRQWusuGeGphRmnNxnjntv2oueU5ET2Ysf1r9/i
NnjnPdhFHRZidG9X5x4OrurB+rWxKerWpiWeEAUaDtoJxleduyEaaDgjQPjiCfAd3hKd58PFfEO+
H+iA0pWjrJY8gINcC4XSJ62ckloHAkjpDYRazQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 22640)
`protect data_block
kOR0M2xKFDcjDIxpgFDW77/WiRUGMO2I6dtiyaxDwJ6ikJ0P8YxbZypDSFdbV2tXAJ0bKQF8oFqJ
m0qOjWkwNZoloxd4qnWMcvHfX2Z5DWsoo4SdWJOCuOy5W88fPkgXg027A5SxPopF1TLrz+avvGc3
2vgvTwTZ/WBpSYlmguGMZTn+ewHe6p9bs6n33tsBjHBNnp7D7nazhvd4Il2ALbW8Jfjb7wpjwwmd
Lxha4Ko0waogjAtWb9AR40o97C3qYn1AqNZIC7bhEdj/HYiKz9GeXvgAoUO0JSeJEEASOKOA0YZU
y/56W5K9r2TuEzkK35h3d0AtTABC+1hl4dWn86imD3a9y8huR+vN1qhJ6OoZBze3Lvowm7LLwKfR
659VHEYOOxToAohTC4vZOPYkYf7un6YiTgpXgKJX2ddlLdW94GY6wvEevQRKx2Kmwk711mN+m7SY
cL8uGB8qV/psEeDxAZkvvphFyVqYyAHNOCyVWjDJJBlD8QWp1pfhEE5wDWSRPwl6WNSttsW4TaZJ
GSlTwuk1p4bLsyXUa3xIGRH6QUoYkUoxzIUfoQEycilK7wGY+78JkQ6a05bhgetcYDyUJNkTJq1i
HT3I1sV2lW8vyM1MfVxGsIx6RGmP0f4+x6gQwcMA3lgtzumFP5pvr2fPgB0G05hAeI476D4YP0Ad
g3UbEiewQQQZLie+p7vQ6+42/bu2Oaz8+9VfcQ8Tb3AvSNQ/8WC9oDAhV1EbHdvvdSxnKadj5b9B
eIQeIBFHf8ynBy5Nm8rbIV43hZ/lWovE6ir4Qj/H1ckAgWD+UwIP/TAxNCks4Gno9V34YO+83RGH
MmYT9jW4YhmY5UqrXFDqwiGqMjexY3pt/3zseRZiA1fG+T1mAlrZp2UrI0TIE0t8oL6gtk/JcIua
cN4H6S3OYRytpJYaYwh+6WS0sO4B4rgTzORpBzKGham29eVaQ+OazK48bajbZkDj+70MtBcAt75f
7AQ1jLN/kg647dt2w6CCObVVgFza+aGdJ71Hi/p43PfQRYDq2BDwE+QNEdgAj02LGoNIVqh4DS6v
KDkLVgJX9ttFN436AmoQ2owoMfylMpzwRK6MeUc6kfK1RaZrnj30/IeBxmgRpHlNrd/hVzMfllJN
kQtkx7vNuS8ZTW6jcreAZZS3fETlFJrtwQUo//rSnNOYXmGNZly7SzMaAalyPXeGoQ+CMCsqD2SP
hqgSFQDBB3/ucSiH1ilXb/xhi6iVIbmOtBaZgSK9BTnskYsaHNpnpi+dU4SkLTIXTWwMz5BIAPUx
TiYyJpVYXRhLAuv+XmSDzZSsMmz/FbxuwQirvxP/YO7jgGXteGzvMjrZtX2Xu2xvuCezj4YtMpJW
6nDWX5aXks1lPbaAqdwFs3wSy7jvP1y1K8TRUB2sWLFQdgbTV5Yvs34mmoZRGVgahcq5PZaXfVFh
Jq7F8yzLyuESFMqdgBX35KGgj3+7E0CPbDfSgNX3chiriNDN90ueb2Yv7gQDlXnYqIZS6gwQOT26
mFXU4UQLQT8yHWk57x1gSfF8E3Gy7QSZZaF6YCQxvfopuSpmNhZSgRR41lLHtfoWLB+DaJLaD6EZ
mX6tmaf5+tcI3YWTYbhWiexZ1GQFWxBCmx9q2TvUsxC7kidw/hUmos/xcY1XTov6wyIYv2iJZk5x
gbDn/tcKTLwGaLBvcDjhuLks24fOsp53GJ8sdtIB3YHwLV/dwT2qHGxriClCk6FuUZIPMsJTE5fP
nqBnqxrAnz2f+s73EUDE2okz5wCwmOkkbZJYWUJIJ7xn5V3kYXjAVQZerxT2bMcLs360wW+IIKBm
ycHNimDCoL9Lo9clyxWb9IjMNaf7PC2LwyCKpi3k+svrPgNvXGwoRoJFaPx/MK5u3hBcj1iHy5W5
nON0kXZPE5njKHpK1XSrrbUOxJGEuhBluf0S8VqDfKi/H+zcw92u3UGxivkIuEzd4sJqyMYT+U10
JRbEcXi5ME0DrmVcvRuEJy79jOYj2WN2/Oc57CuoeaUk/v/8z1y0kmPGAOpUmbfs84eujWHHNwdC
GymiirKGy0QdIORwUTxBDpqtkoASOBpH+ZrMJWg+NDqsRz9K4YthWmIEyBKeIi/dPjR/bX7OsRC7
MF6A3Rx+p5toKNFwK67CD82QOvteaufWzsiF/2wgjpeP4+wDc38Dh0sH4r39OBsx9DdvnLRsYPWB
s40/zK14ZhXVtvpUPOnHBHO7n4DGUbxSr2Auu7KspWG91M5IMLcIRIcSR+daszTsTqWr+rZu3LGk
P1UGK9MZ9w08AmCNxS+QHJEL+kUCMAqrrwYFyBqOxlisJRxisUrPC2svv8wypzcDF6rTg8uIx6/L
CjrsKsaoaz6GMEY1YqnaXLO8DBhN2MyvoJ8xIczU0vcpioEaucmVeDpdb3TtyzJ0KYA/j2+fnUOl
70YvTAA9yTo+ohDQWyuWdXCd9xAZ0Jr2YxgFnRQv6SWxHt0MWKyopCVClyQJx79q6Om5HJSOkMq9
xaO3VrPStKz6c4Jj5vLnavlnR/oANNNY/M4C9cN31dj7fwjwwLaNfgyo4en+/ihOUiHJWrorFGaN
DA+9fdtVu1f8IxqLZoqRpFmca4x1de5ManVEG7sMYGQ+fFkIwbnG8BbMbouBgFz5JJL1cH1uyS1H
TxEysgNL8WEYFU3VuOgcbuKNxkFnkFij25Gl1IZnzbRz4W5jlu4qw3aNOXd+/t9jUnhZ3L9h/zht
+r8YJLVLOAPVo+cv8I0IPds73PWqyyO5tiUGVJehap2CvDXs+aH4BobPTOtOs0U8867i0I/xsuTC
zbInx3J6qkvT2f90rI9lYtzho7K74LvZAuL8N4tuSdT5cIFj5cFPNueex6d5G9ZMY2YqJ/fTNiE4
I7Y+AxVt4R2zkS8Rmv3F1tOcztprrxlFVrCq9JippABJbjhojmLfM4zpzvje1CPPtmoJGck4eFp8
ZugLqVX/wDGj3aqkyimyUo8i/Mlcvrnfgw6cXxln+GTuucVs5I+Hv48fd/CMOdZ0/oH09XfC2jmb
L/OqLdaiXuZDanfNi9BrM/wwfnLEmnH8+PdXfOdV+KUTILhREh07tJxo7w/340ITH5g8LXPv225m
WBcwarrLT9CXSv1CYwkYbCg+G9FLqWY6twLYSjGwtwJjAKcTub76iFZrys4Ki35Q161yVviSZvNG
Z5Heulj3Hy/8ttSIBRBQk95+YeHvZXyXWLon1q+9Li96e7eNXwCfaq4W9z2InMs5qyHCZTEv5cNu
e0fWZZD2HNHfP4ANwJGR6MK7evq7mb3IWUJLgTaLbHjZnxSp0aVYwCfP6We+ig0UNzaT6n+3CF7I
E5AS/iNii/AginMlRm9vn67d6cX5brKQckTpqaVb/hAuJEkAwMGRzD4nFOoSOjWWYBRREmQu/D/7
4R87j1m+JrtmT5UisWnmt3/AtRUpS5nEFRcV22LCtpD3fJ+z91QVFmxBwP/GUBcLtPs2qfkxN3i5
1ZSjfknnVCRoK4GjljxGK4RgbUsi9q5VFGA92JiUrz/Ock+xpSM2F6KMoZ8HrBq1z0vYCm0r0VS8
1hW4F2mLigNfPbzMzSNZRJFKMjMwAu/PA5P+ZCdq6VatrWroBfkcanwGi85drR6E1+4jEnzzvOHM
n3gwgktfjNynZ6BYXj5X/r5ahke3n8BgOdCGFWqgpNlHUl49ggpJFTbkGV8zvLVnCi+agCavsdPk
lUZ/QjdCwteTw80eG0h58+P1uGZUAMkKNCojtwDDQve9LnvW913IM6C5uS+gcljli+9gVEUucZjf
ozYUoQ7v9wI+Rjqw9HWSmWGQBZWHVI8ddZ1HrMAHA0v6w6VsOGf9XYkk60+/I/ZZsQEFaJtMujCr
PW8mbE87Wg/g/sKWpNHgQM6ez3Db3zpjaqxEJ32ax0BEYZonr7GvqEx5AIlnIdcZhCDO8mT8HJMW
vXSR1ZxI5tAJQ/xSjtn3X59z62gd9JnpcriydoDMw74R4O17j2t48DTitR62q5BjZ1/TDY7h8Y8P
WA4sr5B4lbTgfaZ/KRC4sfeMzxSLBxxOsfVHQa6HDS3Ef0QeGF+XxSqtbaFqcU7mDN30emK8Byrb
zOBCIZUrSmzmTEKtSLtucsBwibfPfW/nmF+yq/HIjkFdxXotHkMaTjtmGE1afbATQ8k3Crvo1cZD
0mxezIP3Mst6uKsC5a99fYUPyGUF41DL96/If+WnoXmo1S04+XEJbdpmt6YjDeMepgcZu2sTQRh+
AUjMQrm4VJHzEX66bo0nTJP/G2x9kcspJb+iGKY1xnqWSuO9i7MVf/mhEY+4n43+ScZtjRQthdbo
qa6nIFQjlrZLNoeYiOhwMl9rY6cFwP6e3yXo+IA5TTUkxCz9bbdxb2xCCPg8jriDPpLmnbjbkoiX
m03o97cJ3Xfogw1r+B1FuM3mrehoOZx7LRieBsEaw0CY+oKaXtE0JB8P1VD3f/fQVoWzxFmomnfM
RoKSftT3OvV2z0pO/UnLpuQaRFS2b3QO6kkYWMRN/oS0Ka2l87flNPzlkit+wD9tvwRKKGgXy7O+
HuWkmRnx2Ct/xsW2xy5dhLstEo4PtY6ncTXqIgjZjFWuXqkv3y/Qvi/ciTHgQS2h24Dl8T65cZgY
YE7L2irmdxDrIuJsi/Y1XOZdKIusUjsr4zmUsDy4Htczf6kfAVyyKbwkaK/+z8iQilVeD3BDZnv3
wAFnrCzregmX86HAajTir67EYJfezbfxlHKsFizqV8cEMVIsB01+TztMdyVQy64tjvw6u+CA4Ny5
P/K9w6fSGGQyK4s5ZgqNgDjCP5YnWOlziB/f6PL8xhRHs4RC3lFXM3AppFBqYy2M8UZuNXI3WMc6
zfR6hRmdLA5g4QTtmwBXjIiZQ3o77SUh+aEUT4ZZOUi35vVTbqNaFADGlJYBdeujtkrmTEeodSVm
zwwDIkqVooyiCIOLfeM0UK9v/SfmxGJfSZ6Ve8YQeP8TieZOoVI2q68replILEW90m2cORokRljP
FLhyYf3LcmmPxk+ttCY2KEehupeQcCcsj9Juy4RzV8QPK1NkW9LPraWgXMj5VN6w6yk0bFoCMelN
KIMm8s7vy0HCnmyaQNDrAWmV1KVsLkC5HRv7AsBxLqMBruIYdnuQNJNvkXHFrX62dK/5Hg1qLLki
+VYd5MW9JYMa9P8x1ZqMZ/lFZ51hkq7KxqF/zo+UwjVyqomapWl8QxLPXilIJfeczllEPf6hiyQa
YtoXDA0W0Qj7bjw9LvEXAylL5Bt3n0XmAYrDETt8/0VM9DAlYXScO+Xc1CjSaZ+YJtSFs0E0KSKO
gVVE8ak/k54MX042RYYj7ydE9ZRJ0wyxQkWwsYrla5qQzHSIrzMhT0uCRXAr0yidmUjG4u1kOWrw
GP2R40HkeA9/PC0wVeqmfkf5BAAFspaGbj/2fQNqeZLU9kML2vMA3+KUnvIysGe8eLLoCWB5xVtc
FdN8UikC5nMvItIS0644p+Gnw0x1M7by+vJz9aCtet2u+mD4oKfVTYgwmWeYBRmsRgjboa29g0WF
Gbepol4sN48d9y7Bs3SR6dv1VG/qiDQgDiM5eoc+Fgm/L7Hdjq8t0iTotzR2V95777LFMTGqB6R3
LLkHm1Jsa+E0rt6lg91/Ry023+G7f5FjIdoTPnk7tTGEJQlR/mKGuciWJUraduQL09hVLvvfORV9
B9pd9Md6HIhkJzD1CPXEhrsAFCVRXZuHFKtlD5GYl2yvlH696sslOCLCbQxxkVdMZc8obGU58zt8
a2ZRVcj9rOMPnk6EUUUXdD+ImuSnKAq9NDgFaA0mQ+3/PPVkH2FA7nlgSaomY/fBAjs+nECLfKSf
STotNwTZCRsmbhZLWTbx/9i9pvZ1ilf93roYBX1Dwy+mv0RO9zdorptgDv1UmuGHoLCiBIy6c0Mj
F+w77xY/g1HWPo4hEWIlY8ApN4Z4MHZk23DmVlu68R8r4CPH6gZohwVf+x5DZtc42R6GG/t9kzj4
zaavbONdU13D/MAzDX8kMLdQ5YoicaQ186h1HBKLMxs0sIx4ye9PS6HiP00Ak33RABQYdauM5/A6
xzDWBUCmzAgM68OPxZi4DDUuqH8rNw4j32k6i/1OAfMCW/9W13AqypXseAuBCpNPykmULZYk4xo6
nL/lV7jh9Yd9t17+iuIUMPxlBbGT5agHL6WXFdSbsXwgmveLXrl++9sFZ/b2FSFKnn3jWTa4sFWI
mo8lauCs8LgRwRZZ3DzDwl5/RprYC6u46KRag80pKjp5c9SJZUYzBCqxyPFHvOyrcJFD5g6o9lIv
ZUlqAjIoiIubmcX6sTA+sEnQii0AZVkHCcIrmlObvFnbBas7WEoiRsMYKaT4K1d4/JBvXq0iT553
OMMNTkhJ8BWW454NazCN0BVjmn6IIkPqnP9X0KIfmlXgGGAC6dnXe6YgEgTeBF861zMKQB3VOXg8
nb41uDjIEwVghIUo0+/3k5JoCilh946bKRliWkbOUVe6A2zWy3UrkKauOBuwfY+3E1OF5+kWLxFy
AbFZrIh+rHO2k6ULMTB91gFttcwIxG7Xa6eaG7IqKmIIGdGB36Urws/EFTi7cRf6peTi0HIHwPIh
wRKaajmQOPV3hGzf5bwbJYCy3hEiha1N/wL95xe8L6YLIYKTwI5VuRpVOs0wPC9mEYnziMP4Kp8l
WsxcnF7unTs3SncwtXWX57kQTlHGao/nt8C4AmFItpIJlkwOs8UmW1qj0hwe12i5oyat/WgLnTcl
WdByKsDKZp9M9u1JGcJOeCeg4jib4qVOR7vI/e36c4rIPXt1dyCU3gNjspe+iKrfrRQbUxfaHJvF
KEKJbHHVL876+1tpZJZfD8sJAo2pwMF0IpzmsaPSbvom5JER41c2R0IjpmByfVlScBYB3yzjChGY
TXXX3WA9GfqQc89CR+lSyCADHXCzsm0SnZ7GY3uQcJ7dSQ0utJHpRNQX1ug+K+s+nf7J8F4zCkCu
cWjobyP7g43I1vKOpAK2hP5GvGKxCkKa3NKMYxzFyxvqlqFydpVjxhu2IwSHIv5THexL+XxNH9Xu
WBUxdu+3INZzLN39yngwqrZn8CulRpFDv0tmUIbPt5E5bu3pZ4eaCjzVzrDMFxMINF2o1MrYLXm6
q7f658GCqeBGIUrfO5rcU9n0Qe31pqkXDkr5TdA8wpr5VmB0QdK5pMtxNZ2ec41P/3Drl2NziWuu
7SGX4IXjq1oofMAIapJty2+lWVOVgbDeBX2EIKyFIwOHF+C23+7zoEQEdM0HSv0cImNrA88eRWHc
324MzHkDk2EzJ3iBk5kkqEMLuyCIowRrJPSxlA4gYL1LMPClmxhDYEO2VxGfElBNLzvDB/sY8mLk
libhcVGRs+TBppWx77wTjLGOqP2IKKSWpRNr2WriXeyPRf7EgqfqTx+D8G/1niLBm1jfBGDlSBew
Qmc6KIqQQn/mSNjeVf11KdGsarYlEXNi9Q5yzzv6skriNJkylMZMH5GCTz8oE/SdRUzUMpl8TQLt
o8q0fx+a6+mw0//fzucx9oLEAaLXWgnpv2k+7evoBSqqmySw0dOscCKSbQGCs1/88tXJ3JPOxoFh
UNpzhx9RcGMrFKTA0g8xv6JEv8tP5G6823ynCU9rKb9GyY9b3b431qvS8fUmXhJg7zSXfmRsBiwv
q9wyeZFyGZgyqtcd8zPqej1b4ZBbQhWYgiCWWw7pUOArLcHtIYm/yW0zCCNFN6AxemHeaOMwRr6m
hOQU5h/UYU940U1FfDGqBs4V6qpj/ovtfjzhbMoJ/tszu0tfHQYIDghaYn+Yp5ApAwnfg8ammncO
ONzW5b1fbHrVxqCUjk3DEFnjGEITLZr7g4E250g3laKX6GfdV0AYw9zaKKKxOu9abDKd1kRv/5va
OsIhDd2geIF3SuXrZPBz17SNXqX+gWClLZ8ByqBkDlbEOIIg2o/Yytw+rm61h7C5v3q0XlYrPUxe
QiTZ/Plo0X7k8a6MRQhU9Kc0uQegbsM8BQxHOPjkub6z6g2iXAyJqOc0a/5kQic5BHlfpVzDs7kr
y4gR8QsDTRS6/JXVCAD4S5SdEam4PN0ps07qo+7tfx95679UhJuMhx2th1r1fVa6iVD6qtEE+mTq
ugw3YwuL5I4GSVqlbOW83vFZB9yeUzHiYFXMsj2guAmPq6buwHI5f+IJaVa604vCV79gSulphP6A
ygk10ViX/VqS08CfB9LduGnkjmrL0X7Foqj44D9ssFNdQEnvCNdFI3lqi9mG8P/MKTdXMVTGHy+K
26h2laORadUdr9kwCPmhi8sEWYAPG+iGG1dqtJHYzm88WoUBsIrNjBdtZ7B8hB2yNNHPDNMr2yOe
Nckl6NHlXiGumbhrhyWJ0xlh2qxzXPWgUn+kDcF09Le2slaL0wu0HMmI2db/Jz7OMbiU7/HK0pNH
zHeRIWggd2t93/QnRqZ9z5h1l/pH4t26wXfb0rLesbo4wQ5ndRIng40P3FYMViI0hWuD2JeB1JGX
n5HDnVL7+ODfCg5f9/lnqQoKHGnT+eL/uYinKuul7JPznkWX311vHwDX6sEf7nuFhzbKAWx42uLi
0lSQsnumwcugo50naqh7Upgmlha9HxnjgfFwHJs5BUcZVbDbotPg/0+vtkmXQGakiYn2KEVGIAHb
44vBbdJ6is+hK59VmdRi6H382rwNn+WCaK9ZkQfldgwE4NFz0T/RJz4jbF4v/ZWT36bTV3sjiTII
0KNoXh0oKM8rPhqcKZUGlmtLsaWdqfG8wT9QS31rD6oF2SRG297mprDXK5uHGIkza+AByf3ZecQw
wwq4qylwUt81AKPgk+ic0ASX4DirBigQzyShvRq865J6PtGg+fBYfaB64i6WwAK4DK48s+4ZKWAJ
G0PjYmxwx/H+KT5j06GlUNa8LWQUUBJVwf3skgkiD624go2aaqI+5QhskaH/fpyQOuKfX8zvFlRl
t6guFqnIbSnvIdBKIekk9xRiaQXqXOeh9hKCRZEgKNbQZTg0YBFqOB/WbOvOTBtICOUHX9jSBkHg
+g37ZuqCQN7fTg1fGFyqzbun7rOFEa3hAG6FAF0Z9FEBa5paR0zBHZtH8emTR8QqQ6dy87ef7UTE
TxA2NJPLnTkDmCvhfGiCaKVBfWt7f4wPBVyA0ZOkfRtsUKu7mkOrRkpwX82hpazbFR4MNXha+3Ay
XqpXXBtJbLf56ZWs4bfimhkW4yDc3gXUIRlukcPh4ZPqTkK1UfDXHquvJ4mSKo+YzkpO6Lvy4WqL
hFhoCo+6DfTKtb03gBEJZnYJine3JMNoPT362V7HiJ7Icahe4QN14GcSKhhzrA3Akx/7fhj4NFSg
y02n7WnUkMOyYNhVVD4XwEhoMwNF+CMd/Ny2olhiISqivCj9kxtRbZBkkKpKgl9FOILlF1SnGfvW
elLBzAZRdLa1hevsqTWDhc3zg/Dvy0neBmQIL1Y09KvRmy6KrzIa5kSmZiuydEYmj0OZznlauXA8
le7IC41SB4oTyTpDTcR+pL2KEPNyieIdhqi5BZgFXOmNo9K5cxknoqA0j5pnSC3bVWFbagRoWBqN
BQI8ZkCG4ngpI3V00W1EmTO2wkU3P/7d9Y3VcYGLHIu5QKZ4lsdfPfwi6SOctd07Y4E/8wJkIO6z
38h+MS1/zPUzvGF/U1bhuZBM09BBI7o4HCPzjTpLIcuiDz87KqvqwXekr/shp0mBJJKWks+j1VGB
zuT/uyTqjwwqEMdmvj6sVEnsYS03xg02FeEAMGu+6en2sL/Wg/KxVJPMUNwo3JDdlKIKBEG5yMGK
27OnktkyJQ/uP8mWVSUJthBazK806IG2telPSn2pHBL/C2vWESR/eLhEaLDfirJcXJnO045Opd4n
fFedRYlDj3RntJnSqBoM64BfvlqUFZKH781TWKYF8kEUqNu3Nsm+dTuiaZKOieOvmmiU0qxDIiy7
iQjyLOg9dy0yGcqBBviZHkcC4mNZtEMLNT4ZnB3PhKJq3tPo12rfcN9acAJTftaDhopDXugjl+Cg
OxUGnTiJDnuUD2FA+05iG8cQfjmXHJqKcD8RNzb+Vxzqxaj3UHbhHas6z+/KlbQuW7m1MCg7Ohn5
E6R2cm7Mr7FyfcoNOQXN0plgOG6N5cSf60cJULKcyG5ZJpbG6HwlUOuaau8vUYv9Pmtkt1o9yKB/
z4OPr6fzsfion2qd/bynNAKXemPdKvdWmQMO4rPfE/HJv/hySNZ3C1TEqy1nygV7958sQ9o9/l4A
/zYFLPAx7amJ3BLsELWCf0qd14C9sL42DTwtgp6+7IVTz6ague76RBHWhqca1LY2x3Zh5/a38eph
yQO9aBfaJnAPIj9BBoQXJrbRdePBMdCX7hfRwb8m8Uv3NxLGRpi7NMeaWkF58u9sj8gqpzRIy3gf
1UCzrlYj/M2X5tPynNuyKbne+mqHWu3xfRTEBg3XIKk71ztOwviOgG2D+DsuxyIrlIstp9AH1YI+
4EhsPnaEVXnqMeveqabyHcLMmjO30ZOvg4Uby+0eOsnpHsAa6QgDxJEhPerIFEWLiw4eIksq+Aw6
RE+MgCYogDDI9FbDuj4/8US1BaseUOd9356eQYv7TlOxpJ8AOYiGpWNpOIMP0fdWYz4NyjRY1o4C
qfkC+h9D5J3eUmvlMFITrZ1pvuManBpNavEzfXZZCcdwySbgbma4SlJt6JZe+RBf+nbdTsiN/9c5
XM7v8VZD2cHWCBn6i4dpYGcnAVV46ZYxg0BL1PfMn/aeFKOdDdVXra2romdOuJfo8D2HIeYpl5/p
DsCAHZc50+KIyPGReqqkoHmZ4kwUvcGB/QZDnK4yrdfs75mDRcFTmHwtfuMPjgl9RXNixOo0c/2f
pxXzwIKgb/Xs8FDJIwBYIlqDDhIqwjh4WfI2im0RknXjNVavvN/5iv2PCJ/yUKYEcZJuKxGNbLj3
IIa15JKhH9tigCEschBYTyhAh/fdRSj8hMFOnaQ+1+3LiFBkkrNcLBqH1EOvFf/vswybfYnEj934
U2JaxCZcEAYYIYvM+fcVkxSoeYNX/96gGT0R6R/C49V2TaiLeDOhK6JB+EH4hzXzw7qympbFcPwH
JdVVPR52NSourTQ+Vzj0azgEiekQ/jiLg3gNNLQEm1M1OglF85fndV5zyu+baiOK6UOTMGWQFDet
4pLvzK6NJ+vyGd453OJIc0NJQfi09q5YyUP7p2zDY/WCWV9K8v0Oql16Do2THbbyM1anomoEy/+l
/D75mC7HOcdpWJtiROH+aQvAOrg9xWvynWyXpiy6LAFtSu8itgRN6sGybMFuHUHPt0DIeHUOXL02
pE2qQvvF8tR5DrbpC2y33Fahtd8U8KOT6L9Q1y0z1vtYu4BvHk2xXh74cA4P5W6jI0jSXbYriFmI
r0KXO5+8XCyPa721QH0MFU6zSObVK8vVn9vLchfQZLqqR9TBqgdvgvrqOyTfa0IMPdNJ3pPiO35v
5xdkiPz4V1W+z/ms8s0XH4jqy3Eo3C0mrbV6kkku9Ph9fJTNwb0UtrgCp8V5DPrkx1/VJJ8Z70iU
J44NNZRpdRYhVUnJ1L1gps6OUcvsE5xxGaUV1+e4U49iZeppWQncsqao5fsP/sOeKgx3xvYbQvfj
/CBjEGheaSSyNlRnNHBnw6G3oX9o+sNppGyhNpojI4yzg/kw4b86y7ayd4sabwYxBH0adGJFECJd
TkywJWkeYVR1S1DFo8LNauj+HZ+khB5V15oiz23eiwLVuhcNMAhnPT4TCHBBs4a+xumzqASUCDwA
vnrWnr7jxDuD+iXHTTimamoGRVmH7D3FcI7d4uVI4pix+TovA9WKL+qOlh2NJ8MLipeHOemVLw8o
e5fub4NxIKctX79tIHN7AAdo8DM3OMvuhUjhrFdl1kaDr3ReguH8puhIhZPU3EyUufo9AVaClT/A
8zBV6X0oEZwLGVfcN3jmMcecvhXz7pOOixzpSm70SNUu8LpQ+dzLYlzrAV/mxvMdeAc7pv1rw6bW
Fu5/nWE/nPShhjARWQ7tnxiVuZYZpsFqaFRoMuWaN5z4j7ZP7SRz3F710LFZZsi6b91+WQDmPJxm
+UuJmKo08yROlq8Wy9nTDPdr7c6LO2wUbs9rVZd3aKV/8Fd24ygRBo92wwlZuFq48lT5p28hoaBo
dpcuxwnug6hu8Ezylvngi63MMU3TI0Tv6HmqTaq7jv8KRJs2SfFzSLD+1xrKzf5ppOB+ee24TQ7p
ESsaUgJzDx+s4pbYtAGXXkKhLJbQ6rmAI0LkVKBgnQ47hkVzOqmTlMtQE52Az7JYZVGVVPNVvPmy
4FA/s/RZUNrou5YKaBQuSuSQxzNG9xmKi8wxxiOB44DZPUaM5a/wMTfcgYxg8aqAm0QSgkwaHV0j
5cAE0PFzIsDGoZy3BB3Kv18o+4r+Q3HBQVDTqwQTMgwMiD7zBp0F9fxlvJYcLeZmtpCWhGgFTN25
xDVwwMYXhJoozOzQxzUmpvaPTMCXi/oLpRTrYPYeLtamXGlgnLMck9o+whtQHyxD7EDlYEDy65EY
YE0TQ2OrHc+dO+IKtT20g2sssNiBN81RLAWAmSRl3Q1yG8tAeA1vRDlBHr1agjJRqHLmLZ2t5rjU
3qotboXoT8YlnJ+dUGyfnt/z3ESOfsCBfA77g0bERLjTgYFjyIOZUM4gwPxGkj40OPTHFFXns1gM
vcrJtngPCQTbralDiXpwy3fZhO2VN4I7xG/c7zwf30j0kjcCXNw+eTUdEdLEc4mkv3dUApkU4/PH
YKVc1e8qg5n3MIoox1IV27L7SItQR1WVKqK9GFgf/cJvz2973VEqU0s7Apwg5PL7ats5feIxHsUT
brrkK6FAaT+rQhW+3GPvOY0D0ihAdCBPFrJRyKWVvOTIP1kk/wS9EXJZAJzS4rdzb2soS0JdoRHq
Srg57ocjRH9CO4DqKiPsT0ysi59s6DWJuPGb0tFh+yzEW894OB/D1RWllQa5ZRjjwokLWJ9Ejpb7
Ti+rVCA5RMGaULHFlJXtkjjRrXlPQaxXie/w0evl+IvhuptI/jClnTCQTr930E5G0yrlQAqUh+a6
fodtRB9n5pHXJtsgLd6k/4+iQ20OakNd0uRlX86hanzu7eovDFsR0CyeZoLps80vRedkkZ1GOxBK
X7CpxrYOODzei0agai4mFZfLpwmLX0YNEkzmRHSYth+umDuQLjFeJyU0Zf2f3mWDlMt9HiUm7n1B
PuxMLP5jvPInjC4J86kkasi8Jd5hxp6n6Jt3vjRCzm+jd1Lj88onJ+S4rIYq+IVbawyjC8KoI5F7
XcWf8zAgP0metZZBodnpoDQuB9pnfKQrv331SQG5vevB3f/zQEB/Jzs+YaADOmhj00QLBZtNhrol
rn0o9nAqyZFtXJnkYHAxsNS+4RQAmFAYoFNmZlbEuULVdF7gqlC/GnMDa7igGL5ZvptY8EumGNDO
M83uGJFoydWtRNXm2VIivFFbAxl7cLhDkSnne4Dny8p8hJuJ1tByI00Eyd/WIRik41rFleIHHBsY
PSmHCWiaV7k28rMQ6ZRtfGyVkcvznO68v/xtw02KlXLSbEYDgrqrcci6N3PEZHsy0aqHwq9uDZ+A
7q2EpJsNh/AkWirLA65b+qEbHWUu+K00Nhqe6xhn0pZh2MEM0rveYHqQuYt4r3Vap8n/st1+1JJZ
RUu+h2vytdtJpNqQU346PYbzgcSNhnnGvzBZ/TauuExiRuPSzBLsdad8rUFkPPLrm8mYbjIFz3ii
lnQ6wd1tI7K4TObJQh5BqPo2AhnpWrEdbGIVh0MkgokOPmeMYljOClwLmzZ8mxrk2VSO2+i+ZO0m
nPz96iu1kV+nihbvz9yOe7JKDzlAUpf8v5tYLj9CyUeHdkTK/31mNDpXozu2HvzmipyMh8SWa2Ou
uUnANpUdd8lCxBtKPECaRP0uzZC42DQEftPU5jj7wJYDjsEJ8kgXUXYgL1iELMAbD3TAgR9bVO8p
i6ldTQ11AA4K3G00UJKSMzMFhFG8NmQzQxBsT/rPFDCSc38APBZEPT3EkKzdRbjGf27fAyi9xZJe
mYS0ZjEKcYUQ7wiyT+hxPUNzYx6jxSZLCfIeZ4AkfCiLh+RjOiIHYH00MDm9iOQtZrnhsY+5IoFg
32vNU/74yMWaJFGF4YArxGa51ZXLbd96JWcSfS/2J7LW3bgfX1GIa4nSQ8QzmWeqsiQYWYE0iWp5
m6RSCwplQtzv8vGDujbYvzRJtDfZTJCOHM88OxbWyQk+VbTTv9fjqoU/bpyC7yPHGbQc2YpZbVtO
3VucnOonqZnXR0HzlzbCqQsujg+z98EAb/9x0/ePTEZOTSxHNUQ3qzZGXzAXrW0Kyzw7TJogDaG0
HwrYVJTcMoTl6rxlwEHeSfiVYT5zCBM4g1bOSVc82k2A2W+sFhkkcgwjGcw1Rd6xp5zSeBlgL7Sq
5VxzB50d3/HJXGGkdpqdLeWg/a4VO0i7pnSBPuHUAf211JIsJwweAkqzp3+XbzT8Z2PG9Oq3zwKB
XC3F5JKbjpl63RjRNzbSSJ4cOdrn+zAk9yOuCdMzB2UMujKATxR+tPi/5656obZF2Bf7LIhYsMkT
ME34RFbCHQWEAuqPbJNpfSyW5WzJEgTbWon4ka8ZRXkxr7WAG8n3BIxQfwssKs/uQ04Y8sMNLb2T
kLLGg1liPDMq2s2uThp0Bd6RlgIHFgUDhxsZPqbXb92ptfYtT7pjKixqbMCBU5YMZPaCBaNmTQOd
oq+BFm/js2JvTzF766EhbKV7absPwTULu7tC7gphvILcQlk8tMD0S6xp8nPwtX6hfYkSWj/o9Joy
wr4mDfVNDQeJ3NZMMKvdSDUbYJH5zWF9zP72z2trVzLbmWbh+tR3WYtCz16Z2i+HbU8sMQTlFXLM
UWI5R8zJYQ3SWz9yloObRobVKHckTqiXvkR/Kg9pGZ7uuk3lTuWUQFotXQ4OxxvFfUW+PtvBvA/a
2ZEXPaJRwD6P0XZOajNzJ07yDUKkL2NzSecZHw4JiFVBIw2nktc5I68ao7i7Fj6kpAEfdZ/k4OMv
FnO5qKvES/Ip5bofKpbSH3Jy5He6VEOt4F4L1u66cFeZc7PEwqimgeR8MLu7D8OmObtPXPFY8W66
+tUD23J8r0lmUDSznDWnIUk2JdfTQ/jHFSrhn+UVtY1O+U3wzX9ytMnbbWNDfKeIcH9iO/6MpC30
6FyXdcpsynE6aVX/QQn5yWvR0J3pCSZ9xg5STLG+GIz1iNuGZamrH5GTNFz7DhsoxQ3QHRmDNHME
N3ZB1Ak41ACImJm+Iiq/Jykx34XthQ/ofhpfX5gOtG+sXI0TZdQ7ViqtYBxCqcY1R176899Ve7zp
8waw3dMwp1+14CrOSbAIxER55kDRvSaw3p62HTSjIAcKsmLc/fZ8Q4Zf049SJ4kNBnJ91RgCZUpw
ycaBxc/5d3kIaY4Q2+6E579d2nLSXH7dUYRUiBQ+YUiObEFFIqU1YdC+qpg1e72Tyhg5oMjvyaen
GmymMPmHZh0nzvZl/NF3DA1qBruSrIwnuEO/GVyJoYT8snwJ9hzFwRMHlb+gVaan1mJidKwtjsyn
/eOx7VftSmRh+oT++vtuvZGhRCabSHVG2bGyJFnQ3NVqmU3KnUEZt7A2LOwHZPzfCLkcba1pohOv
3sdv71w7EqhCoxJ+qsLvVZRDavduDg7iYJe7UqHA2OThG6w6n/iRotngv1dE/iy0kh1WAXNvZzjF
3UamiqCCPvYAZ2sQ9y3tXncB0CQG7586lbTPUIwmCKagUPH91cFZzVkMgsWniNBLzzJ3ZwqCmPzE
ngOOIf75mIRnNrRYGa/sEc/4+pMGZAnTFQEr2uwf8EItkIcAZs6dv2hbjzOoYdfTUIZZsEqeQAs5
5pJg6jXRVckWaFv4NiDkw3vmi1M6fjKVUBHyPlbOjQpnBpnwYA9S8c+6tHVB+CWt//5m6oRW2jnT
oICn544FwQ7Iq3nR6bGLk478jVSlbF/sjrqOFsEbEu1XvNTbx/NRnfOprInC2R0QdEErV6VUwRPJ
rZT8/9TzjqBKf4JrNtpsMNaHX5EgXtOv3xWhIkICqsejBa/9cPDy8R4eyB5dfwlb1CZAqHb8Ic71
94aw+noUXoFPVzjY8rKDWwV/5EbrSE5qv2QJedHLsobJPq2NfanL8LEG2C1uGPec1Ln5NGkgX8xW
aBCRIlGqw+dCvde8zZc8z2vhTRY9RCWO0HFiB7U+Uf5bJnDZp0JrPOq0xrixBYUdZXNTJ8rnYuB0
+513MQiUrrXDJgF8nCUnOhH1CJ15ee2TiWSz3R59JS3ark8tV/cXDJJ2IQ4WaMe4+GZbow1/5Xuk
YzFEBB/64cPE7ceUXIWF+QKtLXSQSlq0dT8Lek9J/m56sB1JLi9/I6eZA1fk4026Vw/sODsveV2O
5NFpJ19bFfHnCym/pwM/26hU2PnRzbljRKXE4sChBrY9g9U2smmFYGA/hzP1dlImShg00Z/Cc9t7
ccwWhMKF52TO9t2FTwn0k5ViFQzWXmAMC5hHn1fcHh/Tj3v0J7qzqUTpubEpmdBG3jwJ5v1RSq6K
w2az9M8/s2xSeuOdSLXw9SwIcNFDsInCJ11mR10YZhKs5T6mihlGdfmbx6tEQsfJuCtBQ5bPAJEl
x68F587xp6t77CBal1qqmEfHjNrAPzuF+QAoNHsZjJEV8ZUvPOiE+7zstUN53toq6KsWf93T2YrX
1A7k8HiXwkYz+VjGlbWJEArBlWovtwrJgozmUGXmOeHOcOQ1fLEiEqgB94D3NyJnu7PFKyra+Ftz
9hNH7eZTG2/YCaaM/qVkzs1TzAzbnkpdVNm5AIcZzTy1P2Ue4xZ4zpWlD0hGEMSU6tCH0UadcnIY
kU5k4pJjP5Af3TQGf347Qybl14M6Jh/A+EQUoaRM0vzcSNg5QBi5NS7hATHqwIb89whb50faa5Az
2p7M+SyO9zs412Dk66cfBTH1QH97IKwLrisDIYokpU/2vHpdmHOn3A5J67n23bv24YGoNoHBwuIq
YQwbaVqrIbkLIpbPuO90fIUcQh31mCpju1WZoUjt/h5gJdz57ZIesIEk4z3uXKOeZBPvvaZwz7IS
fxYXt3dTxqveor90fryxk6Utgqyan3SKMSusC5OHSBbkjKFIvzND26GEWTaf1MIXf6Wq+ykyKdTx
6E0mCMkKI2MTVPQ7xgKytd+pqZ5IEFx/C4sGoM98Dyv86siArSvV7qW+9bWKGt9QFnbzL8+yK2aa
Muqp8Wn3WdILEaSMrchf6BLII7NNm3CyCJs6fTKTmNHcXFyXUFPBRFgXZkNncWFlAd1OSLxg0pSv
VMa+jBza56wlEgsNsStrTr/kekkxIHMo216OEeVgZJsbhrub8xfpXCR8sIVf8L+udH6lU6veVOro
HiY2y/Hxn7zrEUwICi34i4QEWSZf8pnywEVqTA2VflRvkIndmXZMOFWU+XPFItv89wcOIplot5nQ
GKqyvTcRpfXHJjx9u4I9+NdoWCqFQTCYCEDBivA4tUbdgKgvJKQ0nPZR26po82BB7QgF+M6BXKa1
42WuNx/xycz+/BkUadohJ/ri0iS8JvO24i97jPh+FVWZ5YgrHDUgRkCDgZZ3JUlIbdNQt0eZMW0M
fPwvEpxZvV68mtG7QQ8nf5MRiCvoRcHZ7L/QXKPWpOeOQxcDZNTrqX0cwdZqYQhnv/bOk3AhDc+Q
Xg4nG9cDuzltZvAvVWeJhXGU1zdLR9ELWpCostdEWso0Np6hjw9x45bbxxN/8LCDuubVaa9oj7gt
PuxbO8ZFgVW1gvbzjjZPvYDhe0ix/MJ5P59ye0lcDDJXMr1spsYNEtYtAVcXj0rFlk17mimqAOyg
IFfO9zo1gv7PhKVyEEFZRD7U6XulnsFJoyxx+AKJFO30xj3YfFfQm03uBCohgOzV+fxwWBR8Tios
ET0AsTzwLwBBB1w/CJTO1Tztoq1gxY+6IzfR384rpQGQcBpX3nn3XPaRWL+bCgd/ZTw0fJGfQOxJ
sml42/aMmHjcH/tWeXlDEGtMkxx2p/uhbmgxcmNRcVmYvZ0JskGsMClc+bsYggv+r1GbUsJi9BlC
XATDSKMuM/qoWaCFDPvGFkLUyXdROU5ESc33w5Inzr33lejJ1OmjKHnGtOXq18WYRvc0ug58ZtCr
3NUiipyLF6ZUMgpTOaKB7hh/ozMxCQ08pIFflbBYT+VeReLjbR1VWD9KLbeaj79KbUR0Bw+o2SZQ
svgqHGCm5hSBuA30d/ZAW5m/csNifELVWWDRK9KubXOoxMpu4JzRuvT4Z9CDC15pQvOOPTeNDnuD
+vNbvjPlhhTDEtbiHiE5E/jr/Q85DsDdNMvPnzVvJWUdGAvTSTpF0vV1pqeztrkGskQkmfe7yW74
V43U41y3NJ8l5dyRrjzpSFuzaBYqrl0vzcnIPkC3YgJJZT37nWTgywjKT+3DwSOyBtOqWPZTzgJk
V3UiEkJn7GRCa6eGzdn7kHsREmkhbQoV1JzwxN+iiI4pHXfmDUct/twkghYGPL0gZyLzgpYaM1hB
WwOkZsHLmR5woIuNn4GZnQrWKXWuvVYeulU36YyiY1Ocyht2eH2I62IMUxf5JxMiY9+DEN4e8T6I
zcESuUxrRTEQ4Y1F5Yl2/NW2vUFtux5PhOgkbmSjEGhPf2i6ENle8+4zg22f2W1NTaPc9kOqTGOZ
rnDtlk/Pgyi2+Is7oQoNDdTfp/zUERqXQbNFaz1neusWhZHsJxcQRPlOj+53mf4ipCLTSMRmG6+m
xwgcbUP1N5gPdGUAbG4sYghDdRfHeyMfEUwrTLW2Ewjgif7V9vxwMP9DkP4V5IqQb5ecjGWrUCUA
8Yg6vw+J20DytrPT07V5YMsRQE+F2smRCSgsjtvfKzdlQ14FHUkfTxNFku1YoBDSUSeSC+6XAz3H
vmLOfUZIsKuScLr3iGgkZe/zZiVVBwUUH76Plg7bAW2FNcNQFKdRVIiuFewNe0+d9nWKzNrcaOTS
I6lNZvMpBnT6jt3sLmYIlLNvB5SBFp5mm7Y/ZdVwGzC5dICX2PoPR8AXOGYh2wXhEQrWnJlSXPdf
GlKx3yY1ygZ9XFLZn5ejYVUgtHN0GOXYSn5P8J/2//rQ2+vY7CGSIobTNJN/07thg9ad2CmiwShA
yam/UNDgEMGyKmaKfTdIlRNr2pEE2LUDaI5nx/sMeZYx6sMoNa6iTNVHLSrtFj635iOGwzVlWVKP
VbZKMEN9KZnEQ8yr9qjLXNV7+wSZYDncB7TflhQhIAnmVQ2PoRHOpT03lo2utwe71cExiO1wxFBD
/TxkzAAeT1vUrMrCo5NjKaF6Dlr1ovbylhujZ9cjkBvW+Ok9WNnVVnWNEQHDeXgLY44suwGmDmKh
O3mAe3LGYHFRdzYr+pEmucMvBA5LOK6lLOJgrloSrTsjkvv7WrnBbmv3U9Wuuysk9N293yavXdaS
T5oAkWEZtjYyWgAN6w5h1w4N4EYo9/GJUmGW8yYSX6ctXN+SMYSR2ckO326A02P18dSe52tEWdMb
eWcXZQzCUKNtLMnIOz8F3F28NURv/XWJem91uD2cKY0JixJe/SqI3HGittTa2/IGFKVkWuviG1cQ
eW2isICqvgeb8AS96yebZUUdfvY3Ix7jp7M87b9y0RpGN/UVnGjqMonb/995yrbsbK4gI7u5sCYY
J9EFgS3lgRXRW+FyD+9XOg9p7TP1U6UXxkiA6mlIivQfZnsJRwfTtG8zRQNIXEoYqDXsgJxgYrvF
mw8CDVD/570yugqqVPS4K4DSJRx3agUzNflXD0zDdMgRFnZ59jxsn+EcaS3nm3X4Xv/nSLcVYTIc
Q/+eSoGfhIAfW2+P80iwTyPQt4vyUNuNd6NZ1KGD3vmvvDAcWMQhbSHLcHz34axrihW3WU0SMgEX
YksW6TKwzuvA7eNRs14FIf6RFRILoZvqDJM8z0vH0T78pxuBGltjhC+NWgU1gTNW6MhFkV3JXeQg
atnmh/MSJWi3G3aNDdPlTNhb62sA7pO0SqzXpRqoTRGbYivFNMU4/l8Q9wvHJbc1mJKx0MDkL3U6
WNw9tLgpcJ8Eki4KDfSw+F80mP1I/555T09oL7+bQK9aptW9quwUS5dVfI+uWX4xgl1QBmt1hK8B
Ibn4WKzLGpmuzTJ/Kse/LdchLwdelUYfbnw9SgFiZNog5HdgRmFh36BwxAWxtHzJm5eE/A53q+Vw
M4JZzUrMpRi0dEVIVaS0CgwZWe3SjP3WqY43INtqRBdQWBnoccbI5U86Bm6i0+auJeXOnmEMIHdV
2Q7DtNOLQGqqKItYv4EDF5vyVwwneseLdl7iCiHKbyDlL10U355HcBoANriDPeW/FWdJY+JagCcn
eGVrBcudH3qjbaBRd1DeRMIW4pShyTs4j0bl0ICAdbrb3AfPS9I0PYKqVCiIaZ+IBglkHYILLrli
IeejrsSQpmP+TU3tzdVqtah0v7ttiudw8t46Gv47mpytmCDebrbD/arTtNL6hzDe3Sv2JJoDbMft
MXYe4ItM+3RvsTcyDNL6CNgUHFjd42gnX1zR0YFtNYmOX4ck9yMQ00PM3AVCcAKdVH8hh9ZTHkZD
w6UwX/PrGbZm7F7u7nViFbv+VShzoWTX4Gd7x1NVJBVvP/80QCM2nZXIM+Cp9MBQrrqgUetKXd9K
ueJ1brW4fR3Jc7spncrH+GyCN4S8hTA7/2mpI7xS1E20Gds28ukY9Q34R/UN0IaJ0kfMKud6UJNa
IomHBtkV0Z3xwBQIgkzyZ9rgNlu0OqPqVKPIlou2C7ubwJXiN8dFoxNfugmWWZhTi+E2oeq6Ciyn
reFPQpTOvETR2rm42Rhy5b1Nw8clbaMo1X1v7j/TXy5WPcX/ijufWQPMuk9RV1s0+T7Lze6i9C25
9dlDlN9Scn5z8K+RuoyWAb1yIvlk/vEnsz4RuX5vUtB52UIfCpp3dYGUgHXKoubFHkKtnnzeTplp
LeyRrkeVJeRmNMg2W2T6TPy264xNvFJpV8dKN94P3nhEkeXR1IiIm3/tjRDSdQZ5/nv9QI/WQ8h8
TEc6vX8IAUBGhRhc+Vi6wNhF42o1DwSk89K9RvgkdNZRGUlvVjeV4RLxc0IEVdQJh2LOl6hGsRsY
q7lU6eQ9KtJQcRKJLTwnsKDp73tqDOdDV6Gaw6BtGw6WX1ge3mEE2pOVhoixollN6J/G6Z4ElNOm
HAFZxp2OiUUlUKjhW/nTlA7V3bNfN940A1EpAtf69nOpxtk9zwB1pJ+Cj2z6bfazZvcl2p0gr1nQ
dLDp29yLCbGtKO22X7A/dqObwqcnRg1X0MkE+ELFiucmTxwuOyQL3bYlnvSFJTIMTgwl1NCzkDiL
IK2px3OkaFI3nHOfHxijY4dk0EHm2mo/MAJVEbViojMYznf9iXAZppxvNdQDn18frUWOU55uV8ba
hi2jU/Yi1vgwd+ciAzcVuji/V+MSh7qufUF8HC7BF9jdLxyrVLh2Om43PrQhwnUrBf9TIW3gWNcr
XLpnajVHlSy0ciAcWB1kkDUcGMuCgxHhljgANgocoNyebiTFcAybAGY3IesI9JI69riI6FrDKv/R
qBXVLa4b+bytLnQ2EnXUwgbIyMX4R55YK3bVRQFWwDJrRFJh/tL31mAj+Retm3tPAm4tvDApdw7y
+HP2WJnRl634lHl+WE2rsAuiGvE9uf1jRCtoIgyWr7HPSSYwdOJIzZgWoUi5KCFYjY/ZxKA15qNc
3lqKwny0+U3b6X/fjzxaVesAmSxUvxSV5FEEo5GT5dEeSFmGzKi3/a218u6hlSPTxaj37us3WkC3
Ta1Q5LHxMhI98kWYuHx3GTnU4lpX7IfBS+Ng7LADkpFhcIwr0GGd/VF2O0ld/xOCwG9FWQphAvAG
D+OqGd2AS5yVJaXClqPzBL7uSKi9CbcJjGBCoChI7scG9w4tjE2hUb2G7cT4TiYjTAyEv8rY9/NM
NK84FUmoeyc89IxEeRg0DGX9BDKTkgNNvpLupQbdUHDJU1nBrLrataOFw2LDBAc3q0TATL5HcuW7
1em/UyUlS57fd5HjugG82RcHzVWZlo+tGBrQjt6IgtE2Z14ye32naW1aBFPpngfBf/SnQuiwsrwp
MbaB/hhXr4fp1Lr6fpW7erElZnjg0xGq8K2v7X0nXjOB4I80fFrqewC566GL+g2dSSTHgbM8IbxN
UffV0wbIamPVcfbidywSoDPxjDkKPodkrE2ewFi0NwhJY83J0koTmX++4WsxZVZz4fUaBs14yaaK
/aH08hY9SpyyXdojWSSbN96Bvb8xPO+J2L/8tysUzBrCcN1aa+wVjxGZKktLHIK6TOVr5jyrcDBi
Dik44rVQltefIynZ20DxKY57AxVuadLGcyvpizMsJEOfXn8sK9ddRbCk+Ge2jTdJFefER8tLD9f1
sV/Zstaxvg9Bx03IXpJMyrY7P3DANoVzlZDLb/yKOD+LEELJYEJWqEgpdqq+nJGCr0EACvNpnK7z
KDXUDdjWXh3oQVSFx5wtUe8X8FOpKAPTFKatrHzmAiFQJPFZ+cMu2u2eE87bIUxrVkDTdAQGffxA
Bjs9zSNnYdDIliSGBShp6rVpewisaD3jf17ajnEKqwHacXCW19XHD167VH06IQU4xICwDcCxcNTK
KJuTMiL0BUnb8OXuBGC46Ibkr8b4jzoTHFEariVRHIbdKmVbwBJWP1Hf5A9qekTOaUyTepuDRwFG
wjGfm06Fz4XXb7X+fxotJxSMO0c0h7caLiHXSOQumtLsKnFE7qaHuCOfV5N/3PalnbM3Rhz887A3
1hfWf+fcmv1G/sz8mUp8HVBAgY81+W769n0XTs9QyE1aBrKmAokn0BBdHvfeVTSp9zqYwZhrccUv
GQa5sz9Ktxjz3yWr6IAUk8jOp2jW9rqbIh5fuNsbOwCS8jpK/tRGbKfSYYaDL59aVUbWAiPtlbHI
SG2vrNknnj0WYrIZk33/Gmw9COv+IU8b1ekAOAxuO8CsdiI1UhJ0/qZphk4ndS7rKJ7tlvJtL1RQ
WZ9QTIavcUH6WexRdtz6QO2HV8Kc9rLzbepTuaBCw8z9zLbsP+eupsFoya9rzrTGbY/THkUlgfLV
blrT0b0E1lOcFID++s6YxwPdiM+icqP25wAicp3U4BeKO+S3AYF46w7W2sTmwua5pDhYnspU6fFw
hzYVZI9B3jkYJ+x0MqlfB/LGxYvanwap+HVDZz/vIg2aJVfN2eoxk1MMY0e4dpUrhOL1qrnXP76E
iZ7HSROqT0a4PVparJ9cxCIbiUPU6xmps4EiwQb4HXKgMTF0dqRpx/Z4EHtpfeZYP29ODB7G3+6n
YwVIRF8nf0s4D/Xg0ArGzJWFamGtP6opqw4AQH/wm1198oOs84oC+Js5+zTNCD6vY5JOsZlwQDVX
yCprsFd8mmGQOqqK9u+OHmGtk+KXAok1RYy7A3wPmrkIef1Vhnfe1EjkuIuhg3RgnIGUxncymZV1
1+4/ZB33im71uhl3p5PHfOhH3ochGv6NDL4mgDIQlpnjtEpuvoKWYy142nkvr2IGnEZYSB32qMyU
PfQmBavwlRCpjuEDCy5JlfTt2BksuoegFUIITx29CKD7/K2mJGGEPx6o/HTTyx1eNxPgBR6pdV5a
u+XfR0HfwCDks+g53NMaALBrDMsHz0+h7gNAOGgYDeFUV4KAIlmIM4yeerin79wyrRqKYe8+WS1R
/IkvM+ditpNeKF+N9nGZg0pFvm9NQIusyyfUUZQu8RvDLJgE5BK4SrQylprL9MXcuwKgPeCs08b3
efVvqIRGtg5AGyDlBRlcony7PFSZDH38Y13R/c76iNqnpdDMcyTdFFtbwBpEAqjaPpQ8nDm1/Ox0
gpnqYP1RU4icEzCjusoI7XDbfGFdUzIbdBt8NeLgnCuq8phB9BE0v70beGfomU0alyPiORNhHalm
eDYn72lDWOyiPeft+JHADz9AdJQQ2wWra3o7W+m7bL4Fus/Opy7amFD+ZlT8qKWP+nV3n9u9uDOX
be/oLUAHnQwK/hANR3Scu/ueCiigW6jR/k1nG4/k3J7gMYF/RpnFI1za2zltszPtPcnABIxSj+2R
9WM1wx9ppSvDHz42KL4yZk0pQ6J8MNjhc2iBNY/WGOuD+K6j6A+AjOrw4c9OgFhqOsZKBzVPcLyI
nFy8XWXSFNTRuh46bdxgMFol0T5PMpxBeUFdZ8/fvDP6jSv7yYbivPXIgBdivSa6FB4dZI0Ji7H0
8gNtIDVFmQ9Mx7OZpwIZnLQMbMFzR/IgoRBPQ+8S0cM14BlBjNcfnBax26Mr+bOjVEOocMQteiOo
eWT82+Dc/pliZZBzGfTrs6IY6k+jwjVx9zvWtbb5HYvVlKO0VMA4tF+RKNlxoSc3eApHyrvF8OgU
MBKPHxw6fZzIwRg2ZhzJvnGFc9lPqecPz00tyGV2s2C036LKDTP2vc6LDSg+eBJ8JzzyNhBL8nWQ
SLM8GFFeczNCCnZdvyWTl2bbSLZ+JyHhbwWAAN5KkBL+nDYGQI2NciJ+FF5G0iqeuLQGfBgCXklJ
1OBjUO800cCeYWeNXzriJsPVA1eVO2wmcvLoqwradD87/2xaL0f4JovQtFlGQWJKf5xPDCGyvkx+
ZG09uL1S8EHNA6sIFG2LSkNluIp55hsvSBwkdLTo4Te9zUA0F/X1hFGXmgYGFmlWNdfkOG3B+51j
/OvS9+PlcwFpuJ9CqVb7xj5BEf44/cP/41La+gXqmWv//0RsiMus+deZZ9v4IZP/cY//WtHGFip3
S5tGMm68iCfZ5BLO4lxofP8z9QWKAwXUN3SHHjUZ27G4av5DHfaP3URA6P2k8Ux7H6UYMrO4Xt7E
ymcLNqQpBoDqWvOoxn8zmVPzX+3piWHOLruAapOBZ/m8HdGW/D8gZF4X19erE1sw4hVdul1nzlPs
WxmUCWKf841zoWZ5CJ+4s4PSxQWy2nR0ikj+u/fUAM/qbaSy8Oe2GPLNWcO9qBvei1ZL3ZNkcDlg
Kg8A1tLwITsMgO55BKJXy8kU502yVEocx6ot1VnV2P1KFBhSchjebymb2yhbfBB5sfF6UoD0nTXc
5ZDrRL9KwfMBuWQrPoHmwcsLPmU10rG1ACZv+L42VDSih24kxRCxY6NwqxdPE0mJYz8VmLsUK350
lCcJKTRo4AYUEZP+ZRu6rmR3iyMZVFqZE3RK1uvoSt1kEVcnEXOyh+gJahxw9JYc19yQSPb5tliP
gmDJUD3mJ6RH5qK5T5Lbmsgtrz49L/FBNgwUn7dE11PvVKbBbwcm1fAo4I3syMJAhSmfQF/THS0f
p0Zqtx9n8sS3Stor24k+MR2jZLMAPiaauhP1Z85N7G8CepQUC0mwEYJjdHX3t8BMBFGqrX3jSVfJ
AtUVXrHin9NlqxgKwIwaTwAIFpnGyJDeZPd2hgtajGOW30Nt21+91/MbXebbYCesVf8GQN4bJlZY
93NpySORCKxSsZrJhkEFvStUyFehstht2YFIYFZo+B9N1Z8X6Z98kCYbkZ5siGfBisxQGNj6A3MX
t2qwudCp2xyfnBnFND4TEgViz0Z1J6zhuqfFrkGFNgQqU0eufYPc0m0pCKLum462L8tDGNuaPJVO
2KkgJpB9Mx6LRpRCkWWoBxHd0Dw+5gnOPBU/dV2fkK7+8jxWW06uB/dTC1CzYxDMizA7MwYpYAeO
aV/aC0FEF7QAWFe5lpPL57ZESIF2zJFu2tr0thI2OCCnyn8YSafM5yB0gibwdge20jEeuIX+fTLX
8qoT2NxWRk/5tFAW1tM3mMUwedQ2sx4c225gaGsPL9J1h8ilB964buxC6rnSJKqFs8XQvQuTEAoC
vrgT9BayiBQ+10HIsOvKm/UlSdIzQ9ZNasw1Qf5oTcznBoZUcPIJFTLFejvkzuQ5+9Oz6WPmxtrR
0EDTAX2iZaYrlQaWrmOXueQ4/59NJiLwu6E3VOeyI0A9Tu+T8rpeSC8ZufkbU2Oa75Ve/0PxhGe+
O4XjCUFaFjqMgj7Bxp423wAvicMTQnQE05Y2UoQ4Amga2rdTTyfLwkJMlVb52u3q6u6cR4BQsz2h
AJ4JQnZ27EN8ZKD2zYuAJIkDd6oYoUpEZC0pYA4WXagCBy6VZ3nNWoJoc1LRxMzveRjCDeNx0vwZ
BA6KnJDXiDaml95gvK+i0sBr5VAdp59RuGMrJI5tFV6UEkFjQV+FSQe9R9lSoaB1b3kUs0BpEWm+
q2QfiIK5U2fvXa3WmYc5zH/ALFFHJhEjQriL9tUrxXVA2v2QCfslsKlU5QlIIxCKaj44nPx/FtQL
mTBXBOxNxZ57TxlNiuTdlC7r2f7aVz2XBwRyNnVsv1a/QU2JnogNaqv6Fb7dEvJaX0RpP2d7ycUT
zhZsT+mtJ0TMtnI4ukKoyDAkRd4qkq5Jb3h+ygTkPzSDYGctOYCdEXBGhQ3Qqj5yd/s/HlevtWrT
nCLLKFAfmdZWioalm+eX2Q97VjM02BRdB4MphmX4Xd2JQjiCeccm6diMUUceGa0U4nTizH/bj4qP
jR6XtsMgEqkEBBdrzqV0M8Q4PXxKdlr9Oj2rtbXnoaMLEZv6o+6gVYojP7oz1ufuF5xMXl0pgJbO
UeymE1QznycrW566MgQxHxGQeVf1eUX5zyl6cNl88xUQNOEFlDjwHnA+CZxFiJPwzDF/SjUOt0Yy
sHvpNwN9mVmA623gve4lQzqHyGAJqtmNHC3+s7poGx/xCCzdO+9ia/tAkO0/rgSgraEDXjRb+ni8
5l3SRFgfg6txpps/Up1KqB2a+ulJlfjVRsGwESXoWU04OLb5h3+hgP8itWNk4/4KcSDLiueUxvK/
EZgAqEzL4AdYa2qsFvlAsJqsSv5NVq3EfqdiAcwErM+jz+6k1ZzDdLyHktsvvwEguAuNdi7m+ygB
Ym45aKPri76ldS4O4ad2mG4EHFV6SzPnR0h0W+idH+S7mW8NRkj3wdM18Q2dy6ldJVD98e0sb8X5
idOOVn1L4eN51mKhqPQ3y610B/6LGyjo8EimbJeJDjc+rfQygjIczeBev4kFmrpRfxALvrLnQAkN
B2UJYsW3bcp5KJLWDXcAZq9toZhNXoWIuOCQIusBbztp6h5wC3uIu/OOL5A6ZErS2IfGWuuZFGiP
YCnsYHgpr8AWupBEMgucHPoRiYDmaq6p1PhDy5fpLsGtQkuPkfOa8m7oQRgG+NlR2RLPCdSvx8Mw
smw7GYaFrI60qCrJ1/Hv90Ku8OsRmArI8DQuBFNxp28V5IxgP7bRHaMl2BD93dadAFr2Kp7gbzIp
xbEug9sCfqa3hs19GjFbwXi+F2E++0qbjDwodcnceFd6DHk6cfEZuZMfN62SgxlpkgaGXlnkr7eJ
LvcOA497bCB4RjXl+w7UzJ70qVmVIn+J/4PLoqXEdLM82UDLpZidt49Q3TnpkpGfZVoJN9B2MoNH
Frl0uXauc6OOBHUClE3XV0p1jOw6CebFLbEYGeLKiSLvEB4tyvjKRVDnsqqbTO9PmqeYIv/6Cm29
nFXjnkRLXwSqww7hCrT9pu4VX+TC9AUCsbk52WqutisUFfrob5D8ymIw3L66UHL2XsUxh+q9QJHE
dvX++S9snDiAgfKLCvhMMiBQLt+QYnkGeSF0BNvcWHpaL5XiDHJ69FiKRjdPXJMht8mYrNsSKIyB
hwdMmkG33zirCR8zx+EpEX8bk0HAKRmk+gkbh+nz3LOLSqdjlvrhMieP+qh5Kvilbh3IDO+bluUM
QWFv/YfGS7FehDCONOokeo41dLPI7cJ07sYXiocKtlBrz9Uu8E11iEe56d6W1ftxl/ZgwhyivTpY
wh8KpHYyWjkqg9L9/yU7RCHzIiunpvpixBsI3bHw+go2I5O4M2uWsV7TBJ+0ysTFFplb1THpwh5M
9QRmKAw39S0bB0h+OnJ3uqFPwjZdIAz/xACeQOcBaC2Q/IDwAfUcn45d052B/buZ70zrEBDYB8NP
awGg50kWYNkY+YXGyXyCzJVXIfC2/CFTOHal5wb2W94ZXcH0LusEDZ9QJswy4u9iYvf4pfEfP4Wt
Z+VnedoqLXxhKFrimaVdI908wneqnkPvN0H6rH1XXqbg1kXGqcuuKlQeTBYIHvSxCCVH39WnmfFC
ifQWVdgYShZgnSlVtcz7Sh06aZocz5OfbQ91FlT1lnOuP59hdfkHMsuOomr44OL2pdF10xS9+BW3
H8PAv4Ewhp2yCxps8sTA3l8KLtP9S2puNn6gQy4dwCBPlALZlP0++ljxzWaAKn/Bjh4VLyeOtDzB
7/zin9Z8ulHewNhVKJ/lhVYKj0b4jw4bepzg6lKe8lF9fRYqR6a5Iq3dmIVgWHMxhEe6T+3Bn/GT
hJuXKXdMh/76mCeiJFcVLz4SCX/IJzBIuWqU9ggPkMn/mii1S7xz+8ACPJX5eQJEAXO7AR/2TCNp
bg9ZiSqam7wf7lQcbIytebB6RzB6+J1YwGo67vuKMgR1chlr7edWY3nNBP1teT8j2Mr/n7q2fTDf
9fqlPyFDJ1H+lqUWQ3Sm5dwjs7IHHUnbgw54+4rOB/nyzHnoPKhqPvJjfCUS0DLb3SH1Rp6BOMV0
+vb1Mk9L60oGXVteeZESZVWmjKd+x0wY7v3VnOC/6ySLscimx2zspr/GGbh4x0vt5W870ed5bj6H
KUcULu/pGQxaUEklJOwGrcnQ1JhR9EisHoM2DsoJArPdT9/Ng8BgEv2UKcmNNXnxgsomouvtF9cz
g5nht/DKJ6VEX8C+rsGHG7GJRZD5dwkO3flPEcW9C0pEQ0e25eEpz+Bb4oW97uNogSyx4JJ0TMQ3
X3b9PKQsmSVrABkPh92TrJCf9waudaq7sLL5cbpw27KnKrRrBfPRDLyIBR5CgLNL4ItewjZKBow1
SYn9HNvaDOixqh8Ul/cWaBmDoG2N4MZADvilFSjgRyJYzeqMz5rnxuJTwg6TWXMtQJQXKGAhahg5
QwutYjsv4TXl+Jr1ORw7LI2uArpXwajVPqtX4Tc3Uxo+Vi/9FNsZ2ODPUYlLUH3XhE9SKzUuqxCA
ThSORbOH5pS2GJmzp98ZpD6A4pGJK5GrdwhfywaElga8Uk+LHVqYoH0v8XgnZxU3VJKpV/HKLxwC
gT2B6ivT/Y1hK45qGHWehB9PvZNHnKAcwJqXiz5zBFELt0yoYKPG8X19ZPwkk0v6TGmducs7AKF7
9KF1f1GVD1KrErTK0b3DjLg0c0SLRk3pFai7OjCQ/Lhm0xe09mZ2R3vzZSkVGxhNaVIF0YlgWE+F
8zWo8A7a2ePwM5/YqqppujsXZmTIVSQ0LBLo/Gc0XnXF8ZfBIati2MGYmrW6Z7x5snKJ0GZ4jSEH
OIJl7v4ZSIuvVXk7s2jJAOgYp2Wv8C7O+4FzcbfgCcscbfRg8BpnnSTEmg4gNDt531gVQIlx18Ow
J8fFrVch6mTGf/so+PWYpJ9kIsfKRB3Yv9+b2X5E+T0+rDY5Yk5MqHwjzGzY4v2ic5MrucvdWWj8
QxfoOwUNIPwSMm2T6JxuoPcg9+CP0i1I17AA0/qbKbPqjrgwOAk64HC6oAIoA1NGJwcK0lBJvK/D
wl44RFEZg+GEriL+TzZlswLZNQm6ylitqJQfl/Ul0KtQ+ZtZocwKy4ZtlPosFm/xEvBeRm45Wab4
ZC/BS2bvm2wxR5MhVaOVvDbmA9xMwpRH+ETl0WHgx/fOMvJptWWfDqQNd1dlGjYHhnsU3A3n6ZbQ
CATF+SfrStJT+9xMbHSDwZ5omDxvPsrGskZiAHmXnXzkJ6wgoOfnBUuWq161yr36F97iKObsRGUc
2KIkpSqJQxwjbHcr1Z3zz4pvH2THfycev4ifNhSY0l1HEOOMht3kXxpe+3ntkVHWrC5JLgaUy9KC
OeWEGICO1YY4xxHvk3LUY4GVjUxsUD6uT544M+pk8gEzNRtsW2R7kwweEqUSvGXJPh/Ke0b7w+A5
3OkUAvpr1haqhvljrruPDpoSBy8fURXsyuwmo23wHRffiTJgNSnDY6zvUozjUhvCVF8wr3zkHw23
5SGSYqRVU3UpyNXXmTEGjbe6Ei5cC3+XoGnJ5QNLug2VEK7Pvr75rVMdmcZona81De3/X1OASAk+
vqV8xj7LwIxl0W+pOyvIS4ekPZIIO1brpTFlrR0DM+1U96ViC3UE1Nl0JoMVGv2bB56Me8p9Lchg
XMO3bEBom/Sm3Wc=
`protect end_protected
