-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
TVcMMdaoWQaLi+W0KaHeqEgrjsIkNL39+zW8Gvri1Gd+URYKHGU056zKmZv1IsyY
iD3ijO1p5iRWlEPlYFf+wbcJZ2bqTHwblZx8QsTW6HWX1ZMGruj2i3HM9w/PeBnI
TKw3HWMA1ofpZMFCvbKRyn8s6JuT/Mpaqpc91/48Wlw=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 111846)

`protect DATA_BLOCK
ilkUKwB1Xncz58fq4iJPTdMCXZ6X3ns629cXszaKEFL5eAZgDLTd90uFglAe+kPf
qff0t7IFQjN7BBy9rEsgIp6RWr2rxnBqeH/gTO/5QFRnoaA7j1aXRf18rkVm9OfD
RZJHgTvQT+GK0ieOV3gcikizzHmBjC3KRpToCEs1I0kP72F60wDtQlSxX3TSS4ju
jSNXQDRRhWdJuyodyTb/VFQMhqU3/tvUEp7oWa7zdOfZZkVNzkd5koR1MUCg3M5F
M9UaowzrQTP+RBn+fSnWZhcIinjVbcJj008pRZJXTpvH+Bd4ZAv+XQpP2Dk/Vizn
Q0HZiv01IYwfx73fE0hcgj5NiZx0bm7R+YhTZA03I7vhwSG+u5PL6+J0CcNnvAGD
fTXvP8UH1W8RHpNEOy7SxxS8VLd5kuJKPXdtKPGDh234j7k0Rl0OXeMxayB3yToL
UMFbd1lo4/W8O5n0ajdOV2nAOwTiNU0agGnA667nU/qxihHGCcI4n/540sPBRd9R
30zOLOTZdzXHJurjTBG+EYTAlLmYOMxEPBvdk4T9pji0Scc6kbD+RjbMX/At3mhi
SjGtS7TDV2F0IyV/usGOYfCGfxVlW67Ea2oOv/WuOAaqpojVM2nySdwhwlQQhWW2
2t/YnxvSZNAk+R+tD4+kQXuuSbK4GTbadxqdKAkCC0afAznDzpDqFKZOLqtsyObn
6SG8mtkkWFeDT9tz7J3x/nDvhypWeZBRpe4n6o7SN6geskOjAzJn12CPbKREiyp2
IgGsrcph8Prn0NWTaItfd3Dt3xcYm5lvd4GW3GIQMZaacGK0AyiYWcSPK+7DcTgP
vXBqb0CDNHiVfeLN5S1EJJrXIzKKka0YLWrESylwzHWcjlilW3zHLcUZILszUZE8
NkFQlBHIq7GRChIFzF5ONGpKBdFoM6fhWPUwnIWrNY1b3pb2KUwF9ccjzcfSs2+o
EO0WvZrWn6w1/UUPeOmCeDxgC30WBSATG7vBqRSh6cTABhb9DgXckLEiV+5e+usq
Wxcuw2LlZj8Fnr3bM7IODmh5bnUduGcLJSO1982aEwmTGEwTf85ay1jePwx08rny
SToybE9sZYRjkmMaijlR+jBFxdAqIlCLpm2hseWJdwbIQvRBZseiFjURk2xaIB32
mDSbLeCa+BWaYV4HsixvpLqk5m1ut2E2B+LK7GbKAbA0ox4GUmkr6+n3MNYbw4K/
7XLfL6HhX1CnxgwQIDJbeuA9EvSL0HbNdszUus15iQ6NJxGRR5nrra+0mVGvrj8B
FEdea806r7dsQwrzzBA2AzxI76wzv+ZAheD5K6h10Xn+N3K3WNF+QwgfzvGgBQZQ
0gkP3MJ/eWIPgdBCijSD3C9Lyl4wGqDtaW+Un9/qtPZI+Rzihd60EzV/zQcopfgi
jXkIQdyg215o5s3VVVCcBpBLt4WM7LqcjBr0YgcAboa512D2ve77fimiCrCYpEwZ
UyIuysdK4c12Lgh9CjbVsG7pzwaEGmluu6tXEDnAAAaHnnMuWgOScZfTojplBl24
sx88KpczkQlHHq5xj8vtQDLzXsfFSqF4UwKA6Z5VikKCl+9Dl6YaOQfpvDpI66cu
NacdpmT5HrytJsevr7kBICvCw6dhLTlsCaGqRTuTkvoDWZc31FYKrlF4KXD6uidn
hkhnNlAP2is2BIG5J3EmRd6xKmtv9eFryePj6xdUCU1N/PyU2Ugg/Z/RvMoR+Si7
CIASsMi3akSChKr0EFcmsFStZiClMteIAKbNMOuJUdr0AS9KC8CJagM+bFhWAHoo
Yp7kzSnHVNaR0fJ1xUvQZ8rt5zhVAo7eBM8uHOo97jCDrjlRFOyrALuX3Hrk7Q26
6gRwjvirlB1TG4ll8g1EhrzUeATx5cokXEZMPeBsZ4iFDcNXBNpqa6WXEoPF4lpl
GOP/LsMHqGz9R/5oSwmvHP9YqV6ib3M1nhM1/fPlqDEwa8ZAUTxqvXU6S1bb/UNq
KxxSPEqsn9nu8jOHgp4Hz8PVMlga57TDDOISX+349ML8giusfvpWXEhj+jceTClD
eREEfRYT00pXrW9Xh28Y8zHtufttWTQ1ODbPDJXdVTjUDf1dv1SWp28yYDh3w07U
r0e5dSF2eeYJ/7uVQuzreQqV3YGBrePAUC+mem7A3o/ojJSCTVGHyOY2yA5PdF0N
ClwuzBuu+QzZ5U3LzzQJzVBqHO1m81BK5Bi58lUbknj/dswnKTc9HJDVqrEM29HR
FyKeEVEhQ1dBqup8gM/cy0tW4RFt+4rtkWQ6+WPEvLE+alfo5+ECdGLlsYujNkha
lV068JqScnIDqmyBvZs9aLsQZTUgynzVh9RHisVuZrFS08GB+HGbdyb4Vy/7PLY+
PcDJyjrfyk+a/bGS/Hg3JZnh+NFTB0cH17zJcOXlA3YG2mPS19YTOGOL5chjYjFM
LBuYt7krU11WSSbPFYSHUb9Sq2mxCJMU8i4uLlL55pXXfLm2v1n4XWsx0oNPkcO6
olz7TRueM9BwQ2k+7qNGHW472gfND/QC74XqbVi2xbumK6EONnCz6sJZq1N7b4v6
Qw/MFpxZF2b/vfvv6Jck59Z0jCivo9TCM5xwC+UCgqZw6oCxrjVl45lOqQlGuq8w
rga39jBHeEchM8NCgCKQ7A63B8CDBKNfWxYRzCKk4CqJT22hf4BXLrOL4o/DfJ4D
7V/oDEQH8i3TYVx33D/ZVsxFTBRhgfuoWwXd2+EJ1rQoVfLSJsviC9/RjZJaJA6H
qaIVjD/a43+mZdhkLsvVzDT/JfoFDnGHuoiENqKh3NiVnSGFCIHPQFw2VV4jGoN3
ATunZGajuJhlyQTPorpWnPZc0ItG4xJam4EJ+Mu7sx8wgViEigWdZJKB2qWXrhx6
c0dv92Uhx8SrXO/Fk2ehsBqznmIYJNuf0WjK28wMWeVY+hAZwAShOHMD2aDy82N1
WMtEDmGg/CLXD9hMFRjNnRy1l5Ny47QE9pC8OCUP6vwZTLyOnynzuus9donhzX8J
kjqtckCYM0GBrbM6F8b3E7vg9VZmThx3nZguQYi9PHj3xhsLDdkGatDaVQKc/BaZ
3ceCRaaMoBVIuOCmnoRkNRPesVbawqLVfPSdQhZhuEFzKNBBjmdA439t1ABWJw0w
Km2o+g3ANBEkLLwmzxoJQGdNItf+zK9r2wlxKT9f2lVWXj6uQiWM+/hFw6CcbJF8
UeqWqC5DK7DS4HQt15HNEoRGBFl34YfdiXLtaY/5OyxmrNA6ghjst0gi4lnTQAT6
bIKl9COVkFWFcA5YPTGUM7l/6PqvqOEdixZluzpGljFi1TmiLFAg8Q1jGp3mwUXp
JB5N/11/2zAQKjhuwTFWHXEYrbp9pic3frEiBhj3Zsw6WQelNkTKwi+Zp6tlr+RW
uW1cYACqVCSdhUchGfCq/YRmV3tZNmxzQ2XBCAz357XMY0JX2uysQ6wYqyhRmD07
ofW2EaAWARiCct7bnxnDcPB7eIdVVjCqDLLGspONKGprhvZCf1lhYp4NkynlxYrw
+PqCQssWTXm/RM+GiKaFUvF4+Ncb8RBcuAlyJRt113Y1HpuSSmBhNQwJ0G47hk61
xmL3mFIWN+qPYt+HDRaoF6Uhd3FfmaGvZPnC50bcx7uC2qQ04jPkrKkdWJPHS4Nw
TsZIbWRlG1ynvS+2dUmdZhnF4Un9h/tYOIC72m8T6M/uHIlg79/dgRKlztSZfC3+
/kuiYjQIEySSVXdX2JFnIbytrd27OQhE9VzIafqu19uMDRgPL+8mPdTr7KO4qB6D
Tu0OnJbXeZyJKgTU6x+6JHGmQJkPex9hRclaGKl1HNDKn69ndHqDxDPpHGoiLVsC
GPhQap0zilMemSKu5ZklSCB5JT/2OgS0nFbDkos4r/JSyyG5AylIoZJvTdR9lMpq
X15u3vl0Qhfg768GjnJSVYdoSdJVDOU5uc0Ab3Am0sOweiCanYhX9Y0a/V8L/CJ3
wnlWsq5XqBz/nVh2WlhJeloLTH1y3liSvDGJfhSYhaGES6b4ZZ/fHeMDAuvGpV4w
NKG8YBDY4YIOuIR4eNZKlWM9jOkUvILAANS91PDT95sitt9wdal3qGbNn1K49nJ0
4y9HeUHr1sFZZSOVcPrmaGXiXFvMamUVqfiE0kVjNB94E+ldeBJRH4xNjda2/HMv
561uyK77agwzGp2+pJeCj6uHfnC7uL49it+nqXGSgCg2z4rRVWDz2wXw6XJ8UE4v
n2oervKB9CuhEhXTwRliqFUIpq64raOzSEaDMjNeGSEvGsvquUgzisXUamWQ35Pl
7eZmBCeEW+jq53LWepBirG4joUg59MXJ2xpBqwUDEMuW+nPQ8JhVvObiA63KuNR1
2QHoUQrt8Owm4AQOgQj+SDb4G9TvTRcAmAhVS/TA6TvedymmGK8keUynrM0XNqJX
pGnFrOUzd82sAf8Zu8cxz24wvpXw88lbZacibZVFS3BRwuW/opCZUcHzusjbZmUr
p8idHg6hiE7UCiSh+yznh6CcUrCA1E1vT8TFko1CoGeAnvQEFbDwMP4S4ApSsrsj
Kj0rHNSfSJMSY7A9M+oEJC3GDnIpjKo/nwgfToOx1uhueRJ5ueL6CbggYkD+bn5U
VtgWmGDtIfxBfxTWBqgKvzYFwxSdnzwKdOEQKbZdH3YJ85tABz/fGbotgLZRYpdO
WK0R98CxP2Q3KffqhdRScb+NjtENfizQNsyJ2ypaDmq6ZemgHBPyxh/7cGnm5lU6
ncnn7vfTiVWS6aI72UE2FxiGWJrkZtS9oT292i1sI0N3hWg0gHueORysDAcHdvvd
iDeYuL4JobCqSBpH73d/nssY+S1bISDIAGjsuuAWJe1I4H9W1fEWp1ewXU/Ug/aT
Cw0feaRFXCITUK0tvxeRyml16JyF32mnaVBdgtklUZTKrW95VVzib8jDE2g4eMB2
c2wajJi91+IHft7gCOdaT7JFWVnz2ZAhwt1qvEb0y2c6IKjsEzdQKqeiduAfI3Bh
FAL8r8GMrj1vPqTwlnR98QiC3GmgkACPV4jORGUHus5O4LpTF6Ve+VMGGSglGqrV
EGYDEBpSdnmhRVTA8DHDzyHomFJacc9YZsyDKjwVE84tqg78QiwcnWz4AI5JUTnK
/s34LLYOTcmGjZcHOYMT6iqVtShFXsn08yNDVjKFCeU1GEsbb1IJslpmEvGfI6xP
85b6w53d5EYLE3m3ON+abLl4rFrup39Cc4p0TX79CKDMARe9PW2sboDXhhTT8Vat
FkBU1ur8gm/0dLLJI1mrGMwgeV/6x9bTR31QSFEFHe8W1R8ArBm+W9sB5JP1L/EV
TBm37OkpL9g1rpSvLI48Ly302J2bJtapauvMMArIDGrj+FS/oGERfBxlrimchPH2
kNI2uxNMCCaV/Gvy9xludP7IdtI8IPb3Yx39IKzTpWPdQoty5/6Uq5nwkUNgT3Xc
MN3IwZXPuvevrIs6jFJRgG2PDM1lzAsyMDKeJPzCbKvqL1c8FKfhCH4OMFYPHR4z
3MGlZPLNTgiZ2DNyrfrMlJUfT22cVKXXcb831U4GZGzd5WBC9aZnjoM9nGlxe+wd
CG4myU+1Qx0CkV5z+/x30nti7KT9xp/hKV8dQighF8gbxR+w3N2GhV7nVpfY3DZ2
dLdIqRqlCit27rTp1R4jWgZySrtgsUwb+aghJ4v1adA9vM17sHATEd0hfclmNc8a
vvnFmmtysvjpCkNGq4/DM0gDac8wCHibkBRcE688APo214wXjN/06QRWGVeE/D4y
s1dTOitJjenO6f0aXy9g1hqOJX7HHN/4ntJ8DiDX30qkkfX0EWSUt36TWMs6zKlJ
JYLUapKimPn9Jm3U5vKY5xhJBJGKDreKwl8Ieyao9d/f5iROWAx82tktIp1d7xKw
x3EhHSDAnXyfU9r8K/iQDQRIthlvgQBoPuVTXJ73wLue4zGrKbF0LxDPkoiL6x/f
2t9CWFdxxibuiHXukG4nIQGDMvIsZVHhoYgkHKuDvoKyXticdPMCst5tVlVVBE05
/KsCBH/BwCXbSk0nBgiG7VJRWa9ujTAqkNKq+uq1F5aDGUN1U2rTDzjiOc5cLdLP
fnxyemBYcSrpLGxHXP4lw+wkm8bNfBTErFkKgeKps/vEKKFG6GymxOjYofFs//sO
zAtw3HXjJquJS/7R3Yu5Ybil11lk11TwuTrQiO7AtvE0fqV+GjBimjZpMyavfDOJ
cd5T4Rm97LeXWLp2RlZcWvXwPZWzXY3XumtpLyyqYkhmu5b61b72Rb4xiZ3E2zht
Hh7lIY5tB4I1QV9LwzUVOnHbquNTNfhz90JNLzyOjXVF6OTBJ2JjJpGatMKzakqH
CGoQ6aEj2sTc+PHsGlIiwjr6wU6SFP+f9HFLrW0p66n8cmrXbUWOH9g4r68xddBf
eRWKOtYKtINmVUgQCIscOYh4IJxuy6zr0mOp+NuT6bm/IgCfaVCQjxUJMmxPf2D+
Gmf4O5j3qR2eHHuukhQ8y7gT4xdWqMsrO678aX7sguC/nl2SssO0w6Xp93YvmRnn
tdAE4JJu6zoABPzbvgCDuZii8dgdE5OGz9zYXI0E9dLYEKyaG6EsGARqMzhy4dMB
3qta+1SACTLdEjzjs6n8KBtI1El/FmVFBGsw7Zp0DhHnZL38dfWxb23YIOCKLZcw
jfZ6uSk4vi7K1qwx841Gj5JtvrZcMWFBcPr5eyUnnbtXGwHiZPvlCwIHmJvsmqBB
jC1NpsILdQHhj/G1aVzw+Py6r7e1Kux0Nc2/p7Id0qGXPuVu/cuJEUCLzBHBgDsQ
1cTeoeX2IkY7HTXO2f2zKCc4ar4bzyM+meXCCh0M3itPNfSp8tRENCe8FYhrrNSm
3nUr0W/oOmECh6a0//XD6LMB3n7AZDLU1GIQ+3qoY2DknuXO2m6CwKj9+x1wtR6k
zF/Ck+1AJQOnRLqjhWiH1I+jzzlqN05Z8nmn155/hPfwX98jWTb0wWdehvLkZSXM
t8WLAnI6yNGN5VUVfbwVf/N1bnMGhCjp0kxK2TxqSP9AtKsvzpyk7ABle/EgKy5U
PN9SPX3aUARo+HfX6sKfFTm5/z0lwnEtfGXectZ5sMg9mHBmxWXYaSFxUPeIL2f3
HpfK8/Z88Qf9GlUjxEWdkXCsb+DBTgezYmMqOwYuTMUyFtfSLgR77biknJMGP+8w
xnr+uT/n1xrlsDmVcCMockmq2F6cEzce95y8TN1wLLlJDlK6JsIui4tgvHFIn2xN
lxMxBGPxKsDd6736VgSETPPXdlQrftFb2Un3nJB6vO6CobfZVZDYb66hnWMdiWvM
5iGnRB33aN5ce7U3gVjGrrfEP6lfjlsAF4ll+paLZIrGfZlyLLOSz4pOvIZPiW+J
8WvN+L18jG95rx9nt4t5iiq0GxWPrwXrif6HLefzs1MnY8PzVq1P/qj0rvrQGmXn
LSqZSCWwC0ioS8y5WgmeZdpGFheb/8TE68n9S+y3+joiP+AjrysqlVlGzUFga7Uv
ihZG00GzK3UztzVyynjtHtPfv4QXOEuiBOGRydhwyCymZrGwoRIVZwV7FVNpsW1R
JuvQLzdgttJa5brgMnoliVq3FNO6N6VxEJRRXcI3XBz5R0znLwc9PiVYOA2iLbah
F/n3E0icIZLrUotxIMomDG7g2i5Qtd8YQi4bWVcB2AOwvHYyB7OIFnKnmzmDd3Ih
7ylXssl19JvrL4LpUCULgAJ8Tr80Oz04JmdUzs4NhAXkcbpC/KArZe1Ju65n6/cb
YMdqIKwcyfz6SIJaQ5VfMCdQPTp3MuSyXkKVlJzMNxQ209i3v2BTBoS1eP6g6uep
w/81nkJwrhqF8eD7gAZShez770mZifcRv3ExsNYjsfMJbG3Tr1SIjmdhy3blNrAt
tlfsbBcQN7Nci+c1O3giZgGLaSZGzYAxjMzWSxb9ghTFX1o81r14nXzTi8NfwpAP
lQaOPdQ4bQkfmkkdD2/Q/3hlryShD997WXufW4hPdAqYjrevb5V1KykjRi3sS7wR
BID+fjkf0uYeNUYfjGC+2zbrzAMWWTTO3thTlH9lhwWZfiKF+NphC07joxbppvnd
ugspKKRCeVm/i8xdZcpHnkmjFFd7pIaq48NMWjwa5iWiXuzoJOduTh4+OUYYTUAy
yoCB1QvxZlrEQIJv7Uf/hthiOWto2qLt88kUx5SWX8Pg0cTX7BxV2TDARE0YA7bn
ymzDthxOkVMaycdmPY6qsr2gsYPRh0ODqwWHGRMNS/HIUpegbJ0lU+gsTBSP0sAJ
btaHX4rjnT9/+Yx17NUDdDAlSiMCjQ9UCqMOrphO/Iyud4i4dC97cxfnXkX/eURZ
pibA35oaWTWDMIwVa/WrKzox9GTAJTBPUdkL9Go6Dk/GHdLNE5TFxsHuXYEsDU0z
Tg1ezyfRQhQV72SpNH6lyxzRL2prl7W6tTYuMb9CvB+IzlUMLzvUO33Lsj4qNSDX
Va1nHr78aN8ey061GYNmoAlyVb77iBCL6ObuSNcepCHe3gAz5fy9gI9802jlHc1/
/3+TvTsrGGJ4GJjA9AlPCsJqhxfpsExRwCiMqH0bmkinAIs4wES5gZWnQSjwT35R
mRgBpXPy/iKKnj+kJYHOMxnnuXelGTkjWUkHGywDhZ93efsbx5toUKTI2P0kFVoC
dB7+Cz9oY+jGurXOGIbNhazI1N+0zHghcW7ocCYeNMmqAOK0xv2wcrg3RIe3Mu0T
hia2xBvhgNUvZh0xHL430FFQQxFq6ss8SPcQFa+tXRA0z7aNnOcbvdQFZZyhWNDp
VPewhFOZ0bXPThecl2o+IYnGc5bcsy7TKLY0LfVOM+z0T2FbSTRFsyW1rswBGAue
jn+O8e97eAXYZSgK/dAGv2r3mIvpsL3uu9eVYhb9VZrAkp7HcwiVKYMzd6DbcJdy
kN5aRmJKPpBx109vcQVl/O1aZZ0RRNXDDjB/lfnjCV6nBU0fVbgledwuMLKDQZ8R
PkB0X77X3edA7S6mlddAsXxObh0OFeWTqLgpIj/ZULucddHFqPKB38aA1nZwzrTv
o35XAHwjM0ck3BcyDITGLSfy7Xj3O0JRtF6DmIQ9qUONW4lR4kchfD7JNWRMIY1m
MVM4pwFsdjFqy8XO9/p8zh/lScSDpOF6CKa6LTuYSueGRTzrLMABFEclPaiDmOKr
YsLf2VM+w9IZIJlZGx7E8IUf1EzT/ckN96GMD/xwUEWmKMOfgFmAQevYeOIAUrkP
Psrcdq+srD/kKmLlpSHHTcKeqiFBXyZkL9VCUgPhPCdKI1826CLXKqmh+G2Zgev0
dq1CTnCnBx0/KPGYgvCflX/81LRuuCqceBCTwDG3k1V+Lv2a4jngLV6yIPoxFG6f
FwVgH0ENVmhUb8Y8p5wf3T0HzM/oErPU+P+JdL87SPn00X9LvRtWDEgnNhEfVACM
rOuDn+WMtXXznp4k+ubiEttcZfeMI3TjzwCkKhDBIa9lidTZuBZtJR2aTnEN/K3t
BV3C62GyqalJ9hrpMRrRe/ivPvNAVdeMFynbRhlBUClNlSAT75ljNe/rT2K1hys7
lB/Bepun53k5WeXcIzZyBdem65HWUwEJlONHOGjjhTrag+sQ4I1dNIJjFrr2rIl5
dGqJYl1SKbtSuCtD6pTf0ojrL9Ptg3BcAPN+KheYWTYvjjhfMyS8nEkYnETasxcR
HgvNAoTo6X7yLkhrqFtIIauHSrHgjSma+B9WTvzI22TXKGBNMRg40EVRZlh8Pydd
X7AEX0GTUW07x/ityD+ZG0oW/LghldcxpZtmvbtY26U1x83Ne+66lyy9bnsb3SUh
Y/FW5ymb3vfPb94c32XHs6ak8x7skPHR61YbqV59Q+UoNC1EErmwGSaQ+CH1jpt+
NTvaDRMKzcqMm9HqOCrba6t9ZSmRKyFQ12MZVaXzQvZ0kFfl1ocTGX4K3xde0PuL
0g6t0UQh1711OvDSdrQANy35oyBttMJ07XtNJTxqZd6IVedbEEpJQulUjaRvMAn6
Gj7opj0ZCHZWP63uvg6KkBaWYqG3bCuqM9oz7VsTOYp43N6i5ZEdlbZa6arLQONk
EIpB3x28QFXXPoOpiuEKmJ4xNdAqReBDnFx2Xq5tiT+/hS51IVfWiMhP9drJndVa
3BSOZ7lW51HxgsmJwUtZf7arpvZbsE/Byp59jjDodL6reuNUS5MXU9QDHAQepASz
Ybfi3TxQKL2G4fI/CLYZvX4Aj8FZZWm/CeNZhtK4uzdkC/N5FbjuRluASSzgfSUU
DR7SjnZBnlbcCH2VUi85+IVJ3AGEP+lLzKgbeThJ8wasBw0uLIOJo4hoZxrBtfY9
nYZc1eGSWGpZ50IbBqROmk8QVriBIbxYXl9d4XKhgn06mxOqqUSZV2AY31ncCy3B
SF4Wi0EiYucctyqa46+r3M+gHyx9ewcVef9FMpEYzKA7DAA2AlH18DG/X8XLHcMa
/OJBwa5RQPc3f0MAesJyqo23SImLeU2ag8aJashF5RS68sj7txSC+FGxuYPburS1
w/949/uZLYxy3b7K5vnX9O5LzVbNYGfIQlt6lkZg3R4IHKnQJ+px1470qduOGCW5
BJhIYUoiKvHrETSlSpy1WF/gos8UmfQvU667+hxjZrGabT+CAwBON21DCGVyrpSn
+/0fkYDjbSV6iuJYkjaJ80SCNQgQn6Wf9nmLsxfPGf8hvrVdPIVt0h/+rtnXPtXV
s0pd21Wg9UVjIdSCOPbBFu2pQq83aWndEIfeh5u3WkY+uJHWRE5HXH4mBKxJwJB3
rmZmhxSs0rMA63paREP1pVse6bAO9MTKmso4iX1WFjFEriWKxn88z/4dM8ux2lvk
w6K4U6w6+dqnPJVkqViDA60DTmojN1Xc2XspHuwJEDlhTPPA0ZnqCNfpMP+AlOv2
F9I6CiMJIQqhBtQmpO39KRp96ckKMzlEVr9qiNUCtdktVSf0b0i+H2Bq+rLHV6s5
J0b7I8dlMq33C/joj2RmJFAgkagWb6lGzHGDzZegF8AxJmX28B71ASFyJtV7kU11
aqlJfN/C+r7rq/A2qIs2+p4bVPCa1TbHqrqFMR7JBPegAp5TXTMOGKTc1Cbv5wpY
xlNgwGzb24aVHF1YSPCwUiRWePSCp9/BVcIv2r7LbSQdDnYH7a2KW6N7HPdSFy72
Rh4WW1TeCT4Lpqkg47ODcaNte5k94BgCxEUDTWm+K4/xRKiYgzwpNo4bT+HZj2TQ
O+dw0goBpxdBpe95N7HTl4kHoiuzhGIM0sGgLdoPhpu+f+muRryYmMcWkcsiu7R6
/0gOwtT9xZ8irp4PG3mFow22R9QuKjrWo8NtODlD4zF2a4PJINrjtOnlgxah96H5
b72wmaN/1DGfABVXQgBsGr17CMxEWsaQ5kvLcFOBCS7845olxC7zMGJLRwLe8hee
ifG5u6y0I++W3Xx+L0B1hvS8fcWnWUp8x05wMCCyC6LRYbhYxxMgtBeh5UITgEWD
zyVtQg+73I12iw6kG815cQAlx3VxnU62vKnXBe6ayfOCLaKvf3Vr8RZV8HRZ7Jnb
meHZD8hv+booh5A1jW+hEHcGB9CsQijf+mGBBiLrVKkgOiLyXxV4vPlGofsnFYfm
OWNb8Hz01fESYh8lYw66iyMuFUPsfnxNL+EjL22ouW48DfK3F8ppI2CQ1KcYMNF5
TrjFuBPjM0hyQJiEtEoDaC1LCjzHa/ysrntK20899uwhUEZ/drXyBShesDqo21Lb
BcYYQMNTBvrUga0+o0pyLR3Lb1VHZ7SRMezQowJta4sJ3/2HRaSDlzQScqLpInGA
NdshM0jdhJzalxRGIIyG+qip1xiGej9FJjlS61JLnbjSx14cFD1JGg1HxaCVd5Qg
2BrgAF+ezUmzoLKPLylyMV66uClSLYpsIDNCw+s125VqlmYrzfsM1IweoSVThOQf
XeOqwnEQWeV2oScbloLtjU4A4z++FHC1yV1kYWugdfsUUKK4b34Z4YemwC28/hZ3
kW5daCjrpYl/BPrwygi8uxzNBc5Z1wbIGwwTnKbQEXBdczB4k5tngrIeutaCY14H
LllH/blhUKYOBBoIjnmyKJEKtihMFPoO8Gp1aYbjPK/d/AknmNIWIfVgwWLfBFWB
WmmIUCipriqd03SzJsXvxR1XOIGq9WQ6PNyZlhm4SKFy7IR43HC0QPNZ0a2nzTuO
TukCnAlUym9eK9bRej/znlwQD6U/97+HsvSHbtTv0rWkF6Y4pVvhbtXGFiHWwFn3
n6aVYfwi21TkAhMZKFHBQqX94dfcIDDen/q+2cKffpnUlH72QN+xIP1qNZ79FH29
zk2AYpr9qIYrn53Gxa16og59fsTGnOvO7LyZzHRschDdKEFiiNbzKC/JuoOiKLIH
wQf3IHjsf2smY9cjmyWzgImQAizjqcK9/IlM04HPiqMwstDFR5I8HtO4TG+OZHP7
ISVN3wV+p9XU5w3EkKWgrvVN7Z2oQ79AAYgrFiB5RGQ/fBCJ+8spzXj3+rQN6Qd0
iVabyrinqs8fhpj9kRtvAduZ5smn5zN7lqtA7JDfYhj/M25dVXUF7Z5+Ob8FGDg0
pdzOVW431CfSceqBsSSlDlLP/y0haGMrYeDdw2ByO3aQ6g0qSWW5FcKQie930gJD
uoOPEEYutakSXurouMiKvXzsQdUgEf+SDvG5pX9aJ5YkpvDipEqSyjp1yPiWZlpk
KaBM5zz9m8WdHnihRw9t/dl/tgyqfrj7Wy2GQi1IhZpwiGTwTfKNh4D9O5fQVpTc
xuFd3bndpuL8PlU9dBeB9HkNRuNkscSnzPj95d++BxqVaRLzOdVxAImWs6Sgyktd
6m/jo25wq21wBxUaPVvJeiZDwnd/bfwBYibaznqtgBVGKhjugXomEerhgivjvnv1
Cwo+DyFWPHEgW+0ur34kTvRproNYAUTjKZ0ba2rUsAEhJnu+hHFZBKArizzgddI2
3LqAUhI8D0AeBRzb0+dwkYeM8giJvcxxt/VUx32TAeoHzcnSH9KiHZeufTHuPrON
g1GkaG7LldwOqR/Z77TQdBXF8dLQg923BsDoTzqf5sgTzPqZm5P92v8If32lbUTY
OVxUusXjh4nnfC6gV3fZioBL6+85kbu6qMEO+ErxfSbp3oODNe6jMcIEOLPu3Goe
ukt+jgH4uo8vpz6mksTnOToDSH0EI1mNdajeRnYviv4oUedcJEQpUvQyEQOB+FSh
2s2nWayu4fG6vRBleJgcsOH1kGuauHmNm/AH34hMniliBHEgJrSBbRPQ05M/pkaa
yyeAIkgLXz09adZX7uVpO1WNIZoeKkXQw1vMuYifqAOTXEZGXrx0UPnGnWKYOL30
rh/367MBmGVpIajRWfwmpW0wnYZg0W3/znGWXnjtfmjwk6UWOPy3C9ulhRuT3knL
uRIg+fkLSu9ei80XGplINnJH+C1TN9vPlOMUvxS549ovdKSkMESpz5pBxOsY+63J
R5zps2FCPjQxlwypNVUKKYj9aDPwgg0vIWeLW1nKnq+dF3SLXN2ciIRN+4JLhHdk
riFQmJjcBehPM8ZEVupICKm2/l4GS1uEhk0qvYsJ85p12SekUPypv1tKP2qOBFN8
YhTpxVXzxosAOlS+ImIgsamIS2tJYuwh9FyYxpfHQ0Hy3Uw8Rr+KVz26T5Fw6Hh+
pAjHU8+vYANm78cvVHTVcle6uQY+SY+P1ZnVP/1Dc72S0+xG8q9Fa0RM/Gah0Ldj
TTpt+CVcKO/1/qSjO5yPx2I8XgPyUmy4Ydm1JgnXrjkqOBWWTyTjs741CMlxS517
YHQyu8roy0db/Pt4dB7h5qminGyyTfshKw9zyL/rr3F/mUGGK4vUcYe26sePyoWR
/97dgwdLrdWyMvix4fCjaNRvquz6N3lbrcH/AGdgZCrDg/DwFnvouw5dOMAmaGgk
RzqUBuvVh+Nz2pbPavhQJ2Yq2YEmobogGsdn4TBz+L1KOJWvOyavhrDabASadyas
ZHdqkgz3LtcEaojnuW+e4JPtBnT3AtWHY135oGcRdAMCwJvee2iyEHa+sI0QhnTB
odrq5lRJro8GzUwiQuMh5912gYsB2Xv0XpjcoA2UMxey7gHQEj9KVNjaRZ3PRmE8
YyYF9isTP5OXHNpPLab+Fn7F19WVns8XZbTQ77oXPEkSGRlESIPn2V5ko0lChjJD
7x4ugoqfrRKthisEpoWWVNeIAPAbxy/Ejb0wEx6PaNwSJng5G2SQ8I4YwQ/ZddEv
nHn5/FYk7h03zd32UFkF/g7Q+/UFHiDaZ86LUY74v/5/W/IUVN5eJum/oS81u2X3
KAsBcnFt6Zoo/oJkVVBjc5LBVec42YKFEKauuOLeozii9oKZ1J7NkZrc2JbTfR7r
mvv6z4dJi7qpXwlNXmqyER8SCoFEGUcrCPh6gJDMBD1pBsOrR+jLIJtcH76FKoqw
tkgzsKIaCxi3vaz+CZhdD2OSrhJc0L4qQ+SZxkg2o7aeXcUJM5MynRlY18N2wD+g
mUpprpjM73o45u4padpj3bbYr9rjrsWwZUSirU8bZR3KrKOxfgw+kfOIf7vfqVX+
h0bIjyJuejCXm1BdrEgWYrOQIoxgaLNy1iFMG6y1wAxUnVAtXLpjmIOFpoa/ZBJR
27J/p5VHiojsLA3HyVdR1x/t9jPchhcp4au1A4CTZthE9vmc4xquQAaztMTY5lTk
QIFNxhhveJdlt4M4wiz0eD53IST9J3MNBhUrsPWaVU+J9MDpl0SXHszWPNuZBpzj
H8iNmYD2eiwIpsFScjHwqKRyvBcJljK7yRpE+GNiZky2Jah7pYNWBsBH2e0oiNTS
ghpvp2H0We7sUVTTEMY1RZ3L2UkwKnNYSSlr4bFAYbtDhipznvvpx4+A3O8aPFr8
BgS8pn6pr7fqzSkanU+EdmvWXgtsgR+cWqrwV3LDS0IkGbvg5PfsQw8pYDKSvR0q
ZIFlq+A4ZOeI0WOsbwUCw0mRT2rhqdn+Xgl9yWrngKvL6Oub6LDPiNtghscz7AEt
IJy4eeVufeIvypk/PlWY3PwNSX+S+Gf744xB1/Lorwnutt1Uaiody3vOl70eu81U
3gqwGfcgdmItzJFHZXumtt4NjruEbZWgRQKjx7o2aEi703jH24VimxaUODNSN06o
Yf7RZnvHKZviVAsyy2OJWSXxhzva6DNEWf8aGQWTcIr7Tz2ceDpJbKxuvDwwtUWv
UNti62zxBlPb9SsNVKQrJ8cQLel5I/3WUG3/3kQwr48pLH5ea7Kb1N7p5zxprN1a
X2bYhhn1LTp0O+tUHhsywrx5mJSwdsNQ4xtZult7rZS1+EW93FBL+7AUJDWh2/76
MNdYxWsb1N0QFyxATOXvtfIB7S/u1mfxh6dhqxJgPimz8Crztnns+suzgk0eY5/z
FKmGW9jSpnI4gcLsHw0/lAVQP9WYD0u83PUDebOSt1aWfc+2LjkzivbcJLjEymqP
isyt4zQBmE34qjTJJ/v5b/tnH1FWKB+DPOp0RySIIUGnLv3iYfr/1m/irsCVGpZR
KgMICu3bAt8MMILKAhh6E5qvL46smIgIvGpHD4dYdclYbRpN67haZgFnZMI138wz
QrusgkL1c0G5ZWp67/AJwFi0LZPuAbJ20nNXeAZmWmipzrA1RxLt6ZEgDf3PKYdk
uIUtcggjI/tZAL7PHZXWZpSEG7xe3/cnYNtNXvnukJ0UklQpvS9xRB+Nwstnjncn
ogVWJk7D2EZsqwlNo+9V4FDMRtgCxRr9taknHSY+It4JYR4w4ZZqpXO0gz/DJDSI
TNVaURT0f1o/uNFmlVuBdPymudov6PH8YaiIvOeograiCctzIeUl0yAE6Tczws/p
HTW9U1ZMBAmDvWqkWNFDHKVQAhPdGEcIe2dLg4ihl+RM4za9wa5wnE/LBbCgbATR
TAJLADPvmoMuwbzVsVLNaD2A6bJG4ah/sWizhRaPCYgoQRL5DQ+o+2M5ZJAsNSXN
LrundCiCzG3fSC/zNkK3IQp9HzwUG1ln/pW3KZ06mo4tXeXkg36EdxRdCut0yuUS
3IMaD61FKyDZ4j/EwSPvrfSOvHrdIhitbu+FWSQMnVSkoyzOvzQiiTQsIhdCOYta
RY0/c1BYazWfXRNGin7EuTYRrqNtP1d+En2SHLAQH33KoOfxfZCO7XiB7/+U9ug8
48XIjk2dN9/jl+Oon2pJvd4e4kP4a9pW8MJgU4796ASM3OpdyOuk27oeb8eVrzbd
TaqW1VIief1yXi+PujrTnSVybOqnKqwxXHavOzYN4ru/oS8TThN04FtkcA9RjUmN
/ZeVBLCSKukvGsPVfaxwkNNrcLjPttZ25qJ0TXrU7k6Y0760BJBUwZ/5Kv55xwyx
Am4FEmOH8mW+pMr47mBXSi1eX8sjPGEs7J0mncD7tLtayzVZeeRmfJCMNxX7so4V
4AhQl+5qg4CpF/an7FDJM1v58s7mi8EnPtBsg/XACIAmRXvLdBnMUxQNrRuvg7zd
yJuXPzcE4Q5JtNbJ5EOsL1b7kO7glljt8PhfEEuEq7pAA23Ary5qlXdUXTbziK9F
C25tPgCUcdvTza98KfgLJ9yQSfJKZ1aS/mCrNyfCo2EILaJUJ94yUbHjAGRV+uYF
0ELesgwbGv06oBIwwI80L9gjLto5jAM+LOHEc/Bk8G7omu57Wp1OGLokWiZPdnqB
dOAa8OtP8cv4tp+UuyaKUSYPDy+xsEaq+z1SHI5CT/R2q9P8dJGR+lCKZSFQs+ac
TjG3+pAQfW2JxSBhEhuK5LVEIsQRsrd2fKs24nSH5lFfIy+WA5dRooFdDFu62A1T
IQWPjMavNuOWXNKcThTD+bbCgW2qVR5jMAS/BBUM/Yw9zXuKEn41C9IhIruhQ7u5
S/aRvR1GxbB5ZLK3VcFs6ViCfd999oLvkeZQUR5ZWQHUenIMTSSdRfNg7fTwApsD
8JqPWuPC/JjeLI0sMbf0RxdmdKeVTjufk2/koCtIkBAQChEoaP5D82t7h9ze/fPh
UwxaJw0rwsLqsIk6ueBAgCmsT28Q6BFEoeJ1wCBFOHds1kjnK2f83X0G2KreYJc6
qwpSNx2vp2oEAsuTVwvmSbsdWbtCwpY/g12x6MT6AYhcxHMwMhCdbkTH+Mh+j/Vr
dDu0GepGSksSxnvPdto/lqOaDwymEZA1m2FsTIy2A8KOUBMhuoWtFvBW3o8haF6i
DN3HZT2+/hVuZIOvRfKLgekYgZbIQ4oy8FosEUJwdoENTonjHXJf7sJRtLXio2Ow
jwV7dZOZ8W4TfXAv9kct/XF9PsOuUTijZc2uOEV2msxehxBhU9P9OgCRPzJlp3S7
extVOmTJy3mifD8HaRdrbX5M42OFpHVagbMdtzlwZP5RVoCEHIgMR2vsXvkA0zme
gFYiRxQraRCvxp8fKjXfVlrw76PMstmZr1UTyS5MrNw11sca8siIeC9t2KOzUN/z
3m/8OKHeZPqeO854ADfPRh2auBXYb1cgJfPl1CD0VBxWFqJ/Gfj4oiTkK4V28dHr
+3hI2YnwPoCqzYCixg5KmJUw3Q3AMQr8+ZnlDKw4mCPeyY5qmiJrlBM8XrFy84LC
swiaaPBwb707jomFiEfb8P73Gz63/jhK0lULEQfomxmd5VyPiJ1wfaxirTV36ysa
8tY07UeunziyfXriX8SdgGzGl/Yz7+9q9NNkX9h7XPATmsKLSxM0X6HZ6N1aa77D
iGzRkJuV8yM26MXlC82f56Hv7QkyKb0i65hDIqUKd1lwuO9NDovzaQSZBxbmZC2O
l9JHIn2eJP9JPnHlmABDnf2uiJWobUgqJ1pY9Rdo5CT7D+qB/3GktIUOWI1VDjmU
0dU5oriJIdMVVDjygPueP+6pSMR0/128b/Y3SOJYiuMRhODZCKEwdYZA00HNZmo1
fu+ONjix+Hh6LlFWhsU4QfaN26izFe21uPoVADdNoDwWTt7X8Yg/YAq5LYFxRatf
nf7RL125ajBMMeEQj4TszE0XS7zK1uWDeUXSCod2kdKv1OEsu+VlNPN7mNHBaYYY
6yIrVmBLC5ik6pKgYKxCScAIkAR9P5V1t4r+GEgIsY9WDcR6aDkGaWgTuWb2kKae
td6jAPVjYVYJ/TFw88vUl/w/JnUhdqroQieTGafIMUldS3dlT65LVE/oid9wjATf
9VBuMXSs6U11yqPE6VOaeiP5LM73zAQFKWUeGuRirPr/IWidvwHghmZzOxCpo/bt
Bhuutrr38/qcg5ejW2+0HZuZrO2eB/nhAzVD6oKCIN+y5tCAAm4hoBTmdJi9HcBM
XYned6IeEtMCU84oHQwrT9/3hO6N/bP9d+qQiL6mD8kYyAkfXQwXFUfxc/e2evnW
DvZDCSaEKXSoa72yae+XYC/l0/36FEsnb40soRgBTJFqKPPdCECYBYg2JofQ/PlL
5iiuXqWYlobwXbj0G7kBOijMU1YgvL6gwKLJRqqKlydLmVMttjWYPMToE/O5BSgM
GmVFfLhWLbpDRs3h6ktagYQHH7dLLt2xLZHxN75c73EshPuJhItgDhWV2TOGhaw2
4/KdUVODAhSnRGWSoa0PEiq0YUwWeiUZS7tWhIT1wd1et+NirVqpiP6/0qs6/UZa
nUbqdtAFXCdYyA+V2mAWHImsT+ifqX0aebZqGT8KKD0HnzMSXUj+DukVBJJrlKip
BXAmd0AJDm+ZLnzsm7xQllnKCxeYBXGRw+8lbyp9D5alLnFNyywgEz8rjC3e5n9r
YC27kjLTFDvGeAnWiNJtY+HHG9h05rNhG+DM6NWez808RvAB7RQ7nRwMoRCL2una
63KKWseeV4pZezfbsieGp+Rsrh9uz+lR6woJfAuwMSAtlpvtIqPvTXaZPPJrtx/1
uSSosb4/LOm5Uvux6SqNUdQGFT5xHoCiXzCCeRph6qGYUxHMUIUh3qnfetughyEC
99La162hsqgqZN4S0/W+4fwedrlvmH/ChJqJXH03t76Afmpv5x2MpozRI3rtiSqG
WeqGqgRXrSx875x6A8us9eZT1TD+YT0UEDZsC6A7uweXGvLWX9K9YUhzmBIIAkxj
02RLv09yMte/gWKGxxV8bxgYV9BqyFBcxwBq46PE6hXf0ZijiBaJB3yap0CMvD7k
0KfijGIXcQmwNotNXbLSKYLVyJE5kqIQhl8n2nOJs1CeHu5EP9SH2h1sMfrHO+8l
aHmokC33rzw7BPdKZ39QCLVtNwmpsUb0J6/PDOXfKtmdvYyGCGolip6CtcFInoVy
72HOg8i+GCQu2hP7MELCX9tjb8S210+PS598hxz3n5+LhBzQO2VV3ZYJLl9RexFY
AzrTMQ06BMXX/+pc2hwysuR+0+Wzo030RLpqvG7x5asssuxFrdit6aBT28KEbkkL
4IkziJzfS5/5/jZR/psiKKxYP0K4ApCBRelY0XyNkVOuwxqqHfzo7PrH3fkxDzK2
BNjpLHIIq7ZrWyk0nQ1YmPSKL0XMgS3GwfEV0524ft2oravoE0f9FXhnnZGYlt4N
JzdObTHV0rTyTOI4GbCxwE1WY6ppF/B55A0CiM5PGJmoMGZRhShGD95u82Vak6qD
z7RfRfGBL8I7VoIAyr6AyyaYwOzOf0J8n3asMNDtaUZvf/aoxLV7CI0roN3x16kO
b9iz+/ZDOq+D/gvSPfnqLOQW/5Vebo1KMjexx4xSurdXUAFCVKlstO0LZJeaUjef
DyvQCg8176rdUkkj3ByHcQInFDv4+RxrCBTpvcH2113J9mN3SEQYE2yg6qJbNGnL
GiE0ezLcMfZeoBhe2h9l0CY+zDhMnQzHOTSWhQXHUj60zvZjLG+7k4ybwn2GT6fT
gIxML/77/vOKvA9uP5XYj8sM9KEE4KNy559wntPYPVpK17aTlvz8UxT3M+lWd3az
IDVkgYvtcXOXbzUf8LegbfKCgy63kefHr9F2bx8yI9Vc/vgLArYuO7iL1WCc2hqk
k12b4BPaNaQyjUPoKNiWaxuoUO3HkS8DJ4pYuEo0YvEnJqaBuw1Pn4dYaZNMjJ7W
RqoSA1+kXh4JixJly/1ORemxTDQSTvqb2STb4EGjw/EwDmk4obJkMnF/5bmfprnx
KVv9UohjmKJenaqQyiqPkxqe9DRozE6lvC31BvNPgMqa1+GQHLdosKvsy3/mgmrk
VA3FERk+tEA3/xDAW1xfbJJ8QE7nxnff/2OB9xWa1sdCtsRewDIxo6yKy5hzDfIT
bHFIC2w9EmM6vmRzDsq6cAYAcxyFnwE77HqhhRxeFVyeMDUahU860WFLOpX4lvSi
MNTbJCBB2QXW6Ukz6FUsG3cseZdR9JZOYJYyvFUJHRUhGRlqx5WZ6s744sRUC9E6
o75h6uG8wK4D/dQJ8cvWu6Xa9Xm57CZ0M5rCgLL/NsnwtdDa9pocr8/u4u9ROlQO
k1RXGQYvYIaZsPJd2/yR7LqK9nccWf3c3jJ2Ci25wxo2tf6v1FPxFUz+bCeTMVbQ
d/9do7HLB2k+g5VgL+SA8k2e1iukqP+or1jLaG93WvPnNPAbDHaNhyBn3t/8eXO3
LGZCX8cCx3MSythnUFu/TWzkjOSJ9F+hk+tO3zm7sFMq9vixD00P1XD0E2T4d4oK
Hzxd5satmMkZWRBnXLn6+ojfapF5/HFS2f6y/6wWVT8962sP1DzdhJZWieu/E+nU
a6BE8ATFoIf38dyaRkydP+Awi1ku3VoUSeIUU+hqV1BvyP9qRPHc7PbrucKGIFo3
Ms72/isR8hfvMZcLvC3d/87CiXZ2wW6r5I3A16Ebs/JyAWwK9dDzOz38jGK5TM6N
Smd6/F0VR8jfeL+mxjkoMprGRbo+r7LCbzq8VyHjmnSJIiQnQofMni++dAEubnce
/VrHCEX4htVa6C/7e894uS9QG2vPd4HHGvJJNPAiSwi4xqOEK0XIZuMlgIflMKcB
+dlfTKs+x3b4nGaK+YxqGFh8eMeUdhcbdPCmSRfPRGRIe8lM0usNGSiGh4sVr3Da
RDRNVN+rVF3AkT2O6iZi6140IuUYorOQB3T7M3wAdaLyLw/PMxZgwPPHw8ky5IF9
6S3fMQtjB262Pj57hd3gdwY4KsWe/48oJ6Sgx8sNtriKdv3KSrM4g4WR6MftSfpx
ttlZztBb6S7xyplUgebzyA54U8NiWhULOSQMHXNUVS1astwgKzsohmPthhPIzqHy
l122oCNz+1myvH2O5cowM4gaWe6igcRSurdqAx7ug08IMmFRzRISONo74e7va5aJ
2VKD8f4hZZxeTW20HnawsfkBt7QhKqYELGZzyLlk6Oa24XA1tGjSnGQqfK8Ss48V
zZ16lYjhVP4iNrxP14yONn3VCcXbiJkXwLzBpUrndKoo0HDDgtHtgB0r3Z/CX2Ch
aDyhhHhxOiGF5CSqSKaX5lS1PNc26m6IWTwdbG097UTD4u6UNsYE8MiTAAekTMHf
/T9eXFN8rWSC4Q2iEuWlwd7viURVSAz3ZvWb114K90L3VSqvrYw2RF8MovVdmZ7T
cKsNhgJoWz4OYTKvDouT4VsG7WtFawvp13GTDbvhUJTzf3l5h8yGCPqCOR8DCns+
R5ZDbxyXGX3Bsn9LTFoqvh6f6BpdWrk2SKfR/FcdSt2GSZ/r+z0W4otYwGF1mbHs
ORGF3GGlaaGASEbX/ck1tsqPt6y/RlsHePoXItu/Qzgv2nTMKkLYD6r1MlD3eCtD
E8O3o4W7dTszaDFeF5gP99cE5HfvK6ADhTifMJS9sKefMqR1zzv7q6k/BkR8eE4v
SggB4E85WgxPdfj9M402DuxDhBgc7JBqCKyjaaH/7Pqqk3H8JHYeUFOmvPPurAsx
r6rBP9T1WM3VfTTyej63uHXfR/X0G0tzKSNFPM1FSU1HAcsVeLOPJnJTLri5UFPC
FDbq/Y5cl5p3kK3riswyUSnng7G+qY1yRHHee+KA0tOgNtOED/JqVADJFJ+lfqrH
Qh/DrkgQHaRAfXexPjdKMM7aieZKxtATwcI5G9NgpdZC18uWyGqMjAq/+Ue5hexA
uZsCr8qta9ojTq9ZB9Y+wcmmM8SqAsT3I982omhsczdNZzzF6caTokAqU1rRnF+y
WMdUu05jZIWPO9WBceM6pHMEiBqv3t0N+sqUb2L422u4C7j+EjICC3yNbvxcAuOS
XsZKdntGJ8GS1dOsqQ9PLFhWhCHwn4vtit6HBQNap8tMyiG/tArT42wgUF+9q6+j
dsNZ5RePnZrlO+rAeahIdY2OUs2nY3hOMxo+gmBqDrgpj4pKqd7ZEXsOl020f52v
ecW+Mv9QHtgSQ+Dq5WJtPB0JUvbqvK7hD7VV9NRVYIfNXjOF5gsaq87n4OMQ6Lfk
jgRg9ySpc7IpAGJwomRdaUhw2D4fceTthcSSlWkouUe9/o4HYe9VMn8hk/RHiYOl
c3cYJIwI5Jg2dBnzT7yw/VzxFFoSWWCIZpqLMDkcBvnjToEr01+eayo4RTteYTGY
Ts0Z9iGOJYzKv3TDQA7pXlHu9WSdBvsyN2WyhAjluPsUA0YBYYvtPeK1+y3fI/Z0
4Od8zpcALhMLtqkeAYohkHXrdFi2Xa/vBUKz0Yjd8QcPNvoretn3uijq1ns75w5l
r+MxzPYPiE0jZtN2WxdN+8WTNcSEVLZV29Cd2ujPS2PNF33YJPi0gl6lmem+H1pO
pxoCZhHUj77vQ4nu6K+B6TykVEZ2QrhOwLhjcL4droZA6AiaWlz5XpD8RjyiwthE
XyGXefh98qCsuImOAoNWMqasNDBC3BzTwUie6smf2QdDfagrDrMvMpTY6WQOOszi
TOZJ45HJeDpVcCF4jr4C2rh5ABZufe8LEBxTdM5wy8ZZ8vpqFV/aF6Lj3NW5mpRY
djDJX7V/gCOhDgHYnCZO/IKgEgGXBb2kJQ+jocaGHxBMmbOWdzCVsBROx3xtTXPc
e2foGLJ3z/MsgRYUos7zW/TJQnGZ8QKzho4LIg0clNJPTyuIK0GAR1clx4lcI1EX
hXyC7YOCIKwWGLikemwUmFNNdHokELCP6bFBr4y2RUzrTN+jFT9HKM3rAUHAUTao
ZgzWROpALXtIKcU3KE3Czh6D7aZntVQuP5Z2pY+RyikSs45+/o979veGps87hPf1
qpVpNsvlxcxs/DfyCmPJ9IjY/fCp4prDk4gTn6dyCJY+lja7PdHaTm/6jz4XeOSg
BftqUT9US/wPWLmTxODv7nJjL3C3FTTFa5z1+Vmb14peQkzfUK0YuZQiF9Ao/WJv
keYYd92WqgI1/CptUjPdluAEBx2PUOOiZFsVlnnFCLA7YK+zSzsCNDrcc9k74p+u
IA66pJeu2D+G9a00tB5lFnmN9JJxMEtUWGkGNWP/ItdQkT9vjXJdZ/XZfq8ebAgn
erHathSI8CZDObnZBvR6xYWqmprFHH9EziBL+x1imGIn8z8w9wPHc4Oi2z3xjgMS
5iBUI+3Ch00BqlULeJTPoBDo33R/dEKg5berkR+dBK6jNMXaZCZPMLC7Sb5QL0/R
dK4+v9BYg8dDo50CgO8D1QSsvnyU8QLYCVH8bbPHqY3LBK2YgYHXy28xitZvKGb0
3NITpJXM9VXlS4Og5+QTFxIuoaIxsY9ou/o5DBS/RHuDKc+42vlAzJEijDRBBZkd
AwOa+EMFiyjW4YwyOzPkbHp/WLTithCaEJs6TrUpVSFE5yLxyB9IJY+uLzUd6edh
cpCOVbQy9vHMMaeuAP1OFTyMp3o10Z/eDT3t8SRx9i90pJfb8J5bgtfg6ELYlg8P
3Zg+2Qd0tqK24PHFEk6X/U68oSn1JDlo6/bkYKiLy3pLixg2+XwgCSctXKigqh31
NDVzWuOxQhIZbqO3NgZt7FeGbwsyTIfPgaW7Re+/iwBuY5NcYNGNOPIQJnjtIB6t
MyOUwoTKRhUcwAhzOAVDgwVyjxmF+2OtrtuVTn7XxzE+9AAXePoXXWXKYZg3abQA
MSwNBDfcYTMmPviRuyPtDLokJ3/QG5AyfHTKvOQ8gs9E7m5t2fXJdnPcxQ+ijZRN
xiMgJNqpXZUw8B0h5kQrXl1ETt29EW6pOyH/VxDCb/VveM7agNMlO+OJVp6SJJD+
yiNgpPZpXBwL+sY4GdyvjZZTa01Z9SsawVTHzrRswOY9BrltrJ+B2IBr3gKKqpjU
G1OxjhUUmc7qEyxB9PbbIYIOmRUO1G7LwaTRWed9G1a45I0r1KO+ytSPiu48paMV
HOfOD4A+xLqc2FP4JOJzlf0FpwiN5vtkM2XO+jLlfyWTTH44HfrPiOHb1gnyWem4
TY/nGwwZL1Fjybm4suaJ6sXBtjy1gtvti28a3//KP6dfukw2CqDKcb91EatdCP3x
UtBcVV8eG9AY2Vb/qOTb9t1kw2eK6NTJdx4ENzZNgNheA4NkXGzEoRcZ2t5NnGd5
bzqNQosrjX7gZ5nmYatL3AA0RG0qsiPwAwRbdz+Vy/mfIKZys8A+MMXDcrmHhmfk
JbdQx6aUJ0siJcLZ/+zOiuuVlrowOmqr/N26buPfGF/7O/Y6eg2VMKdBdIgcjhw2
kZ0S60xhZyxO8uA//sP0JII8L/Ldt4ywNL4kseqiN0PEegafXjvsS2fdJVoyhOWz
NQDUi6ykxKjoLRKQ+vs61wCohFJOEIRJrS+xNG8vP+SUO9t5qb9ouxw2LpUOkyOe
9y50tkhUZ6sfocTfyK6Bvr6faok9JO5DrrwNXFPaVZHlN26bL37plcb29AOPgNRz
J9v4jg3bUHJT06RXfhT29EQm85POBxoT5vYNknIIn/mkoAJm9XGay7q8EWr6FOwt
PHXhnB5G6Gg9R7LduV8/Ez1u82FpW2wS9KydUJZstl01nWg6gbvM4a6wyNen6pvi
Ecarmq8O0lRYSwfsXrYNV+gRwllEf6BPhLHyyKwFydxXXosDfbPRHRl+n85lpY+f
hOMt2uwGOaeJYokh0SQswcmu8exofEDJTIYpZzPhbSlkZJOC0uxb41+m9cgWmZFz
J8RkuARePN20BhH9XLrGcDFl6gY/0GO5UIgAuKursDDd/ZhwUFEFhj4z2x43weR2
WHsaLbRVN49QYg4uerDBK0Bjb2YckUbmDLUGxszLbp1b1dDyLIe91yTi3r/utVrf
veBOM3afEf88uUnjwZ/5fC92qQAA/17PQKx0y0158ctezHoUQgW7RUuIhKZV/PWA
gU5SribwcSre/peTKcKT7WunXR8qzr+7ptZEA/lyiKK5vHtk5ND2LMK6somMAm9X
BAxENSy8tBuVtiFaYIC3q5Bh74Jb1FoBF0DonyRuZc4+z9pFd2QLS9y8v/RG0egJ
WXrYri+u4sTpM77uskO7UNQFFzJh818vKCqtpVnjYkC0WEJGBgDUlPMtaAmFivfv
bjI6JYXzD2X9wTJ+IpUvOlMuOKXGIPIV0ExjtsTxcIueI7bZukTJ0EeCrAWNDpm5
uQoKnXWfEXmc7zK0fD+FnyBVaJ+xLuETDHZSYhv9hBBlB5AmKVp6naksi6rOvNTu
UE7nuoJBLeBh8zFbNbKf458F0SEN1MnqQRQdEmFjXokQ9L5O1jL3RrK7c758dUKO
Id/kOPuUYdb2H3IUp+p3oL2bQAbY3xlp2q8CJtHnJW/zjiM9zU2CrhSe5XLUZhyh
Z0mfpQ0cOq3NBYha5sgjFpJJiJNE8jksRQfpT5De3V5y9NPhO8sCI8Fbwa1zR+ZC
s3ta9qB4YKNQ8pW5W0cUGvm472Sz0RYbV8i2K9JbmwlQwF1zvON9AZgQLum1Cx//
zBxIuWzu/SZml/IJOBYSJo9RcYvjNcAZb7Wl9rb3qJJLCqmtFOY9H8sZtj4O7SCs
JwyWNWEhGyQ+Uhz0HY6xRnLRFfbPJGKNvmGUc2CAMPS6NvRD2A8lJ8HD4dbo5kls
u0S/+59vekoXWIFT+BDfLL+XDwU7kYp4RDeSTlHTofjrJy8iEyaLUnCXJS9LVjHc
tmA//6B4vdHLSfjZvKdC78bTzS+SqOuSz8HY//kKwTG7IJWIN+6Ifca2KpuRR+32
Zecv0FMqaiG8qvlaQFUTEGhtywIY6qgNMlOP1HzXsKLFIbaDLPgRveKCjAxvV+KH
Sq2zT3PuTgZqmlG8XGAWjl9xOwBUOaL90fHO1efhA4KxTwBneZoKG2CTyEqmyDTn
cEZlQFDwrkzYtawPzRnymdk4ILwrz9ZolZtxgNswYoB1VDKpODzzcd2eroZEVnIa
INiliv22wvDkNIfn5ArJ9GPuEnecRPQyfuPLxCc7gMkAgRbr5qQwi6yRJP2GwVGA
0TmYud0gnhDHYUPPWPICJhRUH/2bVttb7xQ3C80bTyf456eIz31GAtabVS0laBiQ
wwAYPCStFi4WwKQcPeipPrWF4zojfz+WdTM8Ajw8akyIxCZLCMucwk5BcFZ4hMop
Wvh9nVCM1KTp6vw/oV+c4a+rErL8L6g/3pcgE0Z7e7hWUB2HIPJJKxLYK+MB609d
14buUwl/jOfpimnbyhQYKc7iKIJ2Mg4X2I8+/hClDdSvVgGgqn5FllPn2AdInlu4
n9IdvkZ/MVSPKNrjunxzXQvvLeoqURIvV+mz9Wh9gz79BJdK25DMdrrtosn2WMG7
+Qku72qJURMA0Nsm/U4XoOOQyXdavpWlKIbzfZD6hQWqyBTz3UiwPW49Ig5tY1va
m2jQyH+iknGZuGBV6ei8TtfQ5lo/uYMNLsxdEAYssePb7lR85bljsfYsIJ0fh0qk
sa8M8cFT0F0kXOFz1JlsrEg/FRyCDw66jsQE4UKMIFaorE+HHDaE+ssCexvOpZu8
PkE79fLJE/pXBhGxllc+RiIDhsStGu/P+KufR57fyNBj0VvfSMyWyOLZtvU6Ijg6
WVDv6WzUOis0J6tG7/9moIZ2EN5CXDcoccvQL1Sni61xzXRJeDIzLwOTa3dzD3+d
rLOf8NRhf0PoVw+xltdPlwTER9YKK9W+M7S0VZTQqBPa3oSJImJP7klftXPcmE3w
03rYEdSw4kfEHhty+a5k6z2nUFCOiC8O78aEdVix2cDlRDrqKXXnrHrMqTadd1Bn
fmYMeXQO4Pl5PiZiqCXc6a9Q3vefTMQTF5ES/afckP7k6I/TbngEwXdtcMqhKsaG
cjl2Mske4/Oc11L7EjnA+zLv8Gboqgp8tiZDxDCNsdsny3U8NKTppQNYysUdyboC
bjcgnitsf6NR0CAj9vRqw+WcshcvcLEJ1LlvNiEPPQAAIkRjDbDkuCama7LxuvzT
lilmbTnXjEbyccdOTyDsriw/jocBmpmngArFzLh2UohdpL5CYgG6vvd6hBLXjXmf
tBV8Ff78yXWq+dhwQlEdHV/aVTQxnh7e+e2V+DjvwT4PDor1F+3VWgElRmZp+Ghx
zGMeQLfaN+QQYqqiR0XRus8MDj7HUw/zoIOb88/XCDAKaQvpZmnZrSS9NPxcKOKu
/RDAAVZ7cErU8FQoD79Ww7Hik9gXEiYEpCMVyD3eyH46+bacAgjuF6S1WMYfwu9e
bf0cPMVJcqVVvsaknkLQ8OOZdfiW1F9zulRCcr4dAHdE8wmF3jBmqSMhwXAHO5Le
Lh4+nGPszM7IUJFULzaaAjhEeheFkFq+yLrXWgyEFtDNr0tuBKCGMnfDyvr4n7j8
zHhxUyJFJ+L8hivh4shqHYw5qCNnZbCj93xC7vNo9tYnvFIy/cjBmeFfbc7bozai
Pe1FYqrVkiRUeegcGonkGGXi36dm0B2h6t+PaNSdf96AC91ANvXJrj87JH/wAyfx
g+7n1QRL6q/kyrRZL12XmTXSQg3ViMFrP+a/AY4dddWj1B8TzsqfLqaYNsip1p5e
YMY/X2N/jIuXnwLjmYFNmeIBYQ7lDIehLIXFC6/TP67orPCF3Btc8PFBskTx02bm
TnC452xkB7VM5bnEc/ZN9s34SOCqF5KCScKctZ8oNhX5Uxk6NW2GAtwG0Pft4WGy
G98Uu1dJGyikc2eesrifAi3HJbdz8QxHDhJGYpsekwj5o4LQfWDOBptXsJ0ziouv
+RxUw3kiVgVeaLWcYNKrqDfwojCWjZmlJ++NnLbonY1QxRj8LQUgq2imKvDnyUTK
ARcWYr2MdLjMMWalBnyy0N5bjl//wKrDtReNWrGjfL22UspRJJK08ihHiac+ZzNd
kIH7hZV+JyF/3a1CL7mkEL+bVDvscORGEpCzVnezXLDbf3lFlAKwHd60C7eeng0J
9MonbyK+PyGCV+rQh88jKMHWu8rUcdaeO4G0NGard0Paqk+Tvn8YIBrjSE9eQWZl
pi0P291t3YR5LtlC0bTzHkmU4wZNZl/3tnFRC/UQO7W1jXw+c//h9ftgogVm7pF+
yXwRQMkauAepgB21/MgcNoVHMOXxD+xV7IyJ5mNp/StlNHKVS1+vWD7lU9b6qP2s
+uGKkbH1eFSeV54KhO0UaiywuNvCL/l8ka7glwtJ6961ofL7zTO9X7xK89yCxe9p
flouUIjiyeXqt/uVUXg4bHfT0uCiA0hDTghnypAHIJPprgWpLuc6Ai14D4LadAfg
oVUTPc+roXRyTYja+6sK35JobH6KjFZm33c3MPbL1wsR3xKyv1t9NmMum4m83bIS
RXeGiIr0A7CtfVifOOFysS0TWzi97nT2lb/WOBHWIcLJ87jRjHiD9AkrdoxmKq4t
AJQpfLMYj94oa7lgbe5ZWrhOlx9prJO7JI1dDLzTU8yYDctaEuf0BkhzFCZlgtVU
/AH3BMeflEeY07M03NNAjD/z3FYO5HzOFvFVPSmMXl2Fk/TBEL6tVrxm6cNLuBl8
av3S/oBM0BqB7mEo4KX5CN26hbKlAAeYeluXfMeDjCBw0JsHmYW4spt76p6DWmlN
Ka/KgdO1bjnwV9yvZC11uz0CmI6pIEO9AEFDuOol+Lt7siGk3HpYdeDJsiXrnJ7Z
QRvpya3jvuJ1aGXfg2YtooataJcSx7IxkRVMIvHii/hn3abdGVjtL8etShlp/3yb
Dpi0+IKvjbZ9gEI5D9yQ/MfWG9ff6j/+7lQcr8RZnA1LC7v6Kz+zzKvpj4Ic/nM0
MNJCeNSgF7H+FJx+NbTsjFUZwF/ueLu85VO/69efD1Upy6KVOi7/LYm9hQQEThlV
KnM4la6g6xYUDXxYHJPRP3mAnMiDFEfyRm399SdzBDJhrO1cmTDnsVxoJJV8f4fq
ic3XvVxWngSWtGmsFRQ1QwpzcWfpsmidGWtnu4g70kAB7dDAW0LkxvrzeCIm2le8
Ag8wscinAp/qHxA9Th/OcHhO9gAUKAhDxX/sdQufn26tT/YyupH5wvHrzOdGO2fc
0xH5AXVA1+zD8++jhxaVxexeIAXy+slXvYT9BFFZAGZx2vtzjofqtH+wy5G/4H/C
AsJ1If5zRuUg82ojYnsOo0vEUCHDcrXYCFg3efuUOV65T7vWIpzSB/kUR6O3F/dA
SWdtfsPNPur7Vi6f26LMMeUwNKRMyZKHJVHNo9s1kvEGHz9hytCVGEH2Imshbby3
thyL4fIoMbU//6Tga65a5nDk68OPxHc9IlIETr9mmKsIMfl1D5v65QCfTVCMqn+a
00ABkp5XuULorLmpaYX++BiMypSkT7dbhRbZPzLELWhQBHp21P+KoIMjzMl2xT27
l6EyVNVk4IlpczLsVxh0VReInjOpoQfmEJ62DX5oqyn+55JGB7/vtCrr4gky+aq9
EAeWjqr5H7aQZSLxmJ2nXDp5N/93Tsb/mEA30FuVmPCnC/Y1LPb5m01AKPawSVTY
wb68jFBsl0sAgVqy7nV17Mqk8C4vjkuORPzW8nLbdAyq/o2DRWeISQh/eU2Aatb4
oNDa06TymK9x4QsG6EAVEvMsz4qIgDHay0b8pmHrTbp91FW4G2V8Y1M0Ayxh+Iom
dwJ1VHJAERN+TWxRZd9lAzDFhfjCE/EoRxlCv7prMImmcJS6bK/hIcuUzpy1FPql
Nucx4is0P1qORdtS73lmtsoUVhyZZdIuoaa6c0Z1bxFEcSjwLYh4VWKiYcezn2MN
hwjHhnbxtguMbZgGENARI0nWE++1alVrtDyXzkZ7h+GlZW6UyH3vCdFcD9x6KroL
0ukNiwUJ12tOHvUgI+OhlJ0negVFvACG4kOkeQzbsHZP9sIrqC4YnEiRNcgMaSO9
SrPIWoC2eqFWLs4MIBvhF1cbR60NVUR4D1aapekfD4QFKKZRKZP8HyAKrBAzfq9t
ISzFSAs3Q5ud52Ai62q9gOPG6sqVtCNdYCEKe3P7rFNK/QZjD0FbzGIkSroIn1ej
g+df9FF/Undh2LLpQRofVePYa90h6v4x8r0P16Hk3KWHqDI0hZJJ+akv7G2IsJRB
n+5bCBkJjO5AhuMcHzhDdPLWYLlqyGqoxzY8JIkAk3RNjht3CxNiUssaKc1Zr+lk
SalaLXmScD5fqTiJumWSt1mBv2fHqLnUyUAuPszO+ajf225jcjRZGdLw3XDadOIh
vIoZ8bV6AjntDO/caKQQo3fff5x0aQc7qRAzxIgj+QS7RZj8V6DifrPO/IH069p7
dQL6C58fg1WP1ZMJ+gzecc5F+woCOFd8AaSzxGnj6cymxR9RGLtX38BXGITVuMKv
sXQsdBPReFfgOfWDYh2oufOw/oN3+tpoSgt6kFdxr/dwD7CRKYmTFTiYe0B2M4qe
UlQgozWbH85PgxlAoKXGCGdxFWM95KIWg32IOVOPB1yBn8RGPlsxZOpPvoC0R8Bi
Y4DDty0+kAS0Hmw6oh2dR5f4We3ow7v9VvfsxWBgREgposYdAm76iDw6q9vIMu+g
imd7COcgNoCzjvDT5NcNaRk9i/iUxltABMa9yLmaRvcHVDTXvMzkzMcKnoRHJr05
V6o4e8iTgyb8gA4gNc3rGRkunWKjSn+Y5own/Nb0m8TS3L6Pvahf3iNoAOGZgDVa
5fMuDRro3Y326rJy79AOb+hzjWrWc+TTno9uwky1RlmVz/010z+qLt0kO/8wQ+A0
HPmwrOd3J2L28acYHfqwTRHpRZdoJ15l9WLgvrUd/iWBB8aB6oi8T3I4hShP42JH
RzkvNetz1br6hiBSQOCvf7a/szOjJei6hrtJ8PkTkcvxaIIwgS0A/fQwhoRiYkM1
t6HCV4bx6LGAkKD4zOQ+hyw0qQ4vedSrWQwRybRtS8MaXbzEoFI9A6MFScKQ3N2Y
7y0i+FHkUVYnf8NCZPDaboyRrtMPr/e7Y7lHb6eZePU07Y4vo/KN0Jo55YOvK6iW
z2FGyFUrzqaNzPzNDnivFoW9U2rTttnayxvqlyXGb+KWulglSKsxq2ss+DFcy1NA
vU4YtmULND7FH2nTInkF+te88XiZcA05ONhUNoDvYynXUiVso5fqACuY+cpF0gyb
ISny/ZVKxtQbEYX6lP4ktzAogI6o0qdqY6P/pzR4WI0XbuOM8g2uj8ruOUCVThBj
tvuthD0ZhbPgNQgAZu2Cdy9x7SF7v6u9DjRfjJno7r1tP7W6hmH773JCkjSi1bGm
uZ1MT4AOlCjH7dQbPB4OGRY/To04895nBojT4Kfe6nJbqbcZy3Dx+YlFrYj4uV5G
81JsvCY1GyDhwFKGA2aBMKkLNVe6QuNvpzetCz7rRRIk8XNDU83FvI094Oa8wTtn
0cy1iIcNxFok7q3t1Wx1UgFeZD1WALmnAK15m7D4VFFwmbEzGrBi26/RrYdfDsCp
zp/WbetY6zsPldmYE10y3oJqW2PT9Zx4SISUgqoUbt5ILRVnu7QiILG3Fa5RuHjQ
kEMd4tobyFWhff+dfLY/+L0o1nXILelpVIipN4Cadf64Yr4yq1NHtNJwKklkSyTU
HU/FOJxh3ue/SccjCnvzovt9uMVKqfAY3fGwdalELhxsYjhuy6O/et6ajRQyTKx5
F18f/eZwdZRz0BlzbzjCDSzPy1x4m3GAgQABmljsGXbxoTcyRNJ8wkzFm46QmwY0
eNUUdLtp+ros0efOWZ8epkzEo+syGW6oBlOHY0K4F6O8SNL4q3MPugxNpMjE1805
Kn9QhBcQeZBqkfg6X30lVkDQJnBlIDuOmgx5zU+uUsRqVShrEV9egw38h83lxDz3
AK+Hw5eDPg15/vpf5/BkiLhXjHdO5kSVhQQn+DU/EHnAASAiD2SxjQUkfdeCj7uv
f1FGvdrOVNbZX7wmM+B3b8bNiBrQyPat8ErJ25s+mlEWyTUzRD916NFZomWcc6Zm
L8uH1gBN5yxNDHBvHOSAoUMgGoaeLVGi4JdvYs6tH0hmG58i1Z1zklER3eFni9L6
IVFWJlonSaPab/g8OV3qzXn5b1NNCiJj5ejUGmETa/M4bZ3pRnrkj51sDROzoMyH
S1WELL7Z4s6yAusjW1pSAZhD00fBNmQ9/Qf7xlM12yKW4x25jn2C6AMGSP6/DGi8
rJrbKEyNa1X6T82a3G709wm4FuA1sn2rqioUXAqwrIe7Ct4oEYInYS/4SdI+wMbz
RKKJKMjoSHQJt2QAqW7PUkZ8j4mg7+jM7JI5oSdVcuzcCuaWN1w4O0j1M5faThW7
IM2wVTsNBnmMYymcmV3leOF9+DDQqwzo4+pqH/jHKV+v7zAL5B+O/J1TfCSpcjhI
NLxy4huCffShufeqxa/MN6sNLiVoyakMGtnuxBoDvopCfv2F01DtT4M8Pmhg9vDW
seMbe+OOVWqt3vEeMS0wwqdC4S6rSDyWljMXLlMSuQR+6COYgOFJcWAbur/0LMaB
shXjNzdj05GiEGT+c4IpPGwgYSeJfVyhtOmhwxic0vuYHrcreJK6yKNbXt9q/3wq
w0pQBTcJ+xFf2AM2/GHEbtoHQ3rt+xXDpes+9nuWcGAWYbxzg72VgSu3DLIl09fs
dmPDdAG0Cd8L0PFd983guYoabemAvbeEiILrKulbE9UG/a+6Vhvhaxf0k7IltKvE
1AS5TOVwC4SXLJ5OAfJvCaWVSUP2FtZ29BmVSfLQrMhaJXHBfMNEohhGHzXaYVy8
7HmX9WEPCzNvRRi8Q3+/osI7eLrbphUlKocjFuHVFA/WhxCSyPdcBa0f3GI3Vwu5
fHtMnNsMptzUSSrhYQXwGh54B8an0y2ONHSxzybk7pWHxe5dUmkBI96siRsaQToS
ONKdoxvPjgd4nY4pIL6/ZChcZ/7bD9PjUZbK5zqPVLyVSv5Yzmd8MMJ9cZEbo/oB
938pSCjldWdEtTeq3kz+I7BjBekX2qIvYO2b38Ix7mjeK97k4XmQOe3HGWFzYS3e
jnJ4vz/qAJumJ81AvVsZN7xmICZvh8W0ZfFNC5yELtFrw4staNSWvjiz56zUwKCV
+WkaI2u1djza05WJvzNfuEo7+KZDvnOUBp2PpHWEx6Rr7C1GVPcHZXQKLqWWehed
LPMD/w+KCy2sCsZ1bhOUOhorPy8p8HZKZ4ZLm85rNPojCardw8VV9oKyq58afKw6
MZl8X7klX0F5npGH2MPb9fNVDiQ52J57FN7FDPlpzUC9ZBcgJdGOftHoXltSQJSr
XsGW9eB/Uihmj2o4WeGGRsm5R3MTIaA/d35i4NQHtDOVWzEYlZyBobgChW/ENvd0
oR0fr+/yNol9itb3YhNiEp8f8dZ4AWoXFe4TiiKbx1NBDQ/8VBKtKvDHT0aaAcni
oRbeD5kzT+4Cu+Rmd63erI4wRJvxVEp84czQMHyqThzAFMgIAAXyUqVehNZJyA5g
NNkzwubWoxUTxFhK1l0XZWVsv9r1RNAM35Pi745wxxLysrB8+Y491l9dogExyvas
2BUoczvG7LyCEOCRNeMWBLdp71d9oX0pwVgEFBCinExfp93CLsWF0fTmPxmr7CF7
by8uKGIoDA/LnIOBnF1eQXGYhnN+TwTHKiA57AP1Y0m17OviKLmlptqRfdwli4q0
gYli1DG85EzUKcUg3VVF6WaU/WdXyyJrqwBYP/AOE2YB9LL1uB9LnWrS2CxJTTbD
sxXD3pnB4Z8wR6/6fbSB3sVZ+zmSLB8x0TEDXg/2wWoCaIPfXCNYJwiAel6Klro2
aq9jZ9Gz0o5eh6Ra31TxYqrS6QVoyG2+NkmMcykFQ3anYqvYjybpfbhATBl+s+YC
D/weU2NkJnHwJO/sqtrdDBG3Wgr1VOENhSNq/j9s9ccfox2OuKhBHBDFqUxorO87
s6AMe02v63EasnDQ4uAX1TKlf1vlS0slVJ4DtuJIUv9cYCFW469UClphG/sADIWs
py9w0S3ldYDLGPFA51pZEyF/OTwjzthg/8O3GapxHycJzvtYYvg2t3rXm6ZWRbw7
Zr3TZ4mekpKNI9yKsebV7Qa1dT1XbNye/bfY+O0cgw68ekUkfCg4a+72G3teo4Bm
aJc59EdBlpsGDs68UrUWviAE8xU6T7EnCPRA5PoQ++TynPljs3s5hdQn+gYGHt3+
eAG6KhJbj5by2ha+Y+3wfnPS/Aj5OuxDtUCsFsTUpSg3p2UnA3UxI3T+Cfo1PSxO
wGh3gZmgyrL2cFJ79BFSIzP2VqxP5XuHAlI0PvcigFrBjErsGPjnqHzyeaeQD4yB
FHuC1jm+Sf06OnxpBkyYBIsEwYO5NWv0zqhlYGzmCE0YQMwN68ijsNCn3nojl8ot
frdMt9PnqdRIYHWix7Qy9Gncu9Y4ALdmVvPGaS7GXRdhcNIteFCsqJi8pk/EX/+L
U79zlvGFY0PuzvvBDoXJAOI61ownZT2wUQFQr88v1CJoddQZtXVtOePTg+FqPA5m
AJ3dpcBaf4rzwrhzz/lHSODZA+2Oo26SU+L7jpTrUYRztzjpOGe69kacr5jNCWp7
XtNrmkbdO1dePuuog92MtBWKRIsh1oUIWC8vlmnZH58LHJcL9pnE04JE4LM/jE7n
pC/ru4sqg7S9nzt+TunWv8koUDbg2E8CWKXb8l+XPxvkg5wqhuJcBP8kuc16oTQi
UysChp667voHgvNd/5I3OMLKyzMaPm02SmGKBvVYshdEBjvesx70YG2ge43SAvVY
j5iBgv6+S1hIFQzhybmCcWqNuMHsDXMiUXNsbyC1CRXQ7dU1LeVxe4O3J4/oVlWp
L4/213NlkO1LkWZ/HkloRhxV0al7ADA9iCe2SVik8cxfnYy1+Q/A9j4DNQCDAyoL
jljtBVA4ty2W8+bPgJSesO9WY4vP/nFaWbWipZap6H+/l9iO+FmyFLfInr1Ukp+q
uotmhgxuFdZtz6y9zN68rH3Mq73Bs8KyOZYgMvYM7+zhWE97Jrh2WMR9Jg7fhMmW
ek4jcYnJXHiBrFy48JVS9pz9G14owzTf3TRGp0y6gagbPBwbsNY5jAHFcSJWk0ag
dnvsfFePf29hg9vxMVlTSuzDA5trfpPJWD+0N0Yiju0GpmEgPDcgBV1RXtk94nvs
G+2HSD7rrFFfGS6yyBMIkL3McXPWDQqKuVahacKjLgrgbEBzL0ufIPuj9vgCFn/E
X+XDrcCJssAd+tHul+UiIRemIlcL29KSbemBWb11p0waAh0DldRpqNf2r9JiLVFX
kDvZuPzKzkgyjFbv6ppeEUz7WB2F3PeXbR031A2QYCUoPpLqV1kmwsIe70TTYd+t
PjgPTxoKREWjSFxsl3dgXP94dPQ/ckL32Zy/CEXtGOqPXA+a9AolWkqenaAF6tLU
KhrgjD2aTYCQRWFo+/rVKa15sU+VuqSvybMbOQsRktn44CktEUMLjPLGRO0Lydul
Gej1bb3vB+3guGT6k37cGxmLNiXCwZIVBFsOkEF2kSXXTT0hIADY1OWN9nom4NfM
yzc3uCVHDFuzPkPsYzlm11pv7QiwQ0SnnbDFen2BoS+0NvHl2gZP7HtnCMGHiBtE
NYgny6l+kFWfAhIJC+I28mBR2cb5cwgR67kOJk+24VodUaVXpTEBb7+E+vAWO4mv
SpFpUWlwZRlTiUDjEHhAzznrWNJekOEqrTSmIeUQJlsW4yl9Q9bqqAgO4wlXUUxP
r2oiSe+1tvwaHnJHBcvVUQJ+k6+moyWAJpOxbiJS0bc0RCeiXnmIqcF4H3q9qGbt
8l4aU3bJ3mGbkhFpih7O2I6g2PcGi/Z38FPzqhqVj3I4eU/vtdfek13rhSqLPB+9
oLDfn5yt72NpHFZ9eedFcSVV17HOMe3PT0s/5CxNZtcrTrL/vf/JRqGvkfRPkAsZ
ibS/AeKKRZJUdIqRsKkfwxo7y3C8spH+X9lRu/SH+gjtAB2XwCHsYNUA16BgoB8U
oDfQxn7aaRhi5YVuudxHdfy7uG4vsljmwHKpWdh7rhQkmvthK3GrfTN2hiS3uWd8
BnkVKjoIxy14KEjljrnVeyfOneHqQ4nB2XPRtIT4raU3yI2bh+EoFKLk8V+0Nlhe
Nfdfj1cNwVgK/n+s7c9PcLuJK2MX4XycWGoNESIN5ZnU0sAAJ9B90GU4Jt7UMicz
kZmMSATNLOtxO3PUxdlnxEmTKRQ0YlzJY3DV2ttwkaUZVkHndJrdHuCdH2TC6HGK
hAgRDeuk9djMd5pNV5qQ9mX+cUxtbmWD9zkRffji6xR+jmsWGT4ObGmd34Gz4uLX
s/gm00FZBF/ZX5TzOhLQF3hbU8W6HCdCyT8bvY0z3GJ4MIsswMQdxbCnV7RTUJ6A
UNaFVXiIcu8jHuPS+KlvsQTw3JFCulUig1BjCDFFpreUEr81VRJKSl6hs9lLrE1m
W1MAey5AUl84JZar/ekn7jfPE6vJcgvaqDSbhNuXRE36wfWGXwPxgjohwSsuVfp/
oFoyFFu3Zyi8dpppHigNVFlH9UP2FWRDWr/420oz0VbvBjHx8DsdFA+R2LJxT6Bt
v9dLNz+u8+pRHp8RM3vTSXL9zVmsTx75juOS1Xvdo4QleWqt8boq+gkcmV6YPjUP
PAj9jNstsX/AsyRD/6uNCjwsLrkkXHwqNF854akWp4qjJgaRyO8T0y/g8uAiEqHX
jloTtwsqdWEvclfdi+KIqUCMZk1Bggd+0KDmgYYAFyK5IT5/H90MzgciiFlsziSL
4oJ4kdFAXr3q9xwkXkUvaIDWOk90WEDZoQV55VzPhGqqOeWn325P5fMMnFpkj4O8
78vNDJZwCY3z6hWMSizJVf0aEJKyMQztN1V11AS4DOy9JwRhzor5aJ64GW5QY1Un
Rv9SPsW4qD6E2sq03FCEdE0eQALSQRHxQUhmlbE53lZXXoVDBeiyCMHkJ4y4spdX
CJ03vtY0z2iIvd54pX1Ng19KTkRXE4BdFHdS2bm8rkPsa+2CwZmjWsYvlD990MaI
zN1/1bCWY5k3kOI9sKR7kf5/FHHyzeTAayiFqeJjP2XFcRTydFyUr0IG8s5iLkmj
oBuR8c4It7gVrgPPmnmFIpV1+iWODTO/bb/78Y7wC+JVQFDzP7QbR9o+sDL5p43c
2okzeclaZ5L691Ye0lWheZ5AuTOEeccuqoeFjsMCALU/SSaXZcDbUM9opYtCgVyZ
VKU0R9/u4JWHPZlQGhHffTE0rhGB3k8+DVDISUWMSrWscd66TsEUq8wz9ibkAcJO
/ltsK8Zhr6ptJDBspJue4q/B42lvGtioC0+03s1hjA4/tOOEDraus5DNJ56+MOxD
21CqY4vsm21L/9vtOqc2QHKJPP2SazCezVYDdOVoDaR+4AJey1DwNN4m8hFJ50W9
NHXcS1tcagJXAjhvQKZZRoW83d88RjeaFIpOqWmnhOos72xXoaAepneY/d0rZ50R
ncZDb+Wi2Kp45m74AZcksk6cnCVTKpPeVm+dxMHCMly1AMcr7ty2n0NmbpJiknQj
jYTRpbVD5fOVcnlz6D9e7Ba8AHrbmR+MOCSQDF/M7OQx9N9Pgc364fT4lT7pPOjr
GrPFyzhc43kLj3xpExdIyVhiplctFe9IepuqdkcWbeg8+TdVqdNjGx8DZ/646bQX
c++ysyvSQCPM3ySCXZfMEfJkkMx7hIESReWdfDWeoCTcJM0F2hIf9bum7blFW0dt
ZI5u+sSonJ8Cdzim4IYsOSzdv+62WEZ/3p53rKjBhlleeUQaNXCBBRPcTu8voGxV
P3Mf0hBAK2R8WpyNiqxrr+LtJgzVA/p/mG9dpgAJzFX4L5JLBcIbFLXmtE8+S55q
mka3xEAqb8NVPgjSRA4xNbnsvE0V/0zNMKQ4aFzF9N0TQAiy48g+SLoqErWvlPi2
Zb/+xt67aKu64kDvH0cjQXljoaOGP6OqXxsO/IaYNclHD/3aVCw93DtezQVjqmI/
B+QXXjn+LjuYghQTgqtDls6dmLqIf9ZFQPrUsajdYKXBdE0YSqzBD5VNoyAUcyrs
9+j+Fn835PCixTsJzKy492PZLG2s5yfM4L9gKx63TIaRl0dFvvu3pmVVSoQRvv0o
vMEBiW7DznMO3/glGkASlzZ9NbeoS1W5NG/3oOeCS8Xv2hlhrzV+XsHjYX9aBiCK
hor1EYNh6qRz0jiqr8BQVEkOXZcKKnOPhk9CdCazH1sbfmvukKv2uhocOa4sDdad
NZLwBN/7TyXyof5rmvA4uhDo88Eu3znScTQgwGpTlX+wxO9Vw/1dEXfI2woIN2G7
XJgpFfTQpTDQe+Rx5UhuEdJUki7qUKGeFkrjOz29vmt8fUwwkpmy83Q88U4oZhAb
Tly7K2lN0VzRe63Ke0WfapmJH2OpiBaiyVEePehND1s2JouQCcgFiEwqsNO+dl3f
qUgB4yLdWJ3E9qceHkrnQrauUBoZ3nHKtvefd6LclP0O6WVdf9YGRKU9t2AjgsvP
7RsIZU5VadWPzySlcwYQc8r6nLbw/wm6MRqkjVTPycvdBakqKs4NyDv5INJjTJpL
579xR7Do0m9UKOwU9N3NaYwyJF1CtKz3gT/2Y3LcH90PuilblGENGx8TzYb0mStS
w5tl8+wv9Y1Bb23FzxgMlI3Q+bZacByzV0u8zOssq29z+rrhsv1L6gI7WEuNHxDv
T4aLwAjVk/DliDDf/bnutzMDgKyCuOa313ertQF28Iko+Hk5sPoBNwgKA/y6Dl1Q
Z77EwP2yWTvLV5rsCY4cPaapJfaikcM1pI6TMKN+P/4MwWw8rAeLP2AIEywGn+V5
hnhTtRvISwSGN/iBW+dkwsOzJTLtrMC5GlFNIahQp811nvBmxv1/L1zEkh+iCNIH
pOR1aom3xZVx5Q7tFKj6Kb09MWhjaI6f6UyfYYdbIhpBYp2UGlB7m3R2TLmsC89S
MdTv4XGkEkEdAkqwZjfitf9gtszzH6dMhKGdobhWqMntCxNp6Y0oforwxkM4UlyO
wGbpkrONgKh0vOmnD3h5jypfbJZwwSXEt7APaiXwJq/oimpX9k3vBdf2h4o1lzhm
mUkQc9TDzO7ErHBpcrpetlQZoKi2898cBij9Js8tnp/BiXu8N3u53uNJVW9rHqme
ULLo6Fa7SQ5YkTxz8U3e5SJ5liPUu7husiSUYTo7BUXOxLNFhU5DGDXES/BSDAYk
ocHQZE/fITeSfnfNHysOUkBrHQKC6H++Kxqb5jGPuGwNKHf1fxOGtG3tSw6QXsvA
rR2C/z3nsbJS2MF9LFshZckHkI6dyMopb1YKskaUyY36q00+4+vB/pzJYk+UJd1u
ydFoatcCikU7jwVnIM42x6AGta4safE63gSBFyfxD0yBKH195nSllvtyp+Knu57f
479rnmIX6Y9jIIoKy1nXr3r37aVnadwHKe4BOtMTmCCbKgxOEZJ7pF3nM4KhUIJc
+6mK3fqju6aPWZ1l76VgkuGqwm3VBBABoFAfIqES4WwTP16OdpLgkgdkXRbCUCWP
r1fM9lkMpiiMM0Z9V7zR1uG5Z3LiMBhbRwSWLfdZQwaeU2HjVrkJ9HSTiLjSxixj
lkfgzN0ve3jY0dpdOnYAeeNGsb2ca1Bu9M3zKyoxkhg8lAxA1INu5DmalJVjFkVV
jCTyrPZE5VJVhZOaLdDx2eGB4bid5YouscTTZII0yfiU/zgX0PhFX/V7z6MtMr/b
UGLYU/Jt97hxyBpUdzoGmgigozqCtAxQIY3eqmk94DwymgejEYu4Nn5yY7JBn8ln
G0/hkZNTx5GNNP4N3AHCZiEdeRIorxT8lIiTVOKiETt3Mb4iCdlYYTRlnZAjwqL6
XIXT1WC/DeO/OcQWOOo16EGh0aeXox4UMZit7UslugoyqhHIkH7cfxvu/O9sC/XV
wAXmD4UvViy7CPj/cHbBOPikBo+JAg9WFIA8qOjDMXRLbGXzdt6mZ69NzpGAo1/J
nXstZmPaaKKRcoSOmNom+NhAnoPQtLxt0wDvgsS5f12h5J5Hh/QWdg33YPtgFXIL
1/9XszQioe9R/B+RG8QkiGX5zVpoOk+6wkwVk9ofZEM+mTC6Dx0GJlp/6WSlTKkR
jYqaIOO+BxzvoTuyP6lRQ78li/vP9AjgGaDMc7geTdHsceEFrqvn5A6/s80HbIhJ
IOQoRbF9og50eEwOiZR/976MLseoCtaU9zVZRFu7wN7c7SZZncvIBvQ2DqKCmKJC
q9krtLQ1zfU+RWzVghauvlX0fWxw4V3Pvw+zmxG8fAXcjmev1aHTuZTGsZh+Y/it
UhNWHnSPErOXKhligoEunPtAXooPuLc7cNoiVy5TwbaT6JgW78kevFDzBBxOV9eW
MWhVAbspHPGL75xXT1g6FjGGjave6sc3/qBtyeF15RzgGEbZkS2Tn59IiAUmSTB2
B14NfVMWgwDp9/Kpfyn+/Pbc8FLIttPF3l8OSNAn7l4rxaspt2wSD2v5A+UpqImE
5jp3IA4+4uJ5V7XgMmZ/hmTR7t9NSj3mgoFMrd+A3SHfcWknEwzr2cvRxa4IKJdw
XPJZv1yh9gP7yjO41NoSuKbvXrdqRM+UCv2mKoXdkftkUx3XEMl9lNqysskPF8Ws
ZF4KWM6bbsInAQ0G2QTHtUJ0baFAe5P1GUNKyUJcsLjooVB28586A3GQ6RqJosR+
VLfKCva3SY+4KBTAVS07k4ytk4tR7qctp/r6MIMaDly0SPZaUb0DFCWLu0mazbmb
FH1ByxaMdVCMjCSMKgVD5bkr2ZTL//TH33rhjP8IAsVeDP52q3vdCkwF1LbgUIbN
wq0WCuk/34RPtwx328E9OPkO7E4nVoG1/zU1dwZZOpMynBV6tgJcQCDKwUii6thZ
a1i6Q3kT/9Xl1gTyJnKwgBKb0CQkor1JGd7LmgB2Qloe1s+fBvbbbpgYffQdDqOL
xm+8/is13+gIK+5ZBbVzIP+yJqh+1MZWHFeSPu2tmGmkWC3rP0xRoJ1+sHZ6ueLT
yLnKf72nxzQvYhtCy5PKIhj+3NyzoYK6FTOVTpJrGKI8fXsWDnXpGKyB6fEPkowS
+Y6wSXxOxp4VLSkURqq/k/+ZMiN7mhOzl2pW/ciFvZeOZ3xw4MGIpp5TDhj1wEXg
NWNHAsPikWw/M7yrKzLzYbSgwN7pOvLOp6gLw6SZ3SkVfk+YmlkFlILFE4nxU4Vc
2VHr867tD+v2bh4EBtBymB/YI+FXYGzHW4vFBAx9/zaMO8c/56nl6EcGQBrVTUOJ
e2oAfYKuUjeDHNmIKGnUprIrpzlk+RqGxOzv36XpWXdNx1IWIbTuDGP/GvabuzgA
YHErPLL7m/AaeJVpW6SOleqlfQhdkum7wVj9kD7aSpJndUrfbpbXj4PL9i2Duzps
Sy7O4WM1Bho+g98Sd6nPow+sZ2ED92Y0ommdqNsmvu1hIYisz2+uOUCe8eneP6ub
w5x2z4NVaInmKttNfyZ4bHlCPAUug5dIkG+9f4QtVB8rgFXJdZZf4z0+4kbjsmbg
ik+b7TdGJXZsRx6CzAuM7a/aLphms9cvXzv9VPpQPXF1qQRz+XRqygvgYJC0Y2Jr
YoMe9/UPwGgVvs1/72RlTwTUKAbCa1jcP97POEMBcWYIdu8PgxyZMOS47qoLSbxi
DmpeT3indM3qlPHI6Jhwv55f0bM/NdTr/+0nRiSQ4fPqrX8OrVLougFVtfuRReII
vS7oHWsDmuCr+/GC3Z89ftiNS/ppDbyDlh4eYjZymkx0xJ0Ub+SEdgiuJaMv5X8T
YqWiOFB2T60S6tPkn3U201hFTPt58D8hOS66aRNgb789yLHAvAWKIfoT0iw//Mh8
2W4WRT/hUfVjNw14smaUYuGkFSzcLGIEtIPuVgeZ1xLKhYmHE1kYfgkkezJsqBW4
Qi+FHE2a91Op49de+B89qmfs8fQb7lEjhWP+ZoPhcUjXaTywnoMI3mVs6Dlvx12h
XK6EMkJv6tW+etgS0GLCKBjREREK2UDE+M3+p1LsyjdF40R4bxCqM4jBNskIFYOR
AaSnL7Ql2p2LGp9CwvIqbQjPl4BW+l3sblYUjAvjRlfNWKZhNXU9aKkj2vLU2ntS
eFKv4X5ZB1S/jOTVC/fcQUUGN03dAopzW7c27jOz/qiFXRyGYAr++UZNyaCp3Ojt
dOqdSIZIbher5toER6sGaOLoeqFvGG/826sfYjJ866kjPVWiqLtuM6StgtF7iZpQ
Cfrp81TwjaaVeCDZ2mHVItLHVFeFzHZx8xtuWH4gv5HhCwstUaUlhsLok/n5uJVU
2A7txmMYkdR8IG0K1ISoFjUGOxLlkDl8vExRHtwNiF8ZqoMflbVVXlu4AkjNCp7O
LwSmTWVqLLwQnOgK9AaUA8MVc5Y8+dut4QrhXlYhj1mQjDZ00hSEhDvhDiQZzKhm
FJehF+fPZ+GOA5fjEmcGHXgI1jeDgt6U9Lho9VhkKmcfQc29GJmlFM7PLZHctKU/
pUq4wRfelBd/Dvp9DolqYtCleGtm97aLjgZvhDx6kedyhJtNnl0/Im0iyHKSHaZp
lzd6SbsbYPP1n2jiim5nsGTZaxb2SNkRJmEV4khj9bHzn17VL70gx/q6Zq4Mc00y
ei5CAKvySLiJGeYUPsCDoQupY9kltU3hi58gZQBCuehaKeNAgivnhSiCEstJM4OO
0Az7IlnN3rUJ4w+Nw1tkrEj0aI5Jp8QxPzftOTFIdZ7Xa1dkFxiaHDBkbfPAb0gw
cZNaUrb7i9mKOZXV4vGkAqPhmwtp+LuWYiI+ZWqgKzC7LgJp4XxCSnh1RwdWn3+k
Xwwh+c4cNrmDn9kBcVmd82b9D8tHbPS9GmqTJwKvawZ4w1Y6DsA5PWYg/b/aZTGd
Y5RszeiJjmY9d7BX5Q6Oga1tqXCL/shagh/LubZZ895gVYm/6xzBdfPDPoS0jca0
LE2WktBitZIe0ApilLCQ+yM0j3y9dqbenzG26q0daSw3PZhdk91h4BkDMpVGqHty
snzzSVdwBUjHDwyZ7r1uOT5RdvhACSfxbEfDj4u1PBFJPmAH61hBSAbyqh9RJ3AZ
iLcsebHWmxgkd5Qch0jYg/2zigH3Stw+/UahV40lJJ3sWOGwLb0kSSOFCPWW253Q
VS9pErpAA6zgFZJaxSJuOjFTsRIxKAeqH635GzqvqpX0D0ld2wF21P9d3X5PjTRK
MYutiLX5ZsmgePyCA1eVHRUQVZ4jUTK83P+a+ca5R1GOSbRr9j76Ta/mnyYiSP78
pU1ptMjoDxCFzJvkHK8KnsvbFlOHNI4g+yrIj2qVhIv8LbcMPOnETCtt9xdOKZuB
OZiIgqydS1OvonC9mdedYT+sKzH081u//Vh5OazlSueycPkKI9FW52xRkbOBIx1C
hEf/yWJbNFXejrmTYwck6oL39jRqolIiZsk7NZjRqSAqbWaVRAYAV700vZieWWO3
DelE5t77i88So1L9B04W2exkOz56KBrMeMUr+A6/Sv5AuQHlkOJEO0dYGTxVipyd
XHNm+kBSEHjLL6RZSp4H4DXFenEgVDDss30Pu2lvV3N6i8OieFYosH73ZKQaWyxQ
2F0tXqOX5gXEVGcu+uRfaM5uT7VKnz3cG+TPEExebh2BpQdeV30TLAJ3AcuHWEan
My+aWx4TRZVnnJz3ot/JsB65fQqTEr+8lHGtlqkGUHIe8ZCFDdK+K07PulE+eJnl
0VtsnI9QMIVBg7WF0IM2Xq7EqmKJ5cmwE0huxC+kwAaq0/QWzL3AWCFONcmx2IZr
MI0E5HqIF46tCijcMGLcBHoJRi2xnD8Umyn8rQJe1hN3SEglGxRg1B0Rqdih/VZl
roIckWL3+y/9OxM4RL8U5gVLffRlhLumA1sATa1rkEvI0XDzTtYWsXX5/Wrysl3M
JhRhscZ0pFc4zq1IH8T4yebWY5gRtfRCs9fCgwFLGF3bB1qhHpFmNjtx1gCHp6U2
wGtXQ1r725gmQ2nOLGiIsCnUG6/ox2Srjcw925cgIoLLEo1guLaQ8XeKXw9kvW7s
wihK1TN/Cw4QXA2gOVQ9YqepSwRklP8YK43vPuedPRu+KTLUHsVSt4kI/wr4Jpwy
EGMJ9eQ73AGEFWJqS28JVdKc3nRIzNgjtdSwrQ19+UqB+Ny/2Dica03MLgbssGmE
yUxkODiD6UOJ06nTv4TUmk6pxlYIQgRlZgSM83DCq0y6mNR/JvrvwX86wZNnjpwz
Kn9GemCFn/i0ZSJ8COJa7ygzcQ6eynsokhVvUE20sSwScrSXLsdytIyWN1fme2qC
4OPsYPKYZhDjKSFIRC3z5/Ge2wDZCYi37Z//dkTMasiJ/ftGiJb8KtepE5VEVmFq
SmoOgRZnl9h5Zp1Acy1SMEwE9UZVqaPDeJ5P9DC2CXzdSCdQBKk/d/9G/c5iOGXl
0tqPyrVi3ls08UjI+b+kHDC7yt722Rohw9LQKqaJtFvPhqFLP5XHjDUpC5rEPMiK
X8UiFMnXWgkbuq690Sit/FeIj+zKaxqQQvDvt29QlzrZPAPpXjkvxD9ARSvAU4up
/qc19Bwu1kv7GfiJvmMIgB7d2oMtgbtz6OqMKJpq66TZgayaCyU0NilFl4mrgt5l
M7tF5iJTJ9+T3RM+WkGY0OkxEPon3AO9VaoDpzX88sCYMyKhbQDNSzDM9Bzu9vib
xEVSpMigHjuAI2q/LjS5z/AesPrXqLm7J9mFQarI5fQqbbbV3TlHrlsxi0GK9XNn
6itHJBxy/hIKhXDvYpnHK2ZlhQs5/yqXVPZI6CnsVLHdHWoXEaJkkoYywZKAjhM/
rVcDss1kUQIdVtyORFiHyfw9lZUdWAElMv5HmLzop6DLjP39/c1s5lkBOfaBKek/
yjh1EE6cmAmtIlgCpkvMvH0S55IYV6p4ObS+Vv9n10ExNrug+Df0cdTuS2hirB14
ZFzEz1nRsNuu95WEMXYxGLnsXwjcWFxDb3sz/lGwRlG2+fdls2iDtMdrkAMgf4LY
JSI9mDRN0ubVIdk9QX3/LevlpZeoroRpq6h2/7QPHhZp2vgpZF9egcUbcn0osqp2
6Jr8Rh4V4aCLsjGq9D4t2vFeaKcxmzANMU+sj42sMtzr69tNZ7lsRIqBy/P99i9Z
T2XYn4Duz5wRiXPCYtcjKiRpjetKwbVsxBB5WAhhkqfALPmapfzyI3Sn6KvKjeo8
Fa86ni7wSViGZ/rtqiKW6nnZuH5a0O9+UrLOY4clOLyU3olhqCNBLqttcQwI39pW
w0025x4Oh/EKPF8xEr4xXB/2J1lP4/x7kZk4BhXcgp+uiZsLktS3wWnYW6UaMgOa
GnabGPu8HIjzHmbUexv6OpWtXQrgG/P0sPO+AUtmLAZDiRt1UFHkBcpiHeczWZnt
qR2S9btT1Ikzh6PI3EVjcsbxR0+OuLqd5fxRqy9zYomjzU7muqKXanGnEjeV7W9z
YlMYqpWHV+tGASWVBBmdp0IzTaOLfvsbXOH2S+sP5nYF6E5bpXn5g8Q6Lsoy4yTx
UIdWJiuVqPnWPwIPAXspC1R8sKidMt5XgX9o11L201zV/05b4a9SJqAoS9JJc/ka
FDiewh63F/ophclZ04/pwhmEjO6hmAZ5A/2uQMPvZ89zyAL5oJHbpisyheFjaezI
qO9d4xYRZswhilwchxDjCddKGO0FHP2XUEV0rVpd2a8RkA13oAj7mh/tP59zYFAD
ofIqeqKSysuYSjLQcLLAhZnpg9V2O6vcxAN+xR/1ibjYeeaKXMruvUT3eN0wCye9
1hssO3LRCqxdnQveol1u17oPuFFaZ32zXY2vabLQ3+MUDz7sBI7eZtTjNZedC0kJ
Dqp6O2oWBx1OMwqataUCvVhRvkiJya5pWAdMuoHTS60fBBW1tmAXoaGvpuoWeBly
7B14TtzKPa2n031MrMvu4WlMNq9uljKuUvwanNRcQkCsshc8F6eEf+Szgs+m864O
tPrMSCsBmr/0qVuOSzGz+itkLA4EkHF+YJFukVYYwug09Z0lW3Of43UVZGcRVtyi
t2WhyVwg6JItWIoKcDiCQKTiESefSBHdXl2zvy42NPHhlSBH3sDVJKaCPZ1h1Ctl
UibXrALQrgX9lv/Y1ScM4selpctV+U1hlKXQ5cPWGD+WnmSVPSLFMVN9luj82A8h
M78GFzcjkHBCmebCvQGnO9wplni8DH6sd62D+wYMwhRXbB3BV1RFXHzbgh6aTX0d
lk2oXcycOtYDx2QzdWMUAVh5w10N2KIliJcRTGaNANeZguiIMeDRD/WzZVwzWmnJ
o4T5QuGl8hz9vrSloXflQgOVbEcLAQ5lMXNGS5zfnBIT5tvYzhoPrTFrWMrKJJzY
aGJiwign6qh25yUh7Q6kjlcTrF21EvI5TqyW7KkCZvvDQkesnroqcwip5YgKS4XL
I7UnygNQYfDEzi/5aWFeZFQEF/bZqFNvN0qvbm5727sAkndZsI3mjmar9IPauSYu
G9Ep7FRsk4A2Qp1Q1J8a0/vMrdMGq9U0s1I7IGEmIkyBv+URGlJhnyY8/F4wDVUu
MYh/82qtZc9UTwd/VWEWonZiIxzGzuygyrB9nN4H2DwAB2d0WNfBwxtK7hPUlQEm
UjSd6wcxH0X2k7Tz9ZIGtekhCOYte/Y4UagYPe4jXPf2oGzmdv4nwys0dEYBn2hh
c4T6aJTTHlnZT5lxr+8pb/YuO4JpIKchUSdoXvON8kUrd6EwKOniX717myn9TOTn
IYeSHUE3tTGqc1trO+roOQGkHxc1D83LDRjX+YEed74CjI6v+7QoIgt2aiGGhzwp
MyrkGSS7dblbg8lHPrL3mzQFLNv0hxrRjI2euBFIJgXbWsAI+jF8IqlVqdFeVTL8
5yK2ycrjQiyS4E8ehWclzYq/1apBcOsLl8uEUsX2Mv2vPR9PF0lG879Jpj48b0a1
UqW2oA7/ln8LX3dJ3PH54OHot2Of3+B+7FAdF69/61pJwkuVGRku29So5XxAopvw
iH3DuoQ71Zipuoycg9NhYN63T6o0EVsrX9UVyrR6UOG2EaV6CTeo9+jk2OyLyXRU
XFOsMH4pjYYkIm+USdGqFPYxnerdiO2HEepLPa0dLDwRfmZHmj7cOq8iBKXQdlAO
ETErRSu2LFrjb/CvL58nmbAb0vRgOXhDjlWJRTWykMmgjNKQBu1HppO3HWkmK8F8
hq2iykzCVjtFJXL1WJ+I1fb5/+FD5BcKzPxaJ8aw4Tf/0ucSbIFu6iuxFVDKF/Ob
KkfbL6h4DgQ6YGXY2HOCHVYCqiZ+yiTOtHoGs2/2MUypPFtKXB4xcJbWEXzw/z63
y1g1JF2Gv8W5/iMuVdkHfofI/vpcxE1mRQA3Dlr/L0+BfKOMw0x1S2TllrxBHdi3
MPguCU0BYQcEnnqA2WrYNYUYs8n6k/u8liBWT3b/t/lKf905EkGY1QNPtDQJ2j0G
B/w6eaGjLtoExVI4Hw1/FrxEMZvp5ldJsxYuKuVk7c6ppHQ0oYGNNq+DQa5UBuRV
84QzudtQfYwdGsDcuXoD9Zb1EZdcqS1xjaJZNTaD+N00ByIMh4XVDzLSOBd6eCNV
DtzUyiroZaVvzJr3MYvskNUl78GzDaLH7oJrH1pOmSdxRmgYY9Y0lrKdCk/iNggf
EMVBdVj1NFgTro5G46FGrg9XpX313DzhmbMzeuh81yU5qSg/e11UMgz8wxxxfG22
+TMs8R8aVa+8yLhcsxD8aA1j4p9eP4uGjHH6wUEOpkqF/RyAKPp5RjPdUAvlrULM
ZoVnAs3JFaXHzOMhTgsaHaCuBoW7Ay00Fb2t5ErhuONVspVOkAtbnUGhhFsUk0dl
sxSAAp1PZ/yj6kvg6418DGQ7Z6/8Y182jcNRXvZh8Scg56wLRXq1yNA2rqmys4Sv
5owS9UKg4EmqovKr7PIg0bEIblH4OVWcIX9K8xUInlcy0fDVCH9XqsXlbZkbb8d4
gndRTMQwFYHik1Sa/rRXV2F7iUd9bgqSpL9lt4LJLhy6nfujUQ6MzrnH7vy2aDs/
t7AGC03puQ9DN8ak0tQmJ6UVhGkxKGXub5vgkdTbGFvf2Hds98Dz1I1hYBBC0Bse
AbiYgxUENnswAqPRZRV9eAC+alLCdl9HuB8A335J86C8xy3GtDdAm77+G7qIkoLn
HSIk2+hMVVOsoSRY5Um5Jz/PjwPRrDIT3ozr2zX0h3Zv8RhWRbghpMniVYiGGSPo
4ZfeyE2eSpwnsLIEbJIKF9tVaVPAkv3t10Hjr9BsVM1xCLxLN0pibsTNV3Ca+X9y
BScHkx/+ktQ6lg55LKoyaOrrktqGk4PYKb9Bm6zaJTL/p2KlHPKfPLrI0qQ6827w
u33+tWEhUnRZs8VhT4TOml/pTUo7jFdK2hdhmllhw4zbuZMEFWK+HGQQLJYKlJEv
3kGhZ0IF+1dtmf7PbzZSN5EQqTcDscdrtCU3OcgkfB6jJojJAh68fmwcNPJCGWj2
lwgnZL6l7Y3651PasUE14RWw3Fz1dnsN8foA7xp/zpMMIW0wx7ZZ6n1eE7nIc6zj
lnnZA0k0HKMjlUQeRpQ57vcbqod+LFUPVWqYaoYbLMNcjIjm0BUVtAnHjWdZCwM+
KJt945shq7r8K//7xEFSJSJqYjaNrIARSE2Fgd9lEQSwdDaI8MyhNU6S3QAjPRHv
i9gR2XCCkNnPsirav+y31rkwgDn1rYF+BELKD26kD7Kl11f1LmKakS04iOULyT2B
sWql5/4SxzF5R68+5EWb95BABilPXdxpHoFvwnoql6rZ6d+5FDeQHIDy7XC+Ph2l
HzVN52G17x4Av63LfRqcIgUGmlxHrbg/rjCh/YeGraULRaRVTjCpYcW2WZvn3BhS
vm5XOzekdFcuN71AHy2Q6SN0AIJ49Vsea4z3MeLir6PO61iMH/Dc0Pr/NdteZ4JT
rZJm6ZquGlEz0WbHVlrroJV1WTo44EEdRHvAUsnQinLET0+CMoZ1l0MfuPdlpvIQ
BNnnhwzGFx681PImwNuIO/0PTNGLHtyOB5SMS5NQhCNzWX8KGAmPaOtPRG9KovmF
qyJfNlD86J3Q3WzI7MvzpfUDt/UpcHbARBxo5GsqBmQjwGBwfjNsoN+36e+VrLjn
rp8sId41DJ/YdNfxM4RzUH9J0WzeHqz+SfLJ4pcpR2qjiWXFErQ6Kdij28LYGxWD
9zCsQz2IE55r+gyeXoOrH7wJWqyN8INHZ/zYtPXn602SkE82IlySlACLnZ49ZpI5
f0g9VHZAhYX79ea+LxP+n7rtEa7IXYRTxjFl7XgVEiS+mpwvoyZ3kbed2WLuYYZz
jowxM6bR2lfNIGU/LSY093PuNI1+qr9lvtwdzp8NlZW35SE99Eu2n8lK4gCdTr2Z
y/YUjKf3cabSGRlDL3yoN0JVCuG7kZx5XGitqIb/wXXNVQTOnPfGicbndvCuDhFh
TCbMO6bU+eHpxejHpfLdU7bZpubtHj3ttLsVOfiSk3cboC4uJgK+RbsGeUZFIcy4
a5g+yZTqFkKgaDo03E+LxGeHGoMP+EcK9HFldhvsBi1eUT3BzGHJPtmh1rQtax5/
5WOZ9INoAji4hhm5FuQONxSAEOwW7FAvT+wmPFAZ6i48vi1NlsnC4sLY6ibqlJUC
H+QBi8vwEBqurRydgDgGp0H15mH78ReY9kTPVyzcc9/GdoH92JrlLAJJ3GfVprv8
2qYCA4nPSXGjIHRcMCySFndXAPAu51kTK/v1we4WX52hUQgFP1kwMXuFf4fiAqo7
A9qrf+S1tQs3s2/2jlRUkraaI+y17Xj2tBPlCHWXkTIqCNKoXV/Z8bzwnGsdy6dw
QbiQzVI5VD8UM9HmZNUj+Z6otqkpH/eUtPM2cdueZuHs1KtPoQwkVcXsciDqymbn
yO46g/30aGLGj3pVpmspaxSggKqqvkjDl7zfO53ao1GAKd6dxn47EIN1CcNTc/d1
V/bIF+01nzFfgV6xdoTTE6zVkWAqeTZaLrhdwylhbqHIedikU40kuDkOwfTGYj9t
xVfVFTy1Khei6B06HaicToCLcxKXrv/e9Y66twhOLeK1E9szKkUKpZcB6+drqWvo
IgMQ4yb+AWNLTqZZnMXC3nzacjN88IfcGoCeQvPe/DiTUQV5n+0yHAxwwUb32/8G
uUlJRf6h5mOsJuDj8N2/A3FJjFB1FOrYQ1VGSi1FqZC1GsxHG5Y+B0AZMU5qRGn0
sLMfAY5IU2CfUnpCOphV3gpgcD2f05fD5ne4Vn9o+5QNXbeDnf1BouxD+4fBVqs7
ojYBDB61dugWZf4ORkAyCNE9e9zdrotzzLtuFH8Z/1ttTCMy/uEXnOmiKb58zRVD
XI7moeAHXcG7udFoycLLA4cH+Y2IOngiLdRNXlHxju0hfTIbP4H/yWRjpbW4YZ9R
0xHlYRKtP7QIdxkeWzSXuK8hHOUGLwHg8IHI3bL42Zjmn9vtsPT/rly+NJxvx2g8
YxBmEK3Fc4xUm+xbOG57fhDHgZI2sbRMWA3C/whJ0A/gpx13EXStQX1lKFQIbsUr
r3sd8SXkJHCFccEWEgDUNpvXID8Kkf0MucIkCRvi03PdnvMwu3ODHTwblqXPRY8s
yPUlc4YhLePCtgpgVEmwOnoO7360hVeJI3IHemsea2ta2YLfr0V0+VC8WuZeTPGh
ovI9sg8PMn3TDbD99AwnrHK9c34NnMFfjmd8UU5+iWx/gSf4E/Ky6TizpLW+n5Tq
PMC9VWv48BeU1jj9YuZOQV3BZ5kglKv8M9pUHsWfcfCBw3+cYEnFuDiI+6/p1YUT
65bkaQmkpvYW4Fzo1ZgpwIX1u2y+RXHjN+uGFQHs/+M0RCRYD0l0KX4fYIEAdPyS
En1smtQe/JLJr3Ar0mMOJTwuNjJ7B6WU280uEAwUMWhTeI39sG/jbPKEe4eERQff
vHM+8CyjA+bNZ0hP2zP7uwylUz/n0RMF8CoEW56gaMlgxkYom5Yjgsyy1WblRFlN
/6Mj5Ks+Zt9ZGoE0wOLdFH42Nf50R+Jwt/i+ZmXj7/jRIZgBx3TP1AUN8cPgdKbP
2CT1Tx+p2dY/Yk2VIyrQeqOD9PKDwLqlD76aF2IpqHEyOkRXpmka3jVxjuH05rAz
2Xe0PbwAVMkRFm5LKOiXmctD+hCcvZqmv0uLWaZvedLb9rizcfuQSw9o/d1Dv2WT
6vc66g9x67BsIf3y7Bz/8WKUHYMYKsvvK93jXiUn86ELrczHuXAf9wfm5NjagCYV
XubXzqj2ZxyhHwovCK9oWyfbXVEwv6g6s8G4B9+bXewG2OS4tUFate67h7TO+F96
e+v9xzWH0rNMZa1jF1xHLAD5lZ86YHKkNfLLSy51iey87sA3qEN5LHqqkV4CmqfI
MdQBqlUWitK9kzmzbEmgT/3yGX6EtyFYMu6UIa+p8bDSjfPZYNDLY4JhnV2j9Rbr
zJEqNY3bmJMSK+46i56pup3UrdOPif0WMbiCMZjuo72xIm4GWgEgGbLHr5QygyUi
IY5pIl6dWnih9z1VHq3s5ZojFzKHRg48hBJwSdB6ypTnjWHWvlDW60ge7CbwdpjS
EB4GXTsuhD5nGpWIsgkPuni2o8ld0oAgj3U6wTsCwh6Fsj5ZFhK+YvUQNU5LsEB2
tWD6Ezb/f/qpzz8h0AAMsCZG/ik7E2qVMI4U2JWXlN6CK1CQIh8xPhVzyag33xEg
C5BVRwHn3qhWzZs8Ik1M3woH+1uHaH8iC7CNO6Epoe/NDf/s/7ISiNw4paWtHVaE
xEaOByjbJBy9IEe4sDjbJuuO7QhYSDaG7Ql/ix1bq5gCIZW72ZkLKegUNwxZEP1z
BahDNYW7rHgDuQyW3PVCWuAcZi0ELXMyIbUZXnuBbvvK7ylDMNtreUFfbTSy/Cb9
33zz7m+IAdcKHYIiGT+LvjnyUzEAH9YfcLOLfyMZWy/nHDdqPYJuqecPgn5ZtSEo
fI+/JX1sYAZvVc5GVFkKzD6k4ldUbTY816R9+47n5rqzGs8MvVltSAyM7kpG66Nz
utAKWpepJS5jSg8LLsFhkbl4xzQQSW1Gr8y0pUqploptbsSUnjv5b1aYp8f7j1u4
vLn387tW1EqEEgrEMd/9YuUpcT/VAQiGgz3/RUTdFXPFnAjpWbIhUG9RlTFmOxtP
KvoWAvZyhqOVFilkUy+o+LtkCwo3ziNq3V0P3oCFPgi82K3hzNeZDtywSePH9lUU
B2SsvB7Q4dNJlU5Ni+NDzOra7B+YWDr/YglDY5cnoYrqrNKcbDhWteGgapiFukyO
CS00aB6b+BFRkz7FN+3G5ICjHkBSP1pyQDWeWsguZH9WNA9d2RGnfGnQFod7W2AD
as1V5of/OQNLtfVHCbi70+GtQKqBQW6H1RFvaR7FWNrYhosCwQ8zy3ur7xxmj9gk
EdqGsJywCjzipY2fDVxBUnI0kixsp367GtGMy0OaYCgHVCjubYTRXJhfnGkx7JId
mlTeDRamDcfA2kjBl3jJFquAXx3ynIHmxNBqCWYLIdQNsCSpTiefEa8KVtX4D8ea
3NBzPgEMVyVH206ozgdIT6ddka/g/+HnrtmA9g5LjeErtDK+7uho8ec6ubr9ceBp
DC070aDEYrS/ffQ3+Bu+xoNAxDbaf7ATLS/iYAWVJf51I5SONipE1NwvlDTSwSjb
7GcJMOYo82uqyhMmj6JUarczRLZy2AEEh5c7+wY3cs5R7mhwJGxVOdZA3bg1rbba
BoF49DyWEhe5ZMr9Q5DpCW06sGLt8UL0peSSWJ6fpEe9QmjITFeIiAwk9Mgudgl/
DTQtW+p9oA8zm+xDhuEp0xt0K+q1af9E9/dk71bOUwPJOzHQcs8M+nVpkICCs7aw
q/1oB9EzkUeB87YE4kISUzFYBW6D1rXLuO0oX+OCdWydyX30oka0svvxvDpEuX25
r9NFGf2szaO9GJo6wOKlqkEZogOAZtwuAWU7xuHs+Umojn8BIEQAr2OLWE+hHI+t
GRgyWXjJgJjJbejkAZmFojkUhnJhxOjldk/DWV7kagBgBp1ITHkYN9zjDiPDAtiR
z/NAEPeRzj7NdQzh3bMjes2yUO8ybsAb/Afx9+IpgKV+voUrtr+q3e3mEXq9E4+K
zxc9jujjsxgwdYuRutufvS9XlbHy5DA9N06MM9oZVcLICBSWjKZkhh0sGNSYmT/I
WN1xUKCS82zyF9YozZv5PviGFXKvCuO3K4MrDHbXHIGIXDJkrS/Uwts9shZ69m1T
AkQmnOczdkZkwXIDz499kVkDMwGL6jmlvu2eRTw4Ohx6Zsj9KyclKze4HvKLgj4p
ocIl49jBUAdC76d8z19bTEASD9ZB5FrIgNnTV9mnEvBijmdjHPL7RwxkSyY3o+Mj
jlWKAp/tx633/l3do897gT3VAtNMr8UDM2UYS4kN/VAoky/snuilVLzqqPBp0Grq
a0wp9nf30+yT9kAej2u8Y+fsIqnVkODKaGkYlI+uFj/iGNiV/yQHEfX8wJJbotna
eeUgAwgcXyDpudZWsxL0jf72bacW9bNoOuSpsouMgx6OEBM+7QPqD37m+vd6U8rV
JQe7+MATpHQ43Kd6OiN6OTMTIAY1rZ4uEQfh7JlzIxrz3lM31vCGAXH2sVFk40/j
mr9TuRtwzrQUIE+7a7R98e18YBjjVfCRJtiwyo6S6Kn37I7iNrk4f7Td35fF7exG
f9LtFqGgQ1UMDnvqxXIs3+3Ug5PnN7sRly83vye+KXEFv6bJGVSXltCaY4TKnXFH
m+XmvyhCWtY0qsrwc88GF3vdJlSAjEotemeWpeb27e61nK69S0UAhL7wCz94MC5P
CDlLQmIQ3su2Q3p5NNU7neXLJF9SOWJtrG1gZnjPVW869EjaTBD2C3rxfTCPDRq/
mK+eHmn16eEwk9iZ6ASPql13Bk/0QUWBERDATMdoNX/GffGyxUU1eNv3QdjHJOR2
LghjB7Rtn0FPlIFf19X+yrAgLQgYTitV/T7CJ9Z3gexCXlvnmhdIM0K2/LRKFHcG
/TRHHBgYvxw3E9JoHXJbYXeADHCTlxZVUhXqoRq0HijmhtwQ7MG0ziKumsk8oMRa
UM7+QyNs1AExRt3rpMGI1B9L3BfNLqEGXP5oJKrTlWlhzRmeT+0cXp5pCRsig9Zk
ctgWpdqDp9qJKAV4K7t02Oyg47fM8jaBkfhXmmzUPTLTnGmz28ZEjZqyoFCIo7an
X3xNFsv/03ti1tPx9MEjEctycFRcxzaFmPkGc6FHm7d0rGR7RiOHajFi6g7CpIlx
j9DJBc6wvTUQhd80qiinJaBaIQCZiahcEUdLdq+icosq4E8tOsYu1d/lMhJ4nvWQ
Z0wiOrJUbus1ms1r2uRdpoQmId6JyhKt/n+gRZog7jEBOCdpQX4amIrPePqSvHkb
CZwCRf9LDXgaMuGXxoDhnP6LOvp3y5PJFvYW6ix4+YSwGPIfm48WKeXfSrkUR0+i
T+dUPdNUROYEr3/bmE+LUB+2h7Ag01ZO1YL688VZ+EHF7fTDAatWA7vhkss69/zU
LDb2RDE/aFy+uT3ck9ozpQNiB7sIn+bZ+lZKZ1eil/QLhJblZcppbehzTtMY1/CP
hpgyv+tGpVW+XAHTxP7vPcP8sLC7rVwjqLuaRCKjTLjt+3oQyD3kM7ciMuxJORw7
s5pNyj+Sh5Kzi+V4c4bzoeOBUnXw0JPhg0Sse50uw+44dQrVgF8iVbR7IGEbwfhC
p4zLoZpjKqrymCScgQoFqVsuo0HmAeIRn/YG9gzgusQ61Q+wZz1i3Yr9rHBuVMWJ
sZk/yTkUuiBU+OreCj48gssAEHyKf2c+l+EM49vf2Jx0TKgnpehMWUR4gAl1MyaJ
1S3hk6hBNLwMSJ4HzJs8Cp7PkOhGaqXSQODxB91sN84ikSiBsBsy0p+ftGB0bN5P
mG0T9bO4mPsTrxPu7XesfxAMnReYlg83BqIfMPeiF3OuhPseLjT40ZJE7nhaXGUp
P5lPHNb0ETuZLkjejP34/eY1Az5PwA6FPC/DxjWJ0UZquyjar/tf+rh3yjQFR90U
c95Xl6g8RreMfpIG/CL0xHD1E9YzZeXL7GMn0FiMesPo0rw+hXcEtnsJ+pFe44nE
LSJgv1F+jVTTakgumLiCunoau4XTOu3hKnjvaob7xkz8/SmKlWCz5KG5tnHxvVPy
IZRa3tply9oNdtf7pgwaKCYgwMM/n61xjs0TOrKx/fDxxd+nG7eW+4SrHKgGywoM
KGWPjnh26zQ4ENdUV+tCHpnb3k9PK9LB2eAq4xjbJ7eOM8pvJp2YkY/lWuXqlYnT
LmOYg1nKoLy2KGTYjVeW17u1gapF+IP0icWDAC2PYqK1ykseelBfBsoWvuEIHymN
XrbkOR321VktUCve/kZPP04Ueem+KRmRwXUxwRKlr9wmcU7uwTh5uZjrSLW3yLZX
zRPjNtPh4a0UHR24TDmFoi8ro/VXMvO3sQtBTA8kbGx6YfjVQ06+g2zrJ8J6rvf4
7cDWbFqWZ8m4S7lPwh3pDkJjNByiw4W2uT1o7V/tpF8IIAFvHchpGA/SviXLE9fP
PT3vVxIru12abbCJr6VR3MqKb1AYZLIb90/VaUXI6EUsb4BkO1zEDx21Ja37QgzM
ljtVTLEqVwLWllhcsE6HldVIu1tw0ffdRPUVlnkUl5/epm775BbnAaeOXpZ0DSRT
pwc8qZddXw0VsvaOlanrsk/qWe0HI9bLtSRNYvNfFNdcKeO0WaIsCzGcMC2ul1Zt
6ARZ1Zu5PWFOteEBnmuH5NzO+0Es2p6uDItI4NOqJH47L5F8/ZYaZIsHAZZTHy7O
aVHlNz9g6t0srvQhaTl78fGK+F3ZCXV8W8FWctZ0NnjgSeutSEWJyslFPyx3ddFX
I82VuhhZvPniStgWpJK2qiCkO+pG83DEijlcH57m3YoNwN7WJxBBWF0jSMlkQ2p/
JJ2QesNm8GnqsJkAjKQDUkHG2IjTXvKOjfXTLzMA69Ql9A5b0mxehlSoLVnzvlCF
uwKsZHilPN9BLFuOTruCFeSUbbn2zviwH8rZCA/YvOYsm7eMtffeWQJbVmK7zx4k
t18hKBr1JJ6Ee2FZhuAEb3a3BclWYQru8mWIA8LIBEZN+biDssPlMUx1WKSVQ/Ta
e3xGjrgYcHTtl+p4rHOyLDsU8o3leibzPopJLTY0MBB2d5ccItmYFq3X2S3H60Me
1A8nYFPc0KLaia8fiPciq6NN6CG8Y3T1C77hbYRnNzXPiWNnfn2/2KfBEqiJGdXe
MaOq62IUHVgNmFTWXqeoCbenSnog56cpruZJrVvVb4uUdo8KahfvMc6crSrDeBZy
YMxp2sH5RgbwngEGZ5f1K5ZQap7MNKyB+v+dnjeRzHCt0EsOQfWZ8ADobg14tlgp
bZxRPXHkBwhfBSIDFQbZWBL+bA8NHHPmYZXuR8jvrQAC0toM3R2KX7LlZlHRWLTD
vpPV28Q6k/Urm+dN/kh2/qrvUGFMLb+kNPErmF0AQneaz4Rc8CVCFyhM8B28U/Cr
LN0zi/Hdit6mNID3JXeSFyICIkqM2I2dF+O8buJ+aO85wkjd2BzDzloH0VMo6dBt
YPB4uBerR4lE7eE2g+ziPwycZB+xuuLKa7NWrolBPUqWZkYCHOkyqiLfB5XzfGlU
hg4Ilx7wbBjR7Vb0wtBrH6e+Q6gEtqDdzjUKFRZ/W+LZ2v+jrX65F2rd4OlU+gfC
OjohKtl31WtyBqK/GoojkDH3SW+GEUo67OLhykbrb2wMN8E27XjI5evQL3OWocLE
9pLrToLaHFhsEmTd4pmnXWA+ml+zVLI3x/T3Zo/YX0YlV1W7QPAPm3Z3xfkbJDa1
m0lgC4rl39ExGdP8S11sysvNp3ojFZ9rCz3zcbt2EFUbd1VHYW1oC5bb/MsBzVa2
Y2i3U0Cs3VLNtticNF9//qWdqiMp5514oTiuAHX09rL/R0SlHZTLh7e36NcliOdd
KWzz4Khum9WqUFk4zb5aOMmoHN5BiGNHd/Bj3lNQ/uDWgFaXn/KS4c682MeHXuio
WxEcIlabEROLRTc8Ib86zv+7j6q57XBWKYGh1H5WSFZvPILYTD0R5i2n+Ue2k59a
oi9oEHqnSI6sC6ai0i6m6vusXfLGuEQdsH8LFBI7SNvndpbw9u1XMg56iihWZ9tk
VpPf4HCj+G7WbCRhpkiYH7PHJdHSDA2Ou2dcuqgt8Y3EwAhDHq0Dr+p868h2m3wj
Szldmkyi+wpQRiOZhbTmjN3bT1TLG7Y+WoGAqsIRPF2ks2P3CmPC2fgSuZO8bo2m
TCkzYUDnKxHQc39GbBLPZYFtVHkxh63zyEhyT+NWBlMgM+961lOiXHoumDqJliNz
7FfjH6jDIfjmz2A1bUIBY6Ym0iFusbfBCNNWpPiifKNHYZYtVTAZ8ko8zoKcTIFJ
OUD3Knci+WMtnXQOPiH6WF4+Ry1y6OR98vTOH5JHsbmAbt6zARs+bdZXNcRsAg83
jjHG8BN6C9m0rmWdexWMvSXXxPMejrqWsBRla7DZDCjUe0x239EFRxMmHcG64ghm
/zAUakQGIRU7qcJJo4/ir9YHFtVnts8tSH4hxhREAXSlM3ZX32CQHTHhqeAhGUjX
2GvYg9qAfMVVTg6k4hLWTMczyBysCGm08JQOjvd803/Eb2U0XzcKCaZFltvT+d9J
ytaCf84ZBi5tzTv/9ynOnVBh/ARE84rfogs6H/Fh/cAgm1EYrOBy/uEAbtUoBf/G
mTphij2ArdbSDeME4YnF613YKObGY4pIkx2OqzqmbSHirYgNYYa0HKCT8hLDXoQy
+v/6NyjutcGPkO3FVjIMsZTEYZYMX1bPCbtVLaNOjD+yCED/CXBsXWCiopQEfV3t
2vJ6tDV34A691gMTG2H1ZVE6M83dVrQTTOxTbWJuvaTLbTnSJjclLhZ4hiYL8Jo7
/V23VPBQRihByRz/LfonqIB36FTtY7KY1/JSEkuMHqHy+w5dvWq4yZ+SDLh7RU9X
2AG6Thsk1JQJCOpbtQ0FOxTIzr0ZzfMcpRW7k5NWyn+yvsZk4VFowiU13KlAUsOc
Qc/P8oy+Y/9ZYLOduAYwfHvtucYoy7im2dDIhLqvIVvzKGDjbtV8cnVLeC77x7a5
nCjMbzICu77Ht7/w7jiqMbFjzr3VUxTzn6HysaqlNVspB+utJFL6i0VOivzpSEd9
ZNFz9fk5sh83ejOavZ+9A5hIwUk0WhYkWL7VqaPavZw9acX8qukZMPc6LAE5fwm/
LBLOiicOMBt1o57ZXfBpoC4mqKo137fiI9ZnTcWYwJKVYV3sgG/TBAKjZPd8ddcO
Hq2Yg8YtUlRVEFeDQbYtA3Ors5jYSEIysyobYkqMJYnElE5+KUq3fJAQsg/iqDWE
BSlE+BSRyAhcTZ8Du2MO4gOaYhDg2Y0/CJYf4WdWjuKdCx0SXF5quW+2AQVigRGn
pASYs9l1YWYDrqg5VfMUMzzcxJ1L0RRz3JVLE9fh3w0+heOp4rLUAv3etUfr1jAT
8ZW4QiLpPiaVd0+6NIHalA7392mcdID5wQcFdmotKD0z6nyLHU6OuR1zKwh9DrLa
t0+YBV0iQ0mRqN7xNtV3KHQDxwNWeBkgZ5s/SvuwC2prFfNKjcNLqQ03D6MXxZiP
3gsEpcm9SNjcO5VRxN/x3Ws18+uhg/wRrnhjF860VjrgOREPSC94cPlwBj06yHGJ
4cpWwIIoY22DsO93WTGFy/KRcAWsjRirC+7n51FqeeAUdIcYVP/uWLwHmeWl8qDp
zb8INBpqL8hChMFXGFA6ytVf/yqLykFSbIu+iblxts60tv+Pc5/eKY+sgw7EQ8b1
XK1NHdOFn/hVo+7WYgiLEc89A8wodjudsXC4wsss3/tse1cB7UMyvMFeGR6S+X05
0U6gdsXZ7lFxzeF1QHRg3fDJlWuVrPVJVhhhuL7tV+XsBnEWKYbcXeYaNfeakf44
gca92bN59z+KvJ/U+xsm/Xs+ifV7PTEx49hZYp9T5rS+Jl/lYpSP82LC+8y/OC2H
kVUCSmKW31UIglTyXXgBpd/gyDOyqkhnmCb8UWxJL8TM7+1bpy4mwOyXCiDRLD3v
KCPatiSzhhoi8quLcwi0wGcp7UujQ/oZmcFXx/Ro7DfY4wweyOT5+vPG89FtmLvo
07t/7f8CrzL85Ar21u90ZsNqdqGJV/azomrQCCR21QeQSwdzRA48fjonXbpYKwi/
2SdAybfnj7cx/92BfEzBaQRzq5Qbw6JA5n06ol+btnjj5ryuAPGSErDRlYaDhjIE
8YbgliJ718AvChtqF8Dtm+B73RCcfc3tjvk6BgE7xwKdj6eNZLLdh8Ns75/2vnQh
48g1RnWYNIOzblS+BPvx0D+/tvOwRH3BP/sudT0FPTNyzoSNezk1A5hnnccMUidl
ZLxiMfh3RVcZCi8ZsZrEP3F3CAiQz0b+H06gpHZFTt5k99QXdzIn2wr0rJuJujeV
Xeu0iw4mHT9cHPRAqOri1Z3a1nKu3Kgm/KVoFhF/WWKZ+PLQ+Nex4p44J4ZA3jKL
42fETxIyhqz9DSVMW2VOQfe0LoJOIpCEz++lIwrBOLe5r+nPs8f2FKmHjk4bpKnV
GM9qdSCOSn+QR4O0JG4k5IflmbU95/2lAAzkud9jMzyS40zNzRli1aOD7mXxq1nD
mn2KdVfP5hUR5hbvA/B1PJQ3AhPc9scs460dNODMyc9aJH2SH/t017bvcDI9aphZ
2cpfNG/ZpNBpsFp9KAAiHrrO9kuKwa8EPxUzhZ9kSJ2KzTOyFQk5C7eW6aSO1oxq
R9eFIb+8N6ZJsaMI3pXMvevc9hgWT5kHbN59i+IIJrTQKTW7QNMYK0VoNu1u/72n
S3zxYdClU0E58l6kD+PVlqCVtMipV0zhousvbRY1aChyT65tKLhbMc/5tWpc9fx9
iYWiFOIBQyc79YO7IHGyNl6OBKduZizZRe5YtL+Xv7uUB6AO3N+4chjQ8AYOKt76
IKhSAJlInDOssj+F+9uH8Unz5JVrG095SIbpS0n1kG2ih5L8V+TTUFnlc7BIqGMV
NjJxrvflK8xatJ3Yt5esdm2mCZ1ensExUIBsNsdBI5puxNILQbDiCYVfIvv3yBP/
wUvcXVDRyhqtQ+7bxUvFfB90k/1AgvXG6euP/CIGJHe+MwVjwOSOkweBE/kWRwKT
zR+WhQq25qJi/ud1QqVIOSDE/MW1DlBYrE79J6YwSyM6i3FcTJQxri765cvg7Y4I
xBaumMBKp/l4c+XDQdjfHB6rt8DIHv7OZFAZtZ9LQAH/RUkYZKReZhCj7tKC68Yd
S2FUFOZ1IOuRel3qScaAOxaLHsMXeBs2PpdqJR228GQF+FEurTPEWKoukutJrjT6
mTT94Z5Ug00Ws9FSm3fxY+8q5meRDLwjEk7N4AuUgbw/yWlCiEYEdmb79cNnOBFx
VVm9YouwJYV9XcB4oXhaVT4cbum55u1NoDXWdwQEao30kSUPyBk2GHafprmZXkgJ
OgKOXA/nqBE0+r6PGOhl/vAlGR4o48xcf5NhzXs/725ku8POUO8mVTysJmIIzBdW
2ohkYUBedR60MyTtp0a7y0aN5+43KeBVtnvEyME3obGAf8Mbpk9exJJM/5MHYB8t
TL0E7JrQe7t/cjX72GmRZL2CJfINx4Y0aPFVNg5vUEs/ON5fFB3HOgR+UPMnjTqF
EgW1hGA37tqZSzjPFrvSmCG6lIcd2VBmtFo3YI1ddncN+Jy0N9VveuKYxSwsADRW
xTcQVbQZfCbNs9eU548Ikspljx1yH4g2nLtxMoRu1SBcpa+Xwze6QE4TIBSG7fCx
4hBADqJijkSTKlMLD7IdwprnbA4QQq4EM5QwJZmpXuIhImsZoPGHGjZ+CVM0nKrq
b3B5rwPqvvHvmvruKz024QKt3udfrzayDgZXEwAg8A78NyenRf4sf1yFs8BzA0v6
q/122d8UXXa/but7u+wS7pX5yz50potXMaZZBEjVhyNxIsGNNBa3m6QCc2ObTJnL
wUS4N85soN377trS+nyoB4h2z45y5epbEEeT1x7J7Xwxyo3UMZrPiQdLnf8MVCLl
Bir2AOYoRxmRV2nTaChtQp58YMfb0SQ8U9FxziKvHbClS3ztfYQabTtNhuE3X+Re
9xxVTvK8OkThn+mYct0HxJohiiGxvRRZ5TKLflY1ZDZbU48ru9ofSJZjW1a46j2H
qxjr/8XWUS+vFyZhKigoQSJI4edzFoaoWax+/i5PKI4milA5aYirqs6eCuBHJrgQ
/Vca+GE7inyYP5qsZ5JoBU+b/Tyhoygbwm4e0gt0Yeah4jsb/rTtshPrRIvFA8m2
T7jWhCVhsrSN1pGJCXSFcclsJfMZ8Udz7krwSawaK5KOq5SYpvXAKBSgYBahpy4Y
RMO4Mu8EkmQSxkdJLq7ArJVpRbJtRRnqtUFIlxQnZ+hNRlRA9FN/F7kdwKpj8kgR
ZUZJ1DxJMxzi5uH1kAlLn0shMNfSJcxrCVQ+HQAdCOWDsQz5aarojdZ7fVnq3qGE
5f1I+pk3j/y0fDWv/6EznAmKcH/IM+xYOg+QeB5U0PVKphQTobfRXe4F1yaBfDGW
lr/SoPfr+2XDdFn5FDyzBr+yb5Ih1hcg6fx9FHYfP4J23MCoF9NptyG3hMaSyL3P
V/D1gdoGQVvYLmsU1WTzTBlR6P+zcxKTQWzoBL4tv+YYIsn9He3xu3B+22mCOMDA
Nb3vGIHKdJwF17F+6ZdqPY7LaVTLqizJem6OT+dZxgVJVcMsSWzBhZ79Nzr6Xp8q
xpREwvqRbqV2XmTKPLDf4XHLkjUSho6Lp5cghsE9ImVaTAOm72MngSK2uS/vVlJq
SJX+utQIUxH3t4KPaW9uUA+BJxlZz9YtkLTwPPSerd8TU0SNMXYYAqYJ7yJydXrM
DMb+xA6UXM0b8OVZbmcNcVGWO9BTuLryWtmmoTXYwOJ866Q+wc9Idjyk1YGyaBaE
QHAg8rMxKVYSHS4f5GuxAUM/EMiYEivjfOeVwPfhycJYj/KndFd4UXOOmp5/BiB4
ZBjUQmg9Z/c0ZwoReGdkYlcxBBPvQBfzJgof85BMV0BQpsdRQ6nMqId/ynBdCa14
JeiExkhzpIhBjDFbGmwAZYJ0NJvM9R5Uxb1AyrrzI/1hVmHyJm9TKM/GbdKH/ZEX
xEvfU+GTLga8cDMhtR+C03C3ezYr874sybQJdH+HjFDcPFc8HDXn86gbBeUpkDvs
+2asiJSqvLzgB3XUCPUVNXBBbi4B4fTjgtD6kTVtWy8JZoDdDpejoY1veJSpxBXM
OV+ih/oBu3OisTRDNbM7g0aNiOak8EBl2n+UtketeLMKGk12Y4P2gom8Rtb0Z1kj
e2SYpYLOSlwiMfXcKlPx0y5aQG1Mg1gA5uxb6+op4KO5jHuPoLCRWTUGrmqhvuJU
YNwHSuR9sxUeJHPKxLe5Dvo3Lg2m87eik8Dqx+1sFyYCfC4y1Z13m2A0LVAS9mM5
sCM2itjo9BBgEPfVUb+9Uku8IKJ7bTIWPVeGTwTyEVbA6g4y82zQUZx7T0Lus3TT
FK8BRd4Ta9w3c/2k4RE78HuZntg+5biQlzlvIpPm5yxFsi9uyEI2Uyqo7R+NrXaG
6XNnfrvps3vJF+t1nDYdValVr5R3UF1K5pB46QprINd5KXDSuFyVFjMplqaNMQqZ
l3WpPrEFmyZh3y5HXoO7VMzDR5wmttg8UtDan4tGsZ4tmijKvvgaBHtUeUddA8w/
cMS9RJdHj8b/mqL+MUIDTLQ8yFmWrsN6u2vDgc6m9GiH2g2aW+9Dxl6rBGSriXfw
bphCubnCsviDzpkdqMz1k0SfADWkQuAGzRKjvKFFJEMSMSCnz5ww+qRfebr3gRWE
KbtMXI07mZZRqH69BoHAKvbQb0tyqcNeXltbz2vWzISRR3CNzBQQF3K6zgFG166j
h/BAJSAyczGft4BQB64kTjcnUJC9MZzDTz/kWrdfAuXPoaynvhx+1ETDA4l5ylw3
dKIgLiBkytHr021C/SrG9nTGRvOeSP6SksklzRL8GtEWvZp7Cl5jE4/SoPdhQbaQ
MDLvE4fzWqTyn7P8Fa+ggL1hBKHUkRvPbtV9kBP7PBvxtGN+oRmGK2S0/PskcREQ
jP+sYe4FcBwxrepe754pQ10HdKN/rV/SMCEc5LN9u9xFRpFwLQqOWj1+ZwmjAEJ2
TVWmmpPvpmxW2X+SppA9bQWwjflVypHNz/kdC1J1OiQE41GNMqhX0TRJd09FtKQH
VkHT27a7XMCixlgBamNrR+GOKesmcachQ+nnTVg24ML1XxIE08SNiNeKAj39Deay
yDfo+B1CoLyyZPuV8j65kHrMAy64HesTkE4ncVPd3HwcdwAdRxjuhe7UH9MVbRMr
sjQg8PKtn0vvBtfFqEZPjzPm3qhx8g0tloOqb4x6c2WdQLq+Al8RF4FVg62FIim3
/6yPVRmOsayEeRy78RRpiJXCEngn/sJ1Opa2yjfsZCizZKgaMmq6AKDcpwIhcWPq
r7HGkzBTWR9THmjuj5CKAZkPk07WyASp80O6wUs49B7roK4bzfjl38Mv+hsHCxe9
36MldaVuHKWTw50HQmxNuxOwtN0YFqmqS/W+lEPM0OhUGd815ORbylSoMxL83Zsm
yalf5exyIe6MTPaiNGxEvLMemlH/B4D9ZkfafQe9tnNjYo/A2kAuNUIo3iEtb+Ru
/TQT10Y2tCIJ5+9Z1JCLUcpHqrPcw8Pdg+CoR+cR2OiBj5fel6Prps9LEJnyRlsp
wK49hdRi04se4PQ9zjvhE7Nt94xaSycPsKVEHTbbCSXRLuQDSgXM/OZEPrMBhvZB
aMR3C1mQiwz7m35Exoekt9tMiVbyYA6oeYR+0Pa8fUmodDU5p0KBYLgg08xkNy4u
mP+rKaMthqSZ3N70vLRi/HTUHpD+oHAFrG1/mjIrc+AXs+UBI/RmZUqLf7xQERnn
qQqXs+jLi9cD7CwI3FjXmO7AMo7Njq+ka6ouMm1o+XiFmQsCn+BWHOiGA14wPSAH
9b37YwOGTSK6sKAJt5B1XjwnomZV6yPPOW+esBvqI7uWwt3hQEaBv+Xe1/psrqMy
XvZ7w5M4buhnc80izu7R+OspGrMRT7On6JCIIeLXuk9dr3fsKw6BJ1Wgf1NyDDU4
qrgLhpXmyoGtnn7tX5QufoTx0gPZOHIgs8dzXGJhDaldHeGwLAWvAYX6qpn6LS+E
Ys3ttQ7gK2JK4JbN56SOs/7AytVamPXWmJUGXhVQU3yUwkekH3loF6LCZYZXUUK9
jwjpKJ8lQVYncj9TazlTysZyHODlYX1/tUyk3N1qRIHtlkr06nUnkMQZQd7iKFs1
NxUauUnuRBysHAj6Y+3DtsG8BYRgSGwydsOD4r8NdNB1LMnS7syWwFVWAWwEn7zs
Pdyj+Q4AWO0MBonXCeQTkbMXkgaXwGn4szI+pclZI2kiwW3mUasmB/Bb8V7RD5QS
BF1arj754Vh2bDb/u2BqtAD4VQVRYyh1FOs118LRPnXBVsM+FYIo7n2b2dQ4rzjL
7Jqss8vECjl6t9RtEz6O+eO4ESBg/hJJrle64hdYVBdQf9N5zzdKL49WSEBFMTG0
CMfj9b4F/ZKPI+2cq7QVLflKZ1iiGaXGcWfN6SjlBr9ZBJBZ/onjLwzdArIaa5cf
e69YWxDcIndftZv5u58IwyBez0/dpisYwo4W5PH5fzWfqzZ5YQGWElf9GFzG/SXK
yQTaeznBIDWDG0wWUgsHiAHYiuCMyri8Voue5pl2Yu4cHpRhEX/jqvX3tqsEan+8
wj2QnJTBcGR7lfYaoDhH+FTHuZABhgDo7JCJqZQ2XtbmWPxT3yMQ2ls5ysjVSOdk
R9EE0KxdTlTnFy3rU1VBr5d/n7TOGlDpmbRMZR/rvlOOsx3eyJX0YzF9bd/3ZtTr
Jg8dgVwpkEH+Nd3QmDcYb7wMmesoP5/CGFrjGT1mK3ahtEQ+xj8fPGz7jHBI5Msd
BkIi7VfMp3bywnwcD46tfW2amBkPZgqojjHqIzwFhu8M1N+QkEr0TOsDXSHrwFdo
Zm7m6TERqoCCtdhZX2RSL7JIGfbEnWE8QijUStY8AFlnnfN+AWM3udSl3u98JK44
yx1UUVzrwV70rIFRE73MIRYQ44KUbnP6ECDbV//7a1jfys/KOBvhPF65NaiRPvn3
46DHqxOfLRICZ8Uji2lTnqvdNe2iO/Dm23YfZPFJ6x30KpSFoLx6VdU+88Azb/oY
nAB4nmNTqWrg7xckWJJT6O9LqaUZUHoxQaeAe6SeeyD4u8WrZu4etn/3oFQfJJm+
GN+XpeqEo64JimdUM4jASDA79kj3n5HkiDmK3Up2M1r7IW91HIb3P9WyQLEePQKZ
L5uoFt6YharJtJYCqEbdowN3hpCo3Zh+wzkdWLu2xixlTnyhDGojK0xYy/IxqAJ9
7sSBml037Il6YOOGCL1WJqYyon4t59ZFh/R+a4iBtzVe7ff3kIXtRX5u91mJu5YY
6nF4BlYAiP4v2/uALF0ln89Uorpmd6mu+XN/CHVSff4+xFKz/d+XBp0+V3QQWvzm
41hGBloT/BgRag/jZ4cI/bmnBQjQEDsh5/fsaXaa+xrlyXuMRXqo5Izsla55IvPH
6BFPAfnm4ItCMZfDkUTDST+QXg0byXj4yt1cik7Kq+bj45xXkJU20Iiw2r/Vdltl
eSgbM1On/5G74if0Gjy4oxZxanWsnP3iadpOjEMmTNksVwgAYvfozxNI7iQTjAnd
eki82gt1qx9ZBAwrC1JxYzFi0E1tYBCDaJE2DArV50nSONWU2hW9qpG6cNmjWZO/
T1oituLVEOvebl2EWN3j6pZSZew/v6NY3TtLOzSg6HrLme6crjIItXY7bEF/X7v3
QwdXteHbTqwpQq2LIDGVGRfLmN6HaTFiXjvNUwHjqRyhGndsy9aH2CiGnuIvrhtQ
QJdmATYYlIyXANLJ3dRYqnDSa2yQtefMi0436sv81OMnTrx7t++bNyAthDi0s19D
bzGEIOKjr3ICPinnqu52kbq7tVIGB7cgY1ma2MmXPcqR9BjzgGpwkIVJOnLEXisT
c/vaLwCse/MKvORlaZEEXK8EFLChFBTIYU4DcqREyZBwu2PQWWEP1dlHCGz4Y4Yc
S7UfTO2uGEHDYopR1Rnmfqq4N7DM3YyAoDVSctpS1rfQ9MNbYNj6AopU3dNmLZ/r
+MUERFXDjw8L1h1t8i1OBCRa1hf5It2HutKVkc4BQb9Bn4fsdJQm7w2rRMKKXUtc
t07kGDgauM2Ak5XYKct6cyL4SMLDSoRCJlH2kwJy0EPHfBN74dCf6p1EJD0KMs3D
UFfpUAjVD3ZRAHA99lPcVyXZPW9NlCZ+qmICFh0JvWzVS6nD+4MhWfCp5/58w5iT
pccprDbM7o0FFrQZeAVUc0Z1fj2ZiZMxZ/HfsnAj5pNJGE8lhnLfQgaBbnomGHS8
oYq/Wo4ByjQixumQWD9Am1Kql3Zj8lqdedt6Ia2ckj14nH3uDqLOQZDpZiq2BeiQ
nIoXcFMMCZLbMYdo1NIDYtsrS1GwezNs9H76nJl7E80W555njtZc9udlUMMmSoES
A1TcnCYux0M08BVH0btyb9wvpu/B6IzKRSlJ04QaF85PQavUe9UxvISxR2mzh7dp
O9iDHhZKmDHUO4AlqYWzCeAL9htWND3d+DP6WB13vKcaGRpuc3M9hXcttugBflbh
BJhkiAQCzxZPQWFV6cbojaAEXJ8L0s9uJsym+ZfUCTugbqnkmVCjyOZKwNbAnysJ
Rh31ROLx+rASLDrcZxLgRUn9nIS+TvareQ9y9cEUJY4lY3eFo8CrhP/NvUMH37Sr
9ktvMr5PeQHiYEOgun/3zP2iRtnlms4pD0hD/hk2AOW7QN8/IbX5IKfSxOtgQMcG
kM7Sq018DhsNCLgoIV74wWVoU4AUHRBX/D+IzLvmkV2vRGLDTmx3ZcXvtYF9Oju/
axHKxu4zd+gTvfOMAo5vStEAIaslm0xBYF/jUXLK2Zn2cqqxsNM2QlkRggX7nyx+
ac2NwPH0DsJLs2zvPg8Ua9Uhmg8vLYdAZubz8rq36zV32nhHk1hE9jl5FpE7MXFU
nl4+OFzAcETQTImBz6hRLkQclFtjY0xVDSub88X0YgVAgzkEsSGv+hcKbFVDMipd
g6zAQATQC9v2jpINTXH6MWFf692weBXeujczP8XVw1AnkkrT95/wEq/WRBHfWm8S
Z8DfykHWAoZKYzkpj4qxLoSZxp14rddUET3BNilJyBtZSrEWg7Sjazo8ZYAKOSYW
Bgjm83JGAC0uJH9IGCCpxvF1M15xhKiTVpWW/N3dteQP7kBwwdTQwgSaFnL34pkD
1UNYeaRuh8Yl/wrlFg/anlIXF60zEJmqV7BN9O4YMJ31B3xwXfiGkJ0PqWvds9+r
BWeiHXu1U/MF7LHryXct6q3U0izBJjDZIwHAIWdHxudQ4Tv8dcZLzXP3/sjWiZu0
bHDlFMwvM5MbzUI78dB4qfgTj0rUjP/CRWyphwntKInzjKKiOtOgRt1KS0dIJBUG
pmWbay76EiLLiVtGuEkclfYYO8oH6K4p40kcZxc47yZw0oiKhdDA77Q/HohDrSh5
EHDNaOxH1tUy+Ycs1nXKyq+n8+A+RzeZdXGOEpfPvibQ5b2WiWaAnZNk1B3Gc48Z
KZvKFYMq8lEk4AUnno9L8ZGmuQTqudg/pRAHADhHitlGcfbeYX9OHY04KK95Yq7+
bq+BBNxi5HrGkKlmgZ18xHiP1SWxiWQImk59OxvDvq+Xyf2k9UhqmRyY/XV4zFH2
uqjunANI0PGuLLKnOkQ4B2ClIp0u0y1xERuB0PUefSz20JvCX9lJwvsaHNF/UoCg
vwGx38Z+AD/Jt3BstzOT+5SKKol0qNxAiLgn9eE5/Ib0oIb5ybxx5+LXtDn74X6w
HJk/CLD09H9flXKbxpLbmxsDerr7u+lPR67d3CFssaFZv9gJR0/1lpmtxi1/5gSO
wkZ/X1Bfyl4Ry0msoGN4e0stLh0wEDlWKlw3Cz9RWgvOU9u/Cs/L/gZx4fz5Fj/U
+3PH6lnnlZEs6wpo7cq0DKjJoQ++CvWNhEYQNFYDdYAN+o1S6RR173nYB1rjfAJt
E+LcV9Yn4+fQArd+nbp9WUkfACOLUjTZUotp4l/dp0t4Lhlour4en9s2T4tHU7x2
JLbveZh/ml62L2mZy/YfgX+VygPcyjSHOlTgKtcZVimkPFvCk1pAL8XcgnB/V8eS
PMCdn4UkoKDiYgSq/1UvXxao6rA77nG+zI107tWA8xuOn90M0SoyPdjQ+ISl6cbS
4EIN7DgiPWdQH+r9L3+S/hvAPpcoeeaZUCMqbdeQRrN6x6ZI1BERHoBQYeaqRnzf
H1Wv7eSPjmVF52P2UlGnywNlMRwm491t36y5QT2P8/t6MkWI8gVPtojjx8magE6k
fVoWE2FSgs/sR4QExQ2WcsM5IBa5gANmRKqe7fYjxX2iiSGATSYD8drCovDhFJHY
cHTtd6ynk2ek8z1Gj+MPJHt6EigoFxXjPhRBw2+ALS2Lqt7G53GOdwIBnoipBhlI
1V9oT+xdIgrXvuMu1iZF0JxP5rbqD1oprpCi7lH+WW7cMFeaj7f59SQbzyYxKe5G
mqCuIQI42O15XiUYLTbN4nW9YMhK1H6axIxkZlY+9LUFob8JVdCBgmudDhE/gPHv
6yLIv9EePcXgyhb6Wh7NdR4QSicnBFKV6gdSl+5UD/K17MQzvuEHHCjeW0jrpVbC
qptKORgwwalWlHmQsowHT1M5M4yUt6tqUih/aaHT7BFdsH+aTdjz9w7oiiNL12lC
rTzE2M6KxrVnORTCajehTI0JBCmHFghvzSVGdDA/UE9LZU3PC5CZluynw4Ky3XOE
2yEqzhm+HENERqrJDYeB7aPBQw9fThcvlyDjZfSvARzhp5czW/uZj8UUrUZH8l3u
oRHVUTqpZC0IyNJWDhfVFP6hMuEwqvAzKHX3pqN8YnZe0vagothS9yyOeMkWMdcA
gJltz4SDyp1XdLSd4590zmK+d/Z5eVVxr37kJQRqL6HLZ0j9VXErNKLqE1eVZ8y9
nRljqZeLaR/vvWR7NeYT113T1Xvam+Zbb7brZ4ReD/TYt7j/u9P0nf9jw9DM9uxb
4IwLdIIVe7juyEMtIV1NXbdcjpWfrj9YtOW+mfdEIWbQwXYPRsnPoJuZdCwDQurq
2Xi2JsMduh+UA+t/E8sYr9iyDHxKG6mm7QH1/oMN5iYLWrFcv0QPYUAOm/Aglu/B
osngIufH0ftEcLyaHXc6637U/kEU0rKbenOV2GUNtLmanXrTabb+X2TNgfm4Hraq
o8vS9ZYKXL1blZoBmBKTmE8TCyD6tYYFzEmABj6rlezarB+m0AoJZEraL1ImDfyT
nysdhWHU+YiZiGWg2Z2ix/Srju2AjPbsOG+A3KT95fNxogyXgpDo9Du7gGi7oZEC
voSpWOMXdHSsIP82WGTdjo7YLHu7+cfZ8UKryxsx7UUbVKWXezn7cMlr2LK/430a
cgC5TRHhNbV9/PDRY8D7wuT9YlDOE+PM6K6XW/PHDhTo2CAvr/Iaa2dDGC90DolT
yQroxrVpeaHo1ZkuwGnV2wKfKzEsRAbUVBLGuc1k2U3RySKLyV/qAJqt+7sobOWw
I2bhdE3at56S43tWOtyh/uSqKBft2mQgKDMVQg3XKa7wgAXr4nZfLNYQEXDtUdIW
i9D/44UxIVV5hEf7/V34JjeKBWDSmG1t+p0jK91wfegwatghc0eIR6XU2gZFbLOP
QWE7mcl2WrRuY1XxzTsqyaxhwcjionInUNaQ7AcqOrcJsuZ9jDGATbInz94Fu8bH
A03OMx3/zPqJ6i04awCjwoSmuoPW8+p8bHajgtyovOE2FJZNPliL8OMciEGxJ44U
EmKAzhXmv6BIBSFMzcDHR07iqxXCHOjO/raUE8cXDyE5F5zGkqqG655bWbtRGlx1
7MPe60T/01eOICYBmAcNpOPxzQXa8Qtxb3H3xOmzQ7qUBvILOZW4A2dDR0jALEGv
DWbC3OBZz3BnrEa6eIytc4a+5Hm90Pjno2xDdzCWafKjkfER1XTzdRPz+AwrV0j8
V1JOeuTDnEdehNvfKg5Yk7exbYVS1lNWgQUvKBcaRdERu2jPcKzovGFCXxao1TFH
8xPwbHZiNihhKZxO+Xu6FTgLnL7liOlDf0AoogAHfY+7gXRuMmJYn6DyVcW0fP9V
8FsAEYNamn6YcWOVPQCM+haW7N07CrcDBwR5E7iLfN39sfeAC6M+ytN78TpG5Vv9
52F8zPQ+Y6bMT0u5C/dXyN5EsDazbeb8lZGhstXTF/HA2uwGrAiU8X3OxfCTjGmJ
Xk6+wrfcVdaOUhIDZg73+lBSK9ZFpvSStJfgHGuNZnCUw/RTSeZBbQR5ahu+j4kk
CihYgtiTdXls02OWo1qH1Jz/y1tshCxS7TUm/CpOShNmnASQLcr2xp3Zz7UJBmTp
Zf7f1kqEJIkKSqFNnAkqpn51ykcTfEGkWp6yEDemnApjW51EmS+i+o+dzLL7CFpm
DCCC2rFLymeewHS1wd2hud+8BheVGkA6sOL9RxhiHqFIVVSxpUEVqUoR7yz2F2RM
lQXPtxt+5jGgtNINGZgrHDUxEeI8nGNTGjk/0EiNI9stMWxJfZW+pWGByWIwPBTL
ZmnstiO3EVSKojaQuhkk/dOO6lCREFGz8JZ4HfM0HwyROjlUQDVzp/xfoOzbRovL
OZR1rQB4KJXEaQnTA2T/7jekpUe6dYmNK77DX+DZv23ll9hXEh17mL8mNKJ4h5P5
PelW93AakM+UXxWGdxxAgsnCrPh8sEToGu2+Cls8KlAeRPtvZyJXlXlkAEgzJmpx
EQDP0EehFTr/OA2POqMYBuxRp51S6fX97PwxVar7jz543KPclQTktQgVJDdGjHyD
CJX9GfsjnakefzrfkVg85uEhxRz/Cd9xZ8FLd91vYceWc5rhh1Q8Y4Ss0Q9Qzxvc
U9A2u7NZ0D5nP1yiBFZ+uzTSGLdVDapBKWEHkA3gSQp5gdkwq6bEBNkKK9nkp1It
qxbJRvn67yLzyNBhyMEkxpEChZtVg90X/keXfRgVaU5v74rwaXlV2ecmUqPiXqce
fGLJn8YXTk6Zi/nFHoMjZB1l7LxfVZ4PkidXoXRGHe5gumK49W/mfxti06zYyUAK
uYicfJzRDFVx0mBphnrtZbW4i4uBEONw+Slqa6wi2TqLAwopvdPMQlcVkxa0JEhp
npZ0KV1gtx1pfUZyviEndwLPBsouqVf7EyOHgwWTZhf0zf7crGLTrWBP0l0o0r26
9zbtrVXwM5PvJCG+g0AiphXAl3hQ/yOrVQYeYWLVbh1VNuRVdAZ0nyknfCu7Ka9n
KTyjTJYp/+OtqaaTTrG3j11EhXuVq2F5awv8FbUGKLnJWCFw9HlGeuvvH4LEI/Tp
M+IQzCQZJP64hcYZqT8l8IXklgfZplGYyTOgVpagslZ4RTsbuoJ2z1t+oEAL9/Vq
9DDGp3N8HorAv9k4DqPtHxZIvM2RCbwwPV0ZZVW6Dt0jcUGdhFZn8w1EJfxH6vx4
Eo+tuBiEHbwXYK0jTistCEOA1NiB8YdNIWr/spN9oi7GoAdhrPXKB/uCnNZj1VHT
+iMUHNN58mcM4VcSKaym1pPlcBbPJkeDlj+V+2i/kin+D/Pw9BuV6LsJkpHLV2rl
DfVX8IlzS3HMcTuUqIlUn4F/HEvSK8GSh1XRo5AhXyabtTOivRn3eG80+sRjejAf
zCQIyIVxcpYlr/2W919kPF5bWoNtKGLlmi1d/kItvsYbfFo29jqo30YflRzI8Ulg
5GW/rtWtJuRQ/crPcoRvp1TzIOicppsrOIt09tSBehGnmcStKe8JSTOTn0Aa/x6p
ACCmIm4BtPq78j7MoQ3qSdqEn/u2jgsZWs5PLs1HhEjUqZrQmneCvrYCwNcAFd6L
YZehf1UL0st/6cBrfRLGSBVNPpCP7ptrJcKDkyiH6Cdj9nnFgZFcsMWvtt4tF0ed
tEJytvr+BlRouM8QZYMhYbRITehifbNQsfzYM4N8ZRIMZUmORdnuR8IxevKtjEHp
4Ng4HAr5huBYu2wbMiltL72uOFZQ86gLtFukG6qtmEdJ7hXZPYx0TXBn3tqAP/4o
IQ6OhPx3KOH9ySmlQ1cEmKykAWTHBUw7GHNxDQEQaYnTftseL8Nv6K1Z4hlIXQ87
bIDoQUWrLll6caICUjgh7TasaB1GxzWjlXx2EykLE3CB3P1tG3+BN19rMEVp8Vtt
qD2K0DucN+dZz7Oi9Ww2pyaFRokTFcNkOpNIWFJJ1hpSncT36eL5UNnah12qfA1U
Q92s6pFuPJVQHTRJ1a80q9hfYI6W3uCUQVlsbASgEugby4UZ0/iFjNb5psnGfmGx
0WHnMvWM2kT+4Dpc8c1QrWO8Z0TTIUC/jz8k4SLh1mc5ucIUVLUJKxP2N7gvCOY0
C1uj5TdiXZwA5+IDEmukAnCU4UMGRiMbEoOejSrtAm+wadMB3heKB8suQ8HfNVlq
cveJB57Gdj8f1BdreqNb0Qul88KE2ce1RXxzX20kd9yvCJW74zXtdtOVTR8pRS5m
pTIx0pUVYSUp4u9o8ZAK1fKxED9uq9x00zxr31rX4QS1zDtWDQEH+rcrVOwVlcY+
NuFt9mu7VVAevwo7ekg0LC4Crv0SSUZ4i1vm/RVMo2HsfCuHMlh80LX1J4ZDWRi5
0IeVWV9olsfTXiDGBQYsJ5ujOeVnLnNeaSSb4Erus28zGu2fYqMo7JbQVv2hrzQ5
DZakX4Jb1kPmbO3f9Euv/3FuiOBbcs/mwy9dNhkrqv7myWW9c5H7Irp8msr9niZl
ovYlsXV2NscWhs1wV8F+gBuWNnPffMUpR3dQBFcv31p+/FFn7zFAVW7wLmRQgpP1
TB56Aod3f32SpK0JiHf/HCFm52jP7V3W8fUjVG8SHpv/eoggFb5Y0RvH1mXikhN0
q1Ircf6bcmM5Hj1O5GYSW4qk2ajHIX+sI97xz0V1pcJcR9cGRidkPpBxmkrf7PIj
lY8lDH5FSGYoTTVm6GTlErip4P9SWfZIKsMSv4ukahgEdZ8jFBIJ+LglvuMYENoo
N3S6VUPvbMDPG8IdfuqsWVMxOVz9l49Wec0Vk94I6clSWsDfMrUwXzp0lbHwitgE
iCecqHV9pleDoJLlHkmvu1ABQnbqn1UlbHwz2rvdLbjoGF2aBzdUw97shAxezjW0
6iEFqTI+3ZT0IEpjOtp2+0ELYDG4PAw6PdMM8jq01WcHEkCNntR9p3dU38YK5D31
W4ms7FWxzlC42dEOKFBMxfM2MgOccDkoVa1eeGhYoNB+56vhebE6DJkooJncMuz2
5zYpz5s0ywyFYp09UN7dR3lAUkY2P64mDSigUOKiC0bX4izDoAeGHBvGV6Jovh1Q
JxUxdWYwFGLpgvdS/2PoP/uoWOEx9TJj5pBCp5hxsIH8fBwFzhMCQWySd3GsdOCi
jG4/v1P/hKvmsHhN+9Gk0plLOiSDA2giTgP/eJym19NVUfDN0Cv8FNvduEeyLtB0
fziXBxZKQpeXjo52PqLrqmyp7wqCyj56JDgUh3JxofcHaFzC2YB0K4ZhNGeeJWNP
6TmMHlhB3BrJPB7nsDYlUrfqznmHteyrZobcD79sKPYSALZRp9y8h3bfy39Ab+xY
aO1PA8hCj6X3y8rKfedm/4qHMAHs5HWIqItUa5cnGkZed7jHlAO7Ww4QwkgfWXfd
K2/4mFwIe9eZoVf4ZFFrlcC2PT0lFNW9s7AeV7LHs6Bd5VktO0UvabswE6FyGMD5
Vutx+wBjMoId3tZ5upRWaoBfBrDjDh7d1T3NPnd1/eXd+1tl65bqp+g1sBk05DaS
MKfkzG7eyrHDQUjAE8CDERZkWdhsZLp2vxzabOGIc6O9cpNvpSpunjwT+vIfAkVV
ahTcXKhjjZa3zjySZww1lJb1lOD4enfKItTlPJIBDAvNHOmKLmD0c51oELJMuxFg
lY1GClZZboM0vlbIsN0iWsSCQ/v+OOivQYiyozi30x2WjIGbZL9jaIafRxAfYdwl
r+bfjWymVXZJLFsVkCnJgcGLAVPevSduuLorESd6P9XyCUb7wQEYDiCGKzQbLo9y
FWtP1M7Dp73EuKstlbbE0gx1UHXezo65o0K/3ITMIYr0yxJMN/gvPE6v5d2Ey7q/
1Tw7iJRl62Rw5x0qChMsNTBdAUlibzY25DCY/ueTMT6aappOiZWDxR4WBXq8ut48
omsbhM+oRJTo7qR+cg1Ep6p3gaGRA/nufEzIsK8OfWMid2K9knfgSuqfrN16Z1fg
/h7eKQeNIyp4Sdm6p+zWEZy4MAPlVpEIPb1FCQUxusbNZu22iQUKMDHk4ZyKkEOI
avIe2SU2vkS/xb+cZJHRE6EkhP5cHvKl5ypSFyF7ioF8vPG2pLuA1N8X4ee5LPs0
sWImmIb4qNHQEUTXBuGjVD1556mt1wD8RqxIPfKPrZriIDA/G3HMAirpHxEtueaF
YODClLSF+Z9BEL/7C2ULeomRe8AxQ+Ygsce8ANHeDklLHJQ2be60D5gok1tDF6Ok
T1NCCDu3BmP0WGLL2HmH/KChkdWAVaHTve4CkFHNKB4ghXMFAS9gl6iqPSDGiafd
EMlvXtKWzZWJ9u1HHKYu3zYtggNQSdGop1Ey0uPpnIJ5LOhRiYq4SmUk09tAFzM6
Iy5xjx0188pVSuB3oR+P/s976ikIhYEH9IsG3HrjgLiGBaTQ+vr6uIPpfHgJk4OH
SgbRLC63lPTtIXXmY+FQ//jGE0tGz1PnoxTkxzkcwi8MDZb8WMZUJC8KO7apGfun
LxM8kUWuLZwSh3Jr3DRQhNsINI0XaRWOQ6PHik+XUtknopm9vHjaU7YcNcaPArI7
lvHP3anxRmhliH1BNfhzZwbCoPZE+tPXtGEaaDKd1a58Pl8p+QfuK+WjC6yBpu8L
XU+zbyv8pNToJNuikEGNrruOUMp3B7OrGjcDXRFtUz6D2KYNp28r3AMQ1M/CtPAw
3F9SZebLuu2NuT0kWIcQhrWLCwNFEE5zoch3SEL2V1rZGkGBPQtjmOHS56zi8YYu
rjsol7NQWmCdj4PZ2jV2A3ovi0ImgiUCuNAD9RZbUUOkVSx/3EUywmNgzSOMjUaz
ciyDwbjeP9XthwPL/vy+CuZukJKy8QRMbc75RVmVT2DWny/zk9yhx7lFh0WZqRES
ehEs/IMxCJGzWN+6NWM+Lw0ixsNYOuO+yivXjcPabtoknVVvvAOsASlejBl8fxmt
ed+62ZJmt00+tF2rmFK98XDpeWVgl4xxX45RjTeIukDjEW0c6HU+onwKVlk/xkgm
1b5W9UAEWjWaV8ClxitWcyxi6Jeg32vfmQCsczKkxyogMJ4WoJoj67SNjFSi5RGJ
f5MQe3+TvFCOJtHCctl4tNxSoqOfIj/WDq5Nes9L3iqXq06+jPvve/rCV4KqAHtO
FQUQr8Ke5zDoqadxiUlUPpOoG0+f4LuCxBxXQZ4wHRAZtCeh8snJzGCH4zYmDLEk
HYwLRjdFcQqw9qq9ktTsnQqneCgBcxj94zUx4emM5h5Agj7WceHLH2SOaicmLwdy
kVAybjCLvlyInJmtga/R64JWIoPNbqcnorrrPX/UXhfbMO4m4ZBaVnYbmH8KWmcO
ODQ1V6/tBNkeSlU+X997MVSNH/QiYMwOahTSmuAVE8BcW0XIEtbMOfXQ2GyubGaW
GKUma4GMkcuxBH+msA6sHDIRk07j+OJAi17cGM+JdponRdns8cX0H4XWIjdZoaZF
f/JY5R4Asex+MOwzSYuxhP93F/aAg+RPwlP46Y6v0JU5V1y2N0p30B2KFo+COVSK
1qCi7II9yBZ0QiTxS0PWhYacTN1KO141OaMXASLfs94pxnJ6woj/v0lKBZMZWIzh
jqiNJpJefceo/RLKLvcE7VS8v+g21pLnEdZD2q7XoLBUVac/N/13IMioKW9e3MZb
mzy25xQ7h8miG31CEO28saAWFedeS63AIOMlIN0zS/at60VPLvvMfdlqkoROVb3j
PTK6PaqD+nzhK//vhVZKpOzc+wr/M7uLI2wXC7Gvfk9lw2Y9SsEYkIXDYN+VNJ+H
5KhJWdjtvfbiBWHxvDWnIa9bXdkhlWwlNr1pBj9HfvFeuOUzWdbc1/eP+55IHCry
H7N9xrXqlT1J1nF4335yycTppWu9B+shc7K73FcuUDJVwgphIU3GaO8wXwCOr9bU
o9D6EOd87qCHcJfFnTjI5Est1NnlKeAU9+Idn71jaMYX/7/SCqAdHbysJjNTYQ1C
qOkoM2HzFsWr8w55n6VHkCRdf1unJu1br1YbcfNsg0pm063qgl+fv3Fuu5Ojcyju
NVronwj+o6/mribJcJN4RYflyd9oDK91zUKKXVUzCxTzBJ/uxp5E0rkEld/0YwCo
2vcVRqTIbGuUyTUGaJRoQTajuw4zxghR/5KJJzpVi4+vp81cs7aQ0WeNmgNKI4fw
RKi/GMCiNHdq9jf2OQchzSi6rUWM8OJ3DMZQ/5sm+0LAYvm36ObITS8k6LC17OAN
frzmncLN+3ncPxDU3psxQTbKRnQWOaYsKNEqxxGRbuPEBCPKhMNuDGWG9CE/EtKS
vdprVjIxwfim82/ek65SkiPLDAt8SqCzjRsivjk7Hj6kd9ikYCRW11xozOBpISZE
wXJGno7p9w87vAk6ePxA/HAL1i8VIlA8j4sL8Gb99rNqSrpPKvW2eOe6GZqBdbtv
qfpfDjbcHduLuzlJs1Ag6x/yy/gu4GRGqTLghVwUDADh294xXnL12fNFM3hRoeRj
+pjOJJY7dlnuCDEDQXb1KxmXEXSEgyg9asNiO4p0hlB6Vn4QI60E9gwoNn9Plyn7
ZdI1glzhbob+uB6lFLSBMCiLuUTPS8mRPx0MUGqJ3zgf17E6ZzDVlL4fFMPgVIQV
t3uJAFuJ4p2RGkiPlp6lBtdEwLaw2PefLwe/E0zOdppYS9geovWXSlWt88elZWtr
m4H8t7LGIVvepBc9Pkwz35eG54mmocCwuJ1qIWm6rcSjwdHlHDcD5HAwAfqRMx12
KcgkSFI39FblnSkp2+3jXxouZvRnbVB5CzCTxIKIuHhDoOu8Uor5FfnHmQo1INCX
Ec7NUmUImIaT6R9I5tuMwNHGqLTz0E5vPeYeRGGEU1l9uwSRs5XjjkEzI1z5GaCo
RVcIXwcrwsMActKM99WIx2ulCkgh06tEdRYntMTlCHg/1uJmI/K+XMiRsBl7nkZH
2zZFd6Ux7Vx/O2o8e9SM+T8QqAC+Dy+bADas6cI4T9aashsLCU4zr0PFItPP9BuX
iUC9iV41QVS3ET8EXiIsXP8JoKXQ7H2VQ9EKGvYSqR9op0uOgzwyCr8AZ94vOyuu
ukve3flreoCoX8fgYvNcPQUSXTfNyI9AUSkKyzqgx8GyDwq8p0wzaptsII1s29nu
/do53TSiSmo39lhOGKwhcvy8nAtbj8vIY/Zu1dZnHZSPEDjx4GZxXuqXec/FS6A7
HDiI98PwLFQLxoqV7bJtzc8QfUzqmIM9+WF74IErehkHVrRunRVuwvS7ZW7S7Mmm
piSqFI7jLKu7Jeh/H3Qg9PK1cmk/BbD39abKBvnwuwkIk8UnKgy6LmouIXYizqYP
Cw5jAqFvlt+u+uVch+bqhOHT6M6nZ6eEgQ4WspV7o6yBnJu35o2nEcUa4keZYb1o
eNm4yLPBIebTRFg//d6Y6/X4NDlFk/JdqAfXo5u58fbgmAbNPV3/nKR6yT6YYdo4
FNuASrJBW7Kt+ISuBdpAmqCBYht6dohOlkZXtU3zsC+YyEHuFl4CNJikcsyFZcs3
7bMfZUd4epF7Ud9qQTid4pRPtXCUmHfARmcy89Dg8Ey1gQprNSmn/jWlVO2OOVLW
nHQHuaH6DSdYoq+jtP4xmio/wvvorf0rrsG/nmTOuJcg5RlEOpHuXFlgqK8L/ktr
roiT1JU674YuNvu9xz//dNWUmjeFyaKPrbitGHiyHFM6sUYoNRdO7iMunWQbf3Mv
Th7zIsEA8bbnk0F/GfU7H0j98ApGBDQNL6YjilyNufxKmqAk8dLKSaOMza6OPy5v
+U+PCy+PX0U6z0TrqxZeFTjp32qXQ2N88/IaVjSzTPZ8QjU7OU8Tzu+qhdrUY8ik
lXaXd5cWZ2p6afnM2gpUNOKo8ZIYFxyC8ybhLMn1MJvnzbiZsGjTp2vnHsjBg63J
d9iFG3g5E0iKwZXNcl+GeopQLh9ETokdmbB9GRnnH9sOrebim6W5y9twzS+lEbCF
g8yWEKD44HIf946LOqbJGU6w85yc1oVxUTfVJUsiVdlQh5rdmOmJ6kjmA9kfNBfZ
Y+k6/S5oHvzW7z6oKrXEDN1+0K+yA0zZvIroJWwGcD7Vxh4wGewKwi+hfj3szMPw
8tSJ3g+WIdnpeDvUQFz4D4j2leReYmalYn5r5csAaobv0lMSC/3E4otAPiKY3Mda
fpIseUNxUMYdjZZEPQWAyTDExru2YzeAJ4Z6Ik6iA2o3zXy7JgFhIknhn4pdopd/
z8o7+qz2BwvhrqFUIm4cnxem9eEIT2dXSG1YPjns7zGu+/HOKotacVqpyFFk+57e
uAGA2+AdXsW54YGvPsz8196aMYcofKDZ1f3ZfJHpGNwsd9uvS3gl5yxkWYqlWpjC
KiSOyfJWeDv/IHCuWuDkiJPC3SFd+B9ayohRConxHWyMQhSwm3qI+jItF7DosCxn
r8qvVyW3AP5A/gyNtg7bpmbFpj9lz5IBX3pncIU9n7s2zZixaz4pp0wFk9zYY2nc
Dvt1+sY1x8XcMzd8vssotrQkjxaqp/JdRrQuZ/rkSnmzjSMH//LCx1mrff82a6JC
qfpAOJGEh8O7dOT2URiq7cfrOCrDTVSlPTfbo5VztAeMcflbUEPCo2pIRH+caznH
XoesHHI2jBfatRAL07Psnp+sQVT9zWuzu/arN8oDSjVhH+1Buy8m609E1GdlbMpq
dYBgaZUKSZ1DXNuz3xbEc4vD3u0bgqz3PCbzoeMC3cLnF9fs5hf3phzQFiUJKyIN
VfAo6S1z7EvR8WImqV4OWUlIWJVWkCz5lWfCoyXqhZUGfhOe+fbSU4WEdkL6iTjb
uvEUOfPcsLE3fSYhsCYbUvDozUV1cpTsWD/bmkR0VQWjF3GuvxHEZRVvY+PwmJ8L
RTvZ2j6w8om2uUFpbq1cUx7HGehZ5M7hg+vXtASHxL9ngmH10QZVCl9aFUKe7b25
grdXXw2t4TkUootpPyjvczeSnkZHH1dX3WMlAQLbMM3h4c+gBK1i1gRl1QYv1smd
D5LNVmXe65XD/N6Yhe48M3obAFiX7eFPY1x2zf37K28UpOjxbKsDNWvtVmV1AL6L
hvtmwEJY2MicO13DIR5x7KX2caCfRP/nxd71Tc24e7grEksZa8gd2HZ8YaCE+Oif
cdXCgIyVmiNO5X6S/c1LAYMvqaJ5fW3nf7UhLdRsuf0WB4c52on+46UFzmzzHo+c
CochUeLAjPez7RBo4oL8kzRens9aYNGq5NdjvsMAGqRNil/bLmJbnJGotL2MfllP
7vD4BMO5ZVFOj14lqpKD7DYa8nocsMOvyqP+/CGrrKakoL4cd1QO/1tY7Z4KTesw
WCcvsD/40lNieWeQv4MKl85Wz2hSOHbGWlYkjNkOBaf5NyC8EScaVrTHDKBd6m2A
LK22l7G/OG+5VQmNd+ydoRyhmGhiXW6srl25nALv4QSO3Fk8HbyW5Ek2PnuUcmFe
wA1Gw9zUjihWvejeZf/qZ619fYh/Q/gaHPTvCWVKOTa1O2jg/6+ZCF6p+YiFUo4c
HSxWQwBDnEvFz3gkuEY7Gf6VqoeVghA13r9/6g3zZW4XDghSX+hKj+Wze90utZ5o
EmR45ZM991Hbdn/fOYPyMcxxvNz2zjyajDqRZxSYN/8Ztje8CGuBbmSodvg27Xw+
5fK/bCOOluRl65EiiQEqKPdRx+85dkdGzsXeGQXSDpHqDt+H7u4p4ERIEQmPUOFJ
vYAd5B5kr5srs+2XLBPORFQ+cS5bsNT1J+U+WfvsAZb+nYHltWy+CB2nYlB9Xz+r
/MAaN86gq42Q95ruqlTOUUFB7FU5mjBA8Q/RGKecOZqDzd7wHAFruF+uR9SFpoNq
Cn2xWubbNx5jDh66sq3h7E1in+BpvlGaKim1zMpaT8gErfH3rQTBATiZtYKeETR4
HjxJU7thn6PiB1ZwTOyrr328bizC54baLEX1WgWinFGcw2IWVVjAJBvGzXw+FTd0
noQPu4MzVB7WT2Il5JrMW8/CFX487mt0dJtzLsHdCLTZQ3FeD0hM7sXZYrIBeQpM
Z5/8BSOASvXwOyV+MiMfZIwbmAXBQmSLTIr1A/YkykmdN+OtSVDekQjpIXEuVz+x
oKixfBQdyinKHSA9fiLsk7UEeL0Gf28pXbXv1OXJ0lO6xwrWT/E4L1nqnxF7Poik
9w621VdIZRI/jbDQ30BQ+VLE3ZBLkvXNvDB/R1XSUt9nWBeD3R54QiIb7lrIvwpG
447HUU2KwRS2Zlc1374c0Bc1yfIxhDFjVwTpISYmTqdWavtSjYCvGvBf/ax+tbjm
7Am0Ys7jjqIvgUnMIm3bdQnCdo4Rng7fHfjqNlwBeTmSnoIV4ZTWKgc4TMrvXqmv
ol11mDGbSOFCKz39fcngYeJL+0I19Cu4MKOs/nMQmd0ov/f6tQFuMHfGI6Fp02hB
TNuGkG83gYw9sLVEx7kfBuQt9rjJG9OZQGXRo63mD2ebJ0imWRHA3asLimvjA3DS
sehJT/TTfoNIIVns4cDD3V3DExbHnN6w/XI5IApi0ZkObHb73xv2VC6wx0Bigr0v
X8FJw8jomYvg5tSlDw8rX7rQd6GHTxCEQoG/GyFvFmIlFHSF8DFvJa7K8gTkoUKj
wwbBpl7Yqr/QcWAKImz4O2ORGGNUIJxl7rcoSFY2WZpFiUYDY/+ovq2tWTtmkxA+
xFC/EJvjdUg/Lo47TwdXTbdMs4LPMjC+p+6+ImEomiZv47iiNPBYCwPVPOqheTDD
FUtJkWlkTZR29GVYeMv07p5aV72yqmZKpS3ftYhwZPXIWaAlAqwi6MyepSy76ED5
gPyG6gPHn03zTVhNaX6+IB4DGqAASPbeOfNyUarlxeBpukV1z8PGDZj9fhE2LpgN
P86wIw9qG56ne0RUlxO3S7JRkf30HOkQ9BFVSVY87YfMRXwYnVfcwoVNOtjUITvV
qnJp8IrpkmJzSgxjVs6+WKa6Jj4JSKJSlanK9IPa92StMUlCOcPo1fMvnPd/j4/h
L+yFdnHeYwUpg+z37B+jLUiv/Le6hu/YXxYsAH9rkgwgRXwTfO57qKVRaITkxN4M
/2AgNR0MZlybzwMbfIPVEuR1+UlHkS2Mszk0sU6HZUUicf8S78n9fCsmd9QZreWk
61xxNw+UYXRe05e0+/VBxmD14dv4VrFO3vc8SIrA8cQ0dpyvIsXEWD9x0Zg0TnQS
+Qd2aC7bkq5UsJoxmHXjVV99jd0d6h0Y3x4JL7c5Pv+2LZAclr/d72yedGVFAidv
gm3d7wBeipgctjU1J6Iivb4dOiiZCgYkvN4keSpPF762FMXmrKY1If6ecaBL0YbL
p36Lm0GK62RsWroeuVr0/71N5ghCvoUromDKQXezOjqtgdPpInKsuVqF9B3pMnlT
VjT3KRqrUqkLi9WlVc9+JWv1lnIo0gLsi5OckpFSiC4ILbCSZkbXbD0bjElfXeT+
yX7s72m3PxmLO5sJ3zV9fM5ZkEe/Gfljaa3cuO827BI21Hl1RzCcPEMr7Hxrslv6
6EkzJ75AP12qMqJEhIHjcKizErCZsfa2dleQmtRIMtUAWFcweYT/WlLdOdNXhb8A
DQC7h0CSPfhNfYtSYz3qXanMVoT42MXisztwko2GooeRqOkIUk3kRZ95RqUkPn1r
nsOX6Rd28dQWiH4qK1YrZhperFrihedsxwPqBfjGsFg3uT9IOBikZwAevh7QN+XZ
piyVNfYdtc3QL2up9hG5iRLElvFJRLtWrgs3nLvvtgIZjcgwsfBDXp7u8OKlE1Gy
lfm5pVhWrF1oUhMpbCCjfFXEPzH3WNFCCPrITYOFP87cUcy1ZT89yjLt2W4MihVC
lpqWXCfwWGW7Z8ZES5Yucq3DrPXxjwBuGiKR0V92mkxw0l1Iv2bKI58FXxvW69zl
GF1JehJocvBdOLhV/Kh0Ab6k3KB2hlGDcZoVmySlA6uzUSZFcHajHMHsVDF+KaWN
HNSlvaIeM2P2+iSrVEg2rJ09SCCIhaXM0g47R7vNBlrw79dnoIBhx7YLs3PZqR3M
f4YhZ52MdzHNomQ7zwNAfBx47nHQdU3gdPdNVT1wpZMbMVsFejZc+wn/ZmiolnXj
jMZPP9jpl2hzA8oIs+EdpIxE8Y9qyeVkGk7wr4nSIYVxFONT1wVp6MAuEB7QR3ao
Hkz5IRxLJuhGqxVhJC0BnYj0ine5Yj9R3pmZ3uty42+9WxIzJxcjrnKadCMd4mRa
lzKa+C0uh7oF8PrmfIBKNm7PLfRzAPXAwtS6Ze1U9suaiyQ6cJivy4cyXdDp3EcH
pLK7JC1pb0lllkw6zKHQwFwq4tTcTsnFZJ4Rtr3ildbRxHAzbRTyaxfDsK99Rmtv
Oy3soUhXoYFy6msw/HBVqYpTciYeGN1Jm7mkedLYfijyYoi40O5EI8qZ30N2Ptuc
qXp5w8Tk5BDuMNHZbMImKzXerOxgLnihIhRp7OJe+46iemk6qdzfx8zL6ravh2GZ
g9PMtYJY6srebqKVS6tOFSlrMG6VRGATQvcfigKeO4/N+9zuvVJcJ8KR4Jyss89y
ey414Hlk111fy6G3t8zw5QRiHgospLOmKNvJbuUtfJ6FTqJc9BhWzG3SJHFZo6uI
KAl2ytm2bkCkvrAuDkUkBuu+StyF7FfVn3rXyMuOtI3YtjUmXKkJl/azEnM8eBMM
nekEaY3H/hnRi4CjQHSVXAo/OPIz950uUKeEk4Nw8rqGIsKJsGfrG7pyi+4YuK+m
gDIfYtXM1euoiSldN31n8I81knElzaVE/R8TMveqHljeF/uj/q/UQECvwcI5isAE
ESUY3OFhte8KbQlhpAvTmKPIAoG2AGcIs/U95dOOFSgjBPh64qGR5P42x/AHxg8J
ncHBuUE3aK/6PkgkZgq44OQS6Jd+bsZCklgVr+ep2sixWUoxzbZ91g1sUX7q7634
GHBPaC8JtbvUUis90N/qW4Ix2/wPsHXRo/2ddVBSWwxsIVwaCumaFs+CDsA5kaPn
r6uN8w+w3IPtDQeM/HPr6Os+KwsZ3ehzaIMTN/ANfEEai3zCBscWARZHxhPhki9x
a8xt8hbyAwzgQGIq0wrM8GFEWbrxH0lhmr8v/5BKBUpSWc14+1MS9kZAQ8NX02gu
Nbe9n4sw/CNK/DbVcxPnTyV3umrwrVm2MaO0l4alwcduLFih/Fl6qM1wwv1OmQDB
0jwgGMszkX19jmnsuihuwgjd5J/mQkne7F1lg0e1sk7eoiQLbASbWX0fyKcYNktT
5sgwMrDSI0qAmH8w35OtQARWIgYcJxjxE69ywtR7NeQyg/DffF5g+ot4zHbgFq1v
kolQym5JbHGPcxyU8Mmo9LXceq8bIrBOif6xvGb+iN1IcZU5hcfRmjBSrfXu2F7v
fpA9iOHwE3kWWIkf0ofdWdbfE1Zebo3S+l2ihO9bAcTWurCBUw9mx8mKgTX9Gpvk
EyYSdLd03sBqpHcVBO4zlrapBHH6ZpuiDQ8WV+cooN1QMvoxduVmtMdDUfhO5sVV
prWVwiwgjBLqeuiw9jgJnJIOFZz6ckiPp3OfY8CVTJoJHYSe3l6biQyihhdmucGG
RtljAOWbYH1FlyvDmuM6DlITJms276nAmykq6VM7qm74A4Y4FNtPve3eTUM844OH
Hd3aS+HdgfZimki/qiqM3by0gqRzE5F9eA3xUtg/J9ZvudK7C3CScA2balYw/ElR
0N3rzxSaOJZ5AvET0myP0cLcIsp2V6b3yZge91rujtg4Nkwmj1d6C32xi6K0fIfg
Ki0ZK5Zo9wEfHiR3eH5cd1AJYtCqJh4Gnh2nbu3QtAqxT7c7nhgBOPJ0H/CZf6Re
+wKGaF5QvNCTX8S7L7m0GpuLzqJYDm1U5H6exL/3xP3mxKv7XykaX2TItEp6Sbl8
TWZHAjR+9Df7r4KeedMUgGmmFNQ85WMqd0WhreyL7twdvXLucl4GsNAb7a5FpoYG
85PUw7EqW8atQiIYaZh7gcHfsbxDfBZtMtwSIUD0TqpYHppxZMYYtvZq8Y3sXhvo
Fskny8sVmx9sIClbWrwJtSmBRiJxcxmvUbAkNwVpJFHZTAHbK4iFeKeIloS+m7La
zSBmjUVJF5ZAlQUwvf5nJTr6N8v52TipjQEGDBG6kduxZgMqthW2MpliFN2Ir28t
26ate/UD4xPLHIygfDaD8bzdAUe/whgc4fRME9ylL7PhzwLgUsW2G7LbwUnUFpMF
Ija72nfKjDiDhoch1ltADFwkcN7gwgioq8a6fnwhyzuXAIC6eU1ngJEvEKIMAE6S
q+aMXbDoCF0fsfXg+ko3bWq8Il2irK/mKp1nI/PowWfQ+xQYSo9JxIZJVMCuAU0v
UCPq1X+LXVz+6V9upVkNx3NF4rxca8k7WaTjoArmAzcvLDDPBPrNa0kHlXCjl6Wy
Tb4gGJTD/uEsK6BFlE5rwPkhmF/EsWV0WSyi8ESjrIsOG+ROTz87Ql1g2Xu1xvdJ
YKgV+ilcdkngBjx3/Lz+ZnuDwuQr6WcM61j0vhrO3yriNCPM2X2l3bM4r4DapKzq
SWy6x53isNo3CQR2oDEWuFVotvlmVe4SKt2OMXki0DQ68aXtwUAeGh7OaspstNmF
dEkoIDSmMghFPqsLLrIB3ofDCeKVbxWHh7lWKtb+NSRr6iylzQwzc1oiAZ4KA1At
i2FeKwode8eeAiJKQuxdG4DsvEiHwHtzwFChlX2w7rqh8480dOR/0R81BG/mhJ5q
VFxH/hX15ba7BapPlvTuvAtF7HyfQhJ6yoGbHd5hISOCcbholLkmPm6aDzpJ8bEh
SSZTPi5t2IpOcljw08ok2hzgqODvCrZnfZRLHPU5Wx58SK4Gt9u+eX0OF9NSrSdY
kT9ESL2/ZW0lP01ocrEtSx+do9Z3a+OUvaDZ2bj9DvBboKeJjR9Ut1tJNykBzi3D
ii6iHYKpTW/FB2uMveod/sCfL1ezYRiMljn4onchKf0byI3XigRys9838TRfqOLT
ruAkobFFrv6Qr2Gk3eNHcZK0SpVq+TxejNM+AILU/gkrAcjUzHMgDoNOXHWyQGh9
YeffixW4yyR99y07XMkPYfohR2C83tOkjs9d4xmL/gLLhi5doD8/6EFHWAQHe6I8
EcbaYd0e/0p5X3/Imtn/xeKhPR1yUOsoEbiX7LgmhQzFxS5+rcKRkhPcY0zub9yp
ETF3ObueLy4oi0mGjS9te3ypAuvXWqYpHeqtVNlpMsyyddNMGz+EiWvBgwp959Ik
MnhJnL45CClrwhw1zS16uJT/U5X23we73s79y/zg1mnKidv0A35BTcbOHMzaViuk
L2mDLeeRccenjddyWwzquog/ST2cn8VG1DaR0xApMY2/LCUIZF8Du6cGoBH3bSTI
oYt/5hgEiFStf775pA+9oZlBYKJNY1YtKclllToCs996lE7u0ApVnKZOC9B7+YCg
3aIbuccF26PMgiMOn5XfMB96kfK3R41tpVTseaYfv3bdz5WdVNYEzsNs4/n4XIXA
i7sELHgcDkA/azTWjVm6Kdk6MZBywTOSoPTkrq0HyBydKabMUIyN8hXUfsabGQpo
jUxwCm+TTapIdSb4Isai84xbExtMYyn5YJKBytOL1xx7G84EX63sccthPxaQUixp
7x4aS+7/PQJ4IeKsoDVICw3Wh7aycMhkRuZlDINYIxtEw7xIB18FfuwsQ2Dkbymp
/TYXf2xjNah68FBuZ2KEX8rnEBZqI9HxSbE0796p6Rr87cBa+NW3inkwHuVeZXEl
dLHYmWl7lD9XMwMTPwPtO/boqWQbpV2bDA0+7A84YkojzL6kbcKLnHKkiYK4YBhf
2m/25J/TbDvrK5je1YO5eekHoH1vY9zhwFrWdhpQmSVhr+XzqcYlGXeZwtuYToCQ
dzArHwaV7PACEhxMKa38YSHbeedJnysmRWNKVH7X5ohm7isD1fI0nboTZEFA+7FA
uNpkVNWHsbfx27st8MXZcdRSXnbLxvxMz0umHCFB1UxL7xzzTprYIx8JFZhpCPLL
eqnGV+sVN8EryJ5KTCuBhTWNVaO1fFI6y4Mf/IuYm/Wd6a3KCX/A0AMTj3ubfc77
2nfPQtSBxMxFBH6LFKXj3nMvouJkFmVG6LuznDM2wyzf75O91OacwanqlqvBgzyU
I39xZutOajv37wCTt6+1ggSc+c0pCj/hQYsLDDhGL3HUlrzweBew90h9W8LeuNyL
WYp/j153aM8WbMjoGVgZPwLpEX1WmJ1/rcyqQmn5wb19AJb1g5n22ojbTQo3nqT5
ALDjcEQ3+JBgm9SgMmal8qplwmgYuxkg797LQmlz4uBhAEoeoXBpm8uiO+5oIph3
2nKArrn+WWL4ZWODG2n3yDATw7d2Utf+rPJ8puri0XBpfXXuSiZ+CAQ4w2CPUv0u
G5dJvqeWT6G4E10cYUqfhzaasBMLRkrmVJrnTMJBqN6/+8SYMCJN4+1DsijAo4BA
SMtZKShN8040B9LEvwtc7+8JHMXmlIDfgwfo7M2Wq49ZbiwVPmc9JYn9MAwHNTkN
M2e2YCnn9V9aGxzIUH+2DvbPFBodUMjVuiqBxJgTewYQiH7tt0AL3fE1dIxZiy/G
hOYLB4XK34EqBsnB9/LIqj1oCqdgK5sMmFWBzCrfo0zqSecTyMlFqS0OhOfNFFLm
CXRVQKNog3s9KvgtREqhEVpp5DPqu67aXVqtDWjF9HEKuzodAtlsrAeF5hFS0Spj
KFkMYs6aj+pzaLqsjlkuLsbn71sObMBhqqhdzbbmPu6Z2pYRMvWbpDjdB8lT6/SM
fDejYPUFPTV/ppfiB3u/0vfbpRQ02WRe/qigRoGYXAyLGZRhAE/9P65XowQyAC8S
XBNXEZet/pPFGju2GHwA7kUVjKERIXay08XCdJUsoAY8lMJgvECW9xSc+9UJkScv
KiEJZeE67pVGBsc6+oni0fAxG/URuMIHcBT8HXhCcmpBFX5f3avEwBbNDC09DPX3
uAgOel8QtnBCwfps6yBlOC54FBkXOHzO/VxFL7pZux9f/Bn8aNeLGR+CxWUgvq5L
NVqserS1DMSA0ycPdIxHRa0HmgU1TA4s2UGDjczYaToDBZoZhCzG3fVStde8f4Mz
jq4BKpFjsxL2REFJhsGbvBSNob1Yft6hkl5k2sneopUZxk22UibqwlcPqep6DdPC
ZZJ4ATREkKkDyWeWSZmO7JsQ0ekPQ7d7NX06cXNHo6Aq5Uvur/Pvc1SchwH+TcjE
36oDZKj7K7AJDdzmrDV6dpfuVtlJXt4vdvrSNirdJFjCdayZMiwn+06PDhuYrv4W
U4GZKEUZRRfjai995X02a7zslQLyuY2ThwUmM/Ra/edVV/h856rI2/wjX2a18HKK
qlSd7dWLbE8MauddbWrhxXMWMCkSLBjPoW3DbFiT9gJ8XCW7SnIwAx7keN8tB7uw
2pVKyQ7LMsHoJagwGiPf+RuIZ7gpbIv/6NkQq921KdR2gp4V+2v8WulprKjM4Z9M
47Cnni442Wm6G1CeYbCJywiS4znywrGEn/DGAIaCKB4XsDYQp8souF933IDpbHwd
SHA79r0BNXmL5kw3cP2krH8RzCfr3iD+XMvPYQUox/1vw7WfDBelOpkNFULUDgIB
mRgy/TXYgIZ0mPwFdlfoZi2BeqyDFvQGfg2EpmCvxKeRPLoDqusVaUg5Zu2UDbHf
CrFa6u9gUd2HaXQnPDe2hbBOWADClTr3JlHopa2J5UOQv/VoFqLpCsR6hfXnUNcf
eZM7PypDUH9RMbTbPc4qSVq7GWe0nyonBtDruLhrhsAg2IBfVdgEGr+p7XMPDaDo
+YEP8JG+OUDWXZUZnT08naLRJuY4xZZiYlp+l/mu+JcZQuf/NObM6LVlQcl0Aadj
0vBseKDasOI1y0UJmsSJoUj38wGcp3ww1Q6tm5s+CQq/JP5xnma7UVG/p+XnSWyZ
9jEf/Qk2I8Tdsuq+8+MDSs+MWHzZB+y2xe0c7v261o95AifWfBsRciV17mN/+Zss
JAyqocySyfSufPUfet00ZG/bH9j2yl++c4J75FQoXtbGEQBukUHQ9nJYFGPqW8xn
aps/fB9TmIC3II218MPYSP/yI2bQFiTPAuHq76v+gf85DlSTmdXOLGRA/9ZaBLgm
jdp3s71TKzAMiRlIv2nuk11GWxqN41LeiyU0S2NzCB7eS0w1M8nuL0hduowQe6K9
4NQFIhpqmddkfGB6DMct9GV05JcL4YcdG4p3hISvJoXCjJwgACbZq3C5V6ZH9KLc
RdjYdqvMwO9xLv+ByWXJItnlth2GG8YNh3307ntpfoTBe7w3xvC/BENyyJN3zRgg
c+/DyXmBuHAJKT6V8ao+ta5LrdsSpM8IDaYeRCdMrW63ugt3odcBg12vhuq1oA/0
JwCfMB7VRdTEdgUEz8SFlm5gwGJvyK92FlyBQ7LosP0UBL/zQIBzBe3j3HR9Yb74
VhPGfFZMW10SfTSQzEuL450m2K3FrQretGMMcujDCHNDqrKMoQMi3A+DVWYCjxxX
1zrFRAdoXMaq7yXFmk6kILMgKV9P8ZNG+nmw+4/Db5UbP6AAMElMr7xj0S6hlmox
svXlqcgRutOZu53sc1xXbe6n42QMs4amtKVus26tkTqftjZRssgVnoGOiopFFPs8
WBVmImVZVIOwqqHkEhiNxXdQ3xEkoC6rhwhE/62vhm4MRmT68O6h7Okweyjc56wg
19oxBkD8e2cMAqTQ5/F4skIsbCBhA+DJXSzF682TpTgjMZa11vTQQfJWCxzCvjNh
atmR1xLSX+ps2Vyq/bkV52ZWOQSpE7GE5pZCj2RKidXpzoaGrQiDqd6xG9vBFRjr
1OPEbfmYDAme16MRdM5bmXfxbl5a9rU6+cVTADN4dsPD0F6Hw8fPxuhNcAU20By4
v5nPn2K8bBactqyvd/5y7rmBe/0uWV98YpvAPeDF0AXSgFdlfC7Py7nVa5Iin+bz
Qn9iA4OatUOJtycDsAiUqlgxZKI+iH+OKQsn+cNfvEylZcjV4x36TugSmFziUQr6
Pruj1EiJiVsA2SXEchLAEvWKvlP9U6jA20a5xavUN6kTpecf8FpjXmzVT95thtqG
8KWss3lw0h8lwubGSkwOXkMWHft/7icCq8KYqzQQvgXe9uL7EFTGaEMIFusISgqY
nmrwSWlg3dtciaF3lBJM1vb0PkdXA8ZdZxF1pSI6SxGwPOKmAaCqvbWwWokpGcRZ
g+Ey1GolWOSHxgBjrifiyVqpYEQp3InpXticXa1PQ7gdbMcuQuL6ea5C4JvZy/OK
NDzKPABGGX6PqUlcgDx5l6cyuzeGci2ACiU773oIRVYfrUnhFmhbZRmUK0tqBY+3
0lowH2HUsnMs58ahB7E87IAaZff4K9CYmlu8/HkkdifHfFxEy+7bY3euVAZwsgGI
VypoF3XG6BKP6VAwjXu9G7eRKiX0HS/RGjhhAj82lUtlTuy/C897cdtTkI5WfwcW
a5v7SJQISQ7kZsAqO4ZHv/D6zBjojNRooY4QAKraLj0yvj5NBlic6Yw4IZv6gm2I
k2Cm+Tzxd0x+jizu6qvF5sbx3U1iVWG8nBWrHy00dGJ6UoANRiOAo0DABejvAqrq
gnQrXfB6LzKgZZIyn9bS7dY6vFC3D4wyPDlgK5wjLVZTUaFaVOyhy1cMdexfqHqa
K94k/YagpevLQeA5w178Wb5cNAkhdcQxMOpnGH0k2rteMlotFAePubYnIYF1uzGL
2S/MuMJvEn7ATjEiwzggUT2jtYn3fEcAnfcPhgGSmZK24DQMh5PT16eM46HukkxH
Zi7iz/eUZ5RNg7mmgm1VN9/4FBYDuBF84oRVoS/p/kjMrA936DJ/PrWLQZZMuyCN
3yJBubj4PVCCK3+tKgV33iomwVWm/1HB+KujSSOr8MZfXlxn9qkay9ZYQObZJ88p
gF3y/YGwFwNIuAS2Bz8E0HhRQfMDmyzh8khNsDdpAYjtlRBVKHLqn/SETpOBYGXI
EXhkku+fP4uWIxLWSD8BoFwE7pyzmrCmPESEJoW4WNbl2L67bibxX0dUr94ZF9eq
b3FOaYe1Ijs5aX0Pgl4I2zeEEMUDMkvUpu/q5alkr6wBMzeDitzjIjK0r6nnfhup
JsWZS9iwKPNy2Nro7a189BvqZTFVdpQZsZUeHb0l9vYuu75dkB0xh+gl8QMe4xgn
gsG9rAuwT6Yene5iPgw6dFVZlDYi99KxO05Toz7YaLqW2hjViZWjpk0z8Wmej7Qu
DO6+wwluDhWjHkBOf5A2THuUG0PzdpFTLLdguKSrNSZqOLK2orqn/AojQmJ0PEIF
KrpdxAHHMB1mXzrVAo02KEr4FaI9rp/z43GkHdIcGXxrZClOOhdCQqfbHR5iBoVX
h9j3g90Vxmh799DDAaXXa/29eAcsPW19Zfh2YyK9apKaS5xY5UhImRUMDmpmw4A1
eSsfgI11I8hNH7fLSUqzwOHJuk0pnNXPvPsaAZu4AjOroqCxId9Rc7yUpw6xVBg8
8xHFxYSNrm3V+jq/wemXsuupzoh2ohOypnOgR0ZkiIrUcyhZFLlkQmSs6kbfDrgA
ilTBpxQCWTlLx2VLg6gJNDIKgvS1GbF5fs0tOZFv0P4kvAtYCIvyH0jYbZWe1Kkm
LKb72SFo1MKU1getYjQsydmJ7LsQ5V+5AYsIV4Hac473258CnGKPurXT2DQOEIbg
iZ8i0jTz97XOxZPDUfzrnwbFjejTLjbbfAGzYnB3/sPqIjUqlYR3iFobWhuva88Z
vzVj+0ib4iPJW+G2VQJ3xpghI914Lzx+JzObOukAQqZav98ZgqXrXgJM42wvI4aG
MN88jgZH0npMHvi6oNQplM6xM8SQRY3r+NxqqjXA6TaGQgRwh35q3jvO0KQnj5RB
fXEkGKNWuAphcj7Y83IFuKvFa2l1lilFS+Lh/0FwxytS754z+9J5bWnm1MeDbXeA
YYpm1zkPNCkWRBS+P4IiTOAdhiHIEvRvotz39hydihvAGNhEdGBoIvpSI3/9G2a8
YTktA3TEbcZGcYI+ye9vPvF9EitZQHdR1Pq7KZruFAOv27Dln4mqA04SHYJlfG/d
XNq31S4QEnyhgJvGDiIrEifCsVcZ4EWEcNKcaijJlCsORRrv5bdTxzH0oGHo2Y/I
MN2fAx1k07gAokKklXUABjLrZqaPx7hzgZh+/gZo85a//zT1P8tGUg33rDnYkQ3c
vRYVNHJGBUbKq4OqWv75OWZKdFuVzIxWSsISzuQpS1Hb1z8aOSGvZZ0gkPHAklv/
/IlYUDLiZZwVPZg2tyfKtDxzFq21lExHsny7aMU+rr2ZuDuK8ycdfgy2lLKznxZ5
rl+NV0aFqFNOL/jqwEBKlZWPv2pEOjeLmDBZMgTdmZGMzEW8BE7e65lAaVk5wcJM
aViBVc6kP+AB4IonHI0Fd4CR4SS4XlY6xlKe7bOTD0HtiEwy7ZLP28bqIH0pwDCa
kYK8sZsiV2BhzYX1ZkfIrGj6sivfDSWAPNLZLZZGV7htZKSaIA7EtO7J5Pq1pilC
wVznhU9JF0gADgwCfvUUZELiUOR/aH03DKl4xB6+4U2/F6Q2GDKW39SeRJHGwuEs
3/45k31lnXhksELq3ib/qoT16Uqa21J+RctRKonHksy+O2tRyftt/Sp7mwWlxp8W
OXx+hsASf5JiM9l4TBhD7g3vd4nmVKNkogEVzgTFIf1swhGbZ7CXBsmyvruL4CQ4
onocJoUrlnpH6er3zuyutdeuV4AeFznXJkplypFpZT6inH/3on7fEu3FeFS/2gFV
d6hv9MMGexKUMLh+ZhSJsqLAyBLXKEBKocc8n1FsrK8NTYtQ2UHmktdGJyCB29xV
u/LKlCaWP74Sr7pknVpcXhU62V9GyMrx4wKuf+bIKzOrfVx/V7EdoTZVWVSStlM+
TpxZK2yutPUMdZbp7MFJhhbMxozAjGeD4oCm0pIQoGgvBnQDT0OIv4UiYXmGXQHR
jfEgOsxwDpLerRXHI5VQoo99/vLMIE7z5iBVUwy1xGzTQJDH909T8Kx3FhekJvo5
zESs+Z+XsCVmCcaE92EUZgd5I7qCyx59pBuLSg6wBLj3a6h4Qc4uWtvi/YITow0F
ziZ+QZyPAZV5vvBW4QOb+SXHwodEilyFV6qDf496QRm8bwhgLrBx6XwzIIkJf7CJ
VCG3/QmHJDg7PMeCsL3OKyDE4yU2khE9247W4p6BwFBxrXBA+f6ZypbCSvJPH7Fp
nKtKj69Vanu7EpytmyKZIxSB6L+uM2USet7l8AMqHj+X3gDzwfsCMYLz1u69Cvls
qratD/q5+FaDqBCweN87T0xm6aaFXhGMJAFjGRh47maTHmRvsg59Cq1DysSV856I
lmrWc/qoqsGkk94S7tvr04VEe/RXTm0Al3cqCcmpcR4cwLShWktGlNkhwHRMPoda
+zux7yUj7OqjduOtWmiVnzl8UR6itDKG3wtQ4K94r0ZoEnonltSM7VgCadybLlmU
PNliCthKXwLKntYXVOqC3dhlYfidBMVy1Q1224LLqzAtiozU08+i8rSkKAtXnBUB
m9RBl6Ws8j1KWgdqfEZvakI9PQZAsdTvqQ69/feh3QGBP+SPTgejXcd/PbJOMbII
srEzDg+gMgXOmMf3sFp3iB8yyHyLB1iCRbCCm5NqutB0wYbD8cpp5P+w3SKfDI9G
rZ/013mzC7dVCsDSPpBdw+ztVxQyT5IQdwRWOdv3qlgTTfJ9F+mcSAHoAdgihWXP
QgR3utmt91MCjfTPWFu83yhmAwyofL4iSvsGnr55/EvhoOMli5UzcqT5NMQndtOW
svaN3leZ4ePs2XZgk6/NcPXvt0ihry7qPME9mmLqXJSlclzAE2ss6ECP8DAZ8+nZ
jw26/SDKJLM37TqbsWdkd5SRZPw/AuI01dTPlTtULnypqrL7fadbbO04mkTW88C1
tEolnlFzZDs50t0509LCN+cqOpcMjELwk4/psKsPOOo4LlhkoHAhfAbbeJk9gnsZ
xYn2bFeNzgBsG5/4kIYoxeifCBFRE3SppzLRVUmS+nRuZmFZ6tzwJdgvmdnhi6Fg
xuveMoVTh56AKgxOWSTSFI6BfuxEsREk9mWfhzuEGW9KQw/0SPQPOmbSbkfMcmGr
YaL16HJyNkuxkrOAo/nN2/RdQDMtzr9lhVQLRbfEEECb7D3PObDhjRbZd/b0fTYV
8IqjTelmVm0IJiPoi9ZZsMexK93W9KQKlZLvdPHPUoHROGhwpWvbBSzPbV6IX2rx
TewxZkuBU1yi+Ssk/ObxLaiyK/cFIVcQ92ZLU2YDtk8lV9CHL2q4wNPgDajYosZZ
YkdvnTGjeOVHkn+EdJeW4Cph2vu7REQSV39rWSt3Tzklk/JwRgg1VNHWCQQx5PyC
m5vimmoCm5Ah1byWqYnKEvsu+TpIVEa5Cmk7LZi0FmmKQR60s1cWoCGdMCKsBZKj
Ao5/+HPxcB8brXviIRJnTpo2+xiULpozmfFBslUJA7Aio3HkD5z6d3vMWXPPUWR5
S4I5V9rGdzQdLFGVRiJsh1tiAEQp5o/FDJIiRuDOY37JiiYYszb1NYRF4TzOnoD0
k/IRG3sZtDX8JZScpcnQ+qBztu2czfQDzw+Q3SfwEtL4VDoGDM8jux9pEQoFnJVi
fZAEojlIGsZzquoBeeexSmy7P5UriCbiwtGhCHHKssEBrHYWh0KRWIeM4X7UmYpJ
OMftOpDRuobfJo+s7NNYHfadOoZi+QZp7q4j94KJYlvGKxAgLvNEDogK8gQZQDmS
lhVsRim99VGpkrmys1rKwRnbYIo+cJCzFadrsCi5sDwkATGORLj3dVKiNJiRKjYM
b0XNq7AeOgw9FMwwBz0+9d4NR+LUn32SRAMCJ9oEx2zs4PW1UtNebVucipOwEzwp
WqqRf2oxCkWvgLr1/dbT9nUsZ2TQ6hQdLQ61F/m33gwS9K00y+cV5ku4UKBHiAxI
Or9KH5jzDHeELzl07o8V/ZoE+Y4MpciBwDM3UiHOa9FQB3s1Ae7AIGfcX4DBBNoj
R/kQIAkiF969LHdCMgPfiYw5uWLuZ7Juf5CI8yMCtEPaXThD9bEQXXaOIaCDlCHK
9KlvRxtRwZr5Mpli/2zt8TqbZtyWxFCzXE/vq8HBkrwJMGSndAaxG6HJhociIkYu
syW3oLQwvLvbzEC0EvxXPwye0TRqjpwLvjypzjVJxkXzVep2Ola/jqgC+x1d5KI/
hx5B2WjjFKWsUjIHqxa5BGpRFPrN8qj0QaLiXq1KwZATzZloJ/Uam34EEhkQBQ6S
p1YbAnx7NgQV7Rao3cQhxMzPzTGUS/GyI+wIfrAscffr/OrYnecrd1lCBUwuQoUy
OH+uegc3NtXFLI4KBukTFKa+1M1/NxGq3HtSVJja6Blc7Znq3NBM/FIdcuvsJosa
7fZyVHtqnfJbNJBv0rPIKXglTTJyEAWF3nnjDqfhwXbZ5e904SrocpcrlQibovmt
HGJcLYl5amLFmDKHeV2KdVVEhapb0gUNggcO4TqfbAlJQXUMxxjnguJCzSgQTTg/
mp6YXlhVGaQvRSYt5fjTTPwkzChtKm6eMdSVWQgGDpycPIl4RTZM06GFM1B5u5Zz
UTEQeLyHspzEqZAed8VD8VT5Mycdkj3YeF4kutrg5AxlIEGqs5SNchsXwVVkCmqx
GkbUAzpTp4lKwVK6jGc36pR8ydu8BbTLitZWd8j2AIV9OdM8ELxeoH0PcGprbFeN
/0S1a3kDK8kqQSJcj3X/5Q3arDl7xyib0ciTRplg1F4u7XAGRL1PZN2irsRqHrp9
38Lwi9sQqBtmf+4Iet91EUdYKGj6hK4EHq1eMG2jSl3zFUZWZq+z4rrxRtmdn02x
dUan0Oi+f9ZD13BjUh2+OHsxf/yjSh06qNMsoC31KnHyYvBrFq4kwLHfUJNNpjiD
YYUZKVFEXOyCR27cX1Jp22X4J/ZaXuLt344bIR3IpNJldK0Oz8x1IWdwPIefPypx
uZc6XfiZVhyjN1POuLl4ohthqEJD8bBQFq7osweXTDg+uNYr42wzdYEoQYIEz5G2
yo35mFtwsS9ewvnRvZdj7Kog9O6I4mprefP9HfsWVsfppsYmhxlLCzffAsLXCeYa
fSB0GBm6cmXt5h4e6RocGn/EXWBiA5QpIZLLrHReVP9qKi590vnOYyF1HK48btrX
1dW8GFC3iXykVYeQOukRwxQUO3s+qFk4EnoqD1GW/Qbmi5tsholz54LBU3iNet1w
q2Z8d2aLxm5vb8FR3uqt45x2ZP1YVW//n4/X5B0IuXUJDReSg95IsHTdq+yHY+ZN
s+ZHLADMxZ1L2ZFTfpmBn6mqAbro8dgQ+U1weifnf4+u+FbNrKM5MRpLAg/YoA2N
kwYpp0lNkaL2lfZltr+V99mlK2Tcoo3FM9Eb7CGqfllsp+Zyi6oET87auHTuQ54R
y+WYN/mk69CMBUhLVn2NFew0Bplq3PXchisBAOYu4cm6+28mzguzHa665FzNgqP6
2dF/7YaO7bdB9YLfaDvC9g7UKoiUUb9wgap+LLdcVIhAol1Clra47PBfBB0ZzLHc
42smlCmWhpLODJTnDlvVcarb0aJZqe077ouZas62csxqsXDJlxBZMHT3HeQ4754q
7c359SMrLUxqNovSJOk9sCriKccDvXxQU/R2c5pZAWvdeQQkypePpFD+jIAFC1Vf
XKcUjEyrzZhvVuD62aGlBLP4tNcks34KX4uNuft3+axxc5QtDI8aD1uXtExlkHel
ZMet1vtv4Qne5rlIddfZg3X5A9PrH7saLzMF/I/TEZ4rdjas7CN6+d4Cy/y5FUrq
+nNowZLG7x7TEZLk+zFdWol3zYWjd3rpj87U5vag39hFGVTZMQkqMTt/oLAqJp4D
CYYiF9ZA1jO3sg6HbE7U5xI3ACcA2r11p6cqRMdw0eUdIPeAcpkPVRk4qHw1pYp6
v+q/THWkcxD/SiapgPk22Wpyh3rmrZFiTUxaWoBsq3RwUtjOfw97Bg/E+86Z3Qa/
2hVauZIXA7taF9qzc5OOUpneIBVPTfojJT5z/6NFsNdIdrG9QtNin5lzMJT1JRAX
aMGUabxOOgFEeLyx3RSRwn1ZQ+dVjWCUmmgzUpdX8lz9zST66omraDTYibDT/FY0
iBH8sW9IsrCwyaQqiuSamAyLtR7k79unduV/j+VT+iaO+XrG+/cl5FzlSE05Gkhy
s3lCPUVlhv67qJShVjrm8Wscwb47Q0ZO/uiEau579rZr+1gObDwppN0A10orfeki
VSPSiH/59F3oJLxxlGptsPQsjdvrM3Bq4HvZ38dU4nnifrPR+67ZR2kEG8pFqQ1r
o8+pHnIxZS3BaCFfWhxzRl8RnmzlOwvXRHywZcJ/RSbVJ+iTvCvVXnV5w72E8t9E
ZHguPa9qeV6CR3cLDCIvn8fkgvHZ84FXDSMZZ3IHmzCqdfok6dGklVebJlbwi7hO
6AThNcSfTX3es12mW9Wo2/RxuHnsMr2/L+G8F8pndG/bYLcuaERRq3xxd+QoEU03
4Sl+7iHdmVyxo2TqPuDcnnF9nmtvkdqq9wal08d3PPeqhJZ5nOytlz3pO+B3hald
8XQK0JejnUo2S38qqRtfTVIuzQtugxYKIR+LSrDrPG6VBed7kaN4Kc3Ql65ByhAp
ah3d+uZBxqZumBFyh3ExddNso1CUmZiVeCCOOCNl8lTZB/KByTu0nm1U7aJ2oBf+
lXoanXb50/67hpcKq7V6HAN0pUSRnT840RhLySIaqdHn5izZagrGaJEtqBWl+qJ9
JXGSN0Zfxb4wtk9/LVzhenEnRA0qq3fRKNqLEHa1qBg2w4cY/Mo0JYRyyFqsbmQ9
xYJw6/7jrIdqpZIQVa8lN46yLE0jq7tghMYu0wjSWlmNqv7WP8ZFzjNZ0yIDsuT7
pdaF7mESIlmhXTzFQQWPalQPpTnvtLZpLLg8MRbNzrtRoyhAgOqHMMOHPHZTAVeb
NFpZ0S+OFi6OsC1SiSGltSGBn3nhTwEchMf7hPYrMUJN72pT9lxxDpQauIqinKum
hRyM7prhQ8SYypZLGNehInAQfMTSCjJI7XPbHwqBTUwSUpAmf8pm2h2WcI0MECes
jgkTWIDMgJ5tSy+hVgx5bJdybVNLhXcHcN7PK14JMg83uvgOu29wp/UUlFJ/u0XD
k7v3LM1S95gOfAPIzwVVdNNH/sesHURwlQOYqIO+tsLD+kIk8OSfSvWi/ztmilLS
3zhATBc6O2HAei/tmDRlbsQ+QJEh/zru5Z18tr/xg6Dn2x+Jy5t43I0BbDnH5pew
ypfKEuawiAdY8MODbcN+hlJtl2IwFVJ7FJPgP0MxoQeU4DJJREAjdNl3dXP8AIVt
R9TcubnFotcMeTA9WC4n7s4v3Ma5QZXYiTjnoL8cucqn3U8riRNXjXAcRBvg0xa9
zNou/87giwcrTSaEaS7l+kpi+GXu/G4HuqZML9lWT5+oz9bYKdq4N0dBbTyzG2bB
6YpY+pY1m4K8DxVFlrE5UhO0uY8bcL63aUY2LWvvprcODT5CS5/8GCDLLbD0pRsC
cuMlxydJDrZ2PEu+zgx8LqISetfhtOiu1kobdU+VhTfEpMkxssfh0k4TrkmWb3mj
WGvOSpND9Gfgy3ps2v1xVu1v3gxu3Trnw7z8hb3btZuTo/MEqEqwOHGENw93FhaE
raG+GCCBiMLULpyKBJmoYOk/oifkMcciqpGnShXREforQBKOZAy2wp3e7PCoV7f8
wLdEL3KIWfHFpLHOfMwQc6NhfWl0To2gbvOfr4/si7D45sZ5gwZEqz6hHNtyGCar
cCubUap+iRQBlV8heHHbzLt9Pv2WnHriUqBbqC7+hscsGj+ZlVf7CesEVSf7Bait
Aw0+1FimiFFdjqmrzS7d1HsQn0utcfH+myANy9THJTAKeM+PxKMb0PxRBRvZrqyD
HFSyOnjNiYBWtjdcqtbn1aJfXQtjkjrQLW9HGpWcwQMQefUFbxkIB3p8hmlu3tlr
z2bn+aTlG5T1yfE79iUofg7DqsYFFUgOBTXkViHHKM0VAHEH+4tblg5sGT4PIrcU
kX0SsquW/O7Rq4gwRf1rwLNbnfYTFp0vwrmGmvBYrYC9mb4YdqUn3KCj/GKVODpO
vONJ1PrAGjgzNJ/vl2jlhRmhQ1PTJ1etZjXie/QUIwRQqbtL/3Ov+X+DiUfeirF/
4EOzD5kJG2XThxrVNnszrock9MXKEFSwIZBaqcKxy7Nn4IzCDcskSnNDKqRFo5ik
88uRc3xz7ocUshsW3I9HtE46HdalIqeBVc2QS2cyRFvSK2Z0WpNLmXpd6YOwVKXT
5PCcGpyBvC2run+a0EKIwrnaYDWYv/lxgvwwLBpm0o7JKWL/TUt0jbLRyLYAM5rY
Gz1opvDS2Ld/ro2mfTvzKouBsSzZiSrwj5eV0oxuikhuPPxXEVYMzSbZ56L9+HAG
mSq5/CBAtP4WJE2IJOPspbTwB8zGG2+QMviI9MGlgIvGzJek8aZTAFSgWUpNtj0e
Xqqm7lvCGce3xWcz2BOWtvxN1SahZbSaLHCSXkBljgefRm4b5XJ3mV9GWF8SvhzE
45SbNwha5MC9NmZiSpgWgPTJMS/RfYQHmWppkxwmuJWznSUvJbt8Q2I2yx/dM8+v
KIe5ay7VIRcRESrARzoGbTjApvbCa54R90vhkT2iOrcIhJP74T8jBoaKsQnu+wXc
h9g+dcmXEpg5xtApqDSBqH9swpEwDoYd48gL27D69TdrdIfshvIdG9FivwnlFLsQ
jvr24ahomK7J+vOn2A4bIP0zYbd17JJ6aGuzUgBUB8NMlt2j3RHmI3UWrWdM4CVS
FFwN2GvGYgZz1MdqDaMBgdAhEkVv7amqsSsLPuPckmvWEfKgVW5jD0dSnEn6vNzd
jDSnpAsCOFtfcqSzBDphOwrSTEu9322z0tFPTk1MFHaeaFPmxWhMpsMuoYG+HZQc
HcQhy4FCwb6xWVsGmPVepqkAHCFWXh9tFgzziiEaVWZGIdFpdbiF8tdOkuFNNYYM
s7TyZLqeCkQuRCZZZ2IdqGgKrnVYFO7H+zMPBpcr/BgDNP/1Atd4gQIw9l+s/j3M
aWkMSguJL7Kg83AnhDiq+sipTOi4uGpRK3WLwIq3kOjnlFXp9WE35qHXrdleiwsD
KfKFYvXy5At4CTjI/Gj3/y3jhLYKme6WdzqO0d43KfGC2PDNf4njmS01zIQIfxwR
bUh+cUP0bFmxaEK7aEzt/djcyPsk2N54cBQ5xxcp1/0YRAT3/1s86S/xdODKIYxT
rM+WtRjRnWai5jTbo2kXfeeClr5FCgGAutATYvQqevwXxQEiiApFhWXI9jLwj07z
AX29tG2WpNc8uz4Eg9tJw3zf0iR4cZwgFZ1Us2gqClUxbt4YZmsHUAPnXlnCNqmn
qCF6uAsptg9whc+9VntKb9ixp5rMqRdYkG+pq2PHqb5nCbMQGZP6MyIsP1UsC1ub
7/Kx94l1NH4nVuToScQtQDau9rx9NCNSEmfnXdJ5M4Gv45BHYd+g8CFpsx3h77g6
w5XI+3dV1zK+TQ4uDapv9YwhtSTgVK5CSPNnxoXN5vPb1LBJ6NZ4anwEzzlEj96L
jWThJ7e8c/pH+iJw5WhJmj+JEJ0KzoREtglI0n9WR0jv6KGo6GibcKsDQ3hoUpBS
vK4MROOVm991j7dxsbK8VYVAYC7/1gE0URTCE0bZ25uOR+aLXEjua5JEQHEh2Sor
GY/41kGTTDGm+9+MZ6/u6SIUZWp7SA7szbsbolkNhbWM0YggSsgZYmP0NpUyBZlM
vgw9Y0gMaCP176I/c2mQHFXwGppd0Tr9Ivf0dPzfMH7KtZMomjnR3oL5TWtAee6X
p6Q0Bn/1n+o+Wngc3AY0xmpi+wh9Ejrz8VPo129b0I/cu52FY6qVvBVAFZOWY+ZB
lqge1nVeD/fdqdUFzlfYz09DKFDbtBOLQQV064AjSRM7LGBC7nnXkMA0f9nIBkF+
1qPHUr2SWBWLS1HvHVOw31T4+MiKyx8jCRPwhiQBk+hb7LweRy0oBTFmajRlXvx7
d8QeYZXX3Z2C0RhIjPyx5+jy6JKskfPaNlYE+v141HGcC7C1IdC1qw01FIDvNboy
xTqxjzxEKp3skvikQeJfx/QMYyFb9PNMyuKdbdrnqG8sTTzmeSOHnT0ehsnmoBTV
tGTJYURGt9m/C2Fpk5XUT8UZLF72JAOcOYSfXDTrcB3zIlhYCmsELq4zBu/nrwm2
270AXIjRVkZKINPxd+stIrHBhXVOQYtr7wXPtwn4LzzOBuDFsRzrqR6s2UTa5CF7
PvXjk9i1upQ6J3hpPbECak2QFAAcGZlal5xToskV/oMzhynD/FSiNWSh47GGkRAp
oqsBgBsW+nnMMTVAJyObkK2sGeH6ndHiS5gS62I272z5Hr+NKCnO44x4u5ZjdfxE
xYtjog7/+qT3th8UP2aV/W4qn0/+FWv70vnePHp3a0t1SOpMIKQmaPlrYJEP6r26
irrZbJvXFuNfRmcDJB41MfRo26ze3DloILUDyjImg9tnnVViQXDFz4FcjkQxLAtP
k1nG3PMSHEqtCWYzo/7rdVQ9SShJGUe+ZfCVRMNv1NjrN7iuAtKjqWXyJMzwW5m4
qrixWFd3Sh0T8ZB9wsptvlVuayL00N2/4ppvf4lYsmk04yYhwvYVcIsR9F1uE34y
1cCiDppmJEjXsz2Y8l6sc5zUoT1Wq9c1PU8rbQAvY3vaRBJGRF7+MuO/DccY0Di0
5x2dQDVUm+I1JGKMrZf8aJrR6IznKCOaaGdJdj7fh8Z2eKftfwUXKbCUcqVjKF3Q
3JWu1i+5Os4JsurbvybEObyCrGWUsx3nyXaWuU4t7DYq1yw082EWyAP7UDqA5iSw
UhWqe7gidZruNnDTI4wqeKDOmOeJ7uulOAvnKWOc0yLpGC0a/TKHuam+ar2BYxVq
u+rGBcYdsAdSSF21DtLv6/NbrLyoKgMDT0UUQMhnOa3DW5Hv8l7Fcqn3wAQ5OdeZ
VTKCA1EKCOdHK9mGqFg3eYH7+9dNsqhTZm98mixxodnPY7HI1sxMRH7e5JjhSV4L
wXSdykp1bkLm8fmmxemyIREm4+2eJeuOFq4teqi3s2QRFXC3in0TceYTHfehEAJ1
oBVsi4/hApXyK/Lw4zAAvYi4N1Kts2UTeKQHCL7erv56XhRykYqL6UqWWX5UFrMV
2BTxxHoH7ehvPJkrViJODw8q0TiaIyliZWYHH49h6vwlehZMPtA+G+erQmfov0Jk
1GgnH9Rw3F95OGKLgPKXXMppd/HMM9Pkk1rpQMxvSdFt3IBOebXlfYnstY0/MkBG
whdsbtGrKqgkCJYlq3Rapme3H9rjlgxjfOfStokGqX2aw5QgEd2naqisJRJ9sMUJ
CLYc3Dwwm6Qtozg1p9X/KXeW8aQhFKu9NF1BxGSCkUOWHmnozH9qm8cIbSVocB73
21gaiXuiETShm26ExOPqqhj+NwuVC2qLwZRCupH4UjlbVzShcLla9F+zBbC2vFPT
5LRi6/zAz1EQeTtlrMU2YMat5pjhCpO/W2T6grnGBq1yW9uZQl9mOd7KbEx9FKs3
bqNVn1SgSTufDMP1I8KN8pDyHwndnCWQVWw+mzFQdN4QshoCTI34n3/326FC6UPK
KtqYqI18RcpBrU+n9A5C+yL8LEvKQnB6DvVo1hrdCDg281KZPEQ3gpIzcE1QbVB5
P3oSQ4w82sW5zLX+5P6JxYNxJKm88BKmt/FsTr+j3SkRVlncZrez2YX+89buZrc+
lXGyOcm3PXJUfwWm7mAMbN9zGmQ7Krp57xRiAi1ip287fp9tNIetcC81EvH+9nqG
PLtY+hOQVpb1o7cGCk04nPIdonhde2oK8YrfdBqHm0tH92wEquWf0aWIQWbgFnUC
rHEQsn/lZBGUNODCfW+0sQRlA1ih0oNL/vs276G4S+EgI5vqkj9EdxcCmSCEGNeA
NLtGikZCm/zBthAMAYgo2QrXPqXhpInlHaS/6rJZZ8dhkh2tZaoFA53kvoGEfhVW
hHgiocYNOucA9a5DF+WEpBVYkOaEW6Hz5wgFtQsOyxUj/RB9NlndJakn86Pb1JJv
3JZ31xwFDDJVm2/DWejLdwe/PY9jhRFN8hQ+SPK95yeDrfkSk2owpaptOs5xDCk6
8G/kI7a9azx2Tlz5vFeCpcJybGISqu6DRA/lb8kKVHVl/s8IkMq4CgpYOYH6iNCw
myFj6irmqfU+Ye5qy5oOsrohWn+AQPblx1617C1siFrsDQyQFl9PvnwJc1OTItJ4
zASR6y+UodHkv48vkRucAy82CiJlWiaVnlxMv2SW5+vUVnlEq4UiMV1xVnzkQ7sl
sNtIKLqZkVjdtQbU5NMSGDXz6HKsvOKJrbDybZKhFBSIqQ0AKpcyC0ybpwGDEO1X
odfHadrn/4CiblE+FuA37o2x2GTTytoNUdFT+5I2UPpeHfMSDygW+rex1isc2A4h
nhSBJ/q0vgU1QmCNkzkOfIzLQUay4GthtTcITKs+bsl2dBLuHkRke8ZurjVwB9/1
xmYNoGSc6RuoVPX6CyRHiIaP6ACABGqIRCHj4pjJ7Yv4LqpuEX1+MdXHHR+6vfIu
sPxdz+LEdctVE2Xs0wJEbqlzXp29RXpgmc1HJN3zWUYtwDdc9ReY1nzA6t5eZmJF
n8s+lLgvh85p402TCGpFMEK5procnQC+WfFjUBl5fv6Dh3Q195XYB9abujfdOHxv
caET6K8XVe+T1KF1uGvcsajpCaEF0aiBGFNefMvF6ucdxCIv0Y3uhEKVHlzBuTlk
5Yg5BBI9hXiB81UtfWg8QI/j6wU3VRQ6DJZvHgkYEXjATuRbRMMW/6XVPfex/wrI
JLSLz3zn9rqGbbHusALq/GhZDtygl99uYnMcnNOE7bF4g1q8rF3mxZruuaqkfWIB
BReZwdePyerxrlLYEzTngpkClIVaQecSoTEYxPORkAPsvriPJ1xZ6eelMsG9kTo3
8jomkEAl58AHMO9UNVNnNT/AglNVzqiNY0fbo1zL1NsZtCAQLI4Sy+f8+z64agqc
3DOpe1RyDjignX5CokGYonNppQivGMhMUiTNnCS6a7CGoaG1qM9wzukA7EcGa1SZ
B3QCuLtGgQ+XBvHOwpySikGGU+x47zq6OSRVn0Jdb4FeaqjO/HB/C3UIp4AxlwEd
F9bueT5PWH1LZhAEcY5O6+VYjTIhLYoI50H99vOFjE7xEXUkhjEk4t9lRK7d64z8
snCkmbBnRbQSrV41yl5TTUmWa5SwQ/OamPEalFo++CgS0rt6wVyuB6CTUUxX0SaI
q/adQG9Wqd28OTSHUpWY3lun+yZEDJLWdqzB+Z8S/bx6d7H1vFw5zh03ji3Qc6a1
IfbN+4Z8aqGYa5t9F29BzPhLDv3vakAy5wIJhokEas5Ju9J/1gHLsG4Q1UxlkmVV
l4kWnGVFSX2dLKQUGdd1fSCHZQmOZb2541Gj2ObuDTOnJ0Yr7fPRcEwYTUkEBtZP
X1aOTmBcMbZZkVqorhMsQmrvG+DXR86dGQncYKx3rq0McVVP7EEQezOLhFpN7sq4
J1To4UP1WKepxl1I4rFg9G34zKX4S2n+MLPVHbBzygRJ8KLSUTPjdeRwfXEzb7r3
nO7X5PGQ/WGoFJvxuKWiiDUqWa2TYvlAy469ArCQDVYGqWybf9sklDfmnMWD73CF
oFlUy8WAe0Ieq5vmIo8il234rBjy9+w0k4n0X8684RYUjilaN7KWh521ieA+Tx9b
DPXg4RI5ndayc2CWBlCQ21rxllstYiNPAEJyCo5GZ8hnrxtcbFJQiFFKz75o+f1Q
YuJmn0ddzqZCHIh1NOSrY1J3CAizAY4+bkC1vjER1moWl7Zj06bmnKKmROcQbHJC
dSrVapAf2BiFUA60pC/hicswF2VeFw80tkD6ZhPcG/ZW30809PCcGIGEtcwsNlSi
PtYeGZVA9T3EYt5YwNNq7vd/4vS5XEut36Q3NB8gEt/S0KdHdtST3elmVPYKQrDV
cK6w78MIrAVO3Z1e1mh/PnphyQxBQP7UHwWjNQWGgf26dS84ewj29trR+NPM+HAt
1n3A2n11IyAHyTcIjN/nMIAFnqvCQuCEG8IkmmnbaHwK5vKkJEY6kTJbnXwU5xSX
gNgHl2mWixv9Bcleuk+pRTosS+JR2ki/Khd6D32/lCViwK4SJWr4UJweCtt5OKnb
Mz98DFz6TG4xV3CKVa38gUjmg9xBqKJhxRM0q59rHLN68VgtfRMjabvT68cRBYjM
SV0SfroLjQeo0VPfSfYTPpNXkltvcNGtHt3EYMnfjhKacvEIPLj+J49xhDWobU6r
oARoxT4lWQYPmy304JKK9b1BfpdAPG9bbwiwQNzgZlprdmJewkHFvmvY0+jD7WNe
YsLLalf1oGHbVokyG7jg+Ky1c8IvxIs1bax1OC0PdBvJpijjEa2xkGyyZSwl0WDW
7wGztDbbhJImj4jZPmo0zkh8bDCK10gd8NbzQ5pyw8XlDJWbSy/7+0bYVwDlafoA
LaCBI1ols/k6Jz8tTzYseL9/ZY/2DchN2pqczkOtLkLCBRdwMO1NEgXBzUyGijRe
6rlbSI1CIyakj7Btrx0fmL9FwcR92GKYzupaf76XjhVoBfZjHWYO91dzj7WfZvpz
PLirJhH7AMMkDUemtQOc9UoZGwuuJ/SEzCFUlKMLvH0SBNBMQmZ+bwVlxrHPqZsU
H9zQvMIbD+Y0RJaxzAITsHRmH071Jbsh+mTFHOdwTPORmLWZW2y26KEF0PcQGjMM
U25Bidt0/OqMwRx4uyyYj9mHl5ou9+aFEg6qehrvNGlvJV/EmCPJDIavNjJ4VLUL
gXSIt4ms1vbK35yIM3gsH5DFKM1qR51+BZj9ZBl0IoIIsGGGAvoFvO2ilw6jhD08
C6GAO9Zf8KoK/YJfRmDP9Rkl4IGJfWLHtc0TzTzMYeGlGIUrJPfbux4jFKtK/rMB
shRQ7S6cNRx2dg6qgsaXhIjkFNf5JQay8pgsBtn9ulEiZw4WKAa4ESenNwpMkWof
4gC41nVcl8/jE2+skRdYcX2jn6m5jLddqaSVGnXAR22sJCszdJjqWcddTiwloo5m
AkHsWV2DUug+kAswVV+PYIzNa0FwF+wecSDU9VRORtWNJTkXpHOTBjIBapo6GypQ
Gw+p9zGLSuH/YrpaZ2KsCdlyr6NVkUpIQHRZHuknstXjCjn42SplkDtYmWvVQ0vf
sT7e7/EU8cEJqulAPvPHF0szVxim19PNyJa57DuQpwsbQ3ckjV7IjOqPiVqKNoIR
WfXv7AlWn4lCKfBnc9XtfFsLAk3mVqxIdwfpWX9VK+PeKiBfYSBVAH7wdo+t+Vrc
q9FkIoSRjSHf0+YXM04QvFX1ZyD1/icYMbUW7QT9pgC7PUyIyE3mGx0gdrrlHQjb
gmaPEmrpB6UD8/2ewvwFt1KfH6/AX0IqeGuNB91vhXHwgjvHMzYL/RilZqFoUVBn
8VGqOaqlA5fL6YX8/32Q6c0Ipjbe3ZBfq0T4C1ml+7h/TJwT7TcDgeJURFi804gx
Q/EUvLnGBRcI56qxmqraoNBZP5vPWxt5rUKzEORvAAZ1na+NCeJCv+2TAHmrBFI9
3f1GcSm+dtWPEAp1D3oDa4a2IdVtSp1Qsc/4O35t9NgEftYYQReOoU6LTF6vaLND
a0o2kjs8QhAkyuLcsG9GjWUBAgR6sAqPM5sklRewQypZ3T2UV5XRtARKe4T5qp9J
PqFzfGMXGQK/b0jdunZbAyq6HSc91yyCpxT36Lx7ZsD2JWMAYhNmtTAM7y3Zt/Yl
DC2L/a3xqu/os6xVFrPnhMiHZA1iV5r/0pQPoCNSLXtVSfUa+OHiITH4s8r/xR6S
whY9D9ld/C+kAKo6eEHeg+7ZJsrHxMyOJlfvuxw1rzK7Spvufu6XDw8LltuEDRdu
4pP6b0zjch/lb8nHnpOghX8nDXAZPRv5P9wuj5Lm9JZY/1axlqup6m1KFCP/PCTj
FYIpQHG04IVAGhU1xgPvONGVCHeO63+vg3nJXp12RuETZDyVdQutZjDP70ZBH4Hk
j6eneXVbrqZmSJDOeGtvxzDixfbEUQuvqQHRWu0vZxRsSr10mfwNM+40pUxVZQjQ
Qoq2blY3U+C6K38k/WByi4jPdU/9w/eb21BgWYThN1lkDtW7WXCzUdIsLt14bcQ4
qW57Yy9YIxPIVVJf7JJphHckkTcm+mrztEo3za5fJ7Gw6GyTP6iOEGhpg2BofMg/
JSY312e8ITWFYHcEIoI8aXHC3jIZVBn31CiDUZgyKgZPnuMSGLaN+gQmXeoGNw+O
/uGtN/Ew3fgeOcZ/6aTA5IwFu0Gn8WesJIUjtP1yB8f9scqiq8WxTR/3ewJ3xveb
/W3Vf+eENCGVzGAHhepZ1xdI3xprQTNQcuBK5hMOQORrP+R1RsT86UFSAquKneIT
d+442k8mrLRXqYXbmffkYXQoSCcjOhOO0m2Y9i5/uWQUhYreHyRMsoHe/QCvMphi
ruaSE6vTw6g+PejaCoZvcQ/PwS94BUwf8MKepKwsp8QXkoi96i0dY6tZJIipWAGU
zywXI2bwraYybNifT9OPFxsE5GCzdIeJPPIj5Dj+xLYreuJ2/9iT3xuEq6NY8UnG
Q+eySLbU0gUCc5WdFJcRsp3LTHLokOh4esEvW99OsFMgG6XQJUUqtBIIZFXfdUNH
GxPdHWpPxwv8H9b0zP03owBRp7OpIUCNZqP3hkxsWl6DF1TW9ezmmJaR4rWTjDqe
LGIIFriHszfFMkMa0+6keV/utOuhRluTEvzYNfgdexWf4jPXTgYbe029qDKl/pb8
ysQf5tjpljML141aJBMLGZGQpasdHxKEHcIJT9MRfyzV004fnZb/mS6nBqMi+Bm3
0jiURl207oH/cFlNLBLZpTq6ry1D63j7dX4cRUZVRW/wBSiY1cShqyXwP9k8Z1aR
B9ZNw3KfSJTotYN2YC7KYOX26E53b6ldTBaiGUaIpqQz9TBidxN+3LORPGGjZaHI
eMLhYbEWnXCq0C0H/npmIvXhJGj6ljQmC3p1v0Coj0tg0cnB813WSdstzFH6JZWq
f/0hJlHCY/z5Nu+9EM7nU4H6BOFQm876qg/JF7qedRsnfisamcRwwHZWeFHC7Bkc
nh1vr3+GqifAyzw0oLi34IyD5S9S8UhtSVHDLzEjboIR4DSVIOpg2kt7rycoEAzd
WP42RoYhutzYlOkLkpk93A51CFTUwdqRASXF4ATcQSJa6a1UnDaKeibpBj7pc/eb
g9KG5sID81XESRM2dpkz9ad8+82do0H3d3fSE9VSg+DAa7ldU7lPzem8aKhCzr89
ss7kqR03CDPXj9iPqfrQ5NBgFcmsisftgGCqvcjFcV8nTN/9VC76GXjH3mgV8LOV
nJgatzy3UY5dn3lUMMqt1HctjtIJmgWXH3v5i7LA+tR0q0qRiEUQmXG3MuDOucT0
MtI56mjGBtdEWMFLozsFVqnVih8ZtpNvt29cpYytAkpmW3GK38ywI0XwieBI+m8N
6+Kmx20G73S7fmrWtAPWb1LdGFZzDwXJxwRFNJ/8AmF5MrfQkmHa7J68JMFQbxHl
mIq1hmmWYTRwJyeNI0+AjCH0nzLxTEBeeteL72lyXZ84opy15VDEYFWvlTaxVmP1
6iYyT5mXQm3GAledqjofZM/QPFNZkdKfDpjSqRJKNfQK57V75limMFiGCOU1T2ad
jg68do/fG03duYT55eChKsBWZZi9PbzNrSJiMfL50FqUrLJMGJl3KkKTekWtqsQb
6vjAwx13M40TyNojtZ8y3z9iHB9c6E0VnJor3jgTxn0DhjSq41xeXQw27kesoe5o
zvV4KdrDjWlM29rPuF2k6LQ48puMMrYrcnZ20/9+Q0hOLQRkmmDShxdEjvvi68rz
/xxjWp1ywN25hsbBQwrWipe/5cgAMC/7QPIjNIbgrt1+uH+zSnHvsTXQ7Q8CRf8Z
AG6Hveh9NoGGv05fhtSwefkiGrcMBsjhxcqdsh0G8ivPR3vtxoBRcYmXRtWc9CZI
hG+hSGg6k+NimhgssBkg1JS3MIhrJLJt4jwZ6JhgHQF4q8XD5utpZtml/75WBdxh
bx5YQ4ViOIIJWgYJappgD0Cx6B2tDvZwgw1jtEdVD0Uy6KTqE5lfeos81h1YQ5+l
C2QqeaZWIn4dcCpPwtuWHj0smtmU2M76RKheWNRjL08hq4xvj+sS7asSnsAXfKwa
8y9cRsJxRSaVOZFuYkcTIVCTAnVg2iiuWhfFlYUSbZRUYO4lvyd2vjl23u+el6q0
KWZY8/CUGW3lHqcd0rC13nUuYKD0YNqttf4uyrcwTGswzVuQjZW5kQHGjAX2l+4V
ZgV4qbc05Uq8rRIobv3i8May0rb4LD/qMvswxkC/aBlEw33bIw2LbIgQqo0G9APr
tX2QOD2A7hJw6/S5aZ34r9d4PndUhv/CBY/eboZPb+SaN2idOJEGYHZQJpXmC4BI
NqGs7D3+G+5PQ4fbj+UnUO9cRTLqhARIfViERtaCBohLhg6eL3vfey23vMpKvYeH
PVodFnVBU7p0f8vu8mtIB5S3gAtyPoH4EIYYWE3n9GuKsNjov7EhGl16Dc85RKm/
zkjumNnulNHm0Jb+MNZSC71WsxAN0mEx5CBgmyz5gVgvMAQgg34wsOuplj+0jfzU
52/X48op4pdvUhjeYkUexvMe8ajFJZYJYWfIuTpPzulnjDQ8n0X/qK71F2R2wPpJ
iuBaPnMbUkctGNfduf5OOA3j9v1WjWZ/aH2o86znDjFF5golUvkoxQ1gpqpgdZEV
LAe2XSlLDBf+npdTaDyEY3JcVMUddJEjw7FuU2YuXCvPM6jQwxCheYZz0Zwf69nr
hxDfLVMQ+5s78oA/PFp6Vy3g2oMohaq0VMPky4L3d+wqFA0fMthqtHSHzu/qqp0L
1n3EELlT9/BwcS+Bd39f9MZbjoiklDHFue02eRILfGXbCqHLbcc//o2WDBCfv0eJ
kkUihUwrFg92G2065Y0E5fiptC4GouTqupf2kxZzML/Yq+6dGJ8PWFyeGppVZGWT
E/hoZ64cNLRBAdA7+cNjPuJFWdlELWVVTCU6oo1t5PbQiwXZwlY19uVQe7uzeCt4
KNdwp7VyndDX+tvEmw8NYxfkcZd6eTOYNl+nm5Ktr0eREKFh8EFsy03zdzl0ejsP
A7aFxF05XEiDVcqg2bCbwNlHgkEapnOsZeq9PkxQnUDk1NxrgvaykBm0XE3/EAhm
sjjkP6C6L/LLUVObIRPLLRsfcqvkFsL6X2KNkXYsoGo2JiioMHjGRLmd9Dz75NWv
4cAIUGDUR+FEpdKs4YLT2EtYwbQzQqsaZv4SO8NkMiuH0cOvyohErjm2lDPT02mV
3s67hCVqY1Zn1LcT0w38bVu95sdtCC+WeagXZv6SjIIrGI38eP/2IADMch+FgOla
ZE0CsKDq84vOXsUXov1z50YB8KDNsS/A+HHXt01BL8pvf/7euegevCjAxWzRnQi3
SS0YjvtlqEddC7LMsilAnB5CLdeEhiFqYxHPo3KoSHn2pm9uGZCS9tQkTwr0nmeE
EjHuXwug2gpxn1ui3Jbp9kPoHvfC/6+8+nuMWrCTR0rd44Z9VCuUDFxgtBOXG5kw
alR9M3++AZx0supCywQCproodsDrC/iGbxAsxMvDY5qIG2PZBK4QSk4O2z7UN9U8
61XcrBMQS3l4K1yt7ibjv5rVAvlj7iagG6prP9FU9oDpiCcRqhk2urxmVFcHFZD3
xKzzbDvP1M0qhKUL/+aaE2PkrDHFyAawgXJ4Aq1IlNnrDyOJ16LQLCeFpAbPAJun
KUEBUAs7zoMNWBMNOSaQ/kprgRWS90V2E3R+5GWQV+iWsDu6F/8JLjr0t17sR8W0
p6g6qP5WcYaHZRmix6Vm68cqkPMkeOGxnrE7qUd8GiR3ObyA8wqDYcWrQ8jRkCE6
wvgLjMg0S4imXhUSdDiRUSF5rivqgp1lXQRpbJZVbNhxqBXllAQAYBjcAlyCFyCm
gWzuMbn/tqJdUEcrG7fRD8vTSpz2q3qsd9vL2OaFY4R/EwtLMoi8xpq4K8dNv21X
lBg8tcMvg4v9BS2m6mhYv+Dg+JNW+u9DZqTByZM/RkTa3eA7ZlMvIJNW1AQvXzZC
iQ2i883qOqPpYMEBJONWtZvG99Spsgg80K5ijQHtuhc/o4jFcjiIhU1qnNbdgtdR
mUakfeVbIOQWIWwZo5aUnnjavjbJ0lzswIjqEX62MPHssCX/IHULmxrrDlbsA2o5
iIk7ADyDZgCz8UTnEAfwLu7QdBiDMJprdv9NpsrJcYe+l0u8++TPQfoXUjdEVKnj
oOnYurpkUsbDH3Regyuonlz80828ivpKtFhfC2Fx44xERIsCnduF3+REl/g66riO
o0FQBf4T/rdjGLP9JXh1pxZotJlQmWeoASeoapoFafUd7ZUVz7zF6C3hX3sO62wc
LCqVjniAuu5S2yqA8DCc1SwtUOVxwRtuBGsL47XH8uSONKVVHY4SR1Aj/ESVRxJ+
wsE1Hj+Ff3ZLCVIdUmrdVVCmsBtdnP4bMJNCb4cqirnyxwOmPYxUxrzHLLch51eg
xrrSvdxRrBGwhw+Upw7EEJM3EV+7wUmVyrvg3cfd29RzVFwpua5qT4sdGwbyA7YI
qHXDph8ZaoIm+0oflhgwgIls+wo5reu45Xe6nqQ+/MipMFqT890Q9e32O2CqQH3J
IWrmulNmqVq2W86TESLHAye4ctwI3B//VFwx2CjMY4YzECFph0xy4sS8ZFV7S9Gk
QgImFpheMdYgXpAQku3JN+OmrMRrExfcw+dm7e2qS3ItlhpHbO/dbkGr7W6Nnv5o
Zd81dWilnU7EXiroghEAyd66pDqB85uFgFtqXMG6rO+Aeu5/R1k40dGZnmkyvxML
LtnmtbSSb6xDXaZZLbGPZg4Z3JvLrQ+Sf2nytCqJQKuHkLW30vUii12tJY2UW3Al
5C9FCBktzYPhMdU0CuA2AuBHRxwvW8xGk9cdsRbm2AV4hkmA7nvTygIrVH746hHB
VrA2upj2ylgJ/UMwUoCjiiOxWOShb4/6BcplyCPMTag8cYfbX7lpDRMK4wGMjsSO
+iSc62U5Si8BwWEnV6ShYM+xz5HEoOyfNEEzaslEZ+45LJDiDka+HjZmjHYBLOxc
4TW+00fuOUWVXNPucWrT4XxmOV78DbB+c5VuXQrmF9SXnpS3vUjtOBpIjR11XnxP
oKN6LZMqT3O5XVT6tEZJIixCYV8RcgaC/K05re3h0DqYBmW2BEyL1nyS5hjhCX1I
S1M1k5btQvbOcRTxFszLxuuSUOq639xt88jJLI1vz6S05ypRu8LZSPl/yzzt07i4
memAaeeIhE49QmuEAqa4rF+84QWw6+Gma2uvZd1WKBK+yEKr2mm8ZUh4O+iW+q/Y
KfcaeG2Pi+/yerIB3tXG9DZozh7ovDCl1kyr8SOmYhijK87bp1IPQs+HEYArP69w
0teefiX78dPhz+CoE9NDQ1FVjySdbW+ZVqPN6DhWR+AZZw5XCNca63GoHM3SVkoI
sX51INLeoU/4dV8SZ7Ou8IUC36kQ3l9UYK2PULc/ApfyB3EDpk85uZpa+7vLHcdk
wa5aKaQdPGKY1cLC8bye2oN57o6/4L29Bec2mkUxuy4UEgTfxoNzRl/+SicEA+YL
Ijne+AQ1EaeRcPvQ0EWCwYCrlJV1YV/nIfxO7GFTQlgJnic2KftvnAFvbEXRvwdy
fQEeZpX+4C4gJtQh/3XmmijhGR2sz6O7M621Ps3/SA9dxkXLUQ4wwH/KUhuWCvJ+
l1X5WuovlTrrJHOC78kdFLkFB2tZS2tbAIhyAU6qxtz/oP2fGxmS6e9gJhJ3Ty0Z
Ao1Hqa6KZrUqVP7T5hPon6lIk6OBxoFYzLrfb2DplRj84CqwdLrU+FeXd2kFyLsB
GZQMdp0NWHPzJbRYq+nFEizY1tcEX6OPZjJqyHD/iCkLPKAg9YoO14uYUVU8ygUp
mKNApc5kl02JEImOfFr/fVk4yzeJzwRDAqC1OAz6ihcanUzVDvIpjwPZbdBfm8/G
yEpP1QE0hHaLIqry9AwGhCZP56amst0YHPshT0/uxSgu9AzEts9hwHlY1FtcZTP1
0h9PoL1ecnvjeoslL9nx/6KY4hbRMMUU5OQHJMRiowJLxPD7GT247/UtWvU9VWfr
OjIwZFXH85Nk1hdgiK2LjuZi8umZ+YOU7HQ2GKwHnfLRneqFYCKzWRt9M02yINLi
u7aN2ZM60tgtqQn3BtSHXd72P4B29sZZh30zgMcs70PdgLOs3HaIj8u86Xpew6/M
U58jQ/6QHKiseNe+/yRvYs3eXuYjvUxg6m/9sZro8T5IsEyYyNIfdnwOt0bRpsoZ
zsjoVcMBJIP3fEWQZqPg8I6/hI8gz/zKtPwHR8fXpWaNJDJ651t+yABXFBijLtRR
U7HuXWV+VsY1q1DbhzN3Kw1f0Tc0fDpNb0v6Vkm3i/rhgz3Lus7RBkS71MNhoEnN
5ai8IqfcNDZtMUHpq4+FBJ0dHwYr5i7HbKFc2jxVpXTqs0QmKp/+EBPKXO+ROZhc
RKmu5+UA4dHPKo6wWmuD56iTeswbQ6vcffFWXRwNOJFEF6pEebvz49eLKWqaPMwP
lUZO6y6LQ4eXWe6B2GWqTEehWoStI2gujosL/JfaV17sP+o9pTY1dhdckaEOLP+t
/1zAXa0xqQTsuV65bsQOmtZg/JLy7gQBl5t6kxb9HswDgFrePik+70swS6JkQ52W
w9JhoZkHLYm/FK7fnYGz0I1wSODBN1udG8Dj1C1u/rZdq5G3o4VRB6EQ7YZ+OnEC
fsUYfnuiF8qL0cX/RblvgokhkKDsXL0EQfLLcRrv1ctCiNa5mu9SgMwSB4o3bsxW
1CqARLWh5nKeKku76ZTzlJ+BfqKELxgD0fxlBIvuDYwNwjDpGWJoIhL06lX+4NtJ
mV47KoHTTqUx9rDkMa3DckJdlti217cJTmogXjVMCMBIWg/EtAGOXC2KUxEq8Sg6
9TDSOHrwpvaVF/SD+nKL/cXs+6KKAn/TTg3nHQxQr96U/N9ldGkoVxcqhetfF0hT
KvrNJ/6ciFOA/vUh+b1YM/OSEO1sEOiq1H0EOt498SGR4tFCRa0zmTyVrgOL0eU0
ney226gCEY/7HOi3Jrrz0S1q/d8TbDDGCb8b8veMeXUEzg4OdMq/ebbudD56kWBV
6Oe2zASwFK24MZC72wSjvnBY1X+1Mnfp9L8NEHXhOBhiFpfkXTufb1ZaOeX/YYoU
iwRb9nnw/VNbWNuv4XSARcQF5OV8P7JE6V2KbqhtorHAGBlqbmLyyoNkSU3JRlyM
idUej9XdWANMUlCoDPnNA7gFX3diLt2kYCqQRG4QU+n7iIkmr0Tafx9NnQAhBNWR
MDkR0wQctgacgLaO0cADmBxcL/AK+TOjJ9t06ObiWFaRugx1QJjXy4yFWUy+oPy4
Ju9TrcptbJelpQUJMO5KLXqswmPvmFuV5ib942EbNFMFTwVVdeT3Ax8K/FaM3U13
aUwC6qKMtcENdr1Y8KSlwFG+W/b8NJGTt9z97tan734Ui1bYyqGtLI3tJGqYnaE7
UnXsmGvl6b5iKxiiYIvA7jGhStYPvDrPt0IPat1ELXdCNVFYEmUI3czneqd0z02I
ueE33aX7ravsPjU71YIv+i+KWvwqBLS/qQg5VJVE78r9gCHxVG8jkkE3atj+AhuD
0v1eN879SCHr4cJOeKA/y+JAZxHZMvxCXY9kAYfWOzwibJf7+4d9Q42mnQUpxlR2
LHJ/FAj4jPJSaRfwqc1lIKDQw8W/0hSZJEdEEY7nKhlLg0d/BBqgYYYZJPsjcIvz
Z5mHB9PX5yef4I4UvkmVjHND1SUnBVzGiVgk3KMx79GiRSOwYpWnMvT8RlcHtXpw
AWPP1F0tVuBkrwksVk901I/f8K6VYTVslemhJFU7OK2KXAHfdzHCj2qeyHJSq5J0
6zNlR8Os34CRoht43B9IgNFlIdm4JlJL+x/Yb/xa1BUofeiozCXlnse6C4AyaqTu
yNyDuDHuU3XSoagfJNsmvWwSiP66FVK/8uaHRN5pTT+A2w2C/Zt+Awuw9TrUh8MB
MclG2uPPd/pp0n+GbAAoH4ALFQ2etWDYKB1NyMGl0FNQTEkaRR1CeRCjrN2W1lz8
JYbhIGi/LejJdE6Xk7/4IrwOwJ8J5h2ydrN/9wtcm5cWWTCrCetlsuP/8CELIA7M
unFcLn52Sbdp3wiC4RkatgzSQW27Ci87zUL0Nzj91EZIIA3N/C5RhE8249GIau7O
YLFr+e3tqdX3jVpf0p4xNkDEIDMCC9DJdXqXnKvpGgTDkJNp4IsuE443rLyh0GBg
m8Ou9v+900/jW9hY3FpspPZVj+X+1PJMWZZXWZ/WzzP70777yAcnniVOWfJEojPW
s0oyFQURvn2+0pR6qPL4Ux0VN6p0ULX5TCiMLOAvqm2D7CPOozLMqApU08P40dQn
j5+ichrAq2iDuF2yhvKC4fl0RO2VJhdY1K8go1lPhhklqsnQf9FoWjBalL1uM7Ub
4t+4WcVgvYUkZ0o10KyVj4kG3BgCFVHeiQG0B7eTbBwOmdSmiaBfCxavXowEj1Vx
9MJB4JNcIUJvsnv5uucg35HsEQ3AlVECw6dkItK9mC6xidbVf9MesH+5+Xz4WjBP
dGWqbBMT1eSH0sTLWsrsGGLU4wmbQ9e9ohULHjpvsq+15Hgjxh+LuUowQoc/tQxq
Omn/Ycusvq6FdgAdDvSitULk12gZAhuUfB9KM8Zj1qktyNJM/HZnosQc1sfd5qsy
fD8tXUIvoIEXfRdyxHaZwH6uMxm7312mDhNgZsRa18poLLCeCcoQjSj2nhFCzOEq
fz4SxM1DQftNtfzFaO/wHeV6YyGVQpJ5ql7MFUBycTkKPd2MBa4+dpoEQn+YslgG
FP7aybPZ4ozbzP7nAh5n1io+yL/RUSgVcVTqQ3+lVNwlns298v5LKM0kSou9sCJ2
YYBHi84D1MgBF8VZys09Pf/bRdqebh05+vr0323Uk23qNH4Cbg6rZLeYY5uAEa+j
UP5lIarvJJBR50pBucHzo0Hsbbidq+vFW19dCqrXbWaeVWTrX+sJOyBBb9TquXKK
nWhZjwndREa6+xMTIlrKLnZwDQ6xZs8jRlAXBKeuvsllsOQh18LWPLiKghQswWgh
xiONJmOfNG1Hkj7ofVzJG2O0vOyjs8FlF06UfyI2e79d7SN5V+tzHZcKFGYVFTUd
GwOnoSRRXP73ikWHponWCLMNxeYRbUdAxfweoe/yLfztPYcWVAFXAul1pXdM8VVi
nAATyC6nubNHW6qOre9Zy/asPnSlJBxT1+KztzZdYPAz7BzO/qjDLCimM3+Bjuc0
ov3S14AKApw+EiGBodsXAjric/zrFHTGfuUObSjxl4F9As2Okjh0FrqzjvR9r1mu
PIaZfgAISSKlxc+LBI4ovYWlpup4I6uEI8+rph58XhrCBXt11npcw8JxnL1knH8x
YIURCUALdMke6KoPTxBP2rHgZEcxwquoPMQc99FF+JyqStrnxFtKX0JzBGqqeQWG
ybe9PGcF+fkZLYgr3dRY2jrBVsXu5/BaiVOkX3YgQScsEYf3CIaEQiDhfSkHaGmR
lMdVhSKLqVbzqnF1fQmLrIbvF+ikz2TwmkToONThCoMl/c9l/qnKzxxSIVE/UV8T
/r9sKr1Sl9GoM7W6AbNhL9hWTCdpXCSpWZXlO2rT2L06LlqL78zIGThX4K9ptSh3
5aByBZMuICs5fvfmXF+HiTYRIC6rj1lnA0i+/G0h69ijGFUzSeucREZVwg7HMd6T
JNbfTCS6tLu8f0ItqH7esapKrxbhnYbhnikG4lha3WCN+8W1ZOwheGhE/eYKKeyd
T52K58cGQsOUx4aal94qvIBpT4vDMJzo68oLXP50Zmpu5DjWN8BLJa9R2VyvENyT
S60KU3Bb3+K1WBP9ks0db7iYI42qdqhpbbayeGs4/ygxcbh7nWo2Bz9XIHZ8LbvZ
A221jrtQunJr2X/uESSQ1yVE1R3oFwRE87rH4+o935L5StjAAWOcQVL4k18ZuG3E
YgVFhEiBsSCVosUuC0NYLe9dAHjwIWqFcA6DcG6GblDOX8eokGKdWP+f+4OY+3up
w0viQpxlUP2pxgIH1g4U/OzJ7xSJwYtT+BK7kilozvgHtO48d3rVGICdkUXCvVE8
L16R1jZutrjn1vNrLCFARGlPqNFc8y5grN56qsdA4cUtQ+LDEqJ3QCiE1H3wZ+Rm
TLeywiVvxdjZVIrW4f3o5I24pSdWa3ibd0La+Af/oYyp59GZx4/YT3a6BUxcFzVj
txOZy5Zt5gpYXM0+Zd/g0/1aVJzhHpwDSx4Mp4LYrkmzC9RM77H/rbeb0J/uYQcZ
S0DNGQx8MfeLp4RZX4uwqV7WXl+Q+eGH5wshoTDheIaTx7r+353VB3EmLgcgfZfr
pO0hhQFO27c3HLeHWhyuDHC0ScNBil8z1deStnKPzzMKkzKoB+BKuWMq4z9xGoYh
BNxoT7RjXg7UZVt/pTqoYEePAEyje0iFtjHbBbTNURifyId97iEDqFtN7ellNvRJ
disMCT8c1OlDR3t0PtJLT92QCYBo5SvGIMnhkfy4dHQoWCzii9xo8yes9fhEtCdG
h3Z7zT+fL3FZubZg+edWBhpKW8rDfT+uc0bH+4xEApicbMNcXCxWQyNyD0T6ClUu
VWpxPjx9DT083LFnnPZih6yl+wn+weDAV2tvA32qBi7rr38++ejtAFBgB/5fdFFH
kaBGY3GxEOBRh047IzzK/cbvp2j9+FgAPfqFHgr2lGqLQMOpXgLMkQRDKyFenSR2
Gfr6DGrEW29pA/wZ7rd/idPovFgkFpNbgGHgtGI8BcWqKZNL7fVCbTWSpWroBXX3
ACPKDZqpOqyy9vnVYO6mte544m1L3s9n9fUoEq8ok3IkT+hbwqf/9iPtmKAqY9e8
XDDAv8SReyaaeAhYFqqAp7F1ho7WAi9OI3dd2r1ueApVWV+upTnwaxuXkpZyW4i2
Q591yaq8T1j278cC+aw+OFf7Bhv2HCeovEaYpSRgR/Rldk6/2ILVVDg7Z6SKvYpH
guWa8X3BxmEsPfqHR+Pz/oMDsukaKRXsMHuLSAhQaamsEtjitI3nRJagkYuvg3O8
8q8zgx7Vo0Cfjogbt7HI4/3S8NjO4WExYXy2VhpBfdAejSSbTs90A24Qp12HUFhN
uZlBPiiszJOmyBuw1c0uDpbq4reneS3cVl1pRvjK+XJEMsczFm6BBImN/+iJcvP/
9b1d6XjtP8kJ0WoawvH4c6hFKV1xZNntfh0bPMSJJW6CdPLVTZHcfUme7z9Bdq4m
q7/Gc3GBUplzWpDYlBhWLfTx8y6dfXEqY4ouZslO+z8IYiag1NYRfNL7miwQaJuf
xhkWg5n5fediXvE28ihrauKrjFWH0rUXK9lAih6JJPRhGzUrqklvWCSDBz7R4swu
+kAy1P/Fql73FFsyuJs7dJdb8ji51FBZ6il5N+/sH+wxmrQsjy+8eaQ85xqrGZIZ
SdxBgu7Sgixrme03+TPe1tJg2j19jAo+fIMA40DCQpl4V9ILYSWUzVLIrCs1+HBi
vg3TKGkcRIgAjKskwKgWrL3RoIHLvLBdC/c797CBX0uU87SnON/FQ0EI7iCf9H0b
1SMbujEvvs6cNvkd6sNgjtfu9OMJqUMZgvVnk18iL2yiJTOTufzKE73TxqZ5nXfk
sVms9EJMLfgUj/2u9j0iwEiR3uQPtDEltQY9yksVwfbxPkq0/uIUAm7w9Qm7EORs
ygihDxaD5uUQko4thq9Nh9QsSxxgkDeIbe6E/HkyrGRZTqJFhBWA7YlcBte+COjL
926e3T0rW0hh20ANyIwBsi9chq/FAYJ1sWDQTP5HPxtQCzK+j1mXeQyHaPNrfQuV
iJizEPm7rUMPOxcPxrwUa8SYRDx6QHqMIPZJfoHeq3HqWZbwuj5hU8N9HQ1lEyvc
92fh5pVX2859Ha+yoxSsnhuXb2F+ijRcaxXPM3QjLrzb5IZ8HOTtpNFPdm63ysBG
WSeDfg/CLYSSk6pFCVGzZmV78GJdeHOTUkJKu+jND3SurPsctpjCst7rHskP8ZBg
NPLk8v1Bcu2VklWBNB8kxCq1OdK+XmLlCFRuaCRmYaE5DKHW6KlOy7ntpFXEB4hM
xH7qg0ES419Nii+bY2EGsCrLTr4D5nl7x/7MrD2+c1o+oIhRYcT6m/4/yRjI1d5b
e+6OvZ6FkFOqGqgQvHOf8On/J98m6Cz+s1wRuM6Q/0cpaT/ZRUxDetWi3fYKijpV
R0D2obLk6QYFtRsgAdChrx+Ol5ywI3C4FNakmIyj/tEm8Kt2pWNEcdeukumIK+C4
oJgD8Blrbq2AEsYax5gc8hoUHX54jDTl3TaVl0zGOeh2OjPt7BxK7NNa+OhcLKJ6
N7Y3eiOZR5dBoJKs6LI2Hhfj3yys48h9KZvsH8QCj83logObtVjH3z5uZ04vn91a
liUugmIvJudGMZjE9+NTj92w7KM4TAu7JmGpxWKIuMOkgIX98EMgJT/gnDmRPsQi
VJcMd3AaO1NVRhGiDrQS0YVhI0uqTAEKczo14dwpc2jUjw2E4VMksD7VwhmpZi61
ITa/XLxKBsGZ7VwBC/a1hCwyLBHsIbFo1QHGm40F+w5Vr5So6+sXUYH/XgW+aDnh
COW981uENuaoNHcpBf+Bv52R4RUvroEEBqa5V1LoW4mjdfGujUZmYKOB15oERf/8
tWHkLylc0dVSOx7Tz2Aok1KbzECmna95JRGTtZi0SSBf0T1aKbg62E7VxaAdtzeY
d/oJIjDdBw/7raaQOOXVE0I6gZ65kFYNNhUuKDol71lCOvn035YvpfwxDcaN8YZP
l0p5cOCqmC08FYgj2//xLCoQmFvb/CVkwF9PmxHvhkxwLaZfMUVtC2NLyptoqQ3X
pwZTpwwgomkS86lNrLG8RutoBgt2MCnceKw29FWpPIRBn9ZeSxZKD+PGgHIzKP6o
2FIqY5FrAc3waKYg+iJqfeUrBJKuKr1HmX2R0hMc+Xj2U9/4zEHRnRDWRU4NyGFI
YKOBT+3GmHT22DIltEEvO8CzMxSgg8nVsqVVSweNpBeM96goLWVItYCukq6Gp0Sh
Y6v6rOvOcBcUhG81zTkMQhSd0X1OZtxJW7G3q+2m+9zkBCPnDHDzhXgu726mXjS8
+lq1gP8biR8gf5oRJzFMFPph9vpe0atHNp/Q2FmPKE5+loeRv9akKJBRCMCQD+85
m5d4J5XKpfoxioK8/s3Wy6T0cRlrgDq45KcyrULxxsZM0VqiqChUq3mWv1cyk0Em
eRcmt9LezZ+4lYBOSYaq3GPvL+DnwrM7Km7xPUDnnbIxb4/fMOxI1PgMH5JdGeY0
ACb56ReDqiJxax50wtAj4mfYPGZK14DTLcjR5/EjHFzuZyhqzMtbUUXvKWjU2aoL
nrgf/5bVpULB8dU6vYLlu99s9gVxwqqopzIyG3Ig0G7uo2fRe1oqLAnxfdBl1n56
LIAiJqirDBP+WC4oeIHNnkAF0QWYpbEXIq+plngl56rmy05hlOHQfP8MFX/SQW8R
ZAywRbUiLSrl/k9rioQKBF+fTc/f2BIl5PWAh5n15zbaJ6sdcq3phiroRC0zbdZ3
7HeskIQTQMQtZH+CM/Rrsug3lareImvjuvwlRIxbPYYWRd9oR1V+v7EZ5Lx373wy
2UWNg382H0myj4F8ygYIn7cNFUuJXIlttYw57r9OPnZmTG97ZBtXr8/JncqDpcFw
+T2atcW3h16SN2x1kYYGxQYraC6j/fmvJwkdFPvSkVMdte6mVKmdgBFU/ZyVl4ol
InwAzI92QC+a/AIXCmPfnT0dfvOgLLMktzaujAY5R60H992+HAimxTs8SATHIyaj
7+XeccsD/JHUdzXji2qXVOEAsUpzB4UbL3ysumPNqRWzTzjrOAyQHwf1wYBbSi9g
U4vvd+AkrP/Yph/wCmkh/cl0CdewtxuVrGwcaKZQxzp1gseprcKD1FMyCPFLbcUa
7KftgEptFiZ3L1M5Fr4+ytfihQtHNA2JZehAXid+3x3vlYf3ZNTn0QDZ8205Z93p
QXdh21OiqK3zDJwEG2FHTqP8jRzhcFlklcmmU1zbej3tJtWEkWqHY3JWX7bWjb5J
0YckoJ+HPUZiH6XZej/b/+39w9fQMW/eKY+rsZ4Cz8doU/IcBszF1g/+ehuOMsXo
oWqyJGxXCNYVKgYyECOVzt0hEpTBAs5AS26Il6mQxD1+kZXaAYucxolIj5GYCjsn
eV7tNm3JFpk+2cgQwl1XJioOM0FkguOcCynEusDGobWeT96r/Mp/DtJsgWZfAxaa
TgXZSr2J5Odi3jyLBv3qwtJ3LGf/fGj7IGiJpGQq+VYWInDQgLmydrOstjSKiV9K
jYQbqKlyIpL+16XWr0/RVF4SyCRoksNOunWTOrzdd0kMG6nWKgmKacTvhQfEg80O
1+WjkuiMsKwh7CYEGHi2mQZ0WTfLYaKpw7w+DrIhufKhI4gvV3i72PYLrD7RuZM+
z4Zx7W5dPQP1DKrqeVnufAZPb15kHmZlex2xFJp9yqHQOM9V2aUHoJ7Y6htt5VTT
OUzP3DSMObDP/VIb25VklPRk8cmWCJ26VVkY61nzHHWwjgKyC9vd5Hlems4Xo+gm
7eKwJ7bZcJQQofFzJDrJwpDDF0Ydu5WOdzNjTxVUXSj1m1+cuAplmIu0W1yKcre/
A62Di6NKsRzd21y8IlZ4ZV/pSIBAG7zbkeMTxanOGQKHrLmfC5wlIClOyx2qbCjm
a3/SGDDO1uCE9yPWxIo5cHC6yktfKnat86NCA6n+39qyhCB5JAXNE9g9S0S7kZle
e589o7hPW24Iga/g7tBN4Ge1Km5KrBZ3MqGdGImC9/7HNd/X4gS8FHef5Tqg0tdK
Y8BbnvsAM/f6AesZMYPfybGtwBdPYzi9WtTHSih17POCAtW/xVYdqGTBv0EkSXaZ
eQku8Zt59jGaO1XpnzQ2kd91f0jXhnxITc3AF1+n8BfLuVlfdWCphDQkqZsfSlhl
1ishY36aoSkZ4SMqqFOsMiwauN+5Z9juquh9C42/iCETuQjGvYle4cfEptaDreuh
Ra40AaQYh9EjkDavEmrC51qGCYIowfCYPJd32NADi+ClpNG5waWycIffV2c1zr2L
F3/Aiq46FhICwMDQX4W6y+YbOCbIuxEV5Og6sDeAaL6LDGT4XzJKWV6t99WTDfKa
DTe4mn6FEVCZZbbvSCQ5y5jOWqcqkGLoifSiBuGuL6wH6RYPXTTrdrlosDqg9IUt
lNtz9zL6kVP72ddnfJjTyXZq5EqGDiPXugl44231IQ+34xdYo7i4rnnmphnm+qeb
5Ao7xv1wKG2cKK4HVn26D5s1/GTHDsDtU+BOB6v8D0i9ab/XCnxUo5RM6+EenkRF
/LHkO2DcsL5yJoI+zWL4DBFuE4VqeoKvpG+1TY9csM+3xVysP+fvt2BHAgjzOSpl
q8zpk+Rk7IXZJr9/8Y2gZR2R4BoQ9dJ1BmSySHvREml0WniQ5+XxYIx+tchQVVrV
oeoYhvyVW8JKDaPTdmkek0Wi2Iaj+KGgDzaFFAxjbXf4RvIy0h+i8offH5yn0m4j
cEgVoehr+/Iy6PXRqivzgxkCuh5I4lKcO5WoBUh6P2blBw0PgEHOL0v8FXTRiiPs
ys/TRfGlf4BNBJMmloZC7h+I/XgPaObQMezOua2PZ1cEe1OVQyOlZH72VO+EtFd2
fDZeRWCDQDsn0WYo4ahbF9jzCH1zuYyRIn3NMO11Ja8jezIVte2nncpZVtjTfWKD
PKOh626xXUsv9orgk/8qouLJjPK6U6uGnG2DdwX7Rc45C79aC/VmyJjn1gdgIvqL
JYbXTqiEFHto5ZeCYxSsYOpzQVW6xuu2t5mO0oghyBpi7QBe4rm4gWez7l3w0ugv
ujiFr6l5om0k1rLwfD6neHzfDo3gWR0z+VJ+CJojX6O9D6id1UCPtMWOgb3o2/0L
T/UQRFqTBlPZpDUk9A79lg0bEI3reEUbAiarzEwJTO7uxDIr5zLFKYQatfYAZCVs
+frwQtr9g7MQM2Gv+rrPy248BtcLC7du9/uoJJWqXy7p+ME97IGQ/iz4ilWQLzE9
nOst6VicSm88Vp8fOyizW2gIeHi4HNonSRphDgmAFJXzShYsYnlCae52NbpqZCaO
cUPlkzEZahTFHsaA5CxJg6S90k5/qM1kvy7sIXgqn3W1FyT0FZ/pjwq8lYsi5X3i
gwCjOuhLDyxKauo84Ap8DPsjv8d5jqj3ySpOOJJV/d7r9g37DnMoJXConBLlp8Fv
pWLNATvoY5w3jM4df9LImWGJ821iNnU+AJw0seAdH0thFJ2dwjyKiZQBDnYGVLjz
aXR5PBB5626F6PiQkUbCXCn9Y6k3Z8so25DIZhSKHthurl2zPIbTeVyOoxY92z+j
n8woa3k54UTJ7iB9YF++55Bt5q7iDnIkJl9SUc9V7J6qkLa8HFVd2Fir+g65h/fX
lFOWWPdD4Tb4ufYQDPPHHg0GlXH/tgT53iJC9kBZERsBEUYxejHdXMPD9MdrttiS
6nsMKrLnZHV9mMykHw4kqt9TBer5gAKR9MIhHx7n9N6Owzep9P1cEvcsmm5u6avO
vFtBGYjNYuwtjDIJEgx4ttAUe3bQW9/2HLvmAlwln5XvJZjVaaVAaCsxFKWG1CLH
Gs5UTrYR0g40A36cDZTuIFylETAyHVf0+uP0MzD2uz5MVxGjL3rWzkwRK8Xl7PCo
A6W6cckzSmxfIuMWu6AMqXyWXnpk/EI9RQ8cEerVgHOfJAVEn9SPZyhje1JPmacn
i8RQXpkZgm0CHoFJUnO00BMTyDbC3QJnaL1CVG4G7Lj+/EG9uZnTRS0NcTjWC2iK
pJr82mpxNjfYx6lMJZP8R6FKyCP+7RQPKDQX2JbBhoJ8YVmkHOp9vtxUgsNDLw7x
9pSm4SgqDhNJw0v9TaNTujp/1UnX9SIJRQ3oaVr/ooKCgAtvCZ7y4KRD5zIv7sYi
lD5W7kRJBcsSRov1fZYEdCt9VRcjNX5hgbsopeBqfhg++qFMPSXooO1HoQPvc1oV
DVMUqB2U4RFjs725Ev1IK4hH2am5Gu4Vg/2XviJBrq08up1kUzy6A8kQS5XxCpQH
wApl+EuRKuQ7Pr079u37vU+4g5j5aCfYDqPkVXHXpJ8zPBsouuH+qVbbOqVz3FXv
fcOUlD49ByerX4qkM3KFvyNL1Sq76bd/l8Q73ybkwu2PIqmkvpwkGEK0T2Z3ptxP
r2OtnDYP6eJU01L1rbgs0yoCELSfu/8WoJzEBjTW4u3I2Edrjim6JhYU7YvAZFZx
U2B8WaDG7fInr5rYftCcf5Oy1TMPV6ZyPLhnAXz18jvGoJt/8Oxe/VoWsCqVbx+l
kWXCkS3TZXN23Hci14545U9xXd7o5bIdxSdIO+yPeE6fbL4/XdaXy0CQbrSek/Ec
hI3JV8PkE7QnCCpykAb46GwHs5rxvPoM88n9JHot5SzJfWa7KhkfYFPdHgfLHlbe
sOE2VzdxooqCVlAO8Ud21puAX8qeSlGBwyNkqkhIDhlEgeUQpxB9IY5++ITe0eyd
e6DkvTMwqCSG/F5huiAJv6ATnxxw3fKqN2MyRkwbD0WxcX+JPHBFTE3clCfhPOg5
knfSyqz8IVgIZD47L3mbAB8mnBT/p5O3F88gZtuOEV7B3s7dANFigil1k31ztcdD
KrhKMbXRPRGb+ErhPktjTD88Juj7LrQ1iy9+GP65um7n8CBdHdThypmyM9xsNZuU
TLXFKBpuZTv4iave0v5K8wLGEp9PXoCfLGLMjF7NP84bNRdZSWJvXXSvRZCqWq8W
XGKZdk3m6YK+O+KREnSfRnYFBTlIFU4mbHEA5l7DUDcC8CboPFNgl0ZkP83WTlzQ
ZsPfxW21GcHFlG2yjfaKmwscvRilfW54H20Q+XT0ltSvrzZ1Tx6X2iuvOAMpH+oo
k3MxHuO2WzETlMcywb0MerJnehqjFBIiKnrG8lWSOquYlpY8/jMMmTkW69x8rIjM
1FthHxgWL49XEpEBT5LWtVSJmncJBmAjtd1aGlYMb05DekXRlxKBcMCl9LNN1pzw
yb9hYki+DDpawlGNkGyO9I0Em/WDkKUJjKKrbMaai8NBsQKsjQy4ztR8ezHVHBEt
x2atT2JlNILvbF3KIBgvleD8g0aa90D1ofb28j/gin9taVbq44CuDs7bJEIT9454
ihDKL736efQ3B16KR2BPAperZ0BKCh/x6R676ajhtq6yTCSXoLZobAIKZXmRahk4
hSSXv949llGhwlLfXvvcmeOXSoSzDZf5KkrbaIbDfc5pW8MDw2ZUebHqyAkSxU2G
gEOkECMy8Jjad6RVyHhsNmtKiF2hiY8T/ecGQHqu5qghtnv4k/BE1LusxWAN6EB/
0cNPJ/+z63rBP0/baYPqlhfPjopedTkDMEkQo7/qA40DWy52+fP7sR6oJA8ZHT+s
Em81GEE29yt1s3IqizuHdQXk2HGc7Ruqzcsj2StxR6Hrc9TVXBkwefv5SLjhnWUm
nyc94iI+eGzp+v+FgR2+no/qMIHwxwbN0HsVDTOMRVlNlucbkFWVAJLWMmbBBM08
ArFV8W9E/X4CE/6M4W1u6V+d5ffaps2DIa4t+O+CN007lucttbcYlrk2oxO9y1Tr
7I8OsHfySLSZZS+Y6fS11TkCtrrobRz3vuhBb6T57dEnUJFrHt49Hnw2OeHE6puc
ahgBPoRIpVlOL26OMJ29CuZziOhh+88M3pAoEOQFEvSIyOWns8a5RSvH5WEu04di
SRtgQKHfeLphgiyt1V8L4GTuEpZeNFeb5NjyO+mbotUgC6VO42NCYmPVGk+G/VPa
PI4s6WvQYMDn1Jdk3shqGdqwJX7uTVFTo/XeXW+ZBpmR1KVSfObPPpN4/GRgFQxb
g3XbwVwIAINxjFMKnvrUyGFfPwTVNVHIz5XdckPYmVAUMy3Rxo80KTwaKq4hk3ml
e2l1qwCCvFKWTuF7ON79mTGT+EWtu04jeH7+YtL92pVgv9XjZyo0qaZzEQWd9CLu
0JVWErLD0RcxevrOlvfJQkGzHSBgz19B6GvXNKeLjYb8sZ66lW9KXXySrkSZWYWx
JTCV71nqylpEpl3IipznextaHUSiRRSxUjpVh/UJ86vT5oVQR4IRWxWM7453Ds8Z
KKD/WlL3S7EAZAR0KSVacxcTBaeVEq+KJuTt2/A7ca8d7x7rAsX6ohHahqiXb3Ar
HRH3ao6D/UhEzXPFxEj67YEh17rtAEvuN566DrYDeylbbIBcPvTlhhEqTzRQz6Kp
iasWjAVF7nPQkVLXKjPwDz+gHC9dpcmpWWBqFTUkm1zJ1+/UnQ3qIVjyE7Iz/w7G
5AUA+778hG9daV9PpkzgQThcS0fXyQn71TpqErapOn4FWluT/f1Y/Ua6Wc+12ycg
Dc9zgbN8Suz+Njc75CbLAiCsx8spIDZiYfBO9sM/kYkaFuZ95ZZBPNg/V1eEogXp
AikwSwH2rKItcy7qBIF6AonlGWA7w9IMNFJmoqtmHPpHCaz1sx4G4Bx71+4Lxf2m
adz6iL3A4mp5XfVB8R7Us+e+hQJVcuOho683NzXhSwz68O5tBkyDngY2o4z9Hpmh
JrNF+ALiytgGFS+bGRk97j6oJY10pCi/5wzEEZoUUErdVuwT5v3Np5f8B3KbQSTk
ozHKanpefoEWO3eFwD7HW9JhzlGDD2QPk9OYD/EXPV4jI7udQZ9K1wgJIISZRRLo
ZnW8pJZkv2DEJyIuxpzFEJTn2iFtklgs1qxkc5pMxrhOThOGj6RfPIPSBB0yvSBe
02YPn5mFZJGat7OsW0vmyzNUNB9a2MvjVz6e7q/WEnd1pQFrEE+rk+JmPUpmC8EM
Xd+270xecLpnF1Wq8AVAL4O1KcBWU5sg4RIeq39lzp2E3ySwsYA8WVmt/4rXb1+q
E5ZB9ewMjOuY+cbsNWhxrMdDHE1I7dozWrzsj7zE55eGcgSehQzgjg43vwRyRugP
XmPhb5G2UKQUrtCobbXF22k5kI5YK4lbDai+GL25U4U1/pqhDlTAGO/gTnaNr+8A
zEikNe7eOmutSztoilCBghtNohL23Vzcw1SRRcg+I2EMY19Jmmr7qn92GvYWJId/
t9hXP8CiBOehvf5pSYtuRggKDmsRpnLbhwCbXZQPMzfnoskjutyv8HEGM1NngQ/+
5/+fdh0BEWI6g7c7oHQ0nL2z0QVtWQJ3+kA8pyfT+zXHM4TM1T3L981XPq6OfNN0
rywYIXjqbMjbMO30z29+7v3Si7bpx4vMygIg2kIau60942XHWRS9veuwPQRCxv1Q
qOfG9XXrEgWgiclBe5wLyqeVMO8Dl1tucxr9ymmgpvz8r4uNj48s7LsIh2Jwwb5I
qVmQipf7mA4aWqEk+F2k+bA+sPl4B9ZNk9Pd+l/rY9hvLBFkNWNsekAQYccQE4dR
FPA/Xagzhy/B8GiOL53jGbbd4TqgMFoz0kSPdOXFEv7Rlp0OloXDxK2HH6l9Q3bf
vCOucZmp8da/tCguQ/FIA7cAUKqcgyiXi4+8aC6uLLfIvRsKxvdvh6/9a3RTBYR3
+1wd3rCFgSy25MQpch1JQT/TXq4V3Dpfef08MsXp/2qJ7zkbXvyFugkw0uf6zt+I
Ocp1mqq0PpmNSk5fXJjzxdYQ/kAe1EYibJCzsSkFuQBc+5ieFgXFq45p62XXyXyf
8AemtPOTZgQQcZXBn3EcHMVJWGPrPhFL8fYR5Zk0AA/mqWRKdlvtIeA9n/IZbhNj
aYL/wa69brDCZXAuDrbn5MJ2V+ykEB8AQd5vCpxMqLcwwAkiUkp/IBD6j+jZCcZS
hptUH/TdgZ5CQXdtvyGcDvTOG5CC7XdlQy6tpd0Nb3stFP5L3cSrgy+lXJzP+0mT
WRm5OZRIkoV4MNvB3kDjTkxS73UsZ+LF7GD9xEfAhU7pbvIlOJlh3mpXFEE9BAcC
SzQNEw7fNbtAEPKywWXzi/uJRsE41N1TtLYrQGVyGZS65lxLlHPftUzj7FS5Y2K5
2i/9ZhoH+YN8cRLp76Frjfol5IIPAKWOkNNqEnfhGZVxR/S4xpN8pAII7yGwXO7c
EWUCoyVUeccvD2Sdx+1kZwKqoO5OSN6vpp5wdiy83X8hAHFfqDGddglSgIRlKABy
ymr3Is653Bp3Ib9qV376SIHac49ico1SAfLbEwW1+sZg3ezCAS4M0+VKaR+fEOwE
vhUJLeNcuU18T9o3YPUa4r3WHKlCUO95CaegXbs20BbAW2CrkEA+vQa7MlVrD+rv
syyxTAxs+8xoOUmvMNSBQtPY9Yq6bzsFzFVqTqE/K48Y2UHJYGyMTicou3ABUeXq
7qZWeEPZo2M/BGrLqEyFgBjPDSmkYMx7vkRJKZYTdFyUdcMK3jzYcC+la0PgIMqa
Huwrh3OmQKxnCJ8AMIL8ZJsvbS608LKCStpmLumC/cWheBDz4scYc0gLoaIfOqac
AgwCQ4GduOON6ndd1Ph38NVHsSnMehtJ9z6i+VDYSuurIcfTGiKAaeeEPh4tk+P6
uBEvAOUnq4icery9HJGbYBQtb5RBj0M6GM0IFo5AjlAenArTqku2Xu58rx53dl/f
Bz0PqjHpLgQkJLPpmpobuQS3Zf9eKLAB6LBTNCOfIM+VJvSqePRf5xQtySedRVWO
MVfDpyiDwsa7eZrYuLbasxOsmiqaksBgEZc/xLLH8KSdIvXurQO7Mc1+admGFEFM
22EFzoGprXL+vjp/b/tM7CmexyZqyPColwpP0LDr9zxYuXqey7Q7Mqonoaii5j64
GkA6DJTdUrrPefh++2tR1r/sVjt+WC9vtoYhCzfODJJEGLrWuIlEDPwv4Y0T2HJk
MUWf6Vg+W4MA/FwPijfcjBEKTMT9H7QSXrPwGQenS9epzszCyze/mFxffMcFecSy
kyXiN833CZfxAj/8oQpNJGMtyAfY0qLvalwfHRaNfx5HuL9/DzZ5SOY5YcIRjv2S
r7hVngtSGp57LD49Bgclffhi+LmmwH1bq0/YmHpglQVDFJGU4DZhGE4thxtzy1cT
jarIXXxh8EElRPN7rb+NNc2Ww9YRE3jfhe6a0ed+UUyLWbvqOG+nkHhvDKcivrOg
UaqOMXBtgTybV1w2g++KLgXcHNugRpvnRzNQHgX04qm1dw0u9KuJ8LdqrdqUdDu3
9mqAsFspM1RvDWUOSAnM9NcnSFEgwDcJnukWWvxZqBYNgELOZxgWStRR4OOW8SCt
xXnHTK2FqjtncYCJT+ueeKya/tWtdrK5HGVSxaXsq6UeRAH23TRVPrIRuiWsNf5k
moQjW+K1ynfUpCeWDee1nfOkcj+2TpAJ5C6IygcJYVe9gtq4VqZG9GNZDnqOICgs
7IrqbpaoN51Axunh1FyNa3ssHm2Bsr2L58oVzKH/meyB6IzyoF7r0a+ad54Sl7An
sGbnEoAe6QCr1qSEz+Wri6ZlfSA6V7RGQn4Qklnxd6UeTLBdd5VI3/N14cOSfgdA
BLF+MFH+8FUb7uSE/WeES+TXcET2MCHUbadgpmGtn7gbQj+q4lxNIQqCvLX7SLrD
wJBuseyCSBYCoU1/RlvnEF4I5SWNqBV9jDQSWOxWRcHqAjuW4SD8V0iRunLwGbR9
RIvGDxiGPKEfqE4O21DEkbn0GaUP+twz8JeBQxWFNPIEMfcsXHxx8rcNaoFte0il
1qZS1fbZrh3vkOu9RSTBYtQoN8qcXP+IWMjPU3AUDU1mrVCQ+QqOe9eHlKlQl56R
TivqHZ2ehQ2hswqZIqs8BAuF8fvQOJkjzzUwlnjohxbdFZjThS4vZQ1qL5DJ7BIS
GeuOxJwVgz3/1s+FXAKt+lNcjqrXJUFyEX5Ra+UKDiRbUfWnczlZaWz17y+AkTu3
lfOZz8mQKqqhOk04hiORa1XbtEiqGzg3D5XLdWLYvCylbe1I+B/ywSe/rmj93in3
H03TX0grXzyKCVxXSnx2I3v7JPv5RMQg/VAO6EwFHfO4gISAWYFVrMQtosPWyjLl
hoG5IaCoY4NEGVFE5tH0g0wGICYp/QbHay4A36jd1aTrrHH7QJmAR2JJzglRb7dh
5SZLBn8FvYjHvPssi8ecvUq+ZMeQxjBVsInll94Gwh9W0mJk5Fv9pMkGQm4ZRQdg
wHStZCw9O/BnRFeXrhzhUQ+V8J7X7YGCklhAXnybnYqgpvnMrbntwJO+nQbBeeAX
NEYIughLa5M/FoRBO3qZVQsEoLVkCuxyYL/JQw4lOvAaDiVpoD7mYUr2C0lhm7q5
ph8uW9J0HubE7SYOSnVpOS8RzuxbwEL5UYj9lRPmdsq5baH8hIJdaYBajuNwrhpN
VzTpPJiI7zPVwrL6dDmUCjhsQPK3Z9deXvOoWvXFoFr9jKikPazpHBVIBlwX36FN
cw1obTmVXh7Rh6kcjUyEk0PC8oj3qa5zRkeE8SS55cq3nolqV2I6Smp62Dam5n1n
Ld9AKmTBWsTgYrPPq93143Mt8j2wKryaVjTiCaqjh0y8Sj+FNKif2vXy+lu/O2Qg
wAkKftFL8H4q6ATQ2ulV13joSiahel5ml6P1AFHI6Pf9S8Df8iluOdsMKHdeMNlB
7J8Y0jomNWMQ6U4YauMTKY5/dLiA0GYyWEryF82hboqVtlHuxvs8tVSCrVYhvdwM
hl8AL7h8f01g52ysCSeXbYaOhc3b93GRaji8Rc/gAMBe5C43avuo97yVshaBDvVi
ACU5RcT8xy0wumVWpDBX0frVxniF6C4utu6mEe2DVw9nL/HYg47dbcAdz7xykQXv
lK/6m7V0rxgVvRTGr6IPtbfs2wx34BA46iFcU2qjV8cEo2YML4oyL+EaafKvSJcE
NzAsv/8z69FDQXvXThoXXV1wC3s0OT/JoaMWoCsSi3QGGk/dg11dywHJj/jaL2oy
lgPkQnKjpvcTkK23KBGUU2wsZ8+PqVVHxRLTpWcYiL73tS2rBZHnQtKVqWDNf0Cd
/2NhNKTHLkaQYrr3NZ1W0Qx3n0I3fqHS4lNyZRAoqdBSRHQsou/V/4jZqpA9COO2
BZP9o+yPsQ2KYyHsPOhbjI/zIPF6aXciLxMy4GOHhSVXIhPIEIAHVDVgEYOUoOrz
D+3yWPXgVPxiltsZxBfo1nYutm4y9DmEgdcMUco8YxDtfMwBuMzh77/ybR2iUJxw
mhIwU1DjV+/1zzPCIziPlP3F8OBsCTKOUwS3M8/2y/FgjFv1Y4J2MmmbXvV1XWXP
vo47L8Z6HR3hA3X8jUXDLwbKHyzU9VDL9/SOshf8Da1VDlbv8MAkL1pivmu3T1CD
0LmoH8gFj48EloKDUkwNl8Q34r1CAD9din+/lBWqG9902xshZdA5OCuP1KD58CYl
rslGZ24UNvqxPo24CPyL4EkojpSIN8D9JJaGl35ZObMB9Qfedy+Dvbqx/em59yl1
WVPqCYF0/K9AuTVDIkcXuivqgMLfFTD0l9T+YQUaK0iam5yr2svYS9Nd7nAXMDSl
GryuxUuL6aj7CtLePFXvbBqCSR8pmhBKMhkINmA3Tj64nzjOMfVF5Rdw+8sMWItb
1eWiC1I//1smfH1il8SPu4eUYU7AN2oBwpcJsTW6cGkUEtE2XPhviWPXCsJpdX0u
r0Pyf3EP5dOP7SrKbrK3M1pPkcd3L5Yfxp5HxcP10pbv6hGpEmrQpwEftlW8YjVz
Z6fBZmtPS1W6QL5YVqEkdfaMgKeN8zc8OwDaaPQCf9bOF5XMrhdS9wHCF0hphZfC
Ie04/jw9CLa8HKaz1fB3PWK23HekB5REysnhl5Bxpx2tjtoKyGoy9+cbKOsDqK1y
BnzHBovoWZKb8iKJrcxm8QOB8vTQfeVMylEtCQd2fjcvvjmssXFVGgSnlv2+PAoP
qewT1p5If3Y5cehkXFk3Uczb4KxRfKbpU7T8JN/tpbJn2q4QSnPcgvTHxaILAyfP
5FOIaGyjFiftkjzf9dtPY5lMgBq7cX+EXUPNYQ7Mh7N9RBwhch0H4+H9YzdEhPfb
Pct320oogDVrJz6/sYK9m+rcqi4kQ28QQBMLk6HxEd3tCo4Uehpm1VLZDDXoY5vf
cgwwCJ+zoNFWy7cw+5++MQ08aCFKCHVn7718fHTiZK6iH82RlszpnE0uT1/TT7DX
/H9pft2aW5qRGtahkvqbnzQM5xSf9fgogyc8NQcf4ZzxuiLcvUqLvf6gxOhN6QLZ
TEzu98p2GKWoziOVYP9xV+fUEV4BpFFzhJoVAJ8vZ11zK+uMdyU3WZ9HQxhR+5lF
FyvnVp3VpDo8xs7Vkt7LL/PnVfCMxkAO23sWpknbWiWnykPwS8z7bVHLzYRkEyHp
oXt1p+1rZPT1MwKEf2hcoSyPIEHA83XmtfVs4cvT9R2ZjRXQFEfwUnUqfCgMhQmo
dRIvLayh3taRaQRRVjuNXld1mhwnU9ze2Vf0ANEpgBaW+EscS21/OwWH2/I+33X9
LrFR111JBp0nwY3ST+CBYuFHCGOzFW3mq0BbBTmqP9boUZ4rwN1zjrO4H6e/kkXo
LJ4Ix/Xn4j4KO+VRphFGoXQ9DNIlh91ACWS6aYriOVSkFFEwLFtpStZjmODnfbiG
Jga0sS5TEw4SAhz0QFQ3ZP2ITYBZpmKuY6L37WB5CoDL7NxnKFTZaNPUMmLJVzhV
V21jB6Ybh4yxrVUvibzA5M7uSWXZ4npI7U+dF+zXTlmjBFY4cMqI7KjT6lNeqXzg
aFbpc/h8r51EAPfsTLws9Wp8ooO8bLBmE9qAcjvFPW3xFQTMZg9/jYytr9IVpXIO
hXwdZhBT7L5h46PCYW0K+PJKj5yGW/QCd8Jk4oPNW23Yx21rVmOyThkKMdPun779
go/gYqYN2GOGUeh4kB9u8TBerkInnPJ1qaiczU/SvgzB/PK9dRpSh79Xt7l0KB6k
LQMVuKRRuV3M8NRbgfO9/FRE+m/fc8/YosxtP8TjwXBpta+tk8tn16Ksl38OwNbV
6HdcTRUbHwJoHOIB6R3rS231gZiV1+lzkzLMbDmtr/DTnJFQv/tRDCe2HR52xFim
tortKOIJ3SiZRgrIqgR4zkoNsgnb95cfrNCwWdJVTa3M0HioeVJqyfpIOw6HTH63
LV1azMzRHmI9ZyY67Mmq2qHt75EwBlsdsmb5ET0wckSS0gMgL1q9zzz1h/n3fxMo
bgIRKrbzZBQE2E57MuXBA7ObcaVd16C7js5qnfssuXN0uEwGpFjZMCs5NLBPf661
a2UPQPvxU8XZYNJopEjln4N3P2tLe3IVfvLex1ImnvQiD7jmN8/8olAUb9s4V6R9
9EL1LW5w8+UebQD4IN1GMDc+O4xolJ50WuUCGeOvpcC66yUevRrZRMjn6y2hReH7
VNcxkKWjmz6SPR1m+UiI9GqjpMu48EJ5v5GnYH7tU5PBvgG7sWXY8ABmbckAktzz
jndMS+oUjL+w/o73t+aD6q4ocAUorYfIKl0AnCID2JxDpAZd7J6yf2Cmf9rUjHdJ
m356CVKJaKszWUecqWCumUe7q8/WkCki+alzZzp2NGfSU1D4volvNpnUQZk0OoZQ
PvyW8Jr6FZXRJl/r86g0oEEaYFoHyb7aSsYQ8OqzpJdtWcGToU6DewD4GoKIQPjc
zG5QGYOrFZgoa5DxSWQULDyy5jUHoQvtCjt+NT7KmxF5Bi9ZBnxVteTUdghk8T0y
0c1ogJE7K0y/M72Va7dujZONfcD/5DhzVUT3hXrHPVyzXntwwgbSj9Pg/s6PqF4i
SUKj1VX3EbMOGAfT/INbV74CpE4ronS3vDNNVKal7S6EffcIT+uZHg9q60LltNlO
VyKKkZb/Qu60KWlThZu/XUXgzJeAlyB0xU1av8giLumJ4kh7um7/CJK9XQ78TjO8
9YXIqbJRO2n6w82dLsfN/rU3sV/8XgjH/Ps/LNsfLN0IAMbxAhCaF6YB0Qq4w47R
NMXJx2mNbFMirYbIFwlpT5NmgPNdLb3dFlCu792wuyeXdH/i8kGh4GArXVEynECr
6yITq3dFKz9Cq+Gi0wNCq2ymImC4dkFOxB8wHVV1YxSNkB15I+FG/uWJrN0BMGj6
nc21zQM0oC8dZ66dxsnGhA8XX9R/fDDwBME31pdhoKqomAIJso5+dlpt12bm7fkh
O5QLdPF5pNNeKQ45ZqLoVaZmVHHyPR8YtYoKigK7aJOKkuM3UYuUXrsDwm+rYV2M
Mu9mT4EvVADUXA2fMdDM7fterceMqSb5x0dK/63fWHfsNlqy8G55Bc/SXxx7qjOW
s9EgZ9KXzVvrPGUdtljfe8QsG+PFLsOKlRXATphZcsnVxM+7kAInbqTn4jEm0eb0
5p3qdDsil4PKHRPleH9qM2B8LdeUBEQ6ycl007sNTLMx45BdxkgwQGKAVNQ8wOUv
UGbnnI6GWMaGujHil3y+4heBK6TZni6goauiTz73+QiTEMfS7QAR1nZUCLOkmFW1
w9fe2iKnckL6QePfWVggTNTWve76tWKdy1kEQJzbqTOTTxuF+9i25+FrXvbzYPvj
LWVL9ua6Rprvw+n0Qpmf0j4bP4jg/5BWMnuEToiQ82Z2MvLjt4PCK7W4Vdp4NrEC
3Qni4jHZBFyyRElBrUvxkoZ6RqnRQn/jTZz4ylJ6y1hZvmZMnodfsarfEAYRn3mz
LFKwyK2LFqy4o9GT3DOTtF3K9xFuKpWraRMiJ1gmw5JF8hUkAKR2aEkhF2FWFvR3
Ns6E7pUu4vohfnMsGoGQfqtYx2kgKMqAZ6ErLDz89cG9UfJUkSA4vDoWVzSIInaD
GaeDedTSX7q8ljIEgbrTLouTkC44y7aZ59xZsDDijj3bA6G81oKzPcgIbYvw0fh/
na3sj41DhHKEOcXJGPz1P1oOYtSn+cSgppBmHTPYNyXjZ6jwBj/e5KM/OR1sXLsx
1v9FL+tuqhEENm0ZUhpoIwyWuDefsaoVaBZkDw+dpbruthU1SeGoaEHGbQMIpdAa
bealshQbN0Jo2d19QIx0Mbbe+NUKDTYZ/hNOTFNHUR5W+rhH1kqeoougXZr7Kskr
FTJWWvCRGVou+geA8PuU/azfUXKj5pMg9Jln97yldK0pYNxZKht1hJIm/9Te6BJq
d1J9b0q+mAHN5LQ90tWOW0XPQnA/WPO9dCQfK3NX13VIFQpjsIzYWnhY/vN7rGKn
NFoakNM5d7aFIhejec6gHrpOnOzR8PDeLPSf+wDoweN3kb48/zmWdgJCoq3IxLt7
G4R9pa5P6WP37f5p4U7olLANzD+dOY4iIc4c9R4XWghe51poKY5m+21gSqGmQwiw
L7RWPS0NoOFMS6qn5ozEE3jea/9mSyXYq0xyfLVUYZomkGhZSTAKSVvG0O+G7vos
vJUGIvoq5n/aUevoJT+FKdB8rjsozGsEHtTLJGDWngqswCHQxUN/6hctCvo+SW1G
U9sdLD6xQ1xXyqnPVcAA41oQHYE6B+L7oVw2dn7dUsycbNSMfyfDqQOAADJudE2u
SvS2F7LmxTzvIqRULCPjhNYKT4RFuUzQgQjLwLFPZI4vyHgkx8OxkvlVphH60CBW
OKxaxARC924uwSIYf5r8gEKEgEEz/T/u+n5CQ5wG5q5T9D8jRaeM0FrkQ0cGHCDg
fMnASSEPqSywEX72WZJ1cRkkHU/aj67cNjUu9P6eJ/XP1GyXxiUSOZ1m/TK1wDQI
vpJTdDzyFaJGS2jyQ217BUSL9uYDbx217GrKlkgmgA87eMJP5pdMTOhaSFj4dSxX
IHiNVcBX5zs3NLb+ElyOiUTwNonC608VF0n43/xKmSY4990VhBWnaFDLDnVadxHy
RiIe2usxRoY4Y1APJBdoq38iY9SJIZxlTQ/k13cyWdVfdj1qvpAOScJzbHZW6dfh
wbIQ6MzsajZdRYukdzLPRWKoRpxTdaBeHZKA6NQT54usQ2MWN7z04KZj0sPAbuQu
/M/udOq9UB4rD3JAy1uwH9VDfwxDmYIUToEgrhB7RRqH2ytEQcsFUxdLlC1OXm1z
kKSPyrrntdy+1OeV+B5dHcn1nGb0YznsfQPhNmcFTGfPcurTscgRJWt/tHKgPS8Q
iCD7k3K3jtz0vdTo0bdn1W96+Mp+DX5aAEiFqKommCRaSQ4lXQDpxzYe4EbKcWk8
C/zxBUL+P2QkV5ggi92c+qaccB5zYVv70eGZ9sP3EG/T7VylorB2fBnK3/st/m4r
0g3YdoOq2SyYi3RhqOUGVz8+jIUlgqodm4pdEgz8r0zT/Xjx2oTj3okKqWPau2Ar
2a7LJqxzOF1U6QKyeYCpS56QMRfHp75G//9TkEioqCJvEllmP50USEJ43vTk2ZZA
Xn+igy0UV1w2TXIjs4U4jUWyE/z0pdhHQRqcPHVm4JzNe0ck1g9DrD5+JgvRy3nl
fxKlPXzG0y+wqOFlD+jWJEqB7GIWqnlteIkuADgA59BxUy2N1qnMDGBnoWEwfXjG
2Fz1rS8VP7Iv9JU7t4GuZwRhcizIFht89c6zi2weFD83EuR52V8R++wAoeuE/IRM
Q0XApGx/Kgfeiv6djKHIAqdQCx24aZJVQESBE1UsrfYBubzWzP9zphoX9iZITVbw
mcrTKdWYEuqYsYNxiBDo/SP6KtCWaxjz9uJAwhtG0AoaJyF1wvafBpCXGHNOtnKX
dI601sSIcM6uk6JhZNSSEhQ4YZLgNMTiFxbWp7M5h7BqE/IXFZBXwlzr384mH/iT
YRgAY9zv8C8jSGFkBZZFdCRHnuMYOwhS7CCVLIEqjpgQ3owqttBwdq8ZoW0favYI
v9x4OS/zQ/mUJSiF5rDtC+N3PvG2v3gFfey6EE4Ocx4M5rt3PykVZb1wgXZUEil3
/XTWSJ0Ki+9iB8/zaVOzxsXfauevU24sV9FQlN3e72lsPptCu0nciu0d1kA8+ftg
Inl5/LyPMBCkfDtT4XOwSR5PBuocahJ4CIuFhSNQaQoAAcMvFwpauLUelrU4fivv
CVWNCCtKPyZaZAD7LpDrM2Ws+nB/B3q4EVtNLqNL93IMyH81wYaCMi+MOlKhMT4r
R41s2uhRi9x0JUIt/0wgJJe1dHUomDGvfjK+BpxVNBoqsGFYQ7RJJqBC3gZUUBv7
2CQOugfompfJuKaLfLZ/nlB4zUV3Z60A35tn9t2sb1gbCy4iKcI5ff+/sz3V6mxS
uD3N8yBtcqu40yAaiZiNzRorzwglEOg33PHlWZTHHtEAyznT7eqPQM2Ohoavi0z1
IgM2J4T+M+Ubiv/X2YEwMpAwA03FrmoEnQ8UcaPRVoQOVaRylKbSUcLDJF8cGJHC
WV5GpE8QfzFjiXLqsS5UaevzUfP0st79SBPp3tQ4Q7sdAnt9DqNiFd11JTd8Dxpv
9HuSwCXiZlZaQ72juzc9SKeA1CjtWkE/WOs7DelgGfPHVdw4/0qmbKX4/3U0fEW2
TzGPFBGrk55Lh+Z2/MeYdfuhkC/qYPgHdv5/1E2LpDZZFMh0fxo/8W7xbUyhvqJ1
+UDL9xGCqgkxjLp/2bFri3C/XAVwPaJwi3fHoQNrns/6P9GpagdpiltkgdxO6PRM
YbZvarOu8WmexV3UQV/J4k8z39XYB3xNVFGW6wAFtiwWj1FEEX6CEXhOo5wxBaJG
KvvSQzjSHVy0vYvVJNCQHnUD1d5SEZLeHqZEFGVJNcSFOSbANE7RT/+D3k4P/jm3
Cl69sb6Kijc0JS7MvYlt2gp+yoMRj+L9gBMG1tLTqxhELSJmFgKr/aWDXHYYzhp/
6dD74y7p79OAMvelfgvGMYZezYTMm36u0CekTv/eSAhnX8b/4uIyZz/zzX1lvPs2
OdxUpYAqVjknG8Ak59IOL4jkB3zc918DXpX1Mf8IKL3KutN0wOEdSGeDZnXs/Vme
0YRsthGq5dQN6MOQCIknyMmgCT598lGXx1GW3ThcOJG3vlLdhyXqp4/ccC8AYn1e
azAQL8JWJcyfLQDOKa35Cn0SyYJHh8I7V2nPSewOwSPs9kNJsOE4O+3WMv0ThtmY
Apz9vcfm7gpmVYps3VZOy05orIXfIH9Whr29EMRVKcp+8CsTdZbWoDKxjgPuymEQ
7PGEeEswEjj96kOVzByRTXHyP3Td/FGcr6CXs6IEe6t39w7tpwp3aT0GE2E/Fd29
vC3k7zR8YKrbqUPeDNNouLhSAEmj8/F1M+A5V488bUHHYYu1ltt/QxsC701bZRTk
UN/3xsQtPrAxaaL7/LEfNdQVT4BnQRmAoTqFUzb8a21SeaqpuLEapG4I1CeSE+cb
JUvpNxfPsoAb7dRujUwb5R5AITGTKzRJe/zbp7YfmPZirKrRbUpGa5ti5RxxKAqM
/YtvWJRpx3/LNzH2JnJvpYA8kRuREpObuBwBDRB7ex08hfL+Ii0+TOORXwcSYahQ
yNHsDFK8YmzHGVIwAp3rVomk5/7PAIlrN9TCDf9s7IGzB6qttCsmwcGQffBorv8f
soOGzoNleqyI96t6Uj5r5uyMX60EMe05m0aESEpVIZeqSNhn3x4Iosky23vFGWj/
0Y9UgJ33yeEr9cYwZmzfwOCdCB7TzMk0SxN8LqloFuZSBr+CYyyelhzuT47UI183
TIRyowFRnjLk2xQ7br2wM6pB956eL1bhRUqNxK+xosC7SGws/JjUQrfhsg99YMhA
17fm9KzN7arPiWi0ayN8YyBgWkeE2IKXWJ8LNPORLS6Cr3eQJi805xCkQb14bMjq
GYUvwqp+Mioe0QKLwVuIeVVo03mPf0p9dXhLH5a/dPUoUxs6EM7sS/ui+2gTtkIn
4hm8uZmOPVmVHKIp3AD5KKnNGQ3gNT3Ew/Mgj+yBz3FYR0fZXgmHhTesgmpGScu5
nT9ivqyalQXWGk5RHCAgHZb0jI7zJndsGtTSEPjbFVPktSGBMp/E/pW0TQYst4Pp
SVbVO4mEKek9yOGFdkrKwHpVKYyxqT1pXZ+sTmrCrbucD3xlwpStE+X0tmNrrfCn
e45EeRk/2JiZiteeJ0gnZiU9pg/PiL6qFFdmtxSnNoQ0tpyhUGbgXewJClpSizYs
PYp8r8UL61IPNQR2Pk5Zd3JbxxZoB1qGLjW4eUwkYn9UuknWzdxKJoZ9Ovi4Xvoj
0TWn1X1abAif96Ujp1NQjKos355HgrN++qbo9bJVdcZ1HyQJDjqz0WZpOtsGKTyB
EODV5S4/2RHHTJPlXF3428Eth+ZIixL6MD/e3/nCujkXqG2+La49PV9Wz8NlmqdY
JZURShMqxiJjkdJK4/ZC7PUk4xWJcKpIWomdBmpdvEG8KIUMm/X+jCW+P2GvpPGY
j9i3pHIYdYgAsIBqx1GEW5+g5Ngs5TBUJ1fJLi2Q9rZkOtaycYhJo3ZWq7CgWXZF
SoM4B0DhNzgyQizkrVwAGGkaxOSZyv39C101/T4x67lO7ZCQdNbQR7L32yX37Jmn
lhHJ8xo+88EX2NsKFvWhu1TUOUgcj/oKSn5QMcXHhzrXSgKmBfjeHUD3uHJ8IxSS
wfEvCd7vmeVIZmPgIQRuTxqt9TzTfuC7VKv9RebmS7s1JjbmmqCuNlJY1EHft2+9
+1qhYqCbnnS/422tYl9yftE+dxBDEb1+g3JRDhgAMXX9/kAZOSSUihRnWPAWi+li
YP5tYI8k23cWcYKGm4rPmCCSVgke2sdhpRFKa27Ns7FdpAO86hndd2viPYRcwkk6
eds1XDpYvRma2W8dpxz1FLFSjAfOG37q0RraTv3WAyeRoa9gKnNDV4dT7ur37e/c
n/erVqJYBNt5cT0C02pKipkXse31mRtdGY244KZMzQS+tgdAT498gubjtM7CXxJH
O+ZXmcRHOzc36vHJACk48A37MA4rlJf5/sYNS6o5APXE3KEo8f8PCfaPvd1xDvdQ
ONdYKN5NMUu6LHpAtMl/0SU5qQNX1KIT2ASnDg14KURq48wmzA4bsazCcjYsV+qP
XXoegCrOZaxoFKKK0xy+X2Pw/vu6pMVAg+Tsqvz+MovHwlMcUfVCozMYpsEyBwos
guee9Dhg9qqj6vAM4xozsYgKPJLv0T/5yHa4B51J5x6AO3eqyC/TeH3+fcCUYARc
rpfQizRZc4ySgQKzGPkcLPNQnSWWKwU6dqWhzARdpC4bRC5LeDf1DPDJ7krEdhK/
AWunH11kHrYWejQIcTxJ7WXxTHx7nAx4oiXIkg+N4xkR3NPE2IoLQZpsEMz98d13
NcHAkzlUHMQrmZQeZ0LAR6sWSmmPFpWcLCV30J64DykeQP3IziJ/wJZDbpYl31jE
G3CkFYnCXOBXFoCLtMWKmRgnGE6/ONnk3iNv7zwSzfOdOmTO8/ITiHTvqXALmIw+
o0qB8Tn4ydyyMWoUDw4SZy4geKsIhFxPj6LcTHbHt5E9eOXV9pT6NaNxQmADYq8R
NrWEI7rr8QEvrycnytd5AbqeQKI1+6eploZYu3vqqZPzZWrwNwZ0sYbDq7vyOF0D
NHMRvsKEwp57YzyinG9q4efiyr12w64xcNmsCDhsOPrxB+eEDEcKrIRbiBoBsKH1
Td8Ip6nPUYqlvCH1VfhP5jaZAbM6GqXs26VOHpnHdQ6CIiC7Z5AQgyIBfzLcODsE
vapIO6dWSMDQK915ihzx/P4gKHANKEL2ngZuMZGmr7x+OujqvoSa/wKBXIvELkb8
vWIjuhIlRi9sxuVwVLmEhq9k05yYG5JzneRZoRZ2EdUDo1JGEOCb5IvpPAle2ECf
QaiEHhkk98O67k7iWB9C54njTrc4SJT/xrfSYyu0kAwvK4N5JDMlDq7QR76zvB+o
b84l3GNUZShJ+std1ZWwyYzRjQijxCsJxHPB2GUrUwDfuk0ZqozNLbcTy9t5vZr4
+7UTJkqb9XuNB/vm91xoSAJRrAK/1991GhrRqmHZl0364vw+U6umcRnBTl7GvvH1
lCHKJ4QFnkLER7nlq0Xif6bAKZHOQHroxZIjyeUXBBUztYtLSoAVXPbuIC504ars
J9chne+Rie6lx65ZtWF8G0TSx2LaxNGo+F/fMzld5O3RReAbZDmZOIvKegvt4YCm
EZW+D2j+VdV4IKLk33MqNAFPXv8ay6XI1Wb+47RmQnDyBM2ZZz3Iq0v4exM1/Cji
4DUOtARDcXFaRQsD4BMtWukc6JbbccOVsBnp+g1GJc8PsgDPUw2QdjhOzSP2363l
9aBQqGoNRFzzuOiyC/HijfJ6gbYlJZzyyExqKgkHBn1yH1CRPUWnSI1cPqk9r//b
9E7ODvwZWBaWY+kogIKJAfer50jzMCHePQc8DcJeQ77eNvUHAbnPQgxROvHsZ63F
sr1WlUUDOhFDbc4lZGZg2xVFajndaWnwAUFGeH64OTnLhXOL6rKaVlsNyiSDw1+r
dEJ3EBRaH0v9BJq3Tkjz0PYpzOddQimvWPf+cbY8aLZSBHxo6ljOweNH3fmLn2nC
3Gm7IxNktX452BE/zfwGb9/JoAkVxU3d3Hzm71WGbKlgM3VOcuUT10zr1Lajizey
8623qeipXAPANNPAW+RpmpF1OnewRgaZGdGlcVIdMH+pkfCk0PgQqiGKnxPrn9ui
F+9n/mMI/WMpB8GrZDJS+owMOau1q+IXxRGQ0n2L9GEy/vfqGtFx+VaMfmyc2mJm
30gLKMJRjmmKQeFAjXQqw2NYi3g3oKWweRYP4edeBVfPwuxLrLhhUZSuZjkz70ot
bC8OVFNnUEvdqoOMM1W7p4vtxWIPh9RN9QIBjVAXW6Lq5yc0s9RzmKbueWHKHujo
O7+YgGRHlnyzRDiBF0HnE2X7wiaIES7tsERXiEnlgDhuyCfBhbb4cpKGaCajC2Ix
fgdxBDWYIRjjBpccHrcTkosxr25eqAwkaUpp7LRjxz0E5+DPehPd+P+DO7ri0j/w
4i1mS7yMf5thmn3YKozOli/XOsvp9v6MGcWTAbxjL7k1ZFkWtVEAOSu1NTWPolnS
Ze8wtME98mrc0YBzEZbKm9jG5W2d2oBvTHj4EJ7XCQy0ednZXu2grxkfi/ZRnEdV
jrdogAoncyg+IXQ+aoJaLoDJyAlYErpyt8xkM22W9cQmpyAppNCAnH/8eceUa8/8
43s3DSjeZeimYdhpwg5Mi/tgQJclwO1IE0RX0IZTMrCcsH2d2bF+sz7f87umvGXR
Cp3TRsWmbB9m865nVxA7fjwcgaUkwUPVSyv9LbGKQ6Vlb0+9Q7fDE/iAk4Itw4w7
jpzY3niEYvyb4YJQco0YscI7LsolozDYVgBO18cYaM+XiGHVt1igFAL6Y1+ZG7eG
d9GpMWuTj5fE0Mu5BxUwy1me/AiV5YHnOP2hMJWnpCn9okeJhC5CN6ypVjjLUPVn
OfFpP+vEm7MAv78aA+UYA3XbRGwoecTIMisYIg8wfrMlAZgriGYcDzBV25Gco+xT
tVOhixb9q3/2R/zzEAkVjrbaqbTaLkkoj8BChDMjaLacoTRFgWsafdv9GY+euwrz
gowUiezfBdBwQ1hD5vkJfZYbHXw7MyithBdXrAP3ugtB4S2DL5RXVDfqSjXgdEUW
6LYmSSLu+5wt/5R7P6cX/JUDZMqcJe3N3UYULxIvXJIad7f/xLGfZS+pwy0QYb1v
ycTATK88czjpv9bQsfG7/jBj4LoMWqeN2eIZd/pnhxo5MRxoaEg8q0iWl2gICv42
H5RJWXolmmYiW0UUk36wcho+rjJWa900YZcOKZvKKpFhs879Qtm/Zrlf1B5qcUa6
EUZR7ZAj7NVk7T0afKHHSFT+WQkD1VPaEM8nIl8fvcms56p4UXNL48yvn9L/yl9x
Y3+URYVIRwxlM9vxmrh8N+AzS8RzK2BpxAbQdQ7CztlWO86hJEYosK4g56mkcGjF
HvxQImkCQMSykDP+viL1WEAPYJ3zSNIXUJgjYp8+isajmDZIPeSw2FFMx8ARWd7v
b35J82bJclCFhGb4Dma1PGaHGZFT5iPMCNjKbQZYfSacWDJPCKm5GA7ejot6MPgC
mhWIljhy39/DGRQ/pZXfO+X3AmHKhLQ2c19LbKM677cCveQfwItuXWK9ieIYK2rT
tVaVM/uejsTX54FC5jY6jC62WY+4MRsso5OlOkTgs8jSiO0+mznK/Kai0V5h155p
xgnjRCA+mx30fYAKV7qVZS3VJdUUQDRL1bWESVKUBYVPSjBTd6BmTeZyByzi7rmx
s9bOc6/yhGh4DBhrFmjQcmZKu3taLrsajgSwVIQvBBQKutdkhxMUFmGsLJy6IxGV
U6DY7DHpO6fOijSvfI04uUDf9+vwD+iu3nhxNOei9L25ZAfB0Jj9HiefPT3jp6+j
EF5dZPfXoqJ3OtuSj4G3omAafzmupl5gMwM4fM8o3j+QP0dEbkF+8O8ExTCgK8kr
fBpEbpqlx6JErjvs6ZrBslYnpMLDKRNWc1m9HwKQVmSSoE7PebegOAhzsfxy6fwT
pcqwF5+0TiPI5eBNTrjzKKZzuq0HXjOBFMCcrn6O92CQ/l7O5W1X039EswzFQfEM
p7hDpmBKyjLFeYuQrxfA15AGMPNeWwyFlDMYs7/l5Dvyh1Z7HZMVJhHzmQUg79G5
cfCElgdb9JXi6vDEHL1FO/Tpvrdi6+rXJZRbaxbhMUOksjRO98xOTIkgpSxOuQv0
Dx2xM8AxDYP2BG5oDulH49eXz5t0Te5Z/zzjc6cB6qye3qLjWY6qw/pQ1hYnInF3
9/Mh1AK3okumsU9U9asaySY/foq7avM+sYuzYgj/VqNxpuI+SEVshA67UATQuiPC
GOVVGlQr0lMKud4uqnDInpDeM/YQr97CqccQQdchUOfAFMbYtRMrEWCPDx0k9ERw
wYnpxoouPhjPa/9lXWc20UOoFgtaccuUqSWDBgJO3K7B13mUTh9C8tpX0ifKaQWc
CIpPdKmjtRX0AqkC9FPv0eHHTL72I0ZJKRbLeFgRjRl6ENrHAHulJXBoUG62OwRW
V1XLohyQelaETNPOgWI+0/JgnLyN6uEDVzu/UE9LFebYYPtoK7trVrXKNM7BtEml
jg28ozSBDBbSVUlAz6PsrHVqAkPIfIivGtXttwS5c6pX95SSB0WJHALLhtDW4Lct
xUlv127eTV5zrGy/id10ucUh6FzgC+N8z2nQDTItFW1N+p3a7b4jnsz0a6icdZNS
hua/YNwUJQI0ViWGV+PNQ56Rx0Onga7v39z5o0gU67/gN+ukeVM+bmgfCHpiiQKe
+YEUqtSe1pyfhej6Q2ADmAftI9hD4a8lo3HW1gVRg1Ahxv89Y6tNFuVjwTM6uG6A
Gu2fFw5VP+gPoVyfj6R9Lbow3uQWqhSsovqgcAGVoZ5qD72QnPQS+bFCob1c2WYU
xv0/CXUxrF0cIq580RCVDGOW83P7KyHtMIea/8CC6x2ffDyh7v7yKsqhU8ElEXFz
sFMx3ewniQ6gZUE9TERRsmLsdkgB40bi5JiVDHsR96EcZRbU8tUmI3dBKLu87Yfr
LnhJq8g+Sa350BGmy8CmXqGc26TxYcmzMsEidyRcX9YaCzJP+BXj9RpE12kz5yAU
FJMN9fomkgZ5iuq5rhMfWMal8QYsnf66F9SdQuq5V5gfgwuLdhCp4ZYpLQlHleqw
1OitKQuEOnrJ0Ip6uoRmVPmw/NOgqCJNknmQhCccEHWwn1l+ZHtUEau9Nforp4yd
HT2LvWOuxTYkdFdPhKY5RWtYJqxN0mxNxvC7GgMjcNxjQuXT/f610Eps8wRMfAjS
7iT7Fo8U0auqlpFCap05TZ339//eyinQ8kPMgY+3fHJQ2N0lqNXwGTiJBts5UZnV
Q9hT9QJtDU/htgiNNB0pQU2DQ2uxxbfavt0KliyogvXZ+4dK6/PRObTrt3hUaFe8
6b5Jj0a63a1pwvpx/YYfzAjf95F0ITDuLUnmPWt1RulqU354iQ4q1nkiDV8JykiR
73YrTcPV93pEw99tVpRh+rjqBN1AZb8FPpt1RJRsfCb1Wmy2ERnC42WiP8R7gcwv
Qgq3dvENLP0ioo2uB/6hZrvbNnl1QACzG7bucd+LonX19DmuqTqi3en+GeUFKYTI
UTPi+59ZQBvS3C+D8EQ84pgjDmfslROa+KE64whkWOJVcgm5Y8TIxpsOFe82Xcxb
PVGO9tTAWlPmDmT4NHyIEm4RX6OzgcTTRohVUcXQuP6m1flQwyvqWAV5L2/lCF1k
S9ntfDxxwMdq/ZtZ+p+o3XGbQFGl4hBowmdoIIXxZItvbDywILXBf4qVEYIo0fvk
5fh+4wKiJ7RuBBiQZw0SuWvuxfUhZNAC3lR9yV4zZ8h63AsUbAovtYXkZdMcz3NX
Hv2HY1xYzNj3NQdAg5ynHh1LdgRrp1v21rb2XtDcNbEcfTKPOeLE3WhjsLTXqKjn
vv3CRtshxRwHJldgoBRpquBcFgUdORbp3ROcxkNfC3+i4/wkqcs9590Li7zBo5l/
daGdMrtyGq7fE11Tnpxy3Xprjk3qJ3JLel/2IZ1DmOljWBg2cLsaRvho7tW1Hj2T
VMwGtaDMQOh7vmh3BcsLw1vMNQ4dVETpIPPtpfQXLkil2c6rFnmPvZRvq79NUNqw
CdBGZg/h1itmsR7Vac5dNRLgqNKkXkrbgKruOFBv1mJsKUhcrVzr1abLYc+YlIxD
jJAcXQmk7JSpQPGlSPOjtKIZ7xLcr4snfKngdwZz9xnBIkMtfHzGqwSbygO/DNVl
XSZC92vCxMSK/QPSlJnw97rUuOeE/hZPRLhdcF4OaI6GTvXcn/Ytzfe15HiuYsKo
GYM7GxX2G1ii9PXu11Y0OXs5H5b+YYNsTxc3VJsMsbMZLySbY1FMx992QsI86JTu
3iVI4eSk/mJhuSKcllS+hOwHFx8AKTPMvuY4BJP5zaSZjwJ2nTKvwlNU3AG/Zvid
qHUyQXbGqeB7hItiaStPimsXN06ZGwevCniRWq4tQp0Xq2UJsdLZCHFNseU3jv7P
J7kyKh135bXut+fR4pYH4JmnDiXiBxYNOe9FatqnFUL5qog/wJSg5vea/ICu4srZ
ZuKtJlVyv1xiNdmF1eM9ALlfGE/Nz1ONza8Mn+2Mu8MUzpPJCuVj9aecnmcu8sGz
5KIeLL9mwa3lmDhr3MIjrypEEWlMCF42btMa9e8iQUlddt/U4OH9Jx+rrZ/uy9T/
y9kSvkrLLt/NGQcDsyWWyCHcJDdChK1ZlYWJlNBFE6Jg2fdz/KZB3q8zm0QGywuE
xdq+EwCz2NhRzPiDbMtenR6L+NAzfHeJgew2ua3e8/exeB31FL363FX7AqNEW/Tj
mjOcE2qzvUECVN6PePNy4KCOpOJNRyfaeEhkK/+pmGfVo9umMU8wO6DJPz/pFcy2
qB8EE88I9otAa4iexFS9O1mEo2Ox7f57G8GCZonRZNTIircG5konhGPJEqkqh/GK
rSpaBi9kHke5xu3ArodHrfxJEKnye4J1T7DUXB7GafYSt/St1TmI1W6IuwJMI7cp
64+IeurkYmmV6E8m7fU4MGD5uyq7RvNnYswsvWg6I5Yaao4ASiKUo3Joz046m6Rx
F4s5qFCx3cFrsf5UKL/Edou+1tG+mcuCEV3uhIQ1ZfsS4kLcczQ5uf8YqkOENhoX
laSzV2mP59M3UZmva/Ceqd+GtSyqulc1tnvIdeUJ5duooUoiE8ar5kEc2bSNT4sH
ymgwmSKyVEEmhIYXrBzEAjqUA4BoE95SHcbiqb3Gz5/h6QZtL3OXETGLifLZDFWj
06IHr/Y4K/LnYHhOv5wYRWFO384S9VCRbe7x7YYstcJPdM+RVS6w3EA+7kc6GxRj
Tay8sNwdThx6rnFQZs4lp/R0S35t6Epl80DpzFlePVIPqBPDxVFLBrv/LKXlNSa1
3JojHbHiNmh8d8x+n55DKsV8baMRVm1obExbNxHrWSmsd/Y5BNjGlIRhnuEEwTkN
s/fxTgRUnEt76EmR5ZxFPhCPZLC3dflQ0pfo43N0FIPuEOgefNmqZf3GzpmouiUS
q3valYgVVa81jbGrIus5O3R1qCElCcf4ar/WsR6+fx65KTRgmsx5p46t8UIbQYAN
uTokG/nDiNUy0eP2YkOZNCvs5bGK37jYhKIRGkWDpLxuxKtVkND/a25CJS3B1LRO
ifZcpiZn/Yy0CnmPJdU35QJrdcN+TzuiMz2UdzPelXsl3/KzmUU+YeC0IojaYBuR
G3IV6xJXvf8O5KcaxqBFE6vS0FcaiptMAaRuwv8JFFJ1T78cau7zIkse8zlUqRKy
cQaLV+2leBs2h1i6FJxgZTN63US/SRsBXEeFWYAbSNc4x/0jJP+4Ou2Gw4RvzdQf
tAYcsdHYswzifQTc2aeLDfiLl5GDYOi27u6K2EvgBO9kvh71pYxTehyue2MujFE/
XVlvHZk93IKRE3LuxINUaYMdHDImBxngxCBmMJzQAM7x+32ChXiQxz5WQ3cJeaFz
g8r2IZntnAGmFRBuLDTirbvYrSqVoPYPJJ/2/zJutAYIfXLWEwDAXOoYD4yFzDOk
xCm2O+nL/mr4LssCxVlkyar7yThAekQZE7GOZfsKAfIlpNbMdtqGXw6xYuNITL4C
IMlbrc1z70YHrKYSaUwJ8wxWfP71a0Ae7/pHqmZI8HRulsxeXfOnRF/h6JfPtL9c
BNSWUshaIg2d1ilKvfg3UDGha9KxVachYyQPcXXstCUPm6TiD49btUrJrKmMJ6N6
FrFJyu7V5NIwxDC006E2Od/dINR4rtkzZ6G7fBXiUu1qrse2p1mXbTkumOP5xmGq
tuBSGFfJU9I0JM422chIdYU7HYur366cPkD0KndCXIu23Tab1HN9S3dC6jkQNNkH
DBx0tSbUOYNdIh+iYtFKAh1IXpnzFVojY3KXRNeOiELb/GBel8pE75M2pP8gmVA8
l6NWW00YhVlVI6bgODleoM9tE3cCLzoOq624+IvTl4AUybK7/e41jpd/p9PQgjwh
IaNuCUSYdYlU5+bap481dOJYkJZpOXwI5JtORdXdcNwHiUjf62h0pEnTga1YfcO1
elkzQPDCK2LlYGQHVDE3RnUn8vQyTF9cvEOGjQId45GepqpZ9vA4GBs+C9TKzNeF
qcw2Qg6i/cLZrL8mCANo0P0y/AWyREykysLidhqN6gTsfciuj7n6o+nJSbSjasBm
WcO2hJApVCxuehBMLRp0+tQeY2EtMM600lX93prGJ0A/eGqFpOheXJbwQgUgdXGN
C1joEsN2Jnli37d5Stsd0Iu0HUO20ptm0EX5qZF7kuwJhnVpRS9o5lmk8WJr+nZ/
STM5X2+ljOluUoVRmoFA4Fxpq8eQ5gqpd/SniM3Qgqz55ij6z0wbNw7oX/Oijn0D
pOqd6/0X59JRf8ri+Jf8dv15NGvoNLhdeb/xBZWmcTlhNfEQDRl3/0N0HZPFfiFT
LrqWWazpvTyeMXr6dMKJvls8dMcFIIZf9MhJHAEyZxNWbdGA0730jAE9Bjsqc+7g
jqOJBzXt8H8gZTEswMRd5DyrjqrK5wt5/OWQbpr5euUkJ6rgaFiD8Bs15jRA4du0
tq9HylHf5MbiO6WJMjcC5oUB4Nc0KMcXwyci6g4DHlR1RrUJnoZsPk6LdSbY0oYJ
MKJgocGblHZVBy0FSC/yfd7+ZJ0l0PewU8B8fj4eKmTGykIX0CD0DrV1elrknreg
Q+5dutrkherPhQnitZZhKEl29HY+PFIhVLkXtQDhliZGqTVhLmwfyeNpL484AXP/
7Xe8Yv2zc+pcoFOHjFFtXksq1HHDKrFi4ELiOSidFLqfxzC1/ktP5i/mZuyLr2rG
hl7g2o938UbcTtvxNieUEZm+bidilt6ENqfwcYUwzSkrcnrfkZ/b8AXIyr7WDqZz
t1gCQZ0XED/VP6dxgeLqc45lnpR4avQUXbAToM8Wp7pJqQvdwV3wijMrQQPYvU6S
HqhgXXeTUbf536SrByS+OYVOH5VqJ2Acag7tDbJdxPhiyteU/7Ega1VXW61w0O1b
jRKHfrMaVsTOfyXkflwLxeZBdULSopKzEY7mWCq3riXzRl8wC76nacId7gAqCEpu
ysLLGdH/P7+EaibsxlZNYfc0FoF+ezkX6oBRoHGWaLyvykuccfMNcy+ijl3PgJjF
L2lea0PPPs2QnTwH4LxKbJxwlJWE4eJB+JB9SQzFaozJ1mhutn9Qb1mrGeQAGr8t
nKyxVqtdeuEsbK4yWd2MyTvT5UyYvu3itJwLacYp0eHb99CUR4eM9WGYTWprq6zi
1Qh9h6BMheYZC+bgzzdyX4i8p9TAzV319BZHJVB+OH5nCN3I2IikcQKjhp4l4C5C
Eh7P6+4nIinbjwRApyhUkpu8tyYFU3kUMZZXbELidgQro6TZu6bNDKOS9JrBuOEY
ktZmVkrtqS4VUVFdHB3QMA7caOo2FVThnDUhvytqD+s+1Tfsnp/Tt8iYZ2lYJHW9
6Y/2ZmOOc+jHhKgPAbC1xXQ3yFxREE04cOFwYRLYySWy0V7qu/69f4ZTDcw1aSDq
5dB6Z6kUVjUwdDvwp0zEgm8sQHPxRnlETgWiin0/rhDRglBzTVUa3uINuFXYeY/v
axbiImP/wtrJ8+lxyYeZxVFdpO8EuYfLnBqzIKsQvWpfWixnqYBpkN7k3xHidrZi
SP1946J962Q/DcvjXNvrj6fWhFHJjWPXxMRzYBnmcQfmoILH12VIG5nJSr9dO+eD
ce9uX4jFqvtj66K24Li1VUaDmNC922xBFQBpZbpI0B18L7Nesn4++iIHW46sktxQ
20oEh4+js2gHUax82jKcPcqjQNDUXzDJOYdC4XJ9pIyXKZqz3kXC2y6oy9x8esud
lACTW8ZVH4Cs14jlJtjfove5z+BGpFbWdbd8HEVI5QKftFbcpOlpbBRn5IIKxVlK
GeyfWrZiB+/f7P32pmvj2Bh54d4BAqjnYk4zEa34rr/A4EubliLx4w4PE1VN9Oiq
8ktjaMNkrrsEVvkaQ4ZI7PzGj+IomC/fNAPgzGsyNlrn+wuyGsVzv9M3y5CZlcIL
CobP34qb6Lii7ryCTYZt2ZnDFMrdfL4O6u+xxp3/Y3A=
`protect END_PROTECTED