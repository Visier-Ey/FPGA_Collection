-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "N-2017.12-SP2-4 -- Oct 23, 2018"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
ckttgoNfNnt3MQ082Bap9Z2Asf8o2xvYz7IXQ08rWKqgYEkRbbvIoETtZXmMZE7e
qZ8BFjDHQ1nuSQu616Mg+8s3A8KdnkXprH68UdwgqXYkQtsAhPXj2c9MN2Y+DuGk
hODCTXpvCxjKANJnvAelXkAGNilD0TwjOPdY/naD8fE=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 44000)
`protect data_block
o/wO1eqZo6V1HTRn2aCuePCW4e6iP730BsyJ8HigKc+9mDCo6SXGKBtbvtbmxLoB
RkNjO1IIW0cHTyxfheNFKYz0Zp5qxz4+fEVZQW30MuS7F2Yc/8seuHA/6TcFOWLK
0h61XQjMZeC5jxzzA1FAAQ/8aHDSEQIfzk4RhhsYQ0b+Or4xFXKNGbI4fe8yuoEG
+ecyE3pMeRsVEOgRvaSecA9u2T+UUVMmK6OjnUA0d7B8zGW0Ela9Gc06BCwST5G9
rU/G5fh4HawhzFFp2vZpa4kJzgQY285htay5DnDPDXnTwFGprM7fv6dXZ1gIMs6w
Z8RFDVsJ7BcUlW/UJlFDabUDELy0CczYbzD7cHfOmWDD8DOhvoxQ6G07fCTMP3Rf
nTbDygGNhEBbxW4DuScXOI3AhVUzCDZOKNlJTahHzKIjfxJhFuN1zohvrB8wNZql
GOdn7cJumf0awfiL6SnYgVtkVL8pO4mRYukpG2leNno33lrPWyxvQ5iu9F/eRIX8
bmGpPDFuzJpuso1YlcCNhHq98JMNMfCuk0YISJccGJGk+yCazmTiH1PG/YwfKiei
ZrZCKuIkRmO8WLaampGEx6MAkXy3FOLzeFdv79vYwLBA3RFl79QzC153otxDdc2o
IXK662n1dEuMwGm1xKvtOAnG5ajIIXHrb+BAGIlLlOnWy7U+6iQOBQYUGzG9hrih
3L4igDDAbifrO7NLelkXUD2qC0wPpxfQeVKb7jQY0M2vL1UezhuyOEDEzudibzWV
y9Nin2igoH1+ePK1JFrjNKeyE5igD/HafRKgZe/1e6HKj6QSukGFd4dIpfQHA+/1
bv61BIl+93lEMMRI95VIZIjWLkJP2iP1qg9eAtv4Bt/c0q26hZ9mvH3XQ660rVcf
hWQHbL62zi1G//jQpJBRgyN9/Q0h+AeaXu8v3GwBTYPlqWTod9cZmMWjod1/sKAD
U0RMYBGFblr2W0Jynyjl7Z12GWmYzsq+sFHZ27h9F6Au0FwQdojKSQO4dCSkgd/d
Ap8/S0kPNko6id4C6RCxss2FFvH+pNDZt+7W6Q1gnxhOEHqu5RVGSUygEHvlfaBU
DMJgO9nw3S4Zxy1C1d9jypjcLt9f4VxX8jBoiMCVrGJdoNi1uRRJ7HJR15qu2BOx
S7WXvUEGg9SO1vTKmdZo3IgsOuA3apmW5eaQqBcJZsA2P9yHwpDE3uWqYMnBiwbP
WOuyKvDS6TeSPDvv0c0nvaAdIH15+XDoDiqeQAveA/SToaheNDwjnbPbiraOKy1V
pH9aBSHqumN/a++yuC2TnS3mF4ycG0XiVt9aquizxlCkhXm+C2eWNX6EFtyH2KU+
BuODyRDtUAHOfFpjWdaYWkikpiGMxDmyTyoC7jGfNr9rHf07UFZk7tyliNzDyQeF
deLparFMjuLP2YB1xULaVpFd2LU0DX0W5i/KaKNtViyb0aBri3xDfF8TpFHRT0Ul
k55qiaGpoVN2/RxB5BcbICuCFBYNfQV+J60Lo2gGZ4HCjmd6IFoKVSN9wqYKN/F7
ynnpK0iLPaQTx6GDyAkLlgJxaKo8QLwNpMLQCZWyeG/WkgrVbEBwqtz2kb9j3qXM
OJqWcUsrPBDLbqJncVtq3E+XQAiLgJ34/+Abs+RnR3kMPlo9j7aZ8wH+nf54E7it
rObWzBZm5jOnBFA3jreQ8oDWZ7ZoznZsgWD6NT2KpYY9zaFQmjFItkPJX+l1phUx
c9V3kmEqGeHAfl+Y6EKMZfPeQ7eFKZPs/Auth94sGY05bJJmYK05pVyi7++kSk9j
l9SYbSA52jTq/e5fyb+XDsCxGfN9BjkmwXK/eKIzC61AAxB+/o17SJ/QEDC0uk/D
fA8vaLC3O7GXBl7fxRwLd+39/J9FJRUyynaj9Y8xGxhsXlMkQKO5PoyMZyd8KMDe
fOCJlLcU6GbEgFPZZdouuRz3aM5aTTPyMrq6nT84U8BB06q6dteO8Bq2JPBbMoBG
swT+r5tkb9UutdpJZFKQwumHLoG631K7fX5Big5O/XGkj51wqZAqOeCm3MLOwteD
A13xH3ZXtnfWLb/qbHpjJm7E4YOxgBa5IqI7gQybFV7Nt2euG13SWfASCHbe61Mz
/n2omeRucbg9XX3QD1LBV5BhaDnCC890KHaWf7wKZcHE1nZZ72XAH/XyXLcPdJjI
iMkX0ONqJmp1hbKKfzpYsmIuOnkL/arFz4e3fxtM8Q+48tQLfWXmrsOeVPOXWnQT
/IceBBiyUPGWk0kkqMIbrXb19oDM6amqBe7P4Tpr7rnukZN3E5kt1K6rwgZp6nBs
vAXGXXupCNjrGIr2LBN0hTGoW9CBcrf7qv3gibJ4jEZWEem5Z7GoZpFsc4o2lDFO
DKvGdyXWXXnyJGBtORPMm+kkr4LdarJPgnLfuCvlcR8bDjiB9PVb6bHrq/p0jeEj
tjv5byqO3vrY+Ol5hkIXNHOXnR5dl8RXyDtcWYrcLans+ANLrBPI22pwU+IiBvTi
ksjKVCHJu6y9HZoi+6ksW8WtnKlCymk71yVNmqbyNDFzhoPyxgNNAI0xYmTyjiJa
+H7vNnCnDdzMsuAK2FRfkFEB8vqSYBqAXIZ5BZgEDcDocLBDwHz4YKIb7JLErt2p
LXI92di80CIfcpRQxFYLWyHSC/mxed2Xt86ujaqqyw9vESNI6kq1qQvt09BXdCWt
e8kVxTX8ewhJo8wxNg5HQknedrbFp4AlRK1xJcnyx331q49iPF2SqeF8Jw1RO4EO
ShLD6RWxAAwh0QWRsxnnE190B6tZIfikGwBGWLB4eyl4J7sdvfx9Zw7ZicpGwpeu
PdLBxcwbNg/Pf17ku6JPtGHvs9JHbCPK9rFxSxvBhtoZiAG95oqtM4HnJgzYFIwF
wKqKRWtY+vlxzp+wju5xiZJcWe8ckw+3Uz1XYh2vIrftYzv6OV/zCshmrlzkAm9y
c83tUt92JO/3K6n8XFpDcrAMiVIuF1r89skV+xKHAgQPV5fOjU+BzKhxZ7czGPk1
xOYzdGZe9KiAD2+diglTVj/bsoFKuHCJ18pukeSfO9DmrqxUmBJJbrYaE5O9UmCe
JnS/ThqKhPRezzXa47ryRKjUHrXvITNiD3FgH7KJjOW1NviPjRnmXTDJRIVcCzWh
TNUGmnSRo1wLEaEznc0d1Tb6+fiz02+01Us+jJ4e7E6bFwSq8q90Ri1LDshe6XwB
W7uGQPy9WYxeSSmWfk/7bMximAnwolIxOsBwH7mvA/AZECGPe4380V3UozQptVBN
QOUb+TDKqNgPAhCGV7Bf4eifB02OuOnS4DkeoPAYURV294eZGv/jQGIVW75CoVH+
yINgAwcWTC8DvqiahVS2xJs6O8KJ9n6LuAB89ZM6DJQ8KaQE4xT21kaBFB+s+add
qpKw2dAK/oaJbN2bmkKvRpk67zTtQdedARAUxUzJOuhE23spO1YE2h5dXFUclRwl
eHNi+WZTnnAh1f3WokcDErK9mu4Hin9calShadRXoJbLrMeImA95u26D1zIJ/00x
TMjgs3ucTGCMsH9ASpzAlE4rpyIRBciqCld9AdMvxbwWTilrXoHa3mSSChTY0EBW
TYsgLMdC3e/3zdLoFiuSTB11QJ5ZegY7QpGmpspeSzN5XQ49+RMTPnZYTgM/qnn9
VfUx8WKxFahqbNBocL863txkqAYQNT1J+28u328zhTo2U2/m/IvEX13E5Qh6o9zl
xywNsHVxUdGxiDnxVu/vFSD9Vel0J0aUvlRMmq/EpdsRZAVVape2+YKp6VMuD3FU
sjj01CIqMuEfadDP8pA1WroUzPfB+2kD/LHhAv+cEQQBpLhRsN9p4l+wdq80aA8Q
NMqX986OfnQe/iiLWybupH7QHgkbtfHKWPMeKTvgYt+6ntybWx3vQS75A4g/IUkO
fG1W2cJz2yWm1m11wNqdYDp6N/7+19R8HpOzMYn8kqububDlQeJq2mMdB2Hm2jsK
wykhqVLpmiMq5ckhupuJ6OMqq9dOWXxxKvQTlps4TkcetK203XZ6kiIF1QTw/RuC
olgnD/NVT0vNONed4YsHl+/AaQ3K5P4wuYoJZsW1ZOFIMFAURKA4eDQ9obcdD/3E
s8vDMT+6kvvk5GJEYC58BGK/1bBGznNrIvBoa6HieXGbIpchCt9SLfsvx7ZzgiWU
rs28gkhqOiYY2t0DwT8ZnC6ZsjajlG6vQPiBmi9fQSMiD6p9j3oR5+tO4iblsf2c
7T+5+efNPho0Uwj6E9VSCWFHHpZ+EsVYorETdVFS7p6tbsGaWt8Zk847orofJ7t7
rsRR1h1aiKXbtTFj0yKPCxkt4JsI4x9GWb0voiqPumUsELzs7z6pk1I/pDMxGFUu
XkPwONXumFZUGtqQ5QsYD7i+gQ0pCG7Aqyctwvr9hDIkksT0hLKIo23TwKC3OrHd
eSNu8XU5jsRYXQrk/hA0Xqte5ggfzzHKx6jhgnLEEVJWCyihFOXziU66sP3ueE3Y
EgUymfJAVrpGAmr0HFpr7teagnBxfOWS2XZk84s6ViQWmvr+15WZcakjzd8wqPhy
kYHJs34+IUXrLSoNsdpWQQWxj0c2++z2YQSL+c2iRt+q1NZZ/rL2ebzS0wRxgCC5
FWzyFa0MFPWRk82SQ/mzW+a0fFXAlN70Kr2BqVXEjDR7sJLfOtwnxlXYx92eOnzT
rDpIKBpPtF2fump3q7GvSBrl9vPjK2J7t0oJ0+bJo2v8DPFPy7CcM1mIAW9U+opi
Kip15aHtRuO1xTLFrtMVjUytQczQy3xgNfx4Rhgd8dtjGCH092av7HL4sy9icQNZ
9+OqTryRTBbmoR7XUtisoO1jsU/SwfCipmUTdnqBHpfvXHQYHvkpqKsZVCqw3GJJ
XXRRN2NC1UCwDLM/8GC0G2f4YtyTF3979gZfcbkYFYPyWv6dB6ckDsOrou1+cg+S
dXBtrQMbAgCF7bJTfGNKRl9VXVgWtajPa2MjSIQNULJ8qMVLviaNnlD/hNnxWffW
38wo5ck1CnvTiWHPE50m/JxypwGG1BXmliJ7BGFPupzAtxLAFl6F4fnZm47oJjLB
jvlRVTQyehbt+Nbf3V9zvHGw0t/CobZGsYe7cyX81c+Qyy1hzYpcX2edQI66YedS
NXd8lJdS344cxV55DaVPOXBDogr1comaJC0i+3JXCHJL1gZtL8up0WA5pv1Z/eH6
QQ1dLsMpODwUAmyx8kupwCmem2a9Aw2n0MPkpRls2l61zHmjGMuxXLhrZ/iqcjVx
7FnJCjqFWBakHIO6l46m5uYJwU+VBkYKfx0VjBL5MQJFNgpQpEIGi+z8fkCU+Fxv
YEhrDfV3sOH5HeP0ABuIxFYqgSzF18OL+hQrxJCZqLrKLwc2516uS28LiZH8bCzn
FleYJ07KIaqNOUqUEDEns9L3NrB+380VGIWUp0rD4yF+AKrWHYWpQi+YUjlgaEpD
ov2XMUuOnnbn1jMDzuz8sv/FKZDMevJFszeWuWU3Y8VcaI+z+4gDOoHmQdQnq0+H
sp9+PNATSAA6MsEso/AWms+OCLCJFrw78rcdOMzeEIA9wVJN9x6USljma/Z4XAYC
NqRfswO2SkgwEr7oI7OSTmOM7+NIoEun1ip2CaOyfSSD7JV6n9xmg8Cla3jWtQzD
tmJ/XkY0XpbiSK06GTCoFOeuq6kFqXWHy4ddQFzQwGvi5tnIat8v7ROL97e68yeE
nUt6SmSBOCcgUhE2O2szN6sEIzstm3oNrfIBDRweifQlvsAwbnBVp002T9v3snVr
QTuc1JMJnSGwgqqi50OAeZKI7hbeXt+EjVPfPZuAOeZaXzgKTbTBVlVd49sksbT1
92emdRlaaVCZAG0nF4Un2jfsIUp9mPSg4hqBetjU+Xhdj+rIFgvArguciIa66Kfx
V8UulevmiJ89CaCqsMbzNCe8gBJLwSLnSdzlk4emtAQ2+CuatCUCQdzNQFsGWbSf
XKNjz2upcj9FVwpjI/M6jrM0oKHeOpVYJZf5Zbarl9vG3hb/+DYcChRHwxq394o2
UitttjH1oO4iUf5ikXuwgErzMZdL4OaHv0jfUGFBL5YYD8bo8htAlNU8+m9Jlmrn
Rd3nKV4KGrKU9RGkmmOEPn6UX7vKjTOk3tcy3OA1uIeTJil+jmnlvGftbpbk5vBy
vPTVAI9qHZHlWOVpSHK8TACBBG4jTEpljneH956gGzO+A7txjH5tw+TswSEi+rPt
zaFZnWU9UGvXqcQ8sSKo0/8dTbpzdMzd7N28QQxNMCETryqE2+6U8ukUh1+6MxL+
Jn7J3wP2+Lp7n8FmZNGHj9/CZ+TmOEce6x3CUhhUmBQjdMGmyn8StjEWUGDQjWjM
fWXsggNTQms2Jqt1qybaaoR3MW37k2lDRDz33Io2ye+FrveRNZpnX3GapbAw4hmH
EOjPZZcVtIUc5za6/XGqA1y+2FSFg5tJB/1VIV4KQBsD0BeAvW3736ZwYo90VDtA
zdUh8BpgSK2jgiPLKDfTzt9cuw1x8oFMvEUf3nDrNjGG7KwZ51W3GeadMg1vx9Qq
BqBaG5FLh2ldsnIcz27wa07P/UpIxEJ7pZfAy2DlLlphA2Dq0CwYelR6pZtkxE8K
zXz+Rayj23TSzAg6Z66IF7s7UstXXnaTs5+vyo63+mMTUgfZJel+i8N4eLNVf7+n
EM0XT0p32MOmBk+V1r4bWnbCi00mht14FapqF6oaeR4xX371oRmYL4Zjxs3d2s+F
BN8w52/UW7s2og8OcfyjK4bpuFDeoveHWBourDzAiYkuuBL2vsMXHHd9sc5TRDxp
d4NDZoGsTi3pjR6jFs4j1eOPLk1wBRqo3cAAbwpTaZTMptl4/A+Sm8q/HdpOFDnO
cdnjoZh9VhGHSd5txP0wmzKkLBukrRnaZkE0De9lw5pMRxP5XReAqdB50sW5c8gX
POXIp6grBZfGq6iZNu5dx8GTiZMGqLSTadnWDKxVHRsnuN9XBJBLfMluU46zLQWZ
rZkbnFKXYJ0KLBCrbJoKpZVN4R8p8Is9Ag8AdBTUwZPmvKBbLatTJ4mkEbeLVwHp
17SOEM5LY33bGcL2ujZA2vXGuzNnjz6kt7QTu6wbYL+4O40H5s3fx2DTsXXsTSai
HGXhFCIjdry97oz7LhWQHhxPj8iKsIVG6hVX3ygyzWcOIl84cv4mgcjd/xtlGpnn
vUuQWP8BPNQtUKsddAiKKyZxEWqg4A+f/xNbOW5BlYBxSu7UHFt4VewmkApbTvEY
tO14G3u+IO5Xc4DpIJ+9nPPnyLfLYqOavwvL6lTQ46YyrQtXsBUiS2HHvoJG8Y9r
+i91kXJOO56OP+6JCJwV+2kZLODH5TL8IpvyydT4pROTMS9nCtSmTkVnZL8PHDER
0FtgqQomu4j/vYKDW47jVhPdcyeczB+Ee9UM/waUrfL2LgfP/I4PBJ2puwppxXtg
vO6oLE6+8wMsHQwR7eF5V+Mqi4hzX/c3vbS/V50MZalI8sn6UosOPYzn70WB0qir
raBPhCZeQgB3KNMsU77bRoxr6+ed2faPICCaecVZUrQCap4I09GbMxsA+OXtKFNV
tazwSr6ensCnyJQu7dgmRrcbmJdw0jA6vgs8T490mKpVUI/2a1lCAKar662pmEVP
jiIw5zMfE1/mQ/yBw7hHCUJAfvSayUmYHEsThRMLtxWs+8hW13KvfvcHtCbHcsky
wZE0wsQJ9T9qRfwIFtbfCE7I905mPwPPFqCSvRlU9eP9w7KcwMLyBmTVrF9ipGoS
6qjsNi+68Qj1NTiKaVvYeNGkHBNPF7y9lBJz6/8vBC0FJoow62ifuXLCPNm/n0IX
DAsg3dUXdGM7ohtCDEi3MvcRZAdXQ+gpxlgJEWjR3NA9OLsKTrByfqp9cDx3twNH
mQX07/XfvHbm8ZPwZ9MHISE3hosCYRuBN47M0W4G2r+56mS1AIHlazsbr6nv2+yQ
2v+Yw5G3Q2LwccQdMgSI+hTT9UH0orFP6ts02Y30s1j8sYzisSB/JRgcjrOxS1xO
put6heuJPc2dxvfMK4MDuiLslNs+ASMbHQXXgfKD4sfITdgN6Tr0rQSjtZE5IeCa
NhgJsMT3QQ1IUDVnkeV3nYhSLT5J6SFXAstr2xRAdiEYJV1WdUFXQbPhi4RRmIUv
i/RG+YuF2748LOryo0ezUGjYE8zFTOyhCKPmOYo3+BhJ+RGOpcbAXROPGAInOag/
FuQ5Vjz+bHpT3aoCLmme8ftGRk2/4qCFncF+fZW7hf0xC+Q6hVDssDhjyMytxCJl
M/DJUK8D+rQ589F42kbV5uBpMT1qIhPFFhWwLrFn5viAzeR8RvWjEQWwSRz78yVO
3mVgKnFbyQ0Ilfc3oZPBuMWkvj8gqykYLjy9NARd9oJceyP5TXmAA5yxDIdOMwgf
ZNOIKC5nvCVI2a8jyUrK9bcsTnhfa2fWUkhppZOyKJWR7Q+b1xhpupaboEGewFwJ
rtGRVaHmzeJB/lnzl2U0U9InWML0toL+4bzhoDsYpEOP3N9a/EHPk98N56Iv12qP
D1SCFqyfgZzCkTRbJpVNZ0N8KL3bovMSvLK2owfgsby2NWqERBjzEitZgPKq3wOV
sGiFz5Nd/lktqr6J7rZPSXXwqnG1sxAiZqBqTDf0JDF9HeukVQYdTRftj2pcjSQv
xWvVgNsxGj7OO9FHVydEOA6xmFtaxi+2LHtElmRyveCGNR4ybSm9QgpsMdHUN7rv
Qaan+gH2ZVcAhzkmwVGnHtjXQL+zLtxh1CdEA4pa1tDlZNG4ZXkUR6O7mRTjaVBk
Prdx2/pMnpOYlE876yJ5UIEMixgf+TVB/VeaV04VZeEoQSROWENgyKEJUapy4e2j
OyvnYK+YdoT5f+0gxFyL7lzFAbYzJlmHxOrQcvQglPWzxv6mznnoV1fcPAW5acV9
Vyz8+JH1uVE9HiXvhWaV9oLQEdDYhe7ugkvSfyr/b+KYUhl+SvjkOLByhc33EH4r
SiqlDjZYbxXsu+xiCffpg6HSQq/XM7Gb7OA3Vjs9UGMdc2Q8LQXYzYpn9YlTewoU
auwdpfd5ejlhboHJHi3UWIgykgUAjYljIlnpig38pqTt336izfTC4ZVIhuYokAxK
oyCEIq4BC/PM98vnLgUQiXqJsk05AF1Jc8txbpmgK+M4assLWuuAtAFtTb5Lb+Gy
239F4GjPyc2k8F8pdeqppYH0jpHKt0HuXS0dcLJ6z/rq3JEUV9Ybd3OBSghK6pCo
TTQCE9wPlSpR8CL/qVy1Lq62LHu4d7IboJqRGH4MvwhExDuXJHCu+gFvJPNRtkmG
r0KqtGhd+q/jh+h9QYEi5DsAsGPNKFi64gyXITgld6qMNl3mkNh2RSoysP4G4FpV
nzDTaPAMoiDZbkD9aNS9CqRihA4UtU2nAgR9IIZuHm8hIu3sMzPspLXTzttIO3H/
0YbUVnGKNPZt5laH1VzRpY1fY6wcuUFt8cpkD5WXOQ16de6xTqOl7lWsmeCECCQD
b36pdSqUSoQIjpGzeXBMQvXKpznJbT5UI+HsBIgIsH5dLe0y1uQr4qmAEkK1FSfB
NPOjRgopYNF1vlY8LDpZxjiuSRCAAHEpKaFepty5KevWtbEPNeetZOh6PpBFjnim
8YTAAUHRBKqCBSdu4iLuu0jZjn3sbsfEfs2oFqtHl43reRCO7953ikb01LEqqXwx
7wH33gmTapOpIC5HGSRY7Ul+TpCFLqRYI5KtXZkLNDhs1HnlVZNfeSioWEMv0lQc
X86DVeKdxilXMAz8FrlPRK6es5qio7Z/cPMTbthE8+jzLCmXlHIPXt/rbnAOUYNl
qZllpqGxifxUDWaTq01uvtmtxuxeIGtyk+l2TURiZZYE/dBPvVosFO+hjlSq1kQ6
wpGKG70y6SIKJIKuJYw+yglYLgf202p3FEeRPle8c6Pi+ZoTGm9a1/MEEyLwIP9D
toIgyrpHBttbKMYMlEqcHiiwfvtNapzAza3bPXQ4oeCekNqpfNUAZglqKYYNnafL
asOiP9Kp66b7HY3LKCx/mfrFO3qZPpqyF/Jb9d6N6SDaYiYc/JsFR07Vz4nYulrM
PFo2JsQ0smSSJLuGGYv1ioTSC5/HdoImt5R4ymo0PbCGwvBy3Iq8oqwgKl9niRWz
EaANvuYKwnGvxBhyznvLv/IQ1NHuL/dnmzWOJwy3WY/IU/qrQ9bhFIW8cRzPe60l
N76bVrTV6ukcUDwLESdRA+8v9R49gBA7ewt4POtgwyNO0tOvPADxkmAujL92BLO/
w/+OXNNMOq3YinuM8igH/0sMQ0XKq+UZVqX/sMqc/vXXzqTBYT5jJu0b+ksJsAS6
sSXw0Zvwczmr+3ZbG7dkxYV76prtz5bhoFX5aVQMxbj+1IKiqyyLamozH4TxNgnP
UNVXDqpzBDuQTb3VjK4tcuF/6HocEu3cx7EomQpAUhjWu03PwdB+FfMcmMvps1Z9
fRY7lB7poxiCsIeLSa8+e93XGGhg2eB40sXQ4K6GPvWQBCJLD1gvsbeRw7L77B+z
c9+aE3Z06vd1J1EGNkFPJcJruPW/VWfzib/Tle1ldmmYqWLdtXfuYiOA22ens49D
Kq2NJS6/bMtTrJ/9Blq0rD1+9eByX6sZUUjzs3ITiZIz+F7FZ18qHXgO0y3rphLv
ba3OU3cM+TzMjU/j4RwPln6hQJT+YVssHuUVZdgH+DQugCS8weUQPAVSBxtJ2L9O
7c9nv/Fhcq1FxBCd7pTDoBO4L9YxP26CsWohFNSO7oasoGNVvm2dRz7gTGFiSVLN
nnpw0Bi4E0ARbWQpCIRwO/yM2X5ALsQ6SpA6nSE0FEERIA10W5ebFzp5Kn/138Ed
gZ89ParOyVdeBoHAwmWCu9b4DyiJzZzOIeylnTGl6DwmoixPKyplGscp6Ap1X7vH
k71rTFy4lbkgXmIDlfguJlLV6kUjS8CIVHPlb8YbLU1CjQqD34d/mC7OqoXHPeox
tVMg8MjajR03+Km2HJ7t5OL2B4fssOQuhn5niB8UMzvfSLjxKmWv6NiFT/x4YMl5
f+jAq5abS2ziCXH+9X1t032mAacQECEnqabCbkXywByK2qUrkm4rN7M6BWAit6EG
x00V+9pUOffT5q0cyNu+0JyJp+whxDKEUOydvMG9OGXmooBxmlfZAdkTwPrPAkxV
sDeH5Aet+7oPxHVxjrwr3g9thDDa1eqdxDWH4r/01089m6D9EDVb6+kRA1N/Uqtt
RPmJ96BOyNzDNYBli4K6m73/6SZkI22xJPxf5+/PF89j4RPk8dMQiRUtX2S6twII
VEzINNe/Htait74yuq2EkWE73uNxrNy3lzSXiWPxt2ur6irEmxoib41354mXbM+R
YC8/s9Dmyc1xVewoZ0pnI3wchW9CqULXyWvFFWs8v2h3CFHT0Dpn010wEQ2iZ/LB
ooAcgxv98A1Pn+N9zbtpW6z1Q+IeFcHN+GYqz5tRj/aPuxnYR/jcu8agK7l1apeZ
GKJdKS8f3Cd2SpaZIJctkXszFLvXtO0DnrGvDSbRsB587e9V+P7f+Ay/yxKJFZbo
L1nGgdjAc2aajvqvZVCU3Kr5MsW9WObwv338LAy3vLmmMu6QZg3IVm/xIomqElWK
tqPwIohQ7Nc4J7XNH90XxQ4aaPEV4Q06/Y6Ni5dlXzCFpbiDMsdAkOOKF0XMLhlR
N5jKjUh295CbkRs2eIJ6hwpnuO+wt3AG1f3lXUeNgTqNjUQWS7exU+OyGhwBr2hV
c+S936JeJI1Qbd47Em9KdkWki4gjZu8q/gcO4CKF8AvWyJu3jSPi1g0KLCst8PRB
RPllipnudTlm4O7AfOGiDpFi2xMKaZO86ffLbO1qFrPLjvH05mHpbnxIgtYer0xP
blvEMUGV/ogWsENZDmhNMsACv/IS8SZj8ibNZHRXrzyd4egU7QX6oVuEu68M2ZbE
DP51Oii+az2hBSW/LET8QPSQvLgnLi4Hv0dwmyiSAlWjLpEUa9U1+UgaXrLNN1nu
kacaRIBMqhw0oy5q3optFoVg2zzEJ4AoaPbCyXhWIotGhN7p0ulrhB23JM1GpyME
OfIxf9rWSsOvTWTlaLpGpK7weigv3FR7TNjGmKWA2NIOfyWtMvBGVJgJSRIWmkzb
3wR82JP8TCin2XG4tzsu/E07AchYgmV+18HUD0nadxxtl0WG+fTcFz04g4+fLNBI
nCseSmul0eeSRaqh89ik/eZjCxBqORKHhJhRwESaG8QwsZgoIWKLyaCl9S6KVwNN
Oa0c0azbMoDwVCttqCafp+zlUxbrQ9t6DOUwK+4dowt9RHg0jeO04ByGidOLXZSW
weFXFs8A/2wLjkZ4rw89PrWxayRIbTik9zZA8MWXuHN6UGQ+JL+u6lW6LPKz2iPF
z3VH6iqHZ5aaK0SgxLBVmzF8iIXNxBu7g6qdw3IzSASwqNsnosWApjacztEFjT1m
p+CMArvXmbV54c+Wm2pxaeejt1/gA2qhkJv6duY3J3nBvHhYDKg3Vqzl2u4ln/se
QveLmnMwHxdlt6atg3TmMSVzPRJ8TmiRG0GVUqRgec6h19+tL0ZPMzN4P6JCA4x+
1e2whwLJod0hedKm8j8OGBmoXU3Ym4mjPpHJ/gmqogXjeJoQkbcWDj4S10IkPELZ
dJPMoirkFpkn8F+fNbqykXvUn11nxS4R8Ze5/JYHOPUWWthRHJH2N12LkWjJopWw
7lrw4BRYqjGztDUAwq+YnhbgI6B3MXdwIJT9XK1PeXUgjahWplzjQHQeYspRz9VJ
79vhrNq3WTJESWSgU5J+M956HrxWK1rl6fHWAmWaNEfWnPdNlmLRq5T5uOOHjN2x
sQptXGB3A6RJIU3aG1Cj8E8+p3d1IXajDY/p8EHSFREcXBFkET0ru6fzVS0z4bfd
vmPdDjZE3bUBGgG47gywKUCdzXKVR+FE4nu/kK6/5QghgNVoMYWDtO3Sf3eQZGTq
hR8t/DyizL3rj3LtGII8HyEG1f2UaYf5efFTmTFIKwoOw2ePDOOcfpGzx50gt/U6
eO7YRIrnjMo21l/Nd5sPkNj8BdGQtLGTCloqEUAOTCqryLgyIYtW6egeNl+H6YbL
Lu+rqaBGDUzK5m1Dxf46YYRzqbLQ1pKInFV8PVzMCmdkj9DFP5KwzhJrH7WTgpUu
rWdFjD0ugxxdrLjbKZsFnv2Z4yCl+BeMSsHhXcV0zZwX4xmzK+femC1BWisG5tER
pKauFNdM4UCwOZe6H8YOj6+V7vpWKVDFFoUbub1w/bUtUbbSlrVs1+MlnGrNaZMG
kEnWiqYdqONKdF3+1JJ36PhSi19X4cAi0Ls9q78T68aBnepdesA76yJ+F2Gyek06
GF/6jPjJHdbc3h7jeGMz6kapDJqbpSOL3Cp4HYaTDtEyHRd01IuvN2CQiMROErSI
Wx4BEKfqahg/UsJI2/BkUfaJegeXuTqkrmui41gIpNQU+dvyfphkqesCnhjNmkqU
oKcf14/zvThte+/43qVmq6XVBAWOfS5Cu0NVa8FklqoIN4bp8pAHknJW9Io5tQAk
zF/PHuMphsI00vjz8hBiRaiRdZxRtUxRWcFSJfQc34JVTtKeGMq2YZitikRkwmy3
uAKTQHsRexRM6xCYLRFvx21Lzih4pEXa5nDBxxfYotYJnrytVjDo1bP6l4/jvh10
TmcXwiT9/gM71lzsp2uVXwEy5Ojv+BFLxfAyaI5OQI857/YhT/TH/j+UPDoEwv9v
YY2tMfNcoqrL34v3O1LTZrE2tM4VK8fx35NtPG8vbdm/5EJyFYdGq+XyPKc8/5YU
ShjxWf0Ps7TvLJ4nyu86sCne3BI0Dt2Gvw6bsNCs/mJwOI8spp6iql/Jx+4Do8mg
mPiBk9yETHGOpBwnQ+fuIY2cPLpT77jOAaPFxRs6vMrQE1Eq6v2L4rkJOZN7i9F8
X20d4HqYjpmIEsLPvZWHxCe8WU8DSLVxXnVBjcPJHZZYi6qkEU5TU0WbB1hVSQ6z
wK1njtbUSGHGUr5ZVSruQttpxL7Tnd41WjkLztXZYWKBGyxk8KyI0Yeijp9UrT/H
sdteBgAf766CEJCpTRFj6K0mHey064Tnx0jH7LfbopitqDZ94GvXSy5ElzcUTic/
LknGtPiDFCiazwKzCKMYLcDWCyh2cUtf698M+VPAMZTPwd/wVzOqBQYiTrXoMw7i
vAXbiJOf94HNXNubQ2key3q7rKbM8l+ev5zetKK4lmCOj1noF2kXv1JgKiss8Dy1
a2q4yzLOXYRe6mUVd7auFykCohGmnhoCKJnrnVTqNOpsCJ4RftYwt6cX8OUuQ4DF
hYFvIPZuAibaz2XcmbXzbXTPS3atktZf5qjoTB4vYv9xN4PlxhGU9qahK4AJVO53
Kaxv2DZ/iBu5VxsqH8ektNPS9xyCJ5IomhVgsttHfADmnc0Bsxa0XSrf4uumqEuw
VpeE7Mg2jGj+NhiaCd2QUVP8OIuyNrs2zZFrGGfggABcq/E/Ju54uH9jxaljsmxS
0F174cGh+m2Ahr+mgL7brphWU5r/vp/DorkIa0CLh1he+hm/tWigBmEPWYaiAgoN
jmMItYpwg0hiiTmcznG1DpaLlhw6rKctyJxybsH0j5+8SMDolgMgvAZkf6EOLdpZ
+BW3f8s3GJBebbo29rNmaJ5XCkzTKZflPVLBER8xrz8UWd+TGwwPTLQ9AKkaXQEy
yjU25SCJ61vVW7ZoCRhtqpDO7WnID7qhumKakT8HEuJYFlQTGH5yKCCcIhrmjwSy
48LsB9jtiIghJdwjKqKx7btAcU+h9FV6lwBzRgDWZ1wll2lBEnFgrVht328WL/mn
l5C9ibQn8fA7PpDxCeFV2mKyJBuoDdVu7tkpVwDi2l7HC1iCKoah+FdQAgSj4rkg
TrFQ4G6j0gSmG2Fcdqg6NVIOyueSeua3MqZA8AVb2Q4cEqDpNdTdzTVHhTv8m76c
OwtgEl/0Q5a29Naes5yvdgu5ShR8mhGnQSbtdwHYg8TH4MsA7d4vIQwT9FIm0azD
qnfEgnWQb0YVyyxFL5BTH8hYCH9eszAtyMV2VzMKAjD6tiWi6QAOO7zK088+v9ri
b8FSutGWTX9sfqO+W7k4lA10isI59QaEgCrwfBzle4Az7bN9jzzgZXLdxlIiilvt
KoW49t4w/CSpJvjmNcFDp0cqWWfXum8d35CZdbgqN4QT2p22SyxIgDBjtS7RFcGU
M2Z+BVQE/oGw8xjvEII5UYFItH5We+4ebsLifqpeamu+LTYkxMHcnxzilFHpVCy0
x9MDsAwzkBg6DPv3V4hVsTR5PZw3fCh+OelU6mOyffTWfSCmZy8ibV8Uhhi+DWeX
HT9utDtxkmcFf2yhWiy54KwHNUmTIg2FO4/7trKVMQJDjIGPxEJNJqLibqY2qN+B
1gFDzmioOJFOht7uWNVm+QK26VLJAF4t0/KmMP6uJjsr70yRj+B5h7A0N/kQGf6I
U0FyR+w3dBoA8x2UmRJBljexnhCVAskfjACkSTGjHmV6YSWE7+/h4wFFQd6BcLFF
9qqSSQSEYDASJjItDDxTxSSlph11GRh2dY8AMgXgHhOiVeSBa6Fi6rEh2xcMu0is
JiComlYACiLnGcSBoRcgsr8gUpo9qmZ5eu2A5MP5/5Z6zbhpqx+trr8+ivZNly38
IV+LgsY1f6oz7y70WMf82HdgloHwHu+CYjtScVUhmNuk3csw/auSeOFGIhK1sqj4
ZZYyMLrxibGYoKUZEHrWXHGr7kZuu79RGo3oEkCJ5Fc9lkuKaGgDDitMv6Y7TOJ7
8VSxIs8s5Bj8qEPbAZSv404Lf04qgcRR/UvVrywfCdRNzw3Fpo1+47CuiesOfDVu
OT8NJy95V+LT50VwYIzCR2ay7CRrC+5BIMaav1i2wi+u+ttZB2Vj7ziGqUJUvEep
M6BmQdVQmmZyzWXYjaeXLYioo0jcKb2CWcVBYTkA2swnRHGrDhTaJli5LAE93Hp0
v5H21yLGtpSJmx0cRIPqcT7988c82poj+tvjG3R0Mt5CmWwW8MJuzu6bnMjkhXQ3
UNTTe2mtkmrMU+8dF7moePDseszM/OKxOCpbxuXYrwQYzAPWcNQFw8KTycLefBZx
LGNOT0pemsmBvqzK2IZyW67ZLksKn+FFPUbFxXUGx9YHlmH3vyq8tw2HmTq8wWJj
XE+cFSSsBZMABC0+pdVUstSHBKLpxgcgroPLpfWmiNYB83HAL83KGi8VFrzm2nkf
kooAqXY96uXJ3l3sHoi0AWktJRhTaei4uDMHijvPgdsrIj4kdinLqjrk/h8HkOpA
ckTPeSgRvTQ62UoJR7NW1ZABQT1ovLaSlMvB7QiwQME3WAS+0Cjvb6Mtk64JtJIt
olqUs10OOWgULavTPQ9m4NOEIIwVruV3kl9Z4+w8gLBRvuYnGzOu9UdhBOtlIqKP
d2MEsXVB6B2xcruLUpvQ1Yrtuh7olobYsXjQ9FvVfWzvjy7ewthpiCrOCnmB1VYw
fk3fLskMFwT9dZ3eBYnnF2W/cI0G/lnst/Dt2jk7h8+SF/FWJXljtjEP8LFrLaa/
DOhzU+CNhqRtcRHEDbzHINNDdIoFTGz3Hgi8hWO1NlClNzvxADvtz30oRXDuTJcO
SPqlmKbKUTUn5/dZjKKsLoXxViCw3w/hOvaRzh3C6YrxxQWcGgbuS1FiI7mDsA2x
rSSaoA5t91m2H54sSZqDoQ8XcAai44WBjU8ervxB4C5CNsodFA6uDbl+qNcRiQXT
AUoan4jrUEVF1TMwlK9+x34lter4pfv9n9oTklJTBbSVCKYzihI/zMZhrydZrREL
m8qPz5yLgk5n9UXxrcVD5WHj+ZfVyoapUKhX0w3o2yRO2/dH+KzmnLggL3qROBEC
Y52xifFk7P+TfxsMEC+/C9K3geepoHc3gUK30fiPAF922Jc3zg6Ya0xaP/Gdb5jx
fKtcdcOz6cVwjaNH9zSH1UboxXqmYL8YR9ZE5jAOG57W0QeywlmcGyrscO8wAPQs
g8x/Z/4gzjwAQgGof+WsEhIhFH1EZZmVjeLldSKds4i9XchRmKwSV3JkmHhR6+tL
1rJsk5INkfm9HF6PMSekKIiDCdmFP4O7gyrJcz6ASiJYgDra9mCVy4KxFzqygZAJ
2S8Con1MwOxppMU3jQn0cG3Gf0riVdoaPRq6TsxcOczs1QkOTnVMz29fgXNXdj/h
WbJ37VjA9WdOZcBpLajB1yI7KwjJRMn+ZFwq2wIUbQouZ6DUOae5IwjMpu09NbfF
a3sCcly85xTPQFe043DFFO9XnkRq/615BhKBJVcSdxCpstYQKIUct1AGxBpvatgD
ge2rhQLO57bZYSGl/6D4j47eb1/B7fRC5TQj9cy0RepkwMqq3/bs1g6kGbnOzx9Q
8DRd/R0doEkA+CbbhflZKMIg3C2sbLDbkrpP3o9sN5bvDZGmkNlySBXHRA/Vg6rA
aSEteB52RAmUk7bM2tbNkmWxcJJ+ogrzhYlKOyH/voUUCrCyCBHS8Ng8uZItJ1J5
OpsLJVTJW61WMEQ1VPjrQy51JtYbpwHcxWprl+3B4vOVS/BYets66To6Ur6h53z+
20lmRJUdM1etevpCGJbpPRk96F+80radzim6+Iw9GvK5kP/zZPgEJbkoMNjeJ4Q1
hYamajPj3ET1rmoAiF9Hmfm4Vl3OoZjL7iGDGxpdP50oIyezrQAj8u4kUVAI6UKm
XTvOT+QbfM2gQuImw6Xu0XCr5fqTzD6UQcLNYB/OUV7IixEb6Yjeh1pBF0Lz0m2C
6mcWySlq4LMUYemNAp9ri+rDTc842qmQpfCMOd0n7724brHoQu+TXm1R+ZT4Gy6O
Ir1LCKS+oE4wmHaS1v1IeKeYBGbAGFukeBR/732J5Rn4d7KJfnQyR9EfAYWhpu8x
3JheMFiNN6dBzHrsEouwFlyhGW2/x5OBgcK17phAhm3/p9kipM+Mhq2Vc+RhVI+P
/6yHqz3MDQT3iN/RqBPhVnLPhDjSvFoT3r7YXR6g3bOY+Z1e0nKs1p5f/2yUBig/
hikTk9obFvKTPOrrojsFtSWrf/FR9oKKwlRyooNE66tZoVWhaOjOBgiswdRYZLW/
x1EnhMjRmiCJUlqWrkrpKjmPanJe0524dHMLsX5MnULaVSlOE58XPWVKXDaI67Ve
S76g6FJA0qlHvyieX7Hrjd4qQTVQs42feIuf39yvulLlZ4V8dT9neHDnWiZqWkBV
0bEeAjWfgbGN8xsxhDfKiuHDg1bEg/Zj6EEoZX6lXl90sHlAw1n6042Ah+zbNdBd
ZHMMLGCE0PwYT6aNzOS9ng2hOyj9EEYP3ka3o+TnQ7ksX1VUWW+EPpBiyzDAE6WT
LIFsp4CkVBJBT0wT+X+pK2jgwSxToCoPmCQkWm5UPFsyUwz6IVPdVAISzRg6qgV8
cD1rrhvV4RxG2g3q/akYTWrJvE/Q0lBulIq8vhOrcT4XfZVrrdcba0chAePSFF7K
fZaccwqXuqS171AGlV+bR7f1LDwSS5YeGSleGdYbYAmG8QD+G4ygc4+z4mDxx9gE
IPwVGEemcoIeToOpvr9OVCPkWq8Cw5QEymOjY5QpD8PnEFv+mYoZYuaLeKMFxla6
o1YoUV18NGPD3huWd7135yU4u6sFjcYsYLMqwJHNwUNL8L148X8k4OtWMoCnPH72
F/85m/C6qfZcTiLI9dVf/EoBZDw/bJEwFMRXtXSOUhLcSVPy7Z4buyF+sjItiymu
KV7fXFh4aLopwhk7z9fFZ8GW131dhjLvGtBB5fG4XqllND9/lPulmhyEX7jqcDU9
CWzYIablAb+ibrLSwo0FlCN7xkErJIDKfmicKJzLjjiP1RFd/rmCuJyBK2A1Nbo6
HHZujKN+rQ2mvFG+XaYoVq7LRIy05lmks36uYQf0BAXerGwKWZxi/c41cWg0NCqU
vb/Vav9RIGAikbKdJIELTL1lGmJDMlamrT51DVT7Y4ZnAD2HVqwDYQtJtFl20hRA
idX25SUq3z33pgL6/2IzDw+da/ysAUdTa2ngSZjzUq8sFHCDsplk5d0aTQMMiPCC
IHg/fLF7Mfi81naCfCenM77TmW9sq1boyz8qaewBYhyLgy05A8EIetmVDhJ3rE2a
0VrXLsNX5b1iNuL1rVnnRAG69KbLB4G86HHCdZLAZ+n/tXDLpNfPHOGXcE2eXN0D
jo/6/yHniTEldW0JY4/yHUYWvDL0oZfcaIfg45zBu18Yvtl0J7zXVkoGUUQBTtXv
lWaCH7fUrqWvPpTIDrz0gMe096H+fP81adRgfGjQfBX1+AD1GOWCbhWM2BCqlEj/
A2hfncYD5ZAU5f2HvOInicNbupq2ZoTjZ1bXYPckqb2DSCLHQkEP29/z+wZpbtT/
TEa8eNfeQ9ptaRpQcq/gmV9ivzeeUMU+txN+iKDBW1Z8lVHDL2GE7f8yd7bFGJbf
dBVzcNMZMo3UCXbDh1nNC7gUfb+KAzc/0FLQibMbjFhbnajVXBEh8uROuiGRxK2+
iv3NKogaRtExLvn/cjse7FgWv/x1CXT6FZTTCOPumNU3aYPeZ1v5kpFkr6GlL8+m
KbXCcv6y6p6znGUKbnmP+VteUNMrXQGRvugTL1tRmauABu9/zndX8fKMHUT5xT4S
XzwHA9UxgiObGA6yKvjwais+VqhiH4TaqoUdEsZVdMxMxzPTcoCfvsl3eUX5x00T
Lor+orUmigVkF/qe62HlphR0WNhXDIMV0JZrS2HZxYM2H+QJd6O9leABfbfM4oj/
hpypBlswVBpmdlyIkhiN8acwTPkDb0bRnmQpUC4qvpmM0rf9/u8COoUSO95eAvde
CDZ3h1tb7T9RoJBgy9JDtL6IGpTJ8/0iRuJZJpcIV2jfOJp2jRks4gKmSqQKvHZE
PnlftJBcYvl/mx3JMcAbsz4gn/R2DqibCl5vejX0ZIzJDOzysDXsp51yOx86YZAG
7iABlyfxAvz7my0FtCly+BBn51U5EBx/lrB3FLacPrNzoYzsEtmIORAvf5OxCedk
J78mS8RzAFGGAcVMoQM+igmFqTUX/1tsAZ/hmuBY/oey+BekAcz+ZODwLcP5nQxs
GFr6eIOtcIBSjQ1DW/CjLuIjzCnPPPEZamY9BZ5Pox66EvYDZm0EL8DsbvYM3HzR
QUcdRXtjeuDs72bYA1t5TobWfM7qL3Di2c+9B8/o4lXwZCiPDJCkuEW2Mmsvkszu
FZBgBLGzI2YPkXedYZ1UYBE7yY3oA6zqYIF9bhYFW1HIQvragIkXyVQmTsZc1Sp3
aoVKJHNCmKo/I9k/4fgwKl/ecr1ISsyDnfyY1MAiWVG+EYLj9LGKrW+78rTPlGFM
2jLFK1OKtqrw2TH9GOQEfPHYp2C1Jr9pyHNhIJdFuzTDLzhqdRMq/DV0y/cgEIfm
Ih7xh8eqPxF8Jej/hdqkLbHLLbmnA8BoCddAerVE4DHmmUxeZVBnLxHbyRaUjXSV
iuEZ+No7azIn45eNr/XXU1dzcX5UnPMOCdBlJjv1/TWwQAXnsUBiwK4P/3LOoIl7
TM0SXdqPaem+JKvk5sKBzYGhUfXG0QdYBSLl4TOsYKkHkkGznXTDKURbguh0yGl1
kMPbuqjSswIH99C1I+/iJCE/PZ2MInvDK7Qn82jDreZdX44kV4JsdB0oYbn8roXD
K6ZITLZhFAo7uZmvMWFq2wg498+Kj2fjShNgICL/WD+9gQ7N0DKgBtqA4AwrzJIF
CGhoKyCWOhCyXXKdd0l//ad6J7WnlqP/Piz5IXp1NG/9ifM1RrQxuzGRELBKGvPe
GitZ/uVjnV8VtmhJgUvc+3ukHNXi9hFyvILZPR4USgrnm+EsLQP9E48bY/KgivKh
DgK3130QCNhR4Gt6Wr9fk6OBnvhhe96JZ7KKOylnOMlZhlv1jHAUzXzJ7OwTu76B
AredXlvp/fpDF7KDuPS6gmUzHF8GHiFlyhRDL1fhPlwO42XEFXc+zhufF4+nttqg
wtZXqNjUyP4xSWzNrfLI/31XRzll45SEkPwIYH8pdiRwv1mzmRdkuXnMyAzytLH7
RTnMZGyTYIANn+rUqFh55SmNwn73mVGK0kk5Dhxzmc09ci1Q+fMGx7pUwmZVMWr3
3CLNk8EfbHz3/CTDeh8qJ/ktNPmc+OUg6MmyDgPm2Yu/ZY8jTddAVnSOIgv/8jZ+
joPrp78mic1ON9hg08yf3eohRyo5NjlCD0Onyb5wvmhliAljkFDMwj0mfFM5urkk
7Fq5fHvRFMCIXQNkQV85n5jdY49Am7G5I4q+3zcsNLPJQmG/jZpSMUDnNLPU0JON
qrFPcfrMTffKLKudKiyRnoixdRkgFhPJmDSx5A8edQTdWyAAnVCGVa36y/gaqCJ/
VtZkYlTHYQuD7rz+uMSzVVYJHoig77wIZ5t85k8qTtI3No1MMecudjtw/AtGa6H1
4QLK7eD+Gcsf5HUZcidLpoO9VAMjuP8/HY+d529timWjOovRXtA1D7nf0Bvzaiu3
zgDhESfRt+81m6mS9/HEiLck2gOfkYnPwEbmDyz7PBUFjSf/J7pZ5B10+Bw//QMN
hWjLGfwQb+p2WeVkufNebGb1uVHLo6rceFHvODSmQbGYQU7QbiP9SGdK7eHwaSp5
U6tEx2vCQT76zfQAk8+j5PYKB8RXZYg5qEEQLERIWVSq65KH/nXB4VzTnyU/Mc1O
WKPJqSDHClulv5yLkiKnxHlxOdZfE7TQG/SXY9WUa6pi6uF5oPgrHyAYmJtJxlmX
AbmtD0iLRZyQ6ySXh55xyN/b8sQMTjbS0QtzhmdStLaBc5oaVZ53ngjopB2h/DRo
aPzbPkYqX5qH2pRK8tZNWIs4uw+6gWnx0NT5TkThZN7DS5Xt+3g0jmzsUumj57De
V6R+phboU/QL0/26donq2Wagxgr0B+j4/kFzi0FIUNk083jgiH3aWO7J9yQfrpH6
ZwaqLtHXZc5CFk4sOdW4VfYEovkXTvElMDA2cEpDPkYI08oLse1ayyb9BFgTgg/0
UfPaHI82JkqWulC1RJdDy/gyCPAlYOjRvifVXczv3RyI6Q+y4pYcI6F7s9mtW1Tk
ltepRsCvHPDYWkvQrJ2mXbBZPMw7MGKtfC8mA1vc94VuPtetLargT7vFSV9A3rRh
6g4acEhJid/9nQXvaZcOLAwbb6CD27x2CL1xkfIBUlDag315/JwnTAOiZDmPdUi0
NHIVLVRYrPnNva6W56Gq0r12IRgo2fTMUOBYTAx8jyrOY8cxqjeuWN0212hAheRz
ZIjTSiYchlqwCtKDBqcXZkxMqCSs2dcA+QzhYFhYnoL8vci2NFzS3a77kbhZclm6
l3GRim4zsUrGQw9Z9zLqRTrDZe7EtRLubSVAkcjXFtxlZP0x15zcUICcqGNL/rw0
E6orCj8o3FFYtZnHOzpf3jdGAnJ43OaGxfYNUt44XsxLXI5eoC3jEZCR+RDz5Jo7
43ZJFUhn0rtlHREsmPi/Ahl15+ZU60kkdRKB/+kbTrsMyUIW59W7X/Lv5onFV0bL
XR6Mw6uNVYSR6jONn5DyLvArvG1V9ZDF0Ql523RmBMOy7P3xXV43VXwUaWwB6OXp
FjKCFNUfp5SqrFafMZQ8EtvjbcopafwjFWbgAhjzsFxDPGMXfR2pdgE/i6NSitNn
zxA2F8A2MG6vdMMi8SKXu2wedJceLk3EektLUrp0yWxeBe5HzTq0i1SgQs6v8XuM
ovBIkNeyOc7S5hOZ65Hvk3R2pPY7a08aHdGOM+jYDv2a3xgR8wGGPYXJaRCTMVY0
nrpvvr3xQVuENkqxkawQInIdtMWXa75DugGMvRlGjhM4yrK5v6LCxmUuup5EyP9u
dewMSAXl9oW60+SDBniky4Wj0DFT81qrEuZNFc69dEqTWd3gM+3FRYpdteteRm+x
ugqewvrq7Yjti+YOE6A4tM+xV5kTMFTCN1e+fssNoUXvcuxzz8Z4c2mlkcg2O0xo
g4Wh21LlleeSQwacUa5/9ZhHUC7qjXsLGeyDLRcNuWKIZx2wHMxp5i8yQfE+wy+Q
4BlextcqBs6PAzMoQDGac61Xj3tBzMrnK3IPpqc96iDchS8+XzisPK3ChfO87nOS
X4na+ENlGA9+4+7bEURcOVwKD1/NAhiHB55xoKnxQ6+Gr4I6Rheu9y7bv4W6Ytap
cPxVeNT808Jf+tib39E27LDkC5eUpBFsoaienunbgog62Dc1Cl08OfGXO6z6DZOE
DdHAbdSOCODdlhc74jCC89wE21xAicvzRYy9QjCZkZRkg2v9g/oliBXsExVy08G0
Gjcunpkoq4bmrlqf+JqfzFeWI8ERGPGsMhHbs1eyK24VJ+v5Tun0QyfTRlvz6I3/
cYRxiky0axlAJnL4Pfhwuxe8vmbdffP7LsY4pLrA00G6aFnW56hPlrx2Uz8X41Pn
DPHqgwo/MFvv47cPxHbImkQFqKkfYJvF5L20XwPWavBYaoTIPGeTcTymASYbNX2l
0Aeo8gJxuZhwcJGganf7n54Hg+fIejQKuurAVVyuDqU6Bv05CdtZsg5Ql2wwPkHW
BuKHsqQ2ZbBcQhkFCtm95bPoPcvCfF9824FRcKuW+PNPeHRuW3xtfy5RPdKXi6oz
NlNJiGpAU78c53I4tSAPG2KRhZxzvlX2xyzRtEbtLWFU0RZjYLdYZK/0eHypPwOY
FbFmd5/trm0a+wOCz/585ZwXMvGLP2qbT2ChoBhEsdRU76URP7xF0c3QVUVDKWWs
r9smN6WVzLMC2QIOM7J0yTKqHdw213EvzaZ4j+03Qyh1hGDPbgwTkGEcL+2YNnG+
HG4gaISR3ctDz7vvWBw29X2cLY627sLUQnagz9Rg4oXQS3JfHfdURoLS6bnilWa4
c8ZevsGlXU8Sg4oaxvBrmfaPAufzg9Co6MK3AcO7aPDIgtOcGF6MdVxlOrzm41a3
96hnhETd/DTKfmkcPu02MpzYSt0aJDmXScmKf73wpjBpC34hmb3xgRy1P1MvOQGF
YzrnoD1+T8h56PHOxNk96GukeWAWZKSNVhG8/GVN2UHHy2v5E3moIem5gWCHRyAj
0lzYfx/Ae6KFNeGzf9pewwbwQZkfxI7/dlrmqXZ3Yq/VHBgmMz3LrHioaqX/g+rc
q2cmMnlcbeE4beErRXIsShqfe40uSMGranEYGO5m9tyQU1ZDpq68I/7Wz0FapQ4U
hUlngmTgVE6z/WWwd3XuOyLPQTmRb1+lQGKYs4x9k6btcHgETsi3agcwaKB7gcnr
eWQKkvMS6i7MXpMV5dlwBx5krgoKf1ZMtG0HImn3xrjg0UfUPWh+/D7KLJIheNNY
t1blSfbyKnOs28V4fdjD6vCUDSXXB6SgJwPZ62ZIEXKRD8unYltEm4dAgDlXLVNP
UdlzOkYrE6X/em3khr7JsxnS/i8SLwH7ten+2xgv7tQpKM0lEbI4oE0DL0qPIcRi
OaG64NUiBenyq+BSxHCFVAIKUARP8xGyK4IhAk5yx5aUqzgisAOc4rufCWII6dHN
RanPEdE2uElrGlZ1n6SopEuXs0D0HaxSTh2m3sDEz++bY3VEmPERXgX9aeemF3Uy
xOkThFnRa1NrwRWSlDHWFfwswv5vRsQbha6lqUB5fSSkjGU0X2iFjT03/2CJrES7
7gljKx5aWu3PkdPggBadmACwCXivCtG4QTqlYlwN30rT5RPIETo8MzrCiUyKxC+w
3FWQIh2pAV/o1mv0Qj+LXog3G0IShUvOKVcKqSvSguhZ/e1RjVpMUPLp8C4+RGEv
C4tZAunjY8sXyHfH9gcpgnJ+c7K+bRjOQFCKm8qqZYNMEHeS4fCi+DsvjAmWP4xs
07j3Va73ztRyO2z2oLyfDIXHSn/ckRNTOcNN+u81BU4Y1tzaAE0PfFY06sLQ8Fi2
LeX0SDXXHCvasdv42DhFc1UQj6Af0It4H0qPfedUNYvVsvzw64VLdOuVIZKTL2bS
Mqm4wunhmdthoj1v+JTRcyJ5CKs3p2wdRT0q2GXMcOT92hZYMJBN0w25Z6N7NIZd
8q/fsFuyGfiIQRc1Lm8UMaUpSfweAxxWhdmVbFDe2Rl7jDO1P7DgB4ztsj4oZWuI
Cl2fTIQDA+xjJhU7EH+90qh4sxySux/EngcV2XDu163v1MKvk8a3QsDUDdNK4i9P
TAmbnlVsdg2FhW45v6EiKtXMbE/8d+7WD/YolYWb/FOfJqlifUtL/iccN/rQFWVH
Hw8SApFRcuVHazLz6rl7Rt6kL4jOYjbMBnqT+mkl/HONLrX5yiFR/W4gzXdkrcRS
pDC3JNvXHdOsetMIHCM9Shke8Ji7xTxyQ8UhPJFJYswzDUwUWuUyaP/epW7UT5Gz
KccNYKiJoWuyWX8sN4gKE6FONbJKXr1z357pUK1LIgj6w/mTMCvwkiOpuul6It0p
Ljq+sSwpv3xxfuFmsKPWUf16yL3qYGBmdVX6Ns+khPRQWjaUwvnLqk1TRI41dzsL
jZ4mS5G43W2a2G2/AFyhzy5e2LOVsJLNg3ggsyQRlDckfQHddM/hQmcwAuLJliFP
Sjs8x20grZs28rjTLz5PQnXuCdZqn39nGtSsNBk0S3L9hwDpooE0mE3F3IdNAs1t
Lns2MBD6uQQwU7PSqqWM8aUYsFOZpBi+rptPGpmlOCEyX+xyNjW9BUM0rL0lE4Kw
SMw86pcpq3WUVb014B2A0U/7cT61S+tj8FbfmRmU/G4oU8BRGhsWwRKEACiqW7Yn
Q8q/opjfoyw/dQhhF0DFRUNtKDJLubw7LJmdIDbx8kW/KbHtSb8NVq35aLDJdl7B
ndSqXVeFO7HeCjPSgUJRjIeiJ4K/yR3ujdFunk4J3ipzZwqD5aqZQbXxa7IIQmPv
KO2M1oi7/mG6NCumhe/tLfc/lra6vxw8HV1z5LhtQSRoZwcQa8WQpvfsyS+ONKzg
9IRTUJ54ZXYTYX4O/G+LsBaAZOJsL/HGYPpqrIPK3Dm1z4wC7ugtzGBW5pFPNejZ
KjcJtznWPcccKjg2QPiNl7xDouER4Jj6qxYLRnv13G6jmwKJ1Zj/I/BDwsL7Ovy1
O+SEDEMH8jvhOTV1cuW5gYetnHUy8R+dtcFzhhpkGrRzhjWf1zMvD0f5m76hQXpx
kPJ+zu1jwYI56SGdrJg0mJ7+ZvYY7aV8QeJkj3jfvefErm+Sx/m56DH3aJQEEU2i
r0oY9QyYm+mQIZ7Ev6ObERXhUwNYICsep2FBNWdEGESBEx7yOJfbHLRmBsa8rLy/
uBpbu9ZyNltRrXkswmE7Ikrp8T2FqvAehd1zk1na5EPD5ZY/G6zBInfv53es2HAS
V3dUtyi7Bc/ohbrp9ecPb5LFhI6CEmsi0asZRzWFs0fM5sygP17ISNVOus6XfAjQ
N4BgPxEE2BOgMCFoXVXXGofwulDuMWMCp5ZFM+BBHwBx8tdv8SALhAa+VKILQvTz
/gwxc90ozZvTy5m7zeZqG1EL54hdaYZ9LliQv3uCqZEjEpu+ltWkvuv8oTid0o8z
0Yv+sJF8T39VeJyLQkN8jfqfivn+1akLfNtbcqzYIYmNRe9kofwyCKToROErCviJ
rSw8ELMQAhkh+dvQfB5+YLfmvDg2cqLCG8TjJh1dnrWSnVcOVHtbUWy+n72xNHiV
e2+oy/JGSt6U0DrE4tR5haNglS/Yfkdlnce0Sw3x6A4txKyUhFJr1H/E7LCRo4G8
aBWgAPNyUHHPnmidPiRPMtP5Wwis55TpYlIZYLVlcOl3YHNmHcilSz0UPe3TTGHn
+zc8qwgo7+GcP0RSx2PsoD08ywZex8yeJ6hqnSbBKIp4v/4+Q4VEoRvAkdSvg8Vm
DKL6r9E3PDzUGLECKZEJIdI90+o/Xma2NX4ufTYPJfstD7MXogYkDIowsvNV2rXj
OXYCkAriJsL0QtlZZG3h5sWMWxR7eIUO/RD74q5R4McaaFppZvWTNqtwouPX3Srm
IpuJAuecI153gTpcCJ7oJYHHCPmFRISgSf4vMHVtK9iSwjs6BNciN27oXxtUqRdn
C66PPhuSFmShLFc6xgLIbM9O65QgEuzFxWKRturMJT/jYZQtVd6kfZKPwFRWwNNk
7GfxPPlByoRg7nBpacNc+9vFHU7wChVDcJLT/WynPHsuD9hyHdfJqTrW+GVAAMc5
L5fDgzCYKRkqYtyNP7gjMfk2BvFzpsnpblZa3EI38jeNupSh7R/0QQ9TMxh1yIXn
PZuPF04mVV/HwyEeR/hQxwLIX3n1p3Jy3skOW30z7padelTACkOoMeYKf0te0rc3
ecn8FJrhZSqUHKCPs2r7gzkirDbcVzpSPPFrebti8hfdAmE82BtxFYwcCF2aoZys
0KXhpqP5KKgToUBkO15LNI9Sla1rLQ2S/PogUbDeqNZ3pQxo3gH330sRAQJ2vMYv
zb4t5WMHZUDAsSzPJ3mdvqdTGei34++SptOKyN4BWmWtYT3FZa0Ccr/wUMrOuQYr
OQGMRl7g9d7EihJWnWBsAquyfzo+qaZzlX8J39NbzADzNjExrkrc8ONDTkpIIw6+
w/TagNWQLMGYtkxZ1ijJ0uVUBPK0i4V15b2vBH0SDMYMa+x2DFSaqAWGum27t+jI
KCRbpwlR6Tw36eZgUtPQ2HPa8GtNUGWy6QUSUMaH759/SvHJfHCgaMERig6mr78F
ldTDJPhIDkFVikCiKf87IyPV/Q8KurOMqiEKLVaft/vdihpfx+ivBSsJVAGc01ek
tHyWHXCh7tLozxMnd/W6pnTDV69uTMWfBFbrsFfOy/q9omMWJ48teWBg27p6sP3M
5xF1s3LgchAeMWOmgTnZrYUJRuNIyVmlkhDT4MsaUV1M1tXhGSetX0YdtvrOCB9h
gBpZ77xOxkJUWXbxBQmbADiXKddWfjX0Mokn+YpJyFglxRAI8oQVxVNF8E55QFY8
1w77nYHVcBy7CS6I3+PBY3gEbiZ4VVsiKY8Wu1YvReCrNsGl1oeRDeg/UNkGr1lV
MGCxC5uLqVsFSoB/6R9y7gfW0i16OrVYBFJXJi+r9eRzLZcSeIPO3QujfPmWYI12
nh6dHpaRSkDi89X4lDd0znE4McQNrfckoJfTsMO/9tF9u+adtvYdvHXl9xnYRV7j
/hDj0G4FYkYh/onO+xvBVUe4lgV0AxX3IeWOcnpIcN11RQ54TKZqHR6Mf6VX48iB
yZI4Z3G/z+f2wuXXXKs5eUji5HV9ozxNTiGZB1s54QruTyOMPZhXSZt3/J2j9mqD
fgy9+/zxj3m6rbNn7bAattFlsioAiLGhM/GPLKoUAZFvYbs3tPhpYXqwwB/9CsiH
WqWjYbcNKummg3UtBTJDCDLzGQk7mTiOFOyiZXoJxKv2BT56aIA4vc+roNmwec1F
XXWTIUQKGN7WCMSNUpw6gUGPF+VYSc77CTBLDDPlvU7xlfoU6KQh9BFVmCDmCOUu
LtrdGeu+jCNTc4NeqddBt8hzHgpWxwlCRoemPiagQ1OuLROMfYIu7/hhgv9pkwdp
/etDDnDgmImi2QKehK4sN1pTxWBZBAxBen0aHOkLXSx043jOJ8VkkoOlmPRpZGOI
voL3G25hGqter8ij9dlc0IfKpoxu3IKDdw6I7uUumoaDaUxciyWLRAmVhTtGgNit
/RpdpslvSGrxY6WhvimiZDrqdK1f/AqtpTvxrHobubnXopU/ezqfRAK/GXR3Ng0Q
lwOsTW1BsnOHRvIsHpLEPHZVG/YVfF5eKJrhPtlxZOnqVtHoq11tsu7rDerdd2sU
x3DLDqq7Uv2yDFaA/fMblEU5sNoLiFK53t+M0/c+NBoFgO8Dr3IPHHH1TkRpavWH
PdmqJhOZ3x0g8B+4pSXw/5KNbzzfd8f2y3fa+iwmrLg0LZI6kXrAi14tb+hkKrfQ
CrkT+ea4AoaKJzQytnitV8fJH8Ga/ytrQcDWngpnYuxk0ucQoZ7KeiYXwDDm7EYa
IxcPbUCR3hWvPKLH71UkNIFPerUOqdc/M+FMiGgnOJt7FpLBw6+sPnVy9BRBMpJ7
x06bcmWrP3KzP4MPkZkyfsC34JEUtONsfeQABRYGYPppLxAX5ZDMG0tUSZ5Rm3G2
yHocIYAlot8F6YXUmHrWw6pc6n7bUs5WSpj6fKhXePgi2XQg+HhP14iPzUQeXMoN
CbmSpJZwBjk14/JXd09e6GxxZ9Xn4PoD2QT5vFcQ2kEKEUNH0B88Y+WAAzqyPLwV
uBTfGO3PSHO275UqSzr7HSvKpSBHKxDzsiUtba5SG4rvFR7O096BOTGOBGVMw+Di
6P1jLpI+FheeC4Ra2fuq0Zn122eYisE20jkY+pHuGipCB2/Cl10tDHzri8ttMl4J
F+HB66dQLmP1fT8MCb/g9N/g8e2Af6hpZuMFV99lt26cE1jkLtVZ7Cr1xmHApJCr
wvtAoNCifi7/qdiP96O1lXab0q9aeLHP1gNxGQgOPb+35nMzfohc202raFtd6hLY
G0sy2QP1peS4IrxrczluRb/UPMqUTiLI4FhMngCg1YyjwE6V4B0i+yJfLbMhJlc3
vwu3zfKNpPRxDSVeHDMNngstIBIj4tuPkPWPmhV5fsITIICbVR0SSQ1nNsONBqN9
mzBelTf825znGl3CE2mza1Ke9QAWbGaeHH3ivkjWafautYbKpLsHYEziR8aeXXjv
i0NFYRhB+1gk3Ry4eMRh/gSCMrPD5wbrSK8nvzy38/+kYQGmcvPuQdUCtxGgUeQJ
KNMpQUnag22glm6bPOfYkodmSW5qbQLWVvRPHlDdK9Yi19zRij2wpYWnAwA7XMGS
rQsURUBJElufv6604WpppkgtXgnmceTY3AM+eHjcujIIJjZEeFkTcmahThmcMJBY
SWZRNFNAs+QC+nXeAByK6oWaNA1BCBtwPA9120tMasHWwA2UQ6nkLUUfj1KEXDRp
R39ZWgvJg3JIpdKhsp8oCKxUbWIQViP8vmGnOMgKmnIG/PLoJW8Qj2nO+bzWWK1I
x9ZmEooUTKdUpQUIzPL22QsjpmiX30zUvlxu98t/cjbWYOGbPANZAtGj9RS/XDk0
6khM7I9ovwsVcGrd9MeJpWIC6OQJvy6+ZmMbn0GxdjqfkoAVeJg5jS2lZRI9ktdu
qN6G2uWuVrfmw1yWMjMP97ERDdi1WSVWouM6p8sNKa6i2WvDJFivLzWDK+Xa+r3l
3pNXoyuPi5mNZcPYZi0TwAk3bwOVtyqlAaGE9kk/WvnaGursAMhoCniyxoskge1U
mNHdTQPIlXDieA3qP1AG9dfD4FoGiw7KP1peOjxA1kHr1qGaJolK5LoSuhgGe/Vz
fSCMMcxt70+eL7ZThF4N/LJIj1AbiWL14FTJgFYPtXyafkI0j4jAh+RD+DSxciYX
8YFObGAMjX3Kh1O4wBeC6xdqOvmAmJwCkriQH1WrSivPWq6oXDV28sp4iTl6lSv/
0YBVGF518C9yjm7HLVOx0ZYGkmLseGhVAkI3sqMmsNIemGyizMNnP5JVHWCVTIj/
LHLqPUZYNxWL16SgGY80jO8K9MDq3NLu5/WmzHgvncfZD8aEyRSxjcx+MvOakStT
cxQ1tusacFxLZOpMke2slQuNXShtsT49GO8/U3HyN9l/MzYx9GVbJ2LtrxZ8ttu7
mhbQ9ydbKVKr+sjq1CszBfoeCsngC7/3EFYGpXBR1PW+1ytWlCmTkNrML369spu/
Kx+NysLqYTgaM/1qM28MMHT9VuUYrsOB+eDHH96ANYLdnbUr+wCeLtCrrNn5Kheq
uNZvY3ApAvknzA0fDJaWd+H5h/3BQFO7ZEGwQeVLqG+UokzwiMPrl2amDu/vBH1/
LnCuW0U1t9jwdhFU//N+dDK23p+Z2G3DWbVWwQRnvjVXup1rwLijXXyKggS09qtL
cUjcOPJ8U9SUZxLFD671JDX8NyIwmgaEyFSlV2hdhdLq7aM3Ct94/a8hhC5EcUMc
DY+u6HIRpVPmHHY1APbGAPiR+W1WLbINFYBDBt6UN8KJRECk0FOOKeFCDpVd/+hP
r27pA5F/oHCADxfxy6K2BagVI/ULeVwuCQhq0vFiC23szYxmfkLxVBSvKGRCqnBb
3tFdzM84yr2/D6xaYXzcpf4AOHOrKqpz+zsWe0dP/rmjR9b//0/7oMGb0O0FGRBp
l9NLozxyIXr1Yer59BWgsBE6LXMJWA95igizYcHj9dIoK+Zrkq+31ixetkE+a8nu
d5qcMBPPXP9mcAR7ji3HQIZqMCrtYhAZc+75ym8eK8Fvm1wXZ094SK3BZ/d/Js/F
WFKO2ut+xwbuzsENSKaMfTHm4kfC+wyB4dIBmRGR1EiXYR+an6Nk+xrR8HruuwZq
AQ8XSMcM3lLhLV1zDoGxKIT8UkRP9/grypQyACA0cZOQDNrt2P8dLEaPeX5slwdV
YeUD4TQ/N+WCPSNglf1hMzt/uHgJiFnrZQF6EMu+s7LOYiLNY6TJI6vGs8KYkkoq
7eelyFwF3+342PlfqariCkmv2N6PoxX1dKq11QrPyNz9CqqleH4mPP4FlplwsliP
5vMrG9sd8vTWKOg5VFP5FPVGK7jgz+k/tn7L1j0d2gOaDYoYNUPdA3KybucbKlAF
H1tPAsPhHLbS3TL2xLweW0oQ8x1X9u6g5aXDOpd1+Qs+s9Qk016vqW7n94pM1fDG
kPpUs/ZHeEAh7EjBwhKt9yAn4MKmcMIlcs4E8l17++j9GATG4uhfC0JxUuPTQb40
vJJu5wBQFi2weXnGuc3CzwuPRnTXCh4D3n9UNPgHFYVlA26dpJw1h5iBAx1W1iXN
aGMAMO8vpl/FthcxairzQTdrn/tYH9g7rfLYDd7QokmF0GEOb6Lv8uc+3r2mLa9f
J/XbUtu/+4nVD1kOxmfTK0l0Re5apn/r9GDTN7oGzV0E3uiLlGZc6ZJuu8YbMgTF
KRI2omQhQNMjBtGWDvHmLr8+2QarCdDY4+L3CTt83x+D4nKCpTqGBGYrsGXBNL5Q
EmDUgUTJS++jt+gywss/w+7HXwzvVqZqscDDPfJOOQvhu7FICLnLQoMzb8iRxRWk
CvACwHCgPfQAr/U3IWQcyNWrU+U6hBykm9LH4+pYYazt9Bwj1jNC9EyVqyv9C3qE
wIVGNhcU4um6IZCxbfiVXIF/JMoAahKeg66/HNJrqTAyN9Gi4YtNTXmsUNBEDFHB
U1awPOGrWrhdAvpFBKdDQSVH0Uww03jwNU8zjHBm+DyyBB4QmV0r0jwNU2ChD49y
L1A4H3ibBOSJA52h1WRYTYY+B9daDaFMcSmuBFk+sbezh/J/4d4tTy5KWOiny42o
94FdXB9vDepf+/K628SwMtoZMNOELRLcHtFgIzx/yXifpoFTaqny43tZO11+Tc4s
qfVJHpRcj2meciB+hqZREqWwUaHwBgieGiSAkTiDuRnZz72t66DfLjJ66L6OBe0V
VKFyqn5jjMGK4elDDUmD+kOcupwdjG6fBxJAIPGev2vEczHSfn7eaJT1zG/mql3Y
FsgLZkW6tVQbB+pSZ62YMHoJCyucskTSpw1sKdgJ4ZFCnWmZqiqC5njs3F7F0wRT
GyFegGrGgilWRBW0HUgXSfm1QB3QzpXsXvhhYlTdZFbtrJYAXs7BBMka0x9TpB4y
XH1bliOeN95JITnv1wIOkVOe90N/XW3QdwaSLYgfIOSKxDSAeejchixb1IPWF8Ho
gg3ecqNT3TFQV6/EwHvLu0RzBNX/lUpBSFRk1J7QUA5/OmLoK/7IErR5midMbpDH
ajFnzNal+Tw8/3wGjnwsLScqQszV1aoF5lF1IC3ZpC8Jm6v3lFW9OT6BHA4lhNsb
wvKgZ5E0Lq8a6Z42DwWwTfbb1VDE4k2BOVHmPBN5yT097mpMiPP5zaVNdKQ74VQ/
iOgn9WTotdFpsjB8dIoEdkxt2YGCodP1Oct9KxJbQIHodU8gNzOib38Jj2Ks5K04
oLTvwvfAdROgTX/Wbut6LS3t88SSTTx+rB6CEwTxdXfw16Ke5tIAbbpd0Bz5qmD+
B16i+olb1XFAq/2j+hKU0ZuUVZfnlBwiV8Upi9O8PKc+qLIyuF2T61lr12sntqx9
AYnN2Nnl7b7D753+L4uUG436hK1CQ1mcv7I7V/01uixqE97t+EZgsx4L/hS5xxum
xDhcm4fFzNMn+scdulLJMql4b9CiQFv81JrRiuA9Dmdk9JSD+ENhVUbF4ULlCTjG
47jQqt2zhQ3rUymKbs1ZzFA3xfNuOFwGpBzsk2EdzM6MxaWSmFCPHsAF6GCRsJ51
3SWeRZ9qqjZ/cJCDcYjyNAuCSyvD0hjlHbCaKcUv4eC7VkhDN/rHhX8fwJYL8HMy
yi3YhhTlG0W/skDxKTxdxtzGA5ex9INCsU2OEFgz1T15ImfF7m1fgZV8gnpsfBZc
0oFOLVBEIRL5L6dOGZioTE/Rpku6dDn9PVLeIxsUlB7E8RYeG0XeMxBEAm706uVL
Ff7TUZh7kcweqX3UR9SLyAV74KR7PBddIe9bE3cmsAmACtka0AfxiSt2PdYtNk3a
5BkShgbF/M5uasNQfdYvq2v1o5LheS8OBW8LmtNBPIFtw1cKviCRrKvc32i/yV14
729NEaUnhIM2nBT6HEyYI9/WoKoBGmmpGllzMe9U00tMFWy43DLLU17F4ycPhdGN
viUNmPTkRiDFTywdFQYy4krMZ0qhxXtaQPbmQ5tbZfWO3mxGcU84wxmmWN/p0Swh
EAB8dGEBDgWnKs685I86Lj69uMrf1LuLGSXixQJY03AITrcyRu1+A0J87J5QfBVf
vdvWFYAQTeUAgrF/sWPs6pNkSgXSoyBUJbmQcjmq9pHFds6RRgvE6mXZs0yJR/Gm
396/RhzMKp/OjCDqTfAzJvG9jH58IB5OkfTM/f4LLaWNT4jJ+OvTaj2aceU8qL6s
QCWvxCQk6hXWxoowkfl5Sv5MJ3lXPG3DDXUvUNg0wC8TtsTg4wDyR1nRf+9cduWU
ghfRe/rmBndH6pVqphXx0hkwKwtDzhsJCASVcwbDibZAhGoEz6bPjvCOg7aOh4UI
V8xhNsUbx/uhXx7vdrdHrS37PnCdIuPT/f84+8ca7nEyOQpGADabQaAEMHRcNDZG
NrwNL0qQeHGlkK6jGYx+t5KyphQ+3jUhLnZfu4JR2kN+RDWJsPoDVqFhyj/o2x2v
Cd19GSMOgMH/2ZW8zOqEq6Ph6rRexmc9Par3HziXGaOXBbwTHfr/VBz6poIWteCr
UYCSJ9kNYG+mJi98X42qTRNZVK3hCWNyqkPN+AijhrkqR09ye4/9YkO1Q/05N0/c
n0qQnLWejt+XDd9/03TmymxpVZP2Ql2gGU16jdBjgo85gRwm3gxjr7/eHgzPscWH
drxJQ4VSOUG9yneWWJwR2rNoih9IXFzP2p/cyYtdxbSvUslMnX64wAPGvbhIuFsz
KlNYt2IG4CWWF+WlgA3AeemtkMxxkXh8WbZZ071f3OPvBDJDjZJ/b1WxAp2DxkzD
NYg77Jvm5tA7Tr2EZvGH0K+A+ExZRuKGwxFnu4kbxzrvY0XqUqplLKJeOWB7dgfE
iMMh0j7Y9RtjhNFWcgfOAcri9G6jMjQfUVr8fs2PaJSmP6K/K4QLVsluQjYfUJVW
vhPBdwMBHu+mA9FBMqlAvyiopEaOlwbQ1BtFD1fu5S7fvl7mW2qyLmHc/FR+cw6A
ctW5hXAMSzTGSj8UP9wYO7s99oQyhwGVzf96tJ0jhqkLd82Zgle1GBxRXEWtmz2U
lPLTxNNBGG8Zot11gvhMTzk066VZOTSslynDbqR9FfKu3W50n/FeVVDKG/4VEHll
vLn2Bcztde5QRhqN5nN8nQdvrtRqPNaza+mlbupAE4NHK1dAsOr15MVwEGptUwOH
L/oOsUZf33fxP7FJtMbayjJBzDnkyPGrlPv7HiP/S9/VlJcLvVaO7HrK1RDuvsr+
pW/tYNb24j2AdjwE7zykAU4xXnU0YZg5QlXjL+YwibsL3Ry24Qyq4V3+GAf6kESR
RPCGgZgBwMBj/CvQyRXaGZgT5DtzfAvFBOXWCFSI8bhNmjv8bjFsUM2eAVqMGwS5
LhkKwqKhHAFz1QLXrK9fByT5FD+ZmOQUG8sXWi7GL2hWhIogYA8wlXOyuwE4xUJM
pyZljbpLOeBbUnaxb31Mf/WBuYAXIIZlVYkx+lC/vPUpbqWfjr2TtJQ9DUC5hOCN
6lui+t7v0/42JVVEm5UIBwi8QbcpgRAGTAAXmV3RwZMkpM88aAQ9xNUdrgS3mOtD
ZggX96ZhN+QMXJZocfsICSgesTH9btXVmofmSRdgMJYDNyp1mRtMJizpkuFhUU0d
yUdsNODD7VmATcEm/96kRYzWLj19V0ZD6kMjaPrPgQUitTFv5vBGb3rxsrGuPr3V
UqTR+g0lQ5paPhBlB18n4dTMRv8QghPaOti7zpd9CPwJqscd4k+OWLLRwIsPJMzx
IOg8DMU98eRFMZ/41D9e/LuJ+4OQyM2rNBhpxoixrKAs4wR2nv4Th3K/e3WO4xbU
SqjAf5N3SHL7UGE+9Die1DHm+5bOZSv+MtTeahkEnl2nkhOOW6HXxQBTYI0yw9LH
CvJrzW30S4433b5l1El4fOhsdrWKpJdAm9y04M2NM8X8PFWQeskBpMRyiTSZjqtZ
bRUuG3ANFLTyhL2enTKb8A8Nf0mgA7GOTzFaA9NwG5YfE0bYCrH1juIHLvvlnv5Q
fYguXvooYyQKqBGTp1eCcqdMDjlX7jhzPVDDk9Sy95N2NWx1gE/SEG22s0XFsuy7
QXJC3DKc7gY4+filQiGzMl8sejFG6iT7jjs3sIKFfJspZJs4DoYxB3/QtlJETk1P
Q3sWx0CrLgbavEwEGlFmPznN5MVaXyMsoQ1ZbWHfHw+90ktTB8cZELy2EE299+Sz
BsysM1GInr4CnQRohDrkdulNZNBxBJYVRSbkbLhFIYJCgAY+taXebVDBKOvKPfas
fO0Blf9DR9ute4t62FCcYWCqQ4400V5X7QPEzk8oo0NT+pVfwXZomERY616n1rK7
/5og9ffvwT+uouSZsDUiBnG//9dyk6l0owFGylt7sHm81emzdzxI4ZIsli5LqEDl
nzrRl8NVc3GO5cz6ACm1+uDNcAmbixgfYTRdFNDjcTmOamK6t3a7qjU1iblqa/yj
7NbfUEpGzxm7Z3TnUfzoOAQxFkWQ2sjK8X63IJsqMnNRo5tTf82MhJecr0D0vQAN
kP7KrivdEDSS8Kzt7QbcbT6Te+mmgtjja4IIMCLwXuCG6cpSrjk+TLo1sUY75X11
K/v4V8q9olw4XBzfyLXa3xx3lDtGZs1M/l5G5GRTsvM1hBRMe2jsRXtNSI1Qi8I3
r8Fh1mJ652qRSYGmC1Rb4qtazXR30XIFotQt21nkoBSmKFSa61Gd0h5TieRLGo9T
eyQ7d7RRBOnp5Rn2hR8lLHFldvE+mfhizAhGImdc8jJZ/H70DmqOtJUwWw6JiqPV
uSR0rkzWPW5zvha+XvSdqYcDXdqEaFgXa8kC9zmJ62CHrzaOMWAtftivQ0CHqghw
SwuLkwRWM5DxDQQr2Ua7XOlHvP9YIcxhhc6cpbgbHPZB8sLJzejuTI/iXlHE0/05
XxuhM02i6VoGHpGAsqKD564vHXZq71+sTmf9fXqpUfPJVcqp7B0BRDM0ScqJOV6W
48z+clamn3Vs1fkaIcKcf+Mu8L+zOMV4bMojzvydVsgYZIUJ2qWql1hKcCOp2r4M
0etcWY5SGBrHEtZznQ1bZwwBZ14SUd9f8vYxih+E9z/K9LLNtEgTHRkQe9LXDvkH
ouvbtrwsBudfU3ARBcMtEWn3+k7RT9YMjoHnWnkOOmd0sUnnU6fURi4ue7obxFJj
I+8C/gqgIOsU1GVJlUy35ImUYLf/ncQlujxf7Z74/V86yzX6/NAxPKZG5pNK7vuM
1KT+GVdWe+Yq/iRux8eL874W5i2dUmrTe1YIWX9i2+RGZyiNIFN/K9lBI7vZygmg
BAnydL/d72CpgbyAMFNwLlMMLxevw+4w/xV1+dGtDcqch0OeJyZM75Ui8Tf/7RSj
IP8urgKqH7xsts8rnS0HrlSCMSlXpa1c/4uyhIDkOzaJMWiCq0sMksHakCQNhr9w
0xpttuPfmS5V3eIhG90TpOWr84Rf/8Y7G5ZUyJyDT/D6d3JyRRP16d2n4wdRZ2Ub
IS7WkeJNt6szLf/fQymDdBzOCk7gmF3B7qhwcjdcuHKdBNyX1GqHe/Vg4p/ksQcT
4Fo2YhffI4UJ9DgptR32ap4hTQ2ajBwDRqOi9SbAf5rHXoYFLZchbt6AL3sWHk4u
7yK76wMmJjPoKSnJ7QYL/XMT/N21o4CLhX8kNdvYeeJpwznqDGoFEiL7rq+4mJ/n
yoQ/xiWAifbMv2je/QYDfBGVVUjyXFbKyMnK6ZoxiwpN+gEByI7L0czWpZ200TFQ
BYsWs8AWD2f0+5ylifmEt574eOhMcL9kg46Wg2uXqihJZHwcsutipu+0kPmhCCWj
CRfEkzDMDn2PyunS4XCfczfEBJFVOlaldIomrXS9kD5IogusKQ57S7gsyGyt5gnz
F2qFeX9We12r9nlmpp9vr7B7FZhjcM5goMPu5cXpTPbpGFxmo7zky+Zf2fykVAUs
IUTaNQtNs54Qjril/UgCPKPqURUbSA/VYdLtKMDbDVdPjZBnI9gaHsyRX3THfw83
P2smKXMEw+NKxMznRMSE4wxkUUarFIdnKMdgy26RfXK9XmLU3o+g0XqQ8UKKPXff
DkaXxb6qrCO5RdTWYbuaRGGrmrNumDpTyvNrPgofpPYbdnEtCJ0PEd7PHo+zArdH
JlJqYohrbNXrvYWAUgkNUtzzGZctxqmVXiuW5gqEKZ9Jpc7hUZ4IJTVe9d1xLa6I
iQ0R6PnGlmzhrFZohjeevjn8k/BSlVSPDz4ANo7xI+rsDvpMC9R3qvDJJThRT+4a
mHcyNz2JqbkYHKeW+8ZVFg5H1JFrclSrCRp7sJc5bQmdYm/SHk8aNuIqcO20fDDG
EsyZYFzZDdS3fP81jBe5T6BNicqlTfK68l5JQV7D88DS4V591VcQ7c/QUz+0k1Vt
uuTbVGuu9xLuEHkLiWkIcQr80h4tEukWgFUJZ7sLu+qGkuTbtfjPmso0PAWWkRaq
M4WOFmhvWqmWjwY6yxPOeKECeYQ0gojrYqMOrcWpPF2BvSIqPO+nr35D5/+rbrwI
97BJt3rEPZkVXsiX1t0Kwj5BP2CXDvnJrr3YcK4CtfnWyw0VNoy1r9Gfv4UfRfYc
A0obiyRDULcdDrfjXyCnGA8pCmCGqLy9LFSw8rW98ngAn1+JDdM1r+ye8/76sVqY
1eAwYfWUsLzOLgmz5ol19SmJe1RPvTIcyeA3no1P8KxnbbJRXDRLKHFSG72twTNm
C3rv+fXflHqtqzIwfIH1nWH7uVECa67oSRgCnQFs12v0TgmbB8PVXVQRDeiL+U+C
IDGJKa/LTY1tnhhjQcXaJwyyeoRIDvb1a391seTqtZvhSidV3d0sPWSeXXlHI9WS
V0w4ikxKxD0i6XU7qKqmcI99zY2AT2uGCL2wrz0ZjVKzf4MBmRhgD1CxqAbCHEIF
T4V7EmKic2AJPr0xmFFRJPFPu200sTMbpGEKOiYelAEZi5Z01fWCZlfx6d0XdE82
K2VMDLqVot6GbePdr6wgQwMQDcu79zc2gwZSb2Wdq3b9ezT3/MLvG2pC4db8ltQX
+lPpzPOKq4gpqlTcb+mLqMbDcqD9fBkslNSCfZ9NHxN4ZI4y08iRN2W5rBPB8PsR
5cAXaTaPQfJsi42+oSDs99ez7mXWDFr1t8ReT9zDlzcKhm44KyBZNQ0QlTwGzmCA
/pvXrQX1hfnrJqmsg9WGZd7L+bZYqIYOfOOrsaqAS0MonnHfBGj5YZav6fGy8YKo
lCxilEf6cRaGcIhZD1KapwBV7KDsGjfjQXRaZRyNfZIGljP3GUjWelXNm+5P5a6d
tFPePDEh5YfyLAIAX0LIFTfRN20wcUMYkeJTj+wzreHr0LY9TIw7ZcJ+PtwlrF17
9phPmYfV0mWGg2AjhBKkvdtzePUmGwrj6Wa3MJkKQ8x+fywJCkLJSbKzNbkZlyLE
wxo+9GLEU29rVu1GKxT/R34nzs+/f8wa+m1jYwGlO/IJvF/gt0eGQ6iiFVS4qYOY
1eKjD4X3Q1hPT6dmedGH5dxFWd/Y0i47gt7gwd1Z5HpEmsw0Ut7i+V/x8JTXwxD5
aYInOSFRzcAWJY7SO0Z7QutIQGv7omffZtCjfVIKO77d/gLD5Kf20Wguq1EGBtNd
onR8ikd0wjldaJhgph8wBMT9S718jyhLdbK3gGSkvE1Gleol+QRIcw7pj/ZdgFd3
oxusd2mZ+/J8KqZlJu2NSJ6HCJJo8Q/KepKJKwk3MEtjAryN1iF/9ZoRS2c7oG9+
3nbCXHMmETxqwIOU/2G7xwhSz+PmaQqQhLN7EmHJ2VFWuvS1AZwpU2OkDuqIzFIY
msYkMxik3SuuAzK+PqSXXjzKJC6oqNOzkRPrgKTdI8nlNc5oRCfcnPkirpS3O8o/
1ajryjnLP/29lPz6593e5PrlXC7mH3k601j8DeK/9rzyki7NcZgI9nq1hXlxI1zr
Hv8ndFMqx0x793rikPjpJOVA7eimWXWgTtOPjt8Y1FSARDs1/6X/y8hcbmOfHGxE
tcD1WZZrkHQK39rCRF1b9/1KfXdQzRWdtWu+GMcabG0yHbH4Clw6suR0ehfdqwrW
zmwWS+Wa0g0bgdBcxPG/zPYqyclXWZ5xGRn25foCdeFxbMeoqsluK3nsi2tAw7Fq
1ZCRR43YzZfcCuTF8bmq322FJSdZNaZ4gzZNuKWp1HJM4MFIZeTsWIR0VccKR100
WRgZuGV7cgEirf2zHgaAaNpjbtqSg4uhtLElV/SWAADl8Fmbue3HBorVNsBq3DCX
DDr/VWqPA8uYe6RY7LzJ1xN1tSbWOg4CiYDVCEbcJLHnCNXHGcdpn+mckRzLP0Zy
7XFpNQq0JR5lh+dGRd3o4Hw9X47sn5TtfHWPMFBvwKmFoC/k3p19LAOopjr+0+OS
RZFBASX3DVejzpur7ys/Fw5elZ70hs1kXldpYUrV0bv/EsqOrIKMcJ8YxCDkWU6i
dV2vpVcTx7qiuATpSLvwb5WiuKccFbFFtYagoJTvc0YpH+jcmRRFoDk/3GSKYQic
b9SAEb3wKb+6DVEDV7F8S1+oJOFrb7pOgNqKwk0ssf30iw+hHoUkM/wtKA7858o7
+HMJKPivkkqvyUqPGvsXayz3OJai7iRb5T0uSgVhX9LSFbLWnyKSXDtfVKN+58XN
JKgd1dVm975xEvaeyjrDuOkMqVIkx/vDYS3q6IpjKe+sPpH4qA6Gbb8b96I8lGfQ
3sQ67eRLbA+Ex6NDetr8YYImGMCWnGyOtVocWBhcINBUYZBiTedg2YHt1GfhJeyH
CnM88UrhGn3a1sYGKVPqKy7mRdyjGBVwjjjuSqa+72pikiwT9zeGJXoXe/LX7wat
btNWJv1q6/4y/kwg2bCuoMP2y2H6CKMbiOMzK5I2fIhkBi5j4bWJem6BIRzEwkFS
SvR0oXoM6cdUKHV6aDCNi7pp7iUWktBkENBhgklYOwZpNrkYaAJ67VnPI/fXjIV9
1cD+Wk62eUB2R3g3rMKs2u3NeJav2xcKowthS0+SBr39CQE/Vx/G30mY7HHAMi3G
eberk5xs2mQvkmv1SRFBuY7hwEQ9AeBaYABakaDcJXSZ0AX0dEuau0d1KTI7alsX
wNjdYTRgQDihs3MYrHjWMQVN15z0tRuDZzkgi10s39AY3rOA1Xz6ctF+/OSJoLCh
fd6XWVCdfUHLPhWPp9dS5IyQjDoNiI4jmuO5m32/ryu3r/IvOZRh95z69HzQXlfa
xqoHAxU2XR8AmRGpWeHXs97ch2kchkwlI8UqRxiiwmHHFkGuPG6UslmiTZojkPzo
3zhe+7JwCwtBLwSPmn80pxia4eiFizuLHytClgvGOf4GtIXTkKDWS9OIU7rggu7M
RVaFY8hsZhgsQT2WYL99BFN1ON5gjhRtbMl5ox8SrSgXtTm++ZqGtMEDQDaQoazK
X3ijduuWLtChVs3sY0MTESVXIsUc+8Ay3kJb9H8z2BIvHATMfYHClsk9sr/GjhBq
5ybMfnLoc1Q8gv9nJGYT/1iRjxPw+71D5fAYuvY7TE4hFfIWhvcJt49fQ2AZ/vOs
qINY/trASgfGXb0dfpWu2JdzxhJy7K1j8iMaL7MBV/KWKdnIVYWcXUXdvwJnlqhj
IgZWb8xLY7E1aObaauUyRRnVvrG7+bLMmtplnuV5aeHQurroSVrdjGkS1ONcoFf6
ATSpOk2GUGCHBgycwggpL05HEK7ZHfLAXjWpg0ExZ0oc+yQ4Hy37Ud7rY9zdX6iU
l/KEFrRMZkC0d+V2sIALC2QrVxNnAwC9w83f871dbLMKZSt50gj6wrBRo+UrEZPZ
yMVsigqm+AL5RChqzxTncPkVmz5dZLOl3XFjsBqhgbP9zjyW727vRQwLxv1m6qIU
bfAtuCuhrwKLkfCR3tFQ3PUljNH8vXjkrM916WjHmCstZyjnpduQ8TboaT36FEfO
JCp8keo8W1JJtOPTALqMiUYYYrdNpmTFnHT5wtquX5xSXqxhH6j5HH437u623L+B
m9zhaKwcK3pGipHHcK14UYkI/NPdYuOzySI9LrYDCkGooS65IamwN/xo4oj7xegx
sOTOFAaobPto5GH4DupcUMaIac7G8WxmyS2TKPo1rYy62jq/tZTfMUNtcjR61Cht
CTccpYy+p7JjRrSYmrBFFDLsAA17rIDaGAGckm8SDrq2rDne1mItLaz+UPAsaQq6
i+x4kfvjLoh91y/zZvUQLXhhTarsbMpSlWRjyOqCuZStwdrLEVKa/TNROU4EbjxN
pcV2TfVlMjBwem6mMCPpB+FfOfycONzILdMZ4QJf4HUInKniaPODDeKDR0Tfcu01
KZxO1a8f+mqDajvjQ1tbBa3ir0DO8OyqVi7UDZH8+4FO8SLs7fw0RD5tHrHe1Jz4
Uta53bi7qjQQZN+af4Bmcb+/O3hQG+Pdns1hz1O0AX9X8wQ32iLkxs56o2Lp/Yf0
33+jvT8OpumJAUCxMizV+s6Kk+V+MLdLGBeRca54M2DzFRN52NeVh6N5Vrew4uoT
O4+RncLDXdegSELT7cDYoP44/bdijRX5mDhxE+usCZfBY7xhi29Gc8xbZmCWup/S
9oXcMNA4gZ3fWZKBD5iHRXyrwyHa1UeC7cGZ9s3ofQ7YqfoN3gFGYQUkWSS1LDUW
NkkqXFOylTgRC8yfnQ3YaDM6awfMTCfeM+xXd4l+7oYyM9O6PvRHU9tTgnXPBtrA
n5w/+Rmwpdg3JgD5ndrVtWgL5IUwjNBiWUynYO4eMheI2cF/oZDvFv0Cdcmr3DTu
0cA3Q3g3Uh1ZYrIqQrGyCvWOMdzey3+guD5V9sj51wCPHDzSJ8kixeO8a8pQ+Gq/
aaIMkNvT3bXu8qEDwMqllo3IdtcDWTxeqQSLCZPgp6izdH9sa/9adARsnOCsNQVv
Hq+BECkiUJTZj2MdqXTiidCLBVEohTPGRa17q4//yKrcv20p4ibphjUN84zaxE8d
oyRwbYpUdY6gmsCXZwJUIqHQD26xD0/nM8Z9lnpTZMgabPnbKKsS7pF5EjsJoe6y
cOzb9UWsC1CC7aIgee/ZuvLUxQtKW6fs6MUvhAgtJvTRlXYB+OSM5RJ0uyhZzELj
bfT6sZLTtvqc7iAaBmObWHkhj2BAbkbHsNeAkiyFcjaY2viluqKIaB6ZYbQEJLDs
iRuCYJlc83Nug5bDU5Iin8RGAcNu+OCAguDliyrxUPADBF05A9Taw8tQT19KPpX4
VVjeL5nnhDcUkciweBUzJWKHyGYv5+2sohS9p3YLlube/0zet8rETB6JqopZXowk
YBwUTJ0EAFBsAUKdRj97jbNgovDwFbChcxtzdeMTwfZF3as15sqAe7rJ2XOvO2zB
/WZ7J492i17j6+MOH+QM+S3A8DxTg9yu/2UmSK5/xWooz6oev4kzlH72iZDXs8ke
STTxNNba4d/0S6U9VFROrwTH+eTFeKWmjlypoeurwFKNSYoBnCBytwoimuRmi0A2
CiK+T+OZ6nUr4KCA73OXs9iuGgjN6b812SkTYL2Q+bHsSQWJ9jRvLoZf46MWR7Lm
Zi7Iqx0+eqPdBdPESvvYhZ5L5nCnzpRVB7fc5pznZ+Pm4EtndcVtqy1vCaCm5j2I
kzUTHjjHXe7fU1hzbpQQVaHfHW/504NbOmtJe7hRcfJq5OSLLk4LQ8ZKuhtUwwbc
75CsYTNgent0xDF+fm/SezOs1CzUl4Blv8yXpn2o6AjusaPL1Rr5bpM1dwg/a+5x
QmDfMzTCJ2zpiAkxGf8FkAzeTgoQqwQkw8BpMeDMeWWn+U+yV5Z/7/UI2m2jfF42
vUTveyiT6umW6wv45FnXRUyNB2JfgpcvVEWOQmmWANGqEDSGg1IikX84mb/4ColY
jm+KwaJYCF8sP8Kdd6f0b1znT5/E/7hWHTKVNVxELs4r1xl/BUt0WIv1mDpr/6aK
wu4Rycg2E0rMM2iKKlRlpJsh3WALiF73lKKcfFmbaV7dDqjCbMOr31zi4IVLmJ50
jAptPGmxEEnm6Wp59L8cr01tAHwJyjYcp+aJUh5nPuVbphtniCBDtrktLWKqZHDT
n5MkXQYhTCkCj40egkTrsUxCsC7rrPlOxrHMo4TzJxz95yvp2xElRyPHmj+COgkO
RovTBLlfdWAcKUR93NdbtxmdJnWt97JsTpKxQN030lGrv0S04HPWgdEJ/TNZU85u
sFFuuE5V3NSRovoL1d6BOOu/l2EMnZxv1g+lcWuPNygZmJXB/DPrMvp5oirwqM3e
+hA9CPMkB/VHu7PeWYK24c8G6nrQtI8hSYtzhGx+HVC3TpuWeeTBiegAzjhonMuk
mNgDpYrr8854UsV/CV8u5qm1hwWsYhWY7UsOQYlUuRf7fJFv742iRr/UfZDDyHj5
7C5hjqotTSuvX+31L0R6O/Sk71CFqBlAweidx7IEHCCE52NatsFomNcAuyrRQIoW
9oZSRPux9QPckAXIf+XRd2vq8qHuqFZVKodpOIFN1rlPVKlxZNOihcOvfWA2ELax
xn478dDxXuHAEgXn53UvBc3va/nWVhgEYg32blQcSbIA6YNiqWK8F1UKMb1O9lkd
UiGylRkXXIWCsYDuiCp2qF8rraYXdlETS6GwswAXHzno4CPMyDtUTTYRKpUxvF/D
Hy/ydz2VA3e8469JO/koMBHf60vuwiDPiBuXXHJy6bvGojh5zcykJm8c1DqpYcMg
G5PLjysZMjMFFrE2vxQDzvLyVmvQd7vg6i8YEkT222pNYqL1FcLC6L1BxErJ0Tee
7l+sjjjk943SukwDKeahZUNsf+j2xsyWUjRoxZX5gE5uB8+wVcvSW2jKBm6meY2e
TKZE31CDRLUPij9/RA9w7Ul5BklIgdl/XAhM6AbkFVI/yCtNQ7sWXjIX8j1C5cl5
Okfau+fCRTi7EV2+LeFShbgbbUwySfwFWm0Fnj4BoDvwSui+8OtuBcwsIQN+Yp/f
6IirPBKJyxo0tga0X+0arRyojo9+zrSxJW1Lakv206wu5zZ5hoby3JOEQUJ/fEsb
2+sN6n5h+theHapggUY//Ay8NQG7ZC9v7CBLUTtspE0RpBPo3r9KXryL0xCcKT3t
Toz/oebHi5HZBBkZHHqnlug53HHtdsiL7Oue7WLQ4Cjn023ZXDi8XMxt8o7a5CuL
m6WTe9Z/v1lB8E5r11hjlsV38+meBEIASIn3tWO12XcAUBcNKD9sSO3DQCVkieH9
ENMUNY1PDa1S/nIgO/J4T0KnCDaQVmR4ilbKanFo1z4Vr3qSAC9xrXdzCKpVcIiu
XmeuSD7iKF4C16tKzgu85VtmrquTFZczSkgViNygSCy0jU7TqRRhwdQzvEAd7Ug3
TeH/4/1KCryOA1s66TYLw8kCBl8fAzZCVfz06+cigSTHANCETKHIGI+jnu38a4VX
z6Z8CwW2JOHlMGtHJct2PDcd7Zd0dzHy2sxoLtwqhWxU6MdahdfMnXY3DwuCCFjy
p+uazVFOR4GkZUxLBfWfS5etOGkLNXv9u+FAYC89hH++EQS1O8fFT3F3nBzXZpE8
1ipNwZl0X2erx+Z8vF2/xx2d7z6p+osoL2vVK+NH943s9367hNOSEr4cnr46x4Jy
70cHzVwWDsmPucRU3fxiF83layh4ImGkkkZHcIrgKt8k89fN7of4H3A6GUe3DYjU
SVd8rHmwyRMQfvPK3vgfbTfB53TZ04cY6CovDfpjIr1UtGx4Yp29M6OHYwYc6ks7
2LxGjG2bNcTWuTBML6EQAYYorcSSxOakIuT6bzsSox781jy1ozMXhFhVT/8p7lw3
OK0Za755AEh+p9WgQfqAsBuxT9m8iYHVxEvyX6HP5P0geAG0Nh4Wtddmsv/D1t/d
UUwJCE0aSqcm4t5RXS9PccbCYtPczM8IEFq+XtJEe7ySeL0pneIW2vZE00LsMU8O
WATjUtbcNOWwSgqkOCf7rVvOqyJclB99nhg7YhTFCCZQDvbRP4x+MpzWko4f2gQS
9M9HzVnGf5dR/4YsydZnvQzaryVsvlo308UmWRj/3P+HboH34X5D+nNsWEzvzMtv
9344CfHQJPF4YU4FsJPbvlY7ypwHhSIZwr1pZe6Y9oSQDQ3np86JzQUPsn4e/wnN
6NqsAch8/42u3ekj9zL6UDohfliEXjdjuVXU0tFmVJL5WRu/rT+R7HGChjO2h2vT
tQ4J6uVVvYE/fhSw0DqmrCxdj4EGIXlxpZoxAYTszy1FsruOIsYCviLBncR3MXRC
D0lhnHeJjuGFCOl7YRJUXV4+lanZFRtO5NY5+a+F3TL5ln8Bec2nAxWTdO/WZPtb
DjbeLwlfcqbm6GRsbTwF6J8QTQehUhlKn5eEHJcm297sW8t7fanGEKFPUI6n60+8
PRCQ21W+4MMiZOGkD31hv5Cjjq7v1AeWaGPsGAl6llzSWQMge142nJ74IYV68lSK
Q1KHVfhqfVOM92iEXulj6Wd8LK2m2IFHoZIRj1/bUgIuM/Po8pT+m5g2Lj4N3MUH
cbVr+8HSmQifIf7S1J7nct7pWfEh8436yEbLmyXMzV0cIMxMXe4x79f5X/R3NsKt
9FzA5QTUzw8YyOTFe7c9Yjr9GEo5aaJZnbILZeAryBvdgnKkQ6BYaw4dbU85qVMG
Y+Dm/YjQBJq21H/DUarSZsrRXHbJDtqAtWQF2cwm3YpeLLkkOZkIXexiSZYRaNhb
hmWpxezCNUylgOjAxbtaUG9Z5U33KgiuYBS0IP+ZSxeXh8aB/ep9pT4k3HWiQH//
35fyP2IM6I6myi5xvSC8b4xqXVXCKP2MYhjoVARcSqBrhoV+O3QK3VsTtGEoymDx
QcKoskMucl08tfvvGkPezu0IhixM9yHTbw2/QeCVZ7WZoYbODmUJ9hCgaFxjXBdu
qWdKs8OLSaU/6mCrHlE0ECd7k/DOaneMYfcCpUrBydBEf8Uxqznxnqg41gzLAp/b
+uC8x3ARSYqfSkHC6x3FuAt4Xavlbjo1bqefBkAIvZIYM/AmwoQxDXFYKMzjyXrP
0A40lBJFrg7txreMw8o9Xs8Fv3juu724HLCaY59xzk9sLa/UU7ix6u4Mp2aTsrR9
LPQwps5Mh03BEJAecpD9qemYe5swhByJawTmw+BFDmiF2F/sws00AfX9yQ//EDwz
PdLAvAh+LTQpc9d3EXKJr3QDZFb2sFo/mDQP4hxbIQUnYun3E2Jsc0ZbB8qx+29g
bxhD2mY4zuhTCyk5/5ugCgoEM1nJw8SctpCr7zCmt839JnI3NnrbL4BP+1fNMsUE
WuoY/3fDkH/VfFivKRiXpL9FkGevPEPaRJnnf48djQ24GV75ZrezBxgLeMrZzUFt
4aIdJ3bktUAaA+NR5ke6a9crj/s7TX1lIefW9xbOATgy+mvBeJSQ6VqzYpfFQHUI
LnQVVL4T7o9z8vvP0Q1FkECizvb1dA/gh4Vl7q1VHdQt0mFvRp5X9j5nd4wrABUS
jXr74Kxh1n3vR9jmT86o2nQIJeLwnE3FoXqKRxzIXGn29/zfdCpTjqjJRFB878DP
3TFaiPX0xZvDO3CDP84rTgrontJZn5dQJJli44DJpZbD9P9lc5oXSvJjtNjBJfle
kuxKyVRPoJioKfx5iqGYRifHdivFBvyOEwQDWY/XJ5y0kxNwTLRoBnasofrGbiHE
xTlReWYPdjx8h6QWnK6nsMkGVJJka5Yr2mhNRPs+TmgyS7Gh1i0OiLd8/xFul6cx
7W3ZrQssw3usLvfJhhioIbazzGECK6Txku9jR/rPa9QWBD4OKXyenpbTpBKd1wCz
NueztrZcmTf8rR+gx2nxpFDlsNlqwt7IwbXkb7YsGRxVtCVW8NGDTYkb6FQhIoQ1
w5/pep/rq5vp2gzkne44Qp2ZBz/o1/1Wl178ZIp1vxAdyHjmqqHbwhvnPOxjUBe/
llGRQNdWA2+RjPDKRAjcc55nRoJ+pzxAy6XpphnY5RjK6QOM54QBw2PVuo6BSNJ2
wUiULKWRiWgSPBemlITuHtqEcJXAVyU5pF9tn9LoWRDbgQxwxac4ClS67xCep873
0hIdAeUER79+G9sPi0asKWvQhdT2iBKauhDGrz1/LaHhFBaVrhdcJ/NQkaBuBQAL
d1Iy6jK2bpluQFJHpj3V4J4p2VyjXFXmVbEY8GJCaFRNsIc4pfBYOL2zHwOXLzbL
nXyuvAU4i3mVgI01IvvL1jfZpQj42uRsP2ZVqtv9jtUCf6Milg3Cb6vy138tvO4j
AX1VbSXLj++IKuGoa9dO9dgwhX63guxD/CKrXt7+16hee9jBKjfsjnGSZpcEjtB/
OoduYIO1TZMkDYI3EKIqqGOW4fyBN+jUf0wzcaeqOEvyRZgv/HmQ0g51tBMSnlAL
wL1FML6lh3ckn9NWqzKc30ski2/xr0XaZU12ws0LzlFmtWVl9GQ7GwPrNVP9HOWp
vPK/C7I16Fy42HGzdUisaFB63S5FWJgJDx4cd2opM5QwLmMW5pipZKTLn5d5MUs9
vxYLMc5IUzmdymZ5nkaLm/U2bOFeBdaX6FAnsT/zxq7bf+aS+kmBqjPnyhRptiMP
UO5jeMGAXS9Q8UCtftt7QjVa8QPvaJtKTMbJ1WmPS6+dgXuJ3mWX2jumi2Ntqfnr
25udW8P8GH+QYYGhi7sP26xHRi7LwjKC3dbbqrL4yBuZn7fxM+ggQYrTf6tVzOBs
lxbhEoVYX5LpSBI3kpMczgHRDXpK6Wl+tqLazR3bfp/odhtFCRHTRn1tDL6+ttdP
0lxLYvdJkp49I01h9dTY46L7wASV+gGOkE9piNWoH7SNLi7PzGaek/ShszIQ2NfO
SpYBNG/CVzoOKNzHUZ4UWbxEGVON0swoxP1yLAu4Gs3vL0UXanqJPvneMWjiVq1t
ihV0P+pVUYVdenGNddZJ+UR6625VxKMHac8yETVWXjNiQYaDOEIciCuJRssxbUai
Ntu7ONPmo1vXG8AZ4482AzfjdnxX/oCOJWoGXa3GoNuN5DYUGEKbm5x0iF+7lT+T
HF3M7W8J7ycfv1DGdWLMyExD6u/77ztPJq1eJKVgHF2WaMzWJPiYtJVxXiKASdtb
EBj7rXwdsSoF68H1R/HkX3YoJUhokh9tcnbH2/MVMYYHFHAVC+xLv7QwtvRQZxnq
bxo1HQVdhHVAfP+pjcyhbuXWnksZsAV8phwp7auFcSjFG2NRnTXsWCK17POSq74T
jrA8jV9XGlzyS8c2CFPmp7FSjgUbAm61liv4ScBjOpQrZsoMCGUTuXpz5D5gjOAk
jhOqHseNpdDgtntkCnKOMdA1NLlPHpL1Q/vMtbTRtni+/QZMZDzNQVy0CQh45K7F
o4gUZ67MqYNRJyl8BvIk7nwD6SYI53YmwR+Nz2aNQxH245OMZUsSyD/tw0azEwC7
WJmwqA6408QjhjenvnmpwJ7RxpadXXILbqGux+tSEVr7qePk6CAnR6tzGJOXOFSB
SRD8cznrj0WGrXaakDcEP8rhwCmeEmWBfAkGze8nnQgi9hpb6zVlrOIKWANfSSfw
9eg1V8gXh8pG8zkhrRHNCtOxJUARAH/Car76DV9CSVQ371qabDMry0tEebg23/C5
I4u5HBAXhqXkhyQDjwXpYGXajPit5V5z+HjqWeBj/+PgWngXKN7achqwrf8Qfx+M
fdeyBjuNOO16kDYBkyiiWaafi7paQaZZLZc32j3r6DURsCZ2vPFT238LXFnLVFhV
+0ShPgRYGaRWhFpW7dGLL0WDXTb65VHtNXlTPY4aLilNkiDgy1vU7MqqDIb1iDpq
M2yM0giSFziTZN9ExAShdW4+nzZheb09Jcu+TrTXMwco6rVd0ZH/knmtuntCNlVY
ZkuNh6flnvbA5ft8szE2R5ug9nJ/Z+VuXM+1dapFboCjeDIvIkj0xymyiVmWwRJI
+/+1j/aguNxqbvCVESFhpJ+rmKnftRnpqRazuIiDjWESCwG+syMmnYlvhOI1467Q
UXH0esBcF969XS6FAVZDEHfUDBuHizHfmSt13vSutGjYI//sAWJE1nzy+6fLxh2H
g/CAhtZfV4bV3hUCx6NR2EwhqrQ1Mv63AIe4y0h09TQXozbX9mo6rsR8fO0RRZbi
SVVyMzipTdLE4vzt870yQOlKlVihEj9/+GyJZ27EA+fGjZdYWNDCUmttmPf+d1f/
bOOqpyvOi+sLlHw9lQfN8fcOQJS0pDWs8LCDWorCRN6lWYOWFY4phxXymHB0fW0i
KXWba+l45h4OGZdCK6JztWb/AIgmMp90aj4hQlHA9uBx9kP9G9pkOmODc427OaHf
Fur95F1tkfL7MGs6QB0BKJHEw2nZYd1Kybtks2hIPUk5M/tdhILZYfkN9EL+99HV
h4EW49ATSvlKTCiNOv6b/xle9HMY0qeoI/e+DcF0UtznmDLtOg1HgjO1BnXIc1xM
wToux5LzxyYVTzvYONdmsZot9XZF29MckyzYvL3YCOB6ygN+KPSY6qr5fgPArUft
SMX+jtXeObeFUB8dSgRGSj4F2+hzAF1C1z9TWR/cAHblcHcSA6R1fqD+XMbC4EMJ
1Z1OI3EqT6+Pi86siQpCLXeEJg+nLieQ4phPiANDg6s+MfCKwKbQh+fUJlkkIxwa
ZLWmR2IFr2zVFjc0FqfMAWbMGd6SB/MIosRy+Wyuj32pcUIzLwLw3gHyg5c101yg
I4EOA1b9qjCbRz6Uzhnpj1K2Qyl6fDk84LZ9NMF6VESO/sibL+LUnHv2KwD3cheW
2evxyCm8zMsXm0niNTkbClQNtfEExTiSY7i5GMmftbrK8KNj5bOUDId20Cdg6+zN
eoaQyRPobr8uRlpDkiGMdEejWPEf5RnSERnBR5BsYEtlpIAT+DVcpKjg51VWd82t
Jdc5R5Ke7vhvke/5t3bGqgHrLzY2XjBHwsbyAc1GgY+O6qWtWms/ipoZN2AUx6AY
pxVbjPjuRoegn5Em/788JNfVpUIheSOhsomO0t2HTwACBlPsK2cfylPcuO/wdWBa
R2uHs97fuJ0DFOMXZJckk4Fvjoh71MgHQcy5/xNro5q95CGtW7lNwHV6sKeO7FPq
Io7j2QpLGJbJAr9I2SkDCnHW4Dbs3tEtSIi8dZVUzertBX7sZSfTdBnSDohnkLGo
lA5+ALKtaCI4RiZAS48wLk9x1EKRosOutKOpWh4pDUdkjGvhRMkSEu/yvKUtfqKC
PX4fYPowNxv9wBd25sXxT8uRqCDLtRCe9LRhN1J4dzHGFf5y2HQF5Kj5NE2/N7pT
hNUG88qxj0PV45QEpHwj4CY7D/wL1K7CYDUmv6YPQ/GPVXL6RP2ZDKiPOlLLYoPi
TfEW6Jmli5zXJXm2/Lrc440K/rGpJxeGx0cKUcHTqxPKkkGm3KNOuV2OKg9YnZfX
fn0hEF1+NZvwcUVa1nZ9jvBIZmuwEbj0YR/+AeTxHbWnqIyFUtEazzbTcaS3sbV3
cUiyxDZOpLoLzr076ehcz3CgI7e8TGnOsP4RVbZF1MZW6jgoNGvwW0zBAm7Yc4If
QSod8qw7C6JfT9RIeOGodtu290zoKWARu3CbRJockWk9k9X6LTUUAf5UGk5MLGhm
VxZ/cmj7gwN0rqOJg87RQ6JbNIhOkCy8GSp5L02WGqUkDYDrMR7zoSH1LT0mqqV6
Syh2rGh5ey6xkC4yIii8F6I3stnert67qEP73A2Amoc8CY8B8cqD+8YB84wvz1Eh
L3OLRxqrNCWk67u6WRb1lEfjMiqwtGyw3LiiUfquAfMzq/oqpbVAaGARNTq+iq2p
MzCU/ypJYE5wIDQatMndEcL5PFMhnSzXQe+NaUxy+Y38lvoTSVLR66ty/yGS4Mpj
dj6Y92ExCgL1/8IxMkKnm3wGJHEO7kwtQAoMX75PE96LU3xLNVGbjHM1KpeWYvx1
tWptf/iqQq9Ba4qTuIi+y4KmenzoLqRgymh1o7LqvCJsMJKYU5Q7aRqDFgwv8h3F
VS8eLN744KE6LorElhA8SE6nq/QcorZ01he2AA32F6o31IKu+h+3lpAR/H09RzBU
gkxTRhpivSFHvAbsXAKsMBaQqbpylBOaPv81q34pu9GcA7yp3QhZUVoQq9JvLpRm
rUdu3tqWo7igy1JWq/nbSsnsnrjiKWVAtaqPqjhZGnO/NTp/nruBiTBqvq+SWt/M
xplNimwfyXwcroheZVgVcPBzAHUsZVhZ6nYLFFiqmCdXpyMPNmd08xOv7Eslvn7D
gp07n/3qDnO/WvPn/4Z+sTIcXJThcHBaOoDEQ7WO0cW0s2VRekXHipd+g1XEejsn
RUVFzKa5sP2bWPO28aC9ofx+NRzRio+634iYLGzE4syKrpXJBltUn1KZGGfeq9Al
RB8JsPr9w0tv5MyBJYdEZK5f0WSC0cuwR1b1tzbIBsQaMLRDZrUPdCcZTmrw1nMv
yPalKE1wz33Ym+a6BWolSKH1Xlynq/cqEcv4eXxcoW3SQ693kbPc/biStNxPNTFC
U8t9rya3d5kWpI2a3EBlmHTNmoTaX3kQLjdi+zj3aZ9wedqPFoMAuIU2VLMP4sOt
HB9buey6ZcFNeFJypTAtGgbS+TAAcrTNrVKcbmY1s8f4uVD8ABXYBN3kVMr8OtgM
w7CcltLJmpiTA1PwulwQTkqCue0E65qLC9Qjf246IN6eBwlfxAs52jzCzmkyOlq1
/naCMWle82M6kJUCOK9hpVIg/rpueqgCgt1LISh2VvahDZ2d6nZQf8OBGymbjXay
91oRws8lzLGBjAsmm0X2buDdssma6uiLzjZafJuK8fTdS3reB7fnvBNyTE9F3fb1
mWozCKeLdLO+Y+LZTyqNI5Isc/uZU507f3OYgPM0o3pox8sPapsIPo1Qb48WXZiT
dWdQbDF6rGCt892l5e5DFupJg0fz6KABWkRnVZI8LVY0XyBJVPcoHsvt1E3QAARZ
68e7wlw7ZxOE/GTj94b3mXexyXTwD/yCTwRwJNNN/+ESJF5tsVlfWpBNaUaSlRzm
tjs+aj1XT+aM8OaFCms0PnmJWgpPqMdaKHPcxcM/cQxTGh+z5RRE3QJBvl0pLfzo
OP97dN1b+HzGWYC0XXQM7XbrdgesPBZE6hNOiT4MmN1rqDdtofXWWNHif/ApxIJe
QX8QahpZVlWx5WR9PE41bBSm//QPnbnI7OpNq+HlSME9UyHcHwbR5OgaWO0TqwWm
KujzSDYAWVtQ5PQbavrd+INDMEqazx8trmxQ+d0CknOVYil8IGS4VOOibo0TAPJF
2Xk1R75CyucjA3sNGaUpwm/oKcompLj5LEWdmG4ZCnuH9kp+0lTq62feIu5SS4+H
cVMC0OQHQ+5ZAA1cK/aCn0z+aALmTYiAdm1HjEYFi3rI/3A+tOL9wcAmpfI1Hle/
SqKZ/kyowl1xuuDCsiulHPFH9kx+lz/CJJo++TFqFdHkBHM+feYATU7/KCExnk6G
g9aMqLwo+rpTDMw6ifFPzW+pVxiXc2hm9KvVuUz1DDNs7uTdfajz3hqhUogp6csf
oYIh6pKTYcjUDqRG3oHqG0rO9GLE6C1W1X274qJm1vhWz4wT0ehV85muXTy0xsPn
efVDRuV/nBviQsiGuupIVebuQfsPvOw9ihuneWNZb1jpBzExonceZrsD9wM60rnO
jOVWNgjQYc3ljVi28h/q/ENE/jS/RykS5XP1uIXrj1HLDdiLBRxENufUsbeV6Y0c
sXXjafh1ibP0Ivqayg8mpb0e8zZcLZanTygBzrV8NC1UMBJCX3B2BQtnUbdAlQxq
DD/O+rkeAmxBTu6O4a9L5DCUg95i7SBSNKK2OrdyR9M03hSPFX+zgWAWPVPedTJG
WSrsQ+HBSMI+xNbG6PB2ZKL/lWtCWKKF2ur8MCXO7f7O5qDGlT7hQ0ELIkVCOIJw
Z6fqLPeXpC2zcmTAgv9Yg+0l2FMxr1AR8YjXo73P8bBs0kA9tABvGwePDwBmkbdr
JJkuMST/7ESqON0Uwoxl8uc0yLIB3ROQ6mtygz/QMdveWEeOCdiSbOzXNIQhy+GT
EGmgV+7S96Byeb9lUOUumf9P82gjJtkEth9fMmn80+1W7nyvEWiw2MEP1ijBGobN
/8F40GisC2OjOlyCor8HcEe5MNZhrY0NSGldLSjZaXfkC4kj1GSGRxw5EzwHTjNw
wqNdRYaBWA35eTLMNIhR81nWRmdffXzrDCH8JhtPdB5Tr68Yqi2cAbTFsNnKxz67
5wh+Th9Vg8n4FLEozpv3TVWlbi3dGzDdebBeDcstjdslQ8GNRUULgQWJGtPqWxZB
4i7B+/TG5usfnJIzcAXdHj+ZNR2z73SVMMn+vkBJMat6rzhuuMYxuKfu74va6olW
uhDMPal43FtLd/M8iXsWXQFa0TVOHezvASERkBQ9Cv56XLpwBsN2cOQXrBQ2v2PN
rXMf38Uwpze/yhoa0aghJqFb9d6kyIcNNl3szb2UOkZ/fXi5ABbcTfYI0946ubTm
h6R59ZZs2gKBXkqqs1Nw1n61SYtVNDFjYMrU9+EYvW0dmOoxe79cJd9MxpqhTMJL
RJ1AWakOKCbmPK+b6KLEEOx+6bqtsA/IJFy5yLelaObgvBJp3M8s6sXwN8vui9g0
weGUxljePlL6iOvNqmR32Lg7G2K3PZGVrgps8PxLKIgjbV2juSjyW3/K522Q6Bn+
4PHdx6atD0lckLSIs4nnynCIp7OGGSNuRPGAve7LqW1oDim4zgivVzHPBtZSc87f
0F2YgBMu6C8hN1ekypIe+G2GKEx9+fN///oeJjItipSON3JBNJX3v/RVC9PZ8RNo
5r2aEPqn3epzAn3MlRsAW2nOKwo8RmElnwOfTeMWI4OQ050zd8XkFrmSmNTrrn+4
Yi+4s25nn09WOHYuAjqecKbCZBU1M490ljuBAC4AsHEPkqhbWZnUD1DFGqDv4SiG
H8oMCUWgHUJFFbUxCWwf5mBm2cg9UC5BttSuFOh1MaLB9Pmkm5POF+d8nw2pOA5U
lvNKRVdCUYcrBZ7NSPtdyERPT+a0qqn6nV0kbSrU7hRuvHbjf1biD5RBjgmOFiAp
ebZmD90HtqXiFYHj+Xlv1Ure6crTZKTn1yYS5FzEH2DD7pa4RydcPujyU3c6l1gY
E5mPHWR1dI7NN+A0oYvmum98koiR+O8ZqOLfQtA7D+8QDPI74lhImCeIWSLAWj5H
PEryTM1eYaAxrE3aqYlabvMZZaCHXLsy34tDM8Rp0FuXc/fp94IzVQi0trkEockN
cW+DFfGxnmvAfnVEwzPrI3iyWDrJoiNiiivcx3YBPwae6PFfqESmMl1mvZEBStWL
f8e+ldr6Yi5tG/6Z/YwI8HsrGmHzOjSvFcf0WpOQzmwc3N5n+Y142c7W4+pQVbTl
JSHzgmGx6od9JpcAuk3QFIyGLJUSGLZ0LE774V1lX1k0muivvcHHjnzNgYT09WyD
XPXbe7oCt5bt5sqf7JUeydqTEJoySMjmTOOCvsk1/ZXxE0TspLln7VpqdxjQGo9n
y45yzjne6D3Rkdn8NrKeyLzMxjFp8JZuhM+GRVpYaaBDR3qA6dAkGQrbJGUhp8hP
8cjTEWqI88CLN4ouT15Vvm+8QpXxJtSuCK+sLeW46mQ5n6QfvjUA9k3uo4XJw6zk
Crib2Ks1qWLHUdVzSaAK8XbQoJXw6P1CRCoJyazDNDvaRMFMFdNYbkEmoEcJLQtV
oxqMw2minx5/XF1wr6O5rbREOCPYdXc7rRAS/cz018xS2CDuz8B59gP5YGqw1rVd
NKfYZMy7ahHKUM8XF79wXMZTsntM8f7pJ0CByZguG/32vU+FLVtwuUproSazo4Dp
Y509z7ZecF3EoJf1UEnLqG2gJW76n+JxQFEbgGwtYrsiIa3/dzaPktKrZp5XFqON
/l5oXq6W3STzV9usWFI1L39Eutl83g9UoIbH3nyZr2xctHAGzc9sb6PF0GcmsUzC
zOqdz9oUlohS/wa6RjRQAQIt8hxgbTDv5wAb/uMvXMUhCicq23mrr+iaWABjRDup
9S05Uuy4sE8LWsII965dYaLV3gBI43SbgWIidT8Lskgx8fK6MW7HUED43DYOdnKQ
fbpxOU1hFnf8yJqrim1Eeew69Yls8iY+Fupuse2UZdWZwjlVCbF0DEHO370+fdcV
mWlI8onm2Z+QNxt/BgaMqKXtwNmrR7RhlHOFco9CDzQwMzxzIMa2PGBXU/lrzgMy
f4Te5WMoAFQguKX9r1lkbOi5tCeAU+x1E2Pl9DfuHdoQiMGxWqbEdNzBZQ6EHqR6
G2Mai7xscGtwSXh3wVoaK3zk1KGMw2M7I2MtExq1qJ6cP8ih1j5/UDls/6lRBF12
+81MZm394l9ryS3177fPP3kJt5nXJAwSdcV2z4AE+U2ZZnqGDE2it9nYqckfgNyv
/NRZtMAWjot1thPPFNoHtJQ61In4mBxO3RYxYgwSlhUX6swX0jcXtfHJgR0b4BsC
0t2rexvye2kpINssrfGAwTg7h2gtJGW5Vysq2GsCLSjYjfAiYg7B3v7JpsHporwA
OYp+d7x4flO4JsVc5E6WX8cnNiad25qhVOau0EruCEVczQkKbuldN2iM3VTUup8Q
dKeqhHwT9Oe2NNf0Ad7uNXBhOTsWGAFsvJsTxp2S41pBKI2cK3jmaHdvI//EGp8+
sqj3I/PGz3/D5oPrI0f6aKfV2Eb16hES/9//+xE+iaq4bLtKP2Z0shoSyusQhY5m
TB4yXFmQEolPyUFVZjEStiBt6T7sk94mKmiDcrt2FuKjWGK99akSyUWUqOnpI2Zv
FXr9tJEv1bLC1/U7RbpTodtGyvssKRG75fMwDweRKWzsyH107oyoWnQpAnjNPWpf
wJmacxdPQKuPytm7ojnwGiAQjLd/eQmc/nl4KmDckYBWeL0cbhwGsUPeUDztUr/x
0ee92cUaqWrovHijM/FBRAJi5W0qM+EYC7BiewJH4Ehu0z0RftANeADXks46pjQX
ZuO60dRUqBufnMBZBRmOw6J3njafzKuJanA/0ipwxUFslNU61/a+iiij6Lsz3w67
jcU5L9iMAykowaepBeVdproa10RjZiplVzuyCvaKD0V/Dlnza9ktz8J+n0kZ0UQ/
2DFBZhLvHAMYesW0p6QsAACSlyypN2borYnnaQ3oqtcTYYMUETV1lYqW0mrx6RTW
ngOczF9+SzBy5ZMJpRGF8128gbLJtiqYBiGqPMkAtaxPfbi7ckM5JdinUYRN9zaN
9lZpch92LRhkOooMmFZQTHzMle88zXTa9HcrFk74lBQj70mK/rVH7OePPp1yqDxt
zU48ibaMGnm2IAoe+KZ7KdITFdywR/b/wUjhojoBW1zwdVNok2Uxcaic9oETF6+a
NUeHjmr/iUTt9OpsqNwitLDbbaIjq4lC8FMikNM9u/ao8HrV8/bcCQWzfE6gcrqc
yK06YAd+SIENJZVZBuQ52/j57RuLKHZQdVKu5Cy6clwF1Wp++7z/1I08a/XT09H9
Vf3BUlYiBfPjZ7U2AIlI5nYDsdr2Z9QwGiLplgTBjdyS0H11oaQRf06Eq0dviCE6
dKGBW0+BZ4A18AF9y44TrF+XWbdfQNi1mk3dvU1tjyfD98yfJ1fBNe26gCqkspC+
+6acutL7l00aUVNakTSBfWmdS0e32a/xspBciTlRVqGurQRj/FGFxQ81oeEV3h3z
wzXPtNxNzRZljYmOJdHdKqK4z+IcbCkBQ3CiTjhfecnbAksOkJf6tAbyPgInJLz/
EMofOx19aHQrsYXYMleNNumHXNTr0SOq2C0noZkdyrWTq0bpoJykOcZRMkMH6MWT
H0mUwpJOHcVpBkkJwLL28ZWaM5HJDQYKKY5uwm2qX/28AP8eX8l4vcUTcig8bXcB
z5gLULIRblAysN/Alt8wzWa2S+CHtq/WxZQM3FoVJMIgVf/Y//sMucRlJCrXxLbC
QRG34xOjyLbjX/w1ur2NhECsLELrtT/y5UBe3APvwAkc7Q4zP9ZgtqWoFUrZGAkn
C6Vx7HI9la63z66u6IGUCI+obV4jtyy7GDxR2WnGW/6/yf5HtGLFCr5PK2S5Ni9C
IK+8avJI/gR+ErdJYGfohWmFTV0dHhbktrRWrSidBimy9C3w76yqS6gXuVK7OIdt
88lH3qLZCjXaqiGnVXDdhKeVWxJrC3uvFXFqUyj7EE0fsbaGiTUw+ySUayUU8f1R
oCsrmpVfGM1YfOiMBVwUbencetOPdJp9CjIvVSkPGxWnGfJbAixP1fa7x3z0ZTRb
lDbLyKJimMnCyVicCIg7X04je+p7F8FcZ3UH5xoZRxDTtw0yurXH/rBI4wl9YqYq
7lWsNyl6bQNSYDxWS6I213tmbdD7Q0A0aY+KGQ8VLZEPPAYMbrP4odSX0le1KnjM
+nVJnp0iZktS9Q3h6IaitrfWigpD0bS9Pmvz5XMmIpax8W3MT8KYeiyZNIJ4MvHL
0+eIfLq9Vi5KNOSF2NjVC8VPYpOoSXM3RfkEYSrD3nVbNcAyP9msGMzbt3LBvrS2
Xz+UE8kyaF5c1v57BEZrTWvB7OHBXKjZ4jNxUuP/C/3Le7scZBmeXwP3t52krXMC
bVjSMHOu+3AeO9/Y6+z0SwKFTB2RoBhvyyyAHEhgI+3wNFe3XRaNW54j3Zsjty4e
QRCCwZ1+88pXr686ejv3L+o4diXpvTZ5zsvFeGjcu3p8GDfJ1bsfRaEKlaiRy5zb
qOnQdntrlRoxWEH2oUYTacC+vrFxNA8jzjbfMcQHcilT9fT2LWbnryNPqOecShHL
g0fQgx0i8DRhSuHGEwvtdxGNedK5TDefHGyIga1sOJVBuExi+Jrt2715BnSlMB/B
8+RGJ+QzBVK1Yx0jbjEH5yLRb1cOCBZwfJBMRP+udUCJTe6n0f0/s785kNCJzj+t
36DQy5+qt4mWpxiC1f7PfIUqxLgqYBXmdhOi6FHUdrqej/E0jmo1E2yZP7A06o+j
BZKfjpS14k+0O3Gy/p8gHx9pNSW8o2dic6XS0XmIg+QnyFvFFeaYWpASIvEE2ajk
kB8AiIrDpRlXp9gjfwson41CaQUV/YnZnrRFNsKWccMQIJP1OWwo6/vAtjKgfyxi
i4IDN8dTETnJ/NZn6dlI6G1yoah0MzP6TaThxF9M3s78JJKRu4CwyXnmImjUjAWY
m0qi3i75YYAlKKffA+qaOPRtYMfbwzc+BwfTXFQu9DE=
`protect end_protected
