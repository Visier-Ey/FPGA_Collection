-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
--pragma protect begin_protected
--pragma protect encrypt_agent="NCPROTECT"
--pragma protect encrypt_agent_info="Encrypted using API"
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
--pragma protect key_method=RSA
--pragma protect key_block
GcXwoiQJxRCDdK5dghUY8AYys7OPvZKrf64jArdreTEG4UAS3LbcfJZbELUf2aR7
dukZuAhl+1mdrfbtHxwQo0FSRqKbGvqOPqzfBRNS2/4e22RQBiudcg3CcdwRJ/JO
qLLs0rEI22Sj+SnxbfEys1Cmr71OTZgT8r23eY040Gkuwb/J6b8/qjolMCBUXKH/
4NgH5p6y8pomZVkDxoWweEtDzBQjdaOrBi1aOXOXDg2JAyUx8pNfj3nQa7qMyePV
nfQshUxVtgKPUlSBRMKr6itd7ka9CcYGrKQ0FQDgnmKoqv0WmqK4MeCJqFozXJ/C
+HNAHptEi976r1irCdsfIA==
--pragma protect end_key_block
--pragma protect digest_block
CqQ9Wme1ZrgksCW8NFAIbOritDE=
--pragma protect end_digest_block
--pragma protect data_block
yK9u6UlkkrjagCRPgIHOTYodoc8EJ5w8FxrmzWKO4HNV6L6F6yBNhfjB0K9q4MRb
m8VyIduRy/XlDyWhD7FDPoI6hxlYWG1ZoZ4PZjwSQDAcqCyko2YymZLcYJdWPiKf
bLN7A8JV00o1aKyG6mGhqdASqwtlEsb1/kugrYGqFWFbGce1iZYZltCv5IQ/9GWl
Zi85W9wNuOb9q1MeYyB3AkDE67Bh1JsZfH+vy26Bq/1Lz9mqUGFaBJtfvJaAaV9C
MSwfhEzc3f9zbMHLHHYADIHmR4ahG1TIhdnEkMqV8mNNe/IMR2GZMCOnXUfcNuCr
bBCX/rqVwjZTZJg9kpqK7nvZENfzs2sicEKkSrPCkqFc+w9ikHtnPFkfTodsO4Ro
porre3KkRMzkeepLqPRLY2t4GperjCtm68bSsvaoqtwG4scmpJAGTTP+PoqjM16l
ZZxZypfxGmSltiNs8DVf97rl04gBma+a5qpbKnsrcKdGvjCkKXUHl9LHox1RSEXt
DdR8gx3HhCJv5NKs6lPR7rof5awuEdXNLPTXwubYjK5cA3L+PjqvW0A2EIeoj01z
fT4PQi9axYZT1Q/qG+YE7v3cRpBS74CborykH1d5KxkTcTfdpBAsBhAivo646uoc
IvulE/2aZuTFdrbOuEfVSsDSP0yJS5QQzhf51rjintOOIgDZDAaymhGQ79b037iw
ii0+jEsl+e4eoiY29cHvgXLqquMkZnoD71aEFadDFFbF01awf2amV1YB0KJ4toNM
vIj+czQpbtugkPz0tuDfkme5CEj7OZqrYPzOMKh2GhA3U6q05dajbkLLFkyd9F32
w/vK3beiGhKvob/bb7DzIjnMR7enh/2Kx1NlWWJ0OKnscYPWtXluF0DscYlNNAei
vgzZCcQTx2OuoK6jYtSrou4J9jrYPPW5QtMPxRD9VDPWGuyOqLGL6ZPVzHvgZs+T
y+02MZfwWQKCp5/jBA9lS7Wf3kWaCK7Il6CneKyo4oTs0L75VFyEqKARY7xhLBTq
FMW0QVTKHzMXlys0kfNX4wsmmxR3/7a2Kyt1mj3ElNp/piSvhilc2kwt1ceRgN5p
pEId0hiEMD2B2YY1A4mdOjVdMNaXspVX+iKENJjaWijrq/WKqxAwFHEgslvGg1qZ
vRegAwNhLO5DvMLNb/B0dcuJqz39/5qvpfNWDF/TqIvqqgsG/E6PaFePw7UpSZ8k
dGqSp5kc5cLvjpkxbb3gKIWWm5ygPhV2fi97NvehddWdiI9qI/neZSRkrWqjwOz2
Rar/tQfeKGK8YZE4tEC2EfCLyEoGg8VoqbhSiogosvmC19jl1edpksfhk2NR1PG9
JjWGncddFAi837F7gUGEGyhLYHLDlgG6mRXTD1oCcHIOEm5X03RbsyhHApDcdVoi
pSXq0QJbleSVREFg72aabALX5OjzqM8BJOBtL42vGPGItpJ+Ry45drsTapJUdTUB
BzUR+u66UdszsVnlHJw13lSnXLJzeK+HuvGdAFIMG8mY3lBUswqcuUDxH9ZQJ2Po
wz54vF4R4OBoCt29HCf+cXYJN1o8zarNAzceyu/vDkurdN9V/T4rGYyMJGdpkxi2
OpceZjchivnUqr0WMdPNMu31mw+WJPH5VnvmbhlAH1m5BpTjoMXotQ8cdc23dGb3
ox9xK67lpdGSZHmHyBYUOROFSfvl5smFDWO7F12gC3g9XaZZP5MiqQbwTGQ2i7qF
lar4K0bdrj4RcIZcVPYOgrb1NGXqyAXWcOp19gfQdrl28Ug5KlG42CKtFEfjPM3h
aETIzjFsE/+TwutrJIQSr66rjRPEg0cJDdDdTcv8gwWylOBgx31TYGCKlkC5zGyO
JS9II8ENvrxl0yoieRpPAJ56IGVyzpzFucZu2HUy1+i7DvSUKgth0sdIANzgXlWv
daDmJPMyfCb0tWyZFwEAS8brLwGSAYON2gz7uNvZqB25NUp/2B4QI4y5/tRawuKL
rP4tUZ/4PxN1DhJrKr/N133389AAip5a2gfz6+t/OuFm9z4Q04Ay2hFEGFL5JyRR
XHbmYvuPo63OAO4BAOqMqKw4BByIqwjDMwEUBa0kSguC+bbbmKLnG2pEfdIVcJg+
WRShioRLeHQkRhmgIgM45+WYBEd4gS5KZdhH/Uhy9Ddi9yDG5HHTvIDtttr298IQ
HiV335HnbkEj/wV2z2qd8OdJi+NGpeB0Ie+wmZtEk4ICl7zWKoppssFqwgeFdgUJ
y7X84wQ8l/pQYq0Bn8TuLft4w7z8YWNoAjfC1my9HZubCTxFN5FEcFhqZRDsuBiy
yMRblgojay1QgwOP88t6al1uVOZbQilVEK7qVzv0mBJ989INzPTwmfaEksN6L46Y
v4Ys7Kk7ojiEQSab6L5/SLX6aqzHvyZn0Rk/3UDDWvKUxfvy9ohVyeohOG6ZESYO
0s1HOgQM9EyPGzpc3vwttDxoxSiuMJalgdeKlUZZPSG27tD3r5DjZaLkMLka/fr1
cWm6Q8Fbpy6i5p5TJj0klPGLOpwmNIxbDnPs2u2CSH4CES5WHBBtJ92Arlof9xHu
MQGnhfZoltKb9KlF9V7/Te+PdrNXfxE5fU6pzIrM8yvhNAE/KraKVzUR1btOVS/I
JFO2bR0SBxvgNCkqy0hBHkYIWuYu+ecVM6adCglJP0//ESSX34aBjcAJBxMPKr1y
0zQuVjkNUGNR9IIr7fLFQgMfklGoAgzfoTqxhKUWb4+uHhoWT1VVXRyDKnlwEvIL
1qWXM8ewlrNx/ZWndWQVCe5orlsBrCM2lHoE5ialqNFeSYkf+Nhc/Jbqoj/QBu4k
dhNXPv0ggx2RU+Ht+VQKhR/lu3IBI0LB71elVgwumfwUwNvbwktDMhG7+gn77Z9K
hQyuqBK/93KvjjmGg9p9M59ZAyr0julxQqWfyVqPPTLMw4JiKlDf/2n2+yqYi4OB
1anCZl/n2WqNH97x/PJEW7TZ0CzqRYh8xswF0+yt3dXBvGAocA8Y1xaNTKZKvBTu
7f74/H+V+gVONhm852sOxMhjOIAh/OTWH504KM9+iExaB1mg8t+fXqEZdYT1wiK0
fdjR8ZXhK+6I8xbRHsToMehhGos4uY4IAyRELxGfTbYZwG4FIE2Ij64fH9z+KZTS
HwbuwamrzSzBwv/VDwWyQobVaYYONMkqG/hKLLQGLeEkr0ScfVupp2gz14ga+39I
rFUcFWJ/LIE6wZkcln/V2jvkQbgba4wl85ZSghX9oU1BNNMq5K4wCODxaUB4/tXG
R3WIaxX/Nr6DgUz9ObKOKVvQ0+a1JBP2WyRf2DsC95cvEcVGfdMSOrgr9ejkZzY9
YUzFDfRjGuCdQ/rcRM3J7xEGS43HDWr0CL7eB8bfwz8HOD1fXXTpOH7nGWkcdwBn
a5mCjIrk34uPBV/G4BN7XoJ5GKjXY2MVmS3rZclSU+OnC3OGh/ycWZ31tfj3vq2r
X9bnfYxNUTM9/J2k2//wNcHPcD3hKCDSqJg6JmaApxp1DivqUe9pkY9yTk75ldV/
aUIDxH592OsH17p5qimyjg4vpOS+5TCmddJq65zuz3NAdZchyeYUlLt5SaMfxiL3
BE1vXm6WqhSXh05DoLEqwxhtuK+BL4LJCP2iesucSjS8nlZ9EXrt7I6760H2WuGj
EbaWzHj0sDXt5vLaY2q0XQny5z6k9N34pd4dWSYMP2MNXOzAcRhgobVgtEslNnVf
oqz8S83jjCi+ORVUDN0w/dq6eECANC8hTahUMCd4X+2tcTCvUCc9McwVtpNycCZ0
IvPuVpk9UUnqxlPN1dQn6T7f9etrVndzXc1tPQllPbrDGmWmWQSRVmGUhgj9Ghqa
e96giUuccfRRX9ndXdrjL+YBgBEb7t00xcJ8ge1wvz6LXulbaoybBMLZcKjWY4Mr
B1g1LzWYMdZeMxCyQxo2JDgf9xz7nA43KXcDFdZipwiyP9yHoc7u6bz34x4sTGln
Nkg0DUPkrkYWpyAmNmxEfTPDmz8qeNVSpTWhmkoqn9mcSdzpmuOW1q0LETxokh3G
pxwTosjL3ZNPcr3+9mCtlKSfde99rm6zY21xD08p6A2FVM/S/wr+Xp2vUxKQ1ktr
kU+WqiaNFIBYr0y4jOjZ3xMKTNAOPE7uc9FQU2OxLWk3BucHrGM6AD4hNl2XnVgO
2pKbGg0V6bdytClipTI0AqmxqbpEHMxTyP33Tu4D1qiln3Hr2sDz0gVnB3JyHPRr
Wgxfh73k1/XhfrrQUcgpLsc+jHljImWgw6MlSnZnvp2dLjRsUljfcZ2I6wZa4W78
qXZRbA7v4qAK7rmf5frT7O7tNuhC0CINKWzrdTd2pJ6L4m1hlKJa+hbzgK+I54eU
Blh+2+rXly2iuezf9R6BNntO34g0g9IEfvjr5vcWoRBAhYtdC5sph6uT19lOoR74
EZh4Nzd9U5DOiVIrsQSnlxoGsLY3mM/si4JCsBP37eVFUIxBB43ZU87liFjfDMRY
jEXn50hGDglC6QzpPwulasbyV44TdNTPfe3wukQHksdkeZi7kNUoudVUnp8LNCWU
SySQRBPYBUR2KjSNM50uzIRNRJJz/rDIjBQQcKejE57IrMvABht8IlrCXbcZYTQh
wNJjZOzM30l2QYoSiOKHRbNTtVhBTfW7RP2r6TeQC8iieoNnUONoYZM4R5KQcHd9
tCKLbBrHwwgOm2eyIk/gNBrMOABnZ53Uu3eKUv1wz2gLcRH0KWa2HcI4enNmG5ly
GYXWctvjPGJPwROlgYYTTzvC8uzuB5FDrl5YjpdbwtwCZqYIjaGLJaY2tSXO/GUk
q0sJM9QJCHnXM5WyEbZPQ/3EPkSvuHp8xK43wIYPGzfTf0IXuiFPtQXZgXavVVjs
rTwXtAMWIN35I8f58aJP381uAbD9ldGevUHN0oMYpUTz+IhwI4d1N+LaZ5tramHr
+YACDYcacX6TSKi8cJcdOUL/jWVJCkM/gZCKIXvQATp3U841bbN/F/ynBXEVsHUU
yjtqdGRlLp3MsB4gNYmMNIzeuJ0VRV2S5aoyLo6NvlD0wq1Koe6j+/MwT/74++9r
yhRXkqniHCLkkqYl1PboRVOiNewreS1ZAcANYywOUuX5Dj+9z03bGHG9MkuYcCH8
lPqnl3I05F1ed8XUhnq2gJsLO9D91fecMRshQn1HcRCyBYkbvhwX+llDYJfClUxY
qH+m2iFV0oqAsfAn4KijxmtXwL1e8Z7WuLWQMjTuy7KmEJJP3qTMYfaxvzNDQpfR
EYDbZqg7dEanDkssQAONmpJmEYyIL4mfW4Ci/WQt7CjFSzYHuYXi08LcS1UECyu5
kVTyIVsifeS/z5dI/fNTTWclh1fD7tXGYhgv3GzqsiP8GcMsBC6Tp4Gzzp7QjRaL
AObmydRGJ8fZ5O0r8nCLaofj/uD9MChFXjCWKc2lNetT70W2UQrimlH0hQ06JvMY
CaxfTOic401bqKaYESMeelJAndc9+b/FU5XqkJQzMjsSvL17s32xI1tgG8WvjwGl
xhtyvbbYtU7xnqirn8fFYdtJSpMffCrqsaZhhiP20F9XWXRjJnRbsNJOC90tFytT
Ip9YS3C4Q3j20B33CGWGnf2sDuxlZBatsKlou2hSijyCTEXhPcMld8fdgxO0rBXy
6nc4QKZD+DuNByxFY+56sH28dhjOxkXfhCSx+dlA0GD5pF4us0Amwx6wF6mvOH8q
aLVUET7vbvFRsmDXMwuiRN7H3/P8rpd59vIQSOedAhlFmcPopX1ciQ34LYpd2Pq0
3sUYbCR6SX5LBy1yWfIX/xK/WIpdahRDx173apfhaReIuE645ClOy86313ZwOpQl
pkVsjvTwM5k+XES1v1+g3sXNuyQ6iw0cgyNFT/EGnKxMbQmFILm1ngytCsIWxXYS
2N3rinPFomvKceyYU27AalH43lsTUs8UY3FRo0FSOALP7+K2NgvIRnLQsPK7O+6V
ZojKr3CZgNf8ga6de3H2HKeyqI70pACBemibsenFUUsrb7j75OY/E3vz3RskiIBY
ngT/vP59pbRDYXpZNai78B06Mo/nxqSzAYBUDqlVursARwPASsCa6KCX1hnrVg/9
C3Fk0B2DYq2Lsgq3Q4/M1vqgh+3maunK7i7MelGJTXjH+nY7kSO94Z72QgPoTujq
2CiK57Uh5jQx+cJA11LBdhuGY3QNudR4p6kZhDUwA30PLm7qytHfqf0i93bQ99rh
U1CxyWgnLoEP/xI2kK0hFU41ic+tDC+0xDrGNWKL7BomAN0ZoPR1CS9pppG93LLY
TzULUq1MAK7+sRG9Jw9bS1rB+VgI7YO2SHEYDIif5IvYh18rlrp4V9+Eo0PgZhue
aEaMy+jhTPXnoc+Dxtx590czvXXPFb8iNZv23FFumvv/Cgx7EhWujkXbjK59xOfi
0gky7jVeab37reWPxzY0THmEa9Yv2NPpyuo6dZO0SnYCJ76ljfim6f0XHOxOrxxF
ITerSjoktlyGzda7yD+G7ocMIZcVYo8feSooJHhV6FUeswvn8ZGLh8S64hVmgQ8u
fjVGV49AwdqRAqdFIR/t3uToVwWL3QHwSUxxpmD53RLFNDczbK04+pzCPMSZg78n
0XW1WzbwaHh5KW8Pc3/HYQmAvooNuKf4kyCTkJa7woUB7v4tF0+CO7kjTjoaL/ak
xfzNnBfHfQsxXdyPFSu8CetXqxIpNkJD61Cm98ZeNZh17j1MahvrsFBQS7kCHnHv
wxLitMFYwrbeBQaPQX9K28phwmmPVYHOvCNpkLDlSXQofEtxYz0JJHZahX1xkJKS
hwbiiy3qJB2IR/g2x+jlSZm6HuKTBtvjQ3w8RLncKvdsk2FFxvFsE2T5FHybhqMc
YikORS0OXlb7a5LKtac3crjKpjXpxMILdk2q+MVcsYaYYFv3+eDpg3YzJcuBhUZX
pQKdMMsZy2LcpDQZ4Gw+BJZGjddaBrDVxBNQFVP05fsKgmM9Y0ejyCA6f4RbD18W
4GFZffKA5J6/sLSkGNQoqJL76PtHnlFZZPQWmcGAfYg+ivZt6otreEyTdswKvqe8
cnPJt996iimkTSS8v5LLl6qNMETPPVtctqqhvBdD/WDVzJhaHUZsDSnVpgO8AWFF
zCYvVAreHyyxp+qPW87e/8bMcfhZFH0kEpgugLHn75YQBmyNkBlN0OA7Baj5a9YE
YmIa5rYZWfGtO0HHBNUG9pxhtHhhBeS56sl+c2mIDXWTTszF/FOHmQdGpnMWqRjJ
w5Vf+frjVhCJv2Mqs35ltMarFMbrOCFjeZRrUBHnDiqwwCQoSw8UClo5IllY4eCv
lQa5XHy/Wo1BU4oQV1jrNwNpakuTAYRt9XEf86/Y5ZqcdoOVI+E8vFrGUmkSuybH
EWfmJYYcoW0hpJ/JD6WSgdkKgwBzWUjSKLyYV7qYMbsKqvb5Yvu5E6/eiG12c8P3
txUU6qnZv6OBhKyCdOwrGoo2Te7h9VSaOVHePwjdcuYQv+Q2TRrChZ1jAOmrfpAa
20njNiz+eUO+Rdx/2AIBcZQ0MUBrT6Z0sc+KNREyIbHwn/Nvm1fXn4zgGmN5DEG+
4fhydLKk3x4bg/tsb2LUkKUd5ysEqv/1Uuj7cO+MyYwxHhVoKYEC0FLkwpqAatE5
hy3hfX8K8tlmnFPMGjAZD6d+BRiMVWiuiNKBGuTYjnJDkvbh3gR86o86UJcNqmHH
lhjVKa0ZBlaZ8a7D639xjv6reXDlwh5x8dmr3yA5vV/pwvzrsR0jT1k3YqXayag1
p7+DP5mtBgczr4Sb5ANMfw==
--pragma protect end_data_block
--pragma protect digest_block
F1ZkEDnwM1CEpbm66BDYoRGQN7c=
--pragma protect end_digest_block
--pragma protect end_protected
