��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F��������n�BJ�F���U�FW9d����T�+�wt3��^��r�q;\��af�י,��9NL���ٴ�[�Z��^��Jy���0�T����l|�x�5#B�o* ��J/�CO������|�)6b,P;����t��ew�u��5�v�u�E�8����R�oIk�����Wb�A1���5��r�5Hڜ �r�n+��MS5��n��þ�|R1��������E�%��0E���;%�6�׸ۈ�6��:�!�#��L�jT�a�S�N�LS�[�&Ϫ���]/��nm� 8K� 7�H�be��
@��1>��?���X�U��&��P4
��J��tz�6�^�O�A��S�������EjS�V�6�$�g)�H!�uA�����.����c:k���:J�G�y�*aio������6M�pʫ��QZkw5~��ΰ <�z���i����Y�T�w-�q$��k�d�V�5i��[�r6t�`?�.�^�v�
��l�;�y/��y6�]*T�۔"N��d�V۬����/S[�B�U��7 a��p~q������~�5�LPؐ�V�T��?*�ؓ�C�r�����	�].o������߽o8+\i+�`K��+darwEi�JI��4?�}͍�<<�,�j��'��u��K�C���=a�X̉��37�Z?�(ȣ�$��Yl\e���=~�Xa��s	 -~����w�N���,v-�xa��$a2��hA$]��g���[\�7�x���{�MO|���1Wc���C��e,m�"��������n�sv4��%-gϨ��hd_�K��f̕�9^T@-h����i��%F�V���Q�%X�q��;�Q��l/��M������Z���ȶ<(a��ك��BXƩ���<�L�q�׼�|3�Ee�w�/*�������pY�V}�hiF¨��}��ro�Iv�A�3zc�ܑwN�8�g���sE>D��*:J���o��Z?������R�:Y�9���Lޫ(�{;{���4����G�Bm�G
o91�5Kc�����'��+��˞AR���w���_�҉��T�
is /J�v�~+cԷ�3*��:�c54Bto�/{v�1oh�:���np�x�������g�E��գ5���~�jO�+�yX��+�2��APn`�}�q :������z"%��R�v�ۆ��v���i�'yU!�$q ��ٺ�$z	&��m�0�QomVP\%ڻrC#���k��K�bt�9か	�}{>����ݑ�s�<���>�O�K���޻~H��%��Mq��N���>�Meo���\ت�5b�U�g<#���:	�a˕/.rJ���1�?*�i�n.�����W��7$���t�x�~��Rj����3� r�Q5�tR�#Y�A��ڻh�z	\�A��ێ�@���7"�D��A�U6y{��"�(cUTB�.ϫ\]�mF�d���~`
_0Ɵ���<���Z#�)������$s��A�pQp�l�%B��P��2��mܗKnjYAA��y6�
�iCߏ��RVS)u�veD��k��Eƣm��ٽ]'d=ހFw$=/�w�׮"�E_$�T�+�M=�R����~Hd���V��8�_�LZ��"� ���h����?263Z�BI�h-lֵ��@0.�e6w&vk/̏	�j[r?t�0:�NAU��r=�ڈAI,�|�Y��ȲP��K�0i�!�� �4u�?Fx
�c����j�<W�dȴ�ōqc ��;�x��m�i+c���M�=�p7m�φ�1�5�_��+����4y̘��' Y�Ä����)P�N�W�o�]������Ա�D�r�	5�G%qC��='���d�� w��PRÍ�%$�qP�׈8D|���ݴaW�Qi	.�zj�s��i����\�҇�S����0��i��v�b�ܿ*$ ��5}��ˇa���Z�Ku�z����u�$}��>U���_��NO���,��
�QV��ݻ�4�\�hx��u2�z��W�%]ڙSt�h��7J�tr��U/�U؞֘��K�D�+%m��W��2�G�&�aw�<�*�M�����ԥ�gj�ݍʓ��zȂVZ1钱�>��۪A��>K���=���8��]1."W�Z�^���>�	��i
��9Y ��VR�0�1�\żV��B�Ԍ���7�\"���kQ!/e��$(,r�EL__$pg�#c��'F=��Yb:�����Ȧ�����P�%ܶnFO���cA�-j��č��7�]��~S�4=�tA�����e݈ە������dbrS�b}�ã���􈒚���S��;$e�H9���V���IǓegx)Ҽ[(b����`��7��6];C+� g����^:)Y���?�H���ډ���L�H l���ۖ�q�d@7�F.���J���x���	�t�Jt�	=K��8��Hr�pf�� s;��}b�"�&V�ΐs�>d��$h�b>m栉
	*�|��l��>��ZZg�3-�r���`/,)/�tt����I{o@��c�(��e��oω�iA�6��5��N#�ʥI�7+��)i����R���@�p���<�hʋ1Жa|+�6�H������C�֠!b=���	��X��;��.�{3#��,�go���Nw�$∡�XL

z�<�h���D���E��^/9S�^��X�<�d����X1�?2��
�d����ܜ_Sa|� n��.�g��(6����dГH#~�xxq�If.���騜�Y�]ܧ�ſQ��V�Jz�x�sC�)`��6��%�5��q"$���qy�C�D|�A�RY�w
21x�g�q{3�~*ؖ:�іI������w�8E�Q'���/j�� �q�*a��BL�߿?��*2�V�
���8Vq��b#c�)��L��p�|�����A!J4@����C�� dj�@�*��'��[�De\�Zyu$P��}y��o&���Z�&�Y}L�r����[)�O��(P��.`
yz7�� 6�����g��ň�X�Hq}F�}$�*u�xb�͛Zͨ �E���9��m�#����_�9
��t��;0���H|�7|3(�L���5y���"��5�n]4je>�L�$HD�����Z�G�V�i�w����`!��Z�Ua���gBq��P8��.�p%V�.�?�/�o���d�8�ɇ�dKJ�X��G�L橵�|g���Y���$�E�<�,H
�!t�m)���jJ=�A���z�fZD[.���G<���!����2��y<��Ji�!k�j|C�aX6�z������9�� [����UwGt��O�����S8�idRi�1��,��������?5��4{u�j�����N���t������FuU�X&1�p'y8�o�2^�ł�z_�( 7��z�Z�R5+褷��F�gT����!a�.E���(�p���T�C�B�
�@#���z�.�$o<��/!�i��l\����k�5.a]��奯�PΓ�E�V��q���7����y?+�n3������W�~���W�������#֏ð�q7Vx��+�E��vov�����k�S�p[�8+�-3��k���+�٢қ ֧CJ�pv��r�*�B��\�|�c�fb�F�D���"\{�&��Hdu���WT�fpd֥x/#������;�`���9q�����u/� �QBlߦ����)���G��Z������(�|�d)����'�/1��<��#�ORVx�-7��:Hݏ����f1���>L> p�*(�_=�+Y���u܇I���=���,����%���<!E���D���}��6��d�M� �i�͔F�q�YV�����,�⩛���߼E����3#\<��Z
iˍo�OY�K�{h�v`���u͇]Lvw�?@� �c裓��Fz�wW���������]#��!N[��)����٥")��:�+@��(�w&Z6�Ԧi�9�i��e��{�+�GtS�.g# {�}�ʩ�,P�:��Q�5������㋪8�"�J'=��%Y���#�"����?���TѸ�7��r�e�G6N��2�S$@7���|.o7fQ�Lo5�w@��>��n���s���6�.x?a!�"/���@e_u�7,P_�M>�姃]%��2�����#)\�����}��v&{VmQ�(��Ҏt��{�/|�w�,�DX픠�*-��fx�_�@1��m�fX@7��؉ۭ)��9��>c��YN�KJ�>�m�\��VB�(���ϧ�}Oy-�tٛ�]���C��Rb��Y��E^�*�`V:^�'L?�=o�ܟ`^)������\�8���� ��	�r(s ъ�d�&�%��62��g�+E�L��S7:�兽��J-�R@��Q`��c
~~~�����l�@ 8l._�*O:�K�n2�0a�u�0K�G�C�1��l`��H� K�t-�����]f%g>�eh7=�?�Oz�� K�E�L.DZ�	��5�6�s $*܂o��É0t�X�~�����ݮ�f�˿�dD!Pr|#� 5����U��I�\�0Y�o0vh�˕Ů��j�S�	�`=���ؐg��E��X{J�_p��+�C�@�����_�~����Y��9����V�^"�,������=ʍ_$�Z�ޜ[͢7y$��u~���N�9�}�u�Y�!w[���6fG�E]1�>����������׮d,���{%T���,m累e��&s�xQy��k\��"�\�u�ٚ[��h�-�I�`a	����YE���R��O��fw�>/�A��L�ʕ��Z�:�\FF�ڍ��t�ѝ�`vfa�	(��߽!qX6�Z{��b�}�苦'�j3����W��c�z�X@���G��I��,�g� ����E[=y�i�G��R"��̨y��wxcR]��Ѽi� ��$��p-�B&9Oc}�,阶+r�T}sA��nd��47��b.�bD�Ǭ�������桉�1�|��ˏ����F�8,�3u|a��r���_��1�?�p*����Q�T~�\�+2�������+�;k��l�՚��v >|����u����0#Q�ޱ�N�v�f�K������Py����H%-�p�5����cy�ϒ~^ê��0��mn�Ǹ�Q��b�o�(��l3ZѺ^�ê	(��3ql�'&O'�;�%����K�4�΂x@7��hTi��6hލּ�i���c:�u�i����{9�t�����=��!�5{�N�o��3x����B0JYOQ�ޕzs���=,�C�y�}IO��|F1��`j�Y�[���5�2�@僗�}��D�]�ǂJ��ӳ��;��&�3��>��[ (�4�,��;>����Y��JJ��)*�L�[�D�����#ra0Q�{ļ�v3d�?��4���T�N�8��à�*%<��2%��`�gъ�j6s��L>o��_��K����	�lB�Q�����ZB7%�8�<I��h\�G�e��,���`��Ռ�<feA����W=��e�/�hP��n;R�D)�'��
��҂V}�\�� z\���Q�?��[����<_��Z�j=!�E���N.�U_�J<>3��U���Ԧގt]2Ђ2L V�\�d|Ϲ��mɠNY9�U��`T4|^.$.�i3&E��� vt��#�[�O,(<�|y9�Ң��Χ,��R�������7��ne�=]\5`��Bp�	w�$�5��׺�V/��}�����\�a�����-��FW�xӚ}� �/Q�	<�e-c?ӳ[���,4Bbr��<|�Xɰ��BQ������v�9��*����m#�*9E���y�.TzTDWw�"_Ƃ�c�9V��������5O_t�c�J��.y*���Jr���#��ҏ��a)��r>*�s�N��'uq_*Əֈ��.<	��[�q�ۆ�o�oB�Ir��h���hN�Uy����ď�}�S�Df��a�P�ȏ&v��z.X�Z��I}-���5ݘ2?N�=3o7r�ϏKR#i�?W����ûT�|~n���e�M���6W�fn+MY�f��h��B(�ȴ�F@s7��P�;���]m"r1�U�g�Ul>��粸�ܾ��&�/�L���(�Q}���xpucI9XzM�}��������+~�|�D|�����L7�j��	}��qP]HB�DǇ:�[*C�������D�^  �(Me���˗��Db6G�������,�_cb_��;�'K�Q��,WB��WjA��~5g^���x�D[-�CϐT#�-sKѭ=�bÝ�����h�	�")0D�	���63Ɗ�L�V�!����@U�w�/g��pNjY�KTٴ�fׇ�pDV'բq�G�!𕒽�#��d�ڵtO��{i�����sz���c�
��1yq���Ʃu��v���h@-bw�ɯ�a�3������G<G�T����A�
!+�39Mk<��E�)"�. m�7�܍
x^����*RN�@
B������d(�[�d�$�v݆K(�Jp��� ��7wѤ{��uc"Gc���[��|���\q�v	m�N�s\�į��?j4�P<P�:������kr���j�T�cBu�AL�/��X#8��#dc��P/w]�����a���c�r�~5#~R�'q�.����1��[���d�^ɄkI�����6a�GM}��f��:[��3�˪B+��7�1��R�Rc�a�N਎�k���/&�P@{l��"��}X!3G+�
;n�IIM9�f�>��fY�g�K}*e���l�������rr�$���TE��f	��+뇓I
���H��{�ά���XT����y�2ˀ�("$���nA9�p�t���R�b�<�B�*��H9�`|9½�mu�*�mF�+�Kr��^���i�Nm�'L揭5lB+���+����Fb�3Ǥ�D����ՠ��/N[Xck�/W�{^9�v�1#�&� *���@��3MZ�]W"y�.�ʵXY��f����fA��Ed�0�_���dA�,�St���U9^��Jڐ��n_ߕ��@6�^�Ъ���*�K)��Pz�\�*P"�;�,�u�Jť���,�v��W�ss�����OE���~ٚ!�>F<�/�N�V�r=~f���c���c/���æ؆
b�.|MYC�%`���605c(�&K-S�3�L� vf����ιG���B%^/�N#ӳ��d.��dJ�n֫�[XY���Q�=ژ�Pb�$��J�Z�u<yr*Æ���6�Vv;v�ӊ���"�Ę��F�pK9���_��秔�����H|����(�y]��{8N����h�8ΐ;�&�+[Oݱ�P����Ĩ���~�^ˋ<�먈�<��NG�f��g�(���?��x5���k��&fV ~.c��� ���O�#��8
��q"��6D��F9l�%���������@��8������u�\/�X�u��E1PkX�~2	h�o����^�_�L�PLR�5����R�>4zu�I�8�*/g|�%ڒ�N����]P+���vw��H������jz�\�ܯ�[1�E�X�|Z߳vs�VbJ�<=��x��U��^��S
�mq��+��#B�����1�&��f]�����\�19�ʿ0=6rRm�W��f�Vn��d�<'�U!��_����+�,��^YU��>HP�����uN��E�B����]��׋kW�Ӈ�p�콎]�Y�v�7K�1����Q�Ƹ�YC4d0�Yȧ��p�5��A��2��~?�=�(�-:H{n�l��B��מ�wW����Ӥh\2��]�Y��	��2qK򑷽�x���
��t?���a�^�9}!A?w6B+,<qD
�f-�4��xA�܊϶�Ӣ�p�.�Lp9����>�;������h�5s�m(���l��o[���4Td�?�(��k����Ƹ��	F��/��&�X�͙Y�&w�^!ty��>�wV���{BxyAu��
L��-��T�Z_���I�u٤(6��f��%P�҄4�}LO��$;@����������%�-������@[�yU:ق�%g-�S�Y�XC�v��3m�}Ӗ�u
��CS>���ѢM�ǯȕ#{9�D����̙�V�`) b.��m9�s"ǣ�^���_G���֧4m��r���� �Z���F$fVȍk���ܣ�.����<�K{����3'D@c������Fߛ*j��νb�=�O@j�ܱ��0��4Ek4��,v��r��?���� ���Ɩ{��������P�ͼ�@��>S#�u���]vĤ!��W������ϒ��z��%��n�B�z5}Y{w`�][��D-�t��[6)A�-I�9�J"�С�	���D
����*��M�x���Uoh���!n\���c���W��6��C���`��r$���l�����R��Ƞ�fv۸ɷD�Y)Xk��ؒ�c8w��G�5��d~��ρ���l\�<!�x���f�9/Y������gp�?w icS\�\	�Z��g����(Tz �r�~ˊeiN`%qrw�+p���'����My��^hv����Y��N�����M��]I�1��F�?�Y,����[5��C;�
���K�ɳl�ۣ]��z��p���� ��P�!'�|��d��P9C4ڗ��w>�cR�Ϲ1��_cr!F�)p��ņ��Sw�|e�'|r��9)iF�)��>�NL}G����`s�arq1ٛ]5t�;F)N|��h����#��BA�&qK�C��xx���dT��o�ffQ@0x�>ڂ�>�t����[1�+=.�A� N�G*_)nw~�f�j���)��ى�9d��>���i��gg}A��e��l�9D$���k�鏒CU��5�憊+E�#Ѝ_��G(	!,"�m�e����uJg�L��_T'��>t���h�O܈�h����� B����kIy9�y�>�CO��m�7O�r�	x����, e�=��9������)����W�	rLU�ء��k�c ��H� �4��J�>����Aax�i�8:TZai���l��