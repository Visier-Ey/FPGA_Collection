��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���Z��?��1*w�k\�d��T6�c�u�����B��E�7�<g���Ԏ���ΠM�0.���������b����53��&t90�$AQz5���*Y�,�w����R";݉aޝ060����pa_拓^d唱�/h+�<��4�3)�j-�d$��H�_ZE��ƌ��R��l�����h�B��>�L&�P��r�!��*67���t����F
'�U�����T�!�:�}:��s�W�+�-�|5�d�K�F���䳤���ARB�i�J6~w2�B�Kؾɩ�k��!�Q��j(��;H�D�|?�ޚ��Mڐ��j�bBR�ʬR�JZ�4��D�%2`v��R�L�}b��� i#5�4��AH�t�Hji��/�^���%�+�[���6�X�E����h�R���K�%S5�r�TN߂�j`�-G8��0�hu"X4)���JP���i/Yg���p���`��vi�!=4ҲTvs~<ג�iq��:�Qh��$�� v����O�mT�[W�1r�S�y�eJ��ܤ!���e�Bi)�M[�m�!�6E8�#0V%K06�L��u�h��鉼��(6H��J�q�ګ��[�]WzPdOV&���C��TXdUQ�Q�k��d�ϖ���֕ꭿ����=1&�zD���7�ۥV���(�� ��V���:4u��G�X����r����0�_��(�B�HJk����dGi��nc+eMA��[	*�L��tm��� ׂ��8�{��>y]�N	�)ֲ?@�	h���?.0怕�hmx(��rb?c<��g(%��#��Ɍ��]�j��憤o�(W���=b\Y��CI��+R���TC�7����-ݗ�N�,o����|���jYQ[|�0�qih��^�mY��J�C�ɈHܫ~yw��s�g��Ѫ�ťV�i��7�O�L�����{��`Σo)WRDd���A����D�15r�!�[��
=mPh�-��k���=	4��riQ�h���w����,9��A�S��N�������ux��6�7E�<�ζ���2���]cJFz�E�3/<�н{�����i%�;� ���ϖ�
���7���?h���Z��6�Յ֓	W�?�֐����;�KNe�_1��
����&N���fTf���cxEGbI
�HH6PxAu��!���+�K\q7�DN;�`/�T�#����Tu�Y��\a�sC�?��|��?2B�����B�Av�y_Вk�Y$��`H�TFI��_;6(殃j��2��m-���[@�'��a֗/J�`����KTOuׄ���u���	�m	c�}�hYк̧cU�~=����g�&)���Z��B�6�la(�NlԿ����g��u��x�,WIȿ^t����nl�.�0S��hA�d������P�?�S��>��n����h3YK��5��["��R�Q�o�O�2�MF�6}s�����gzJN�m�ފ��+2K�,�� !�![,���z��N2��em�#<�/�*�njA-Ī��u�[� 프��l:�&��W�3f���;�vS�X��h�ú]��e�࢖�j��mU�5[�/��S�еA�'.W��ΔLj6' ��4u���jbA�H~����e���q�bo c���È�_�$^ʱ�
�.\�wW�9_G��������45�~���?�V#u�o%��� eL�ݖ��^h�D���a�p5�U�?]�n.%�h,[���T���q^C>�ef�B}CN��^��_��vS��h��e��B��v_5�B(hT�J�ՖT��mDf��I'�����Z�&���K7�?繲N�O� +�l�Զ[M1�����dΙ�{���v3B&[}K�瞿�':,�v5�,�[D�L�f�{��v��K��1�n���j�k'�(����ѐd,e(_��
r��1��[6�
��s(�1�dX[�F��$��^���vy/�]�F8O}��,��ޝ�{u,	�#�&�(��n��ub�|��_̓a���q�~����o��?���ⳑ�}�S�28�OI��	�o�6ӽ>�J�a��WkB�����?���ӌz�"�D K�XkB�i񪬲U'���ձ��6��&��ղQ8x����У��}�E(�#  ������[`����էCP�0�5�<�^�5u��锃������q7YO���B�+4���(%���
E��/��)6[EX�ٺ���o!���}<�e�5��mV�uJT,ؕǄ�����)���>\")���Q+*`�����r��U���,��p�oh�,��u�T?�f�qސL�~��O=Gˋ��5z���+R�u�8zU3��;:|��*��Cws�<H�ɀ�"l�X��Q"�2� a���j�p��he|�J�?�K��*\��U%�IY����ߕW�ʹ�c�[��N����D�\�_F� �wi/tzP�"�<�/��\��;^��P��<���*8����4�����5������#OΩ p4�\n��Z����F��1C�ѳX��C�0����O`�t�n�˃�G��X��C<��d����z��߰,SZ���IBD��j#Β���r35��{��LPP!)�䜫�<��w04;(7�.O��-������=��B����3B�f��Ԑ#Ӵ�
�W{Ήs�S~�u_