-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
--pragma protect begin_protected
--pragma protect encrypt_agent="NCPROTECT"
--pragma protect encrypt_agent_info="Encrypted using API"
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
--pragma protect key_method=RSA
--pragma protect key_block
gpKVcN+khLmBitTr2/N7VtVP7xP4L5GAsvqyXQFu/wlL5fJwazg4jluoBSUas1lF
I91NxXTY9c8HxOAVIaw9OtQElEFXOjsXzBi3tEr3n8vsVAsbwB31sPMytymorG/H
avFIxAGGooz7lAJIXHrZlurCVhRjdTMQMSc2qaoJOe3Rcffx+vXuYhYP01H1wz3I
m3IkxAaWzK+pMt5mvNkbjSDUBmMFgd/gQ5WHhd+t5rhJxkkNyj3v21JKq+UERwfo
YGgwGnAsycI80FGPPpWHDsrrHheyMG+atD+8uAMyoYkvums/OGwk2hZ2rzM82arx
w8ycyUU6kggnralVmHnzyg==
--pragma protect end_key_block
--pragma protect digest_block
0WbH27LKZmgvlgUDTqyH8oceL2s=
--pragma protect end_digest_block
--pragma protect data_block
FTRivN93vhCre59qVmylTwQFIA0yCpPNvhi5vXfe08dI4TpRsqAbKlSV07vCpecn
bUqDva/bM0sdQvKZZvycF+wAc5JZXbCS0oWk3A+5hrkLNmTvsdEmo5uQwaB+wG0s
UbetKCANzyxIUovyPEh7EhQwTqfFleY+IJNneeBiUdSgcqix57UJm9dkjryRWOJM
/DNAOZkj3lfZAoRGPwzdMlC//wn2Q1LHmfe84dYDS6+J2Cb6oPMgTX86sXGHzgn8
pynyWw471CJjCcfmFi2XNGqY3C2SMiPTkMfz1eB7dqlYNcL1DWpTioDxN+o7X5Bz
CBdPqe1wkyO9BuPL50r3erxumGuaMWvIZeSrTXnxROfPs89YfCDvQ+eZ+2ulgfLf
Gni5HUx4jDcogsXtJHORAXnvzf4N7DMVX1iPd+2/5XqB7PZyUejz05rV/yERvizE
0gptKM4YOsEKXWgEevtGgCbJTogw77LRBYT0VU20mUR/RpXG8HWrdUKq2AGGS3Pr
+TXXzJMEBkTVkAB4tR4f+txHOuyAfilSzjEsK5q4Jyt0VT2mWCBSSR4qiyDYurGF
Ly2LBtcpHmtVzH3zEthAJClS+cCazNBDeyB0oEnM99R6IgdDVQ3YTegsl++hS8tR
FCKgt2EWFIr/hmJYR5us+QaPG0xNPsb0LDPU1eDBWHWMvUGp6JAm6sE7mi80VDpL
841r6X8txKffuMbRS7fs1gk8r4SnjbpOhFesk3RUeLP7A8y54t/TUOUSFIuKOc0r
qTbx/riAFKgGnX1+KhmA/ikZIpQ0ky7Kzmzbo4gBLkQRZEwADOLTiCou/OifKRjG
YFgrtaIdS6iFeYoOJgCAOE9TmWEBF/CcGzGgeFccLV8nc+0431QKZB0J3BUF08J2
YTeU3SzISiWCz37+n7G9NvUB69puwV67a8O1Y3F9rHiqLZIyOoYSzSh6AJmCI2EF
Bt9/gXi3A1OvzG4Cp8DHPOYBPb47sfTPjz62wzy3OP2UzZZwAwVg86AUjA5Pl9e9
GNZV5ocC7WF6QRbwJPZOWlVQWivPy4t68y0/nNSdY7pgzBN21PUNYsvWK7meZwSh
naEVkPmPsqPwyz1xXTGOBCff5JZo22ogqxb1oULB0BK+4tFiSrObzBCctJjXt+AU
5Rmo/y/UIOu0cK7l25Y7rnNsMX+cHN3p6ZhcyIfOr79Pq7NbCCJPc3pH1WBDumZQ
hbj9mawj1Hf0U+rb/9xOwU5GPNkHR84zmTK93xR3YzLqR0nDTwNNoPzPA5gLr8+o
HUuhWfg+BQYvnKfxvG/3bGiWnmvmRtLX6t7c7QOLiSNWJqF0B9Nu6WCbIVQx28uN
bgmCkdPZxWaqcarnKTRi2eL5QouoY31gfRb1FqvyhTBDsgtszzzR2kqsANobo5Uk
e1dIuHuNTdpCHM5Vgl74+MKSFjAhXGVtfk6f8ZshdqN8aRdWv0USNo7SgLtHvCAg
4ABLaEdrX75+07fVm6znGzMQGb9ZYr7CfYPddjPrIgB9NyhK/hMtUXKjKUxCVofR
jTOK4f/hbLbPIkrFL4xost5AWEataLz1CK6Y8dh+gRvjmD574bRm2lLPuT3AlE0D
NvCGkNUMu6IBhrA1L7tBKRTXuJ0ZBFA5oqKm/3HRgu+uvhzmIi0nKnt3oipVMe/F
YyKPxhM9DITfQCZlFQEu7AuK6fWhpxgSzDjLvm2BpkSxx47opFkUvRrz8KxQI731
KHhIeCnamF+Ix3sM23KUlR3OTSQhm0NMlqeSRxRYnWU/jAsaeedPqWoaqicgJENN
nQOR/stLRY2kA55yWTvmUSoMaYPxAH1WECB5e0dZ0u99sISgwIKnotTewDCqjdaN
fcSL6qaGj0lvp3tM9/V+p4FurwzJdH0gB1mYeOPbPxjaTL7fPFwGaMn+MiAx1gZz
HsK/OMChNedYaBYKyjPE2i01U+8PYQjixOMTi1w8z6Kn9dnv0lypDuU+pAkJzYW3
BN/7xgf7aYGctr5tk8us05R9FQr239CTJFjpVpc6qCOGAZP+EZevn8J6vqpwHd8H
Kp2/AMFDvR6FpH9QPbjbs1QHRfBzi/dHPdLN/lgzCNq4GgNDIx84LDoLiEm58SBz
tjt/wAXC+stoKXoI/CpSqSxBOICMKJwPbnSluCOpD3IywsRehl0F/R6f9IBMnutM
CEMeF8kQY4cognYrsTp7HAtbVCQPS0VQd0txYHqSyppWyboFlASZZsklwjYia+KV
KAjs6Xu7iFXQ6T627yet7VAAWWKaG1z+GGWVLhb6AapjOtpn7dZCSrPUY9b675vJ
U2GyiBlzDG6dBsFTGhWJhcx1ska/UU3RP8yfPWI0+DKYlOiITTggzHBLMcKNudXO
rnZE9OsGnn4oO4OjzvpenwHKOXn52qVNIc7uBGGoTKf5R7pgovZVx1umZh3MaTeS
BAlDq4gAQxxSrlwfFRDAEu7jHcbR1Jd7M46MWJYZczmi7nM+j9L5xuaI/lb8p2GW
teEY0AS07eNqsT+f2Dwc5p7zhs/Z3FDTMxo1r6ogxcV6bcMY/DzUzJDeMRqtVXKm
8Gd9QPdjRlW1pfD8uTbsKTZ6C9NJO6v1HNV+8rEF5auLchUyfEds/v0faOl9S/kY
Mn8II4U3cwqC2DLFxUhqN8ZIFRX0cZRvSJLMmQLjzt5xLQLelymW1wHLDBsVkVBR
YmJ2pclnIzwgTfqOP1qlGz9OUHly59dEmvusG9amzNN1L5DgIt6tpJnbKR+eAhfh
xTv5vdh50+fRLw/SFQo2BPVDBqTebdWhU9D85Xl9GVJgPP4flNPht+viXF5uCqfw
hj2sk7pfMw6fdrG0D4fpmUkCyniEUZCOD9qqOTWHHXCvHd0w5K/pWzusiOiai3u1
MTmDVqX+sXAU0DH6gtw43wnkewK9x6Vbvr0QTml22ellYgmLiBMzW4V6FDHD29II
4DpeIL5+WyUAnShvd3rfCEK7rC5rpu9YGRmc8AkdLwRZfZMtncLK//jgb148u8d9
zD6wVSVs30yLkXUj91vmGD30Oqdzvn646ghU0J3bQtjvcxSlph2qYuhb8o9RSp0i
d65RUWRzMehgxQNGfPU3sqBYckK85j31BqRFQhGez4diCl6bOeog8fPdk4CJ8IsJ
4pOKK6CsD/lo1n2VvKD/ouIm6MtuzIywAFdpMHWtNrH+ZnkMA6gJytUp66/XdgWC
qhPjqMWMvwFKG14jqVH6592U3/bEnchB/Q1bF02MKzPEkLEkQRyMupIllPNCPvFo
QzyWGM0HDB/VVRxFT2Kf94+8F+lB9KE0RXW9wTR37XIU6jFqlcYbAtORkpCWIwWX
c54LFVwnqVc5Yqlkt8j8tSkIGNWDVpAp7jAdTUsSgbtdJH4V+BlhXd0JOr045Imw
DV/bv09MIUD3epUSkmK22cXsTEItCnOiW+7GiNaBmlLS0Muq/A/5qhvE/zVXUApS
8QjBxePxva8dGdnXDjdk8h/yTIt4LL7eoaK6EBv+AOcUs6511mB1bbWYK8pNTKoV
o6Mh9giDegDmszLlulmQLqRbH4uqwOAcLPkxlhZ4BYkSZSnuY6s1xIjYgpnmFKnM
aktDAp+3ull/4pUHMIA+SlxkBEkLMTrIiMzvDzwX/TBrbjuzZEN1+XzPeQveGO+2
/+88ycbFyTjbEj8FFk58xRKdF6YV0MY3TfQJT6/zhLOInbA90DtIE3btgVGAXARU
OmfaKBZyQKPgh6KAmiJdtFpGt/avvr1KZVM/MCm8ydRtCMzfqT8dANjfrpi785rA
PMCdV2RRDOJyVwZZSucFmqeLKT6re5LTrgJc4NVZG2lpg7s77cicjr7yy7GjLgcx
P81SIfyRBSqA95MFL8UTiaNkTPpUYTxrO04HLuRsgyHsQXVbBSgDxVjgnmfzADwP
KYhP1XU7c234zrO0krRJw/9y4RggfZxbowbkNO6wEPixlnW40gAbQGGUomDabtwA
xz+AOPhWdg9bK70p2fvouZRsn68oP+0KYjTnp48ZGHydBRBNw0JoCDdkiSKJ1yFC
jU6MRbS325opiFpDte1snNCFZANlUJ3+a0+Zk9hhga/tTeHK0Z/EQm/B0WMrOiyO
Uo85RkWoDzqqpWHEaxsEJd+R+yREYBd/QPWsfr2uj9+sMwc1dtqrF+K7AORL30Gf
DVZLKtBTy3Eu8ZQ56klW2D7IXh3OtgnfmiRJSJ3qUeIRGc/z+uSMIKdDJCTJWUi5
IcV7hGAxpQXuGGzbHWTLUf37WmuRZvoyx0XDSWbPEvviNvGq2enbIMcGs6N64A4Y
FEvaMfjmjjHGVTghp1t9OVmYfHQny3lg2rMvd0Te3SHvi9qLGv21YJ5ejb5PZk6/
FYyl7k0vt5oeMV5AtBAMUe+VQSouCnJX2pcjy5y5LBoH++6QTUFFb5M7uwBFA7si
BDaq1hpNTsAcEdCYSZu7tNMWMjKhOuvKtgJgkFtpfE5kRrwOmKu3UExfdroJ3h1n
EnOMOu4W0iagYpN08O78mSmblXYSdBgKp7ehrWh6Xv6DpDtpOl7z1GiraufW1CyS
97DAN/JPZ8S+qFAoj5zKno5X4F0PjkoWohStUVYMDoRmqEmrrqWYlLhkts31l5X4
aWA5RELxRu09bkiaWr29fHnLwmMabYQeP9Y0GatXgIDRTpETu+3eDF1Y0n3l+2PS
Wzl715IC1SO1CXqiB30FTzA3ItGHQnimwq+tKTemsOyH5MNQWqYHWi8M+NI5j9c+
d7/T6iM5DAsF5aFhbjXDt1ulVMcVE8HJYsmQgClMUWBDmxFkPT217ZfZ0GhHdBoo
v2B8DSfB9TkVAlx0VFHVFjhzEWatBKxmo/7fq9rr55rBeeKG+r2WmSXD/tbg4Q1l
LvE4b5seVnPAEKdIEvWNYgL1H9zt1piaD5/aesj58PHFsv/00z0KEGycZEAjL5p1
WEIkmVdbsm1UU6JJM0Ullk6ODkeKl177tsmZzaIbPPzN/oXmuy0NgHMH3sU/Az28
/9g8fRENcajUpM+wrGllELu85jF9//oVCaoLmPsXjDXb3aG25TbUqgsAmX1gWxDC
glYcZGn6viWoMqNi32ccibTPg/mdGfKmCHtpQrrxcIqtHWuhZRwu80mCI4ry0k3J
VLdz3LVgBwBIaiP/DrKO38YK1rr8GUa2byEwzcsVuvGRS6M0DRbkouiMIZIyf8fH
TJtCaieOSCWQ7nDhm7PZijeEwJ7/jGAAc/OP9r9LTn2vXYXfNIX/15hx1PvWnEKi
Q7N1z2t/zxOGsu9IodtEpVsCF15VMxQNanU11iVTsqk98Zg8aahJqWCbASska8pF
V0irn/7/YcIiMFXxAYIqWSfVTFMQ6yoqB2qoWojAZgjZjE7nM/snJYbBqukxOeCz
n4h8+Bh+W6wClnvUAja4CFBdLtqq5CsV6eem4zlNDgPp1olGdVbJQ2qmIgOybbV/
3Tft/fCPtorQJ5T351n26Y0odzXmV7M30H1o+gDwUx3JKldwfOXJKSQCXYHXMPGv
Zwlz7g3AdShHJnvpTIzCqS0P+4tkMnwXnry3Im3c63XVvb7eBBjQu7kdXe4j2gzg
KrvIk/n85jXvpDhxLxn0Ww3hhF+qnjbz2BxF3zr8kMUpuR/Xh0t/XjvA0IHCgYrg
a/aMIDdpx1RLRR+a6XieTDOZL5f0d687FtMjxogojvLbD1cuS0uPPXh/TvVW2eSu
mExzn+9Z5SgAgQqhordyFDGcq1nXMjR/SQVOliIx7XP4ETKda222i5r50S2kjrHO
Q1Zr6OhInlTyCuqGaIZucEZv8KmhgyO6+j5o5PFy3K7nI5wwSjIY07DhJhL0nJOk
P7gxQYWIFLmlCNt4x/NMkCF3kLHbbdECeUglLMcmHZ9CSE49Z92Co6oqi718E0ha
n5505y/I7ZkQasnTSHNZHjxjM5TThcMog8Cxpk4YpcX3z5jPKRFh9rPxom24l9Ot
4g1uHlCfhR8MP+ZWXEVqjW8uwhEXMHXvQ2Ntx9raH6dBs9ZfPmX8lCZt2MZmFpn6
aA2dJoOE7RNuzrKuStBEd54/cEUcE3oRC5eIt5d8bzeVZQA6StRwOIuG5+pyAIaV
n9Xnhrc2AZnpBhhK8WUeoMCr1MKv800X2liHbqWZHdoq4xXyySWxrp5yH+NAgMZ8
nb19Qm5SAx1R4wwZOLkEKP/bzEMlaU349Xt0WbaSytrdjXznGC7pfhda8LDEAJwZ
wdz6n3GKOy+sYu71MT3OycJwBznahtUhy9RZ97GlFIsw/83qYGvGlNSfGUGuShnt
/1SfzXRdG7spDTTRF7OFzAQn/KfB+RnIcyJICVKeqMklY1slvkIIkqsNnBdkY+n5
MQ0DEbtSh5kvMiJll9LeUpv0FnoY65avtrWPZyZcA3Lr7+EvZYO2TSBesOx6/qX5
Zrz8IUNZMpf9FccGoC01lcT+cepAOcK9MVlmhYtYkfXcUMKPmG7MisKQwKtI1r5h
LpFCinrw538w8Q4tWsJR45B8IYzumSoH1sohJukvAE+jhD43IrVyO6kkU/bzRsFX
+LK0rHgj0pChyvaDY6tMlEjVBLeXNt02hkr4yanAaYM3iMQCIY/jQh77ZybgP2LT
EM78j1PHOdopO4muVeekMrdUJwJsOp7cwlrjev+7HIv20mUGuns1l5w+CmtO14rw
jKtqei9zF32J8ckMe9xiavq+v58Pw31fScvTsFGoV/eUBYjztua/Xq80khBzuJEq
8A5L6uI5r7XryVdKtkxI7/Da8Zksj19cuRwy1qmMpGKKOtZ6tgDg9JhRnx55wBWZ
Gk6fd0DuVi0E6nkr0Hw837vz3tkt2NhQzNA+iUdBsrFZiKmDWn39pUuYCA+pELIq
9MbckXaxjNYyIN+bb0aSyCiUToeB5iLfi5Grsrh4Y9kbcUisk17kpNlFjQCZPDxE
d+F5a+MkLuV+W5wrOMQKONSP7fHGtEzU4tAHoAi/YnevHnuf5Mrx5LOyJNSifJk1
XxLBehIKto5gfuUkzhuZbb06XhgLEjCSFdJvfY/RS5wxt+VaRk9TJf3HqonFLeWT
eZZBps7tnccqJQ7bR59QcG0L2WIoV3Aaw8L3Ovkh3t+3rlYQC1tI9cKp8hC0ena8
iu3RblDgpTTS3Ya5SmQr41ycc9IXvN13fUihqG1CT23cD70oqO8eCPm2+uOzTsMa
VYOwGRx4X9Aop9k5FvJCwILjItFfS0kFWuqFL+4+MqY/YpTfMLbk6DMjbdDaFY6f
HmZCni3VyQbtkz0+RA77UbaIkvXoV6xTl10BfzsVtffe7XMD/6Kzg59xJUaq3xEx
Pg49DxXiRuSagVuIWko6b3x7Mx6et44y4z46wfRHo4l6FHls8iF+2Tkp6lLK4enr
vCPm/eyNJPZo5nziocB+5vOtN7rPUtPXu5YKxO4+kkaNzxDbFwcoTU/hhTL4ly/0
C7w9tAtkqMWPQ8iz09UtJw21iQq4OiWKvmdWOC1S2jqB0xyncNMd/Y0YmAfuA8dN
eg9gzvv/XKPRTZyvUdjgqQic35cm3Fq4Hhw+nWylNyEEho8TqooX9DM0xB00ZISS
Fq8paTaReWIdoYQtIUZG8pBBjH4bBBHkpX9OXwI5zdhF8HXe3tvfHJwV+swqhNKS
ZG5CRJxvJA4INz5I579AFd6FEskBOhDS9GCtlNTao/UKpwgBAyOtLCVrtr1/2xp1
uUsP8DLRACF5x/Tqocu67BlULJeN/ycyQPDSGXxhADkg8xHQp+ybRj1hsEuJDiLi
CZghYN7nsoKR8sEDo9G2M7MgWs1mr3qL1my3AlDo1/g9mU6WDzwGt96t4tInxiq+
Mc+nUXRfI5ubYKKpWLnZBMFdfXjUviJLAqUvRPO0VbiDIT2ggl45ZvvXzZG/i3DG
a9NNsHeM2jAvE6CdAnsxsRXa/E6TUgQOmTnComfZSPCdQooDQzVPYIfQaeR4RdVz
/u7FlhUrpZsyMpfJsGUFOu8E4getpoAvS7a0EE7Gdx3vnLN5BBDZ9WLPHg3Wp7SW
84h54vwChJbx7JyXdeNCR0bwwkULiNjZC4fePnNH60nKXRgTVgLyXSaD2XquMjDv
F0MbuFsF46bLAADuldbb2qgdkQvqXp8Q52A0euHg4HCtf1xFykkmJj+KHcR8lIFH
cwK/J1MJDrN5Ahn2c+OdrMOpZ4EDpLk7l9yJcvjfQB1gFeInATejprULtneXAbNp
8k6OXBOf6DJu0/1RHnQZMEyFrs9WkADXjtydqSJhOQFlapyR+bsstW0fmXW5hmx0
GI8zbUQFwvOLiHl5Iaxxckh+u1iC/oEnQhrJxd+txgYimOzF9j4h4H1gnK12KDGV
JlOwtWWiOBtB1Gsu419Z41WB/9O7F05xVdZj+xD22Drl8AvYvkl9tKLtaDeFzvyq
HwZEIWJvlJvCggvHERPiAETtQtJIpLypKqeDu9xZ2JhruB+HOmQ3rBihoY3lmw2j
jnvLR4Wy6Cp2dtceKkvthrjlI5+O++uR406LrUMwt8tPkrwyXPa4dSaPKORcDQiJ
1BmvcW5nk8esK0LabJOmIr5bRMPyFMWB4+7l2RNipX6zlRNw/oI1J3CexA7+aDrc
Ofo+mQ0xCMDx96cxGnnnTY9kzsMXO1Mr/13xWzy7p/ZgFuV1x607sgMwlgYDdnnZ
GzL4Q1eBN4Ma6OwLnHkK0OEiN3IqT3lsRG0oqefnJZrWGhNw7ao+rO84LVL8orCT
omi6hqxI/L0Qoef9qf7AvWeRc70sxjLJOzVqGmntMT17VLFS1Npr3cZdCQZ1m3vL
p0Nip9zX1QZes8oG8Ji1+zGEQRHBEhnBa9E+PfKWLWUiniuykJ/qQ4zVs/8PLVRz
4H64mtOoahTf1Rci3+rUPTwVPVlyAidgAAyAaK597NiQ/4jWc73XvUOa8FIRgLA3
NS8CMaeJg1Z8pi5sHlDrCZWzyS/ZxOdj/2M6LvFcR78Wkk3e0MGMND7XuDyf1PFH
piIy1lpHxvInGUc1KALxmL8TE23U1rRT3SMf2q3+C/W1tomk1elYNkMqVejSv67E
wMk2r3vYGyke2ZIR1plQip0Ka4qkO8N17QWwVtQEFH1pFAHkY6vizW1cUnIDs0Gg
GeS1/yyDExzGGE8LfHy+RY6CbOfvsri3dwgdjdgPnZeNaqeZJYIh4uBGf7qKCO6o
vNA8/+/SX8aSZ/UtZfVNjbE/G0Udq9uXwLLJfLFIsyAGzTITEYNrFdafHx5R5j13
6/O8yCOCm6UUV+uEXJqLKTpEj2FBnsx/MAtI4Rk68oJcVrmKP4gpRwe7ZCNMT0Hu
7A9DsVIyHD32/Lza/1WgZLxXJnkf9RlO0JrWleE2bl7yfw1bdHwILUr2fpkyq2IR
O5b8BKAnhjwwQi+yUt+x6Sqlw/YGcxNyC0SMsXfJ2A9rt1zNGJxfrbF6iVaqt5WG
mF5kycyq7LLKUX5287teZ23NNltyYWBU7mlt0+2s0Lu58SWRf29XeNyK+Y6HMDvq
+eglEJ1aPawJvFf6Hv7kTr1P7/B57tOxbwONoi7PH12SBBoRAFMUlWI+RBZ1B99N
3jwNSnCAd+UJxIbzhiY4WOoia0zdDN38Df226gDT5qZogHG5Vzu90SJMkR85KQPI
pdGAlW6UhzWJz2zL+kNVaEi2McNgzfZsLJsJhMHamwzrKHAAhes4QN5xm+LH3RMC
thE2Sa67BfaengPM/FsRi3L8uCKkJgFzkgXdMYWBawk47ibfTxGtW2NlVl2MOvTw
n6ubq3mbR/LhF7OEhaEoQZpTPXPMSIersciJpbVmiBo1G0GrG1j02kor48hHs2fD
EV9OpBOsk6jZ/Qsbj96sG692PbriMjZo2DhVr9otSexKpjWKjwqCx+0Fx9/GeM4q
4M16/JVTlI/QIuQ360XdN/HiUW4vMZA3imZn7UMg1u6/EoI/pFnuSkJl8NIAnH+J
0C6wM+J2I2jbI5QtxpBhEvFko0F4y/e7OHHiiv4chosbCUCotIi68BVbA5bhlAEt
L5E9jK7lM01sMMhFiJk6FB4OUShdZk7r/EmOSNLUfkUlH6GW5wv5HwZwEuSD9KO6
ArPOqDbZ2s7TIVpcDTquFRf+xNXdMPi7JtH+PCPOPMf5b7o7+u8iSdOlgphHTfJc
rV4UzzUE8LgrwFrdaKZ/81F2L61sn+Ne8InfdDvQrqxMH3+eEGZRjbcJngVAg2gc
s0/qb2oLiQfj6Okk9OvC57n3A2tWxKUWGXc8gb9QlLZBUd9WSkmFrbfkTpmb2B1Z
tCS+SlA8ClNJ98nobwvRYo0desER2q1u265M6/oiaho8OMTMt9SH1C8Ttswy/2Ao
LstyqmulybPzMdwcG13gZiv/qPBGWaJtYJb8w7D7I1Q+NzBrClk80BzHGGmA8pjY
PbXXmEiB7eIjAGd6ObpYglMwb6UAR0VcvniqxOJhJzjqGNl+oiYHnVq/i+NQdumt
Q/4xnbuaN2TNgtK18uN2MexRyC/zI65003B6zbEUvjc4bPiTbvgE1m6al0CNiBX3
RYoO4x6gq4SxGjMcO0AvAZn1yC4ZGK2Bus78wD2332DRYwu/Qeek1kvSwpmzZNPX
70jhThFmq0lQBqvVYl0srzI40b/yaYt0LPfUEr3agxBexLya4rbnCjmVWrebV33m
RtwjzuhiYFfjTpGmnKYUOs7HeVgVD7a42uDmLlVa/1xbHh/hWgy67PjYn7v0Qldg
lxWdjLVUgaD6uBVXJAN1wtwTKrakcRNAQzAah8tH5g0Mts5I1Ip5eBetRCmPmDE7
t6NHRm15mxL9Yjx630/kURW9/a9XZQQFY7yO4HUCsnkeWLmmWCKvycM6aVIqApmI
7ZDRs6V3HhQ1OTgebz/0JS9CeMRqFIxhoeYTMCRcztZCPyG4SoIpMPrK5jrJ/Lr3
2pwZmAesIKFK4BgYGnJ/KZRwSAxSP91hni75wRTbImMPL1xeeq6qUYj6o6fLYDcz
cZ2ffjMlVh6zHPuqgL26YzYHRBt/MPqqt96+xQ+YjieVxq4+IVEWev8zKIL82qNr
--pragma protect end_data_block
--pragma protect digest_block
wVVsGSCllEnLbih4B4nKnx3tICI=
--pragma protect end_digest_block
--pragma protect end_protected
