��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F��������n�BJ�F���U�FW9d����T�+�wt3��^��r�q;\��af�י,��9NL���ٴ�[�Z��^��Jy���0�T����l|�x�5#B�o* ��J/�CO������|�)6b,P;����t��ew�u��5�v�u�E�8����R�oIk�����Wb�A1���5��r�5Hڜ �r�n+��MS5��n��þ�|R1��������E�%��0E���;%�6�׸ۈ�6��:�!�#��L�jT�a�S�N�LS�[�&Ϫ���]/��nm� 8K� 7�H�be��
@��1>��?���X�U��&��P4
��J��tz�6�^�O�A��S�������EjS�V�6�$�g)�H!�uA�����.����c:k���:J�G�y�*aio������6M�pʫ��QZkw5~��ΰ <�z���i����Y�T�w-�q$��k�d�V�5i��[�r6t�`?�.�^�v�
��l�;�y/��y6�]*T�۔"N��d�V۬����/S[�B�U��7 a��p~q������~�5�LPؐ�V�T��?*�ؓ�C�r�����	�].o������߽o8+\i+�`K��+darwEi�JI��4?�}͍�<<�,�j��'��u��K�C���=a�X̉��37�Z?�(ȣ�$��Yl\e���=~�Xa��s	 -~����w�N���,v-�xa��$a2��hA$]��g���[\�7�x���{�MO|���1Wc���C��e,m�"��$�O��
	��M_O�~���jCL�"����V��P�h�Jm�_E��HaT0CS��&�L1<LJ�ګg 9Tp���N�Hm�}r�NBa<��9����-L��s�/�ap6@^߇T��!�3��`�[�� [ݭ��O�>F��� ���&�	��A�A��.V�Sk^�%�M������P ���v׮���w���>��!S��'ho)�mRv��� �=ß��;��!�����=-�F�'��-��$N�9_Ta}u�~-����jL�(�s{1�Cy������[9o{':�����C� \�(��Z�`U����;į�n	��o:�5Y��uU�b�Q��+�IY��,��[����M�&����&��D��G���.^7�L���l��թ��)w�<�癀$E��o+�q������ͳ�q/�K��:z�j\�w�i���S����t.�j���g+���˫`^8�e�Y��|�>�}���#ݩ�x�"���:M3e ��4E-��NuwE��5�Wo֫��;J�AMHː�����R��nEԧPJ�z�֒`C�@�@�#`z�y`�p��B^'eU�-�_'k��z!~5���H%g���)˔\dS����*��y�C	�x�9�(���T##T��F7W�Y-��
Rn �Ruk��S��� ���Phݑ|��fi�Mu��סW����\�0G+�{��k���s���)GTc����?�j��>=��:��g^�Q.�3�� ���-n^�S�/����^*o��^��]���f	�֣Q��l�W����
p%#8ҋ.*��ݞ����J�����B�gG��(��4�`h��<f�:*~�P��naۜ��6���}�><8R���M�0�x�[wTq:�3c_��/:.�S|#R|���Fx����Mɹ�ٽ��ƙHv���eQ�VR�B�Z!�[u��޴�0�)����N���M%	Û�PJ�\��?X.?:�����A�r��P ���!�<u��+)x�9���l�� f��{J���w&�^�>"QWl��D�������嵖����f{�ar�fb��_����̀N�p��u�O���>���3:G�~��H���X
�;&����6�aO$J�;}��t�4���� ���r����3ymmȒ%�*~8r�;=d�ճ�j��~�D�+Wy]��"ϻ�GĻc���4��5�ͮ�A@�Ɋ��CLyWKh�pa�{1ppY�_�'v+�Cg����M��-�ְxu8�
ܙ��)}k��*L���:	���_8h\4��"'$nd/j̈́u�N�`'š��3��.��sZjCC˺�����G�@G����n��+V��@����i/Z
�?n���ʼn�B�(6V���������ae�:�1�w�Vd�Op�r�M��8��]Vyҏ������������$��Ņz���e�Rv��QH��w��3��2;4_��� �A�'�q�MS�]#|��C�_; ���gu����ۑ:�B	`)� ��oT���8��gdd(��SE;�F��!��/�;sB���q6�"չ�!�Ӷ(����đT��_ cdH�7і�O50	%��X�wKX��wY�]��*yF�x�E�zW6�X	�m���7���1ș!�	�\h*�S��+3��"�^?��dE�P�U9V��
LKq��~,;;�e��������(�0O𥖒4�y�)Gȣ5�t�j��`�B�����F f��]i�/S�Θ�7ahC�4�}��H\�ͫ��J�ͷ���߰�N�D���^6�;$�=VS��uh�#o���#.�ھ�c�s�V�, �V�AD7_�t�i0X����ф�1 ��v�Q���o,��-E�Nc<��OJ	w[a��w�1/?�l	�g>�bmy�c92�����+���G�����w��~�0ÖP��@�7L�(�$�{V
ph)s	�L�[z�gj�7�m4:
�=v4�;�W��np� |h�7��37�f���C�w"�˥�}����=��wM4P�"cH>L�C��s�)�P�0��,���������e�-3���������z��t#9,bz��l-,j$T
Z��?y���Qa��Q�S�f��X�h�0�L�{14qR��8�8F<�n�T�=1Ԍ;�vG��<��
c������A���Y�|m�}��+Æ()ox�\��τ�����|��0m�5��*J���������s"���X9u̌ 3�z'�-1����qg�zDw.K�����*t�7!�}��κR��#���`8��wR+�Lc(��/ܣ��M���r�S���<�+��)RϹ�1W��2$h����nl�����4mH�A��X:U��*,%��V5�!�7�K����N �aݒ�f��)�a�|��[W�@���0�N��̲g�b�+�~B�A��r<��!�k��������Ͻ]�Tm�kl�K��뗣�*��m$8p-Ÿ�&��Q��S���hЈ�ƅ#��#ϋ�Ϗr����q������e�djS~Ɂ�k��ݜ���Hm�:bP1mB���EBƞ�T��.�ī��w�*%�E��PMOY�TX�]Ʒ��L_�2&��	L|�Vbv
v��4�<_�pC`N~bvS.�p��?�������N���~�a��w�ի�L�G�T���M�ƴ959�@t &7�c*)�qi0ة	�����|�چ�$�7��AI���K[;��F���x����"ʸ�DK)��m�/��x�:�鯐�i��MҦb�����ﺁ��Pl)}&�(�}moNl�7��a��x;���s�&�4O��7�-�r��₡�{��8yEr�y�L�er?�H�|�(7�t ��������~7s�Ovh�z2�G~;7!)�Q-��jx�P����O�CAHPȨǲAn�(w?b��F���9�N�/�g1m�w|����Kl(�ۏ>�<&M�5$�x�>x�`�$����H��0�=YT<��@�h��{?;�����p��=��1+��c��R�p]\�hﾦɑ�( �0Z|��$gCI9��J�M��5�(/L��,����H�۱+:�Ҙ��_����H�dR�������_��Y��:R�*J�(4�#Z#G������q�Q�,+����j���B��W�zL�2�� �ʼ���i��g�g�y���"<�v��	P��6��*_��sVt4��W�F�@�m����/�$����YhGT������#������d�L|�Y�w�����%��b04��Y��DR�[*W ˫,�K��H%M%��o�� ��� �V<V7��7��Wc�;���ǁ65��Ї�0-Q�8i�P��n��Ӛ\�$Ǚf��Lg���s{5^�ǉid$�l�9ϝ?�+{��?Q�"��Z`�c�+�)�t��m_K������Bz⭼s�LMD���M��յA��+	jBb�MRӛ(F���D�\��ޗ�(��U�4M����!��ƫbv�d��>ܞj��M�	 g^��W���(R�%�`�q�A�֣����R�ihz�s9$�S3��19�ی�~�V�Ԉ��*��D{;�vSC�i1{n��s�����b�?!�Rq�Rw�zU���������J���*sR�s�%1����1�oCGfe߰4�m�p�G�B�!�O��	�v:����/#�5����VeF�J�#,B����d��JB%�l�̈́�0���zq���E� 8�[�`Q.�q��Jl��6�Kg��{7��f/���+ �ʅr2��S��f�"�� �AL"���h�Ä>�+Z}$c��� {��k��������T�:��	�{`T��~����ѕ�r<��{�?�[�ڸ1)�1E�5'V��4����CK9ܞt<�N�J^��I�Th,���~��L*�+m縤��}�~��B��)Ɲ�����+����dI[�	6 ��}i.���d�j3�M�-���;�-h�=v~5DHA���ZhD��n/��kxC������V�a���T�[K�ћD~ӳ�m����D3�k��e�!�-J_���;]����^��̹�l\ǣ|��<L�J��#��#1x������)u0���~w�܌F8 �1#����'r��y��6�s�*���4�w �E2p陀�bL��y�Ń��,CCt��_�U�K�Ʉ�]C$�4�}��2��h^r��grȷ>���ۊt&���:��{ly%�}�����'���̖���G�<� �/9����%���?�A;�s�vJщ��զ�>G��������eٌ�A�i+��|����h����k<T�Zl2T����q�=�X�3J3O�wW�	��"T�=s5S����J�:��;96kIV��ϝH8x�0Ora0.�;�څU����7��L�w*��/�~���wu��"�)��Y�N�;�����oI��_O�Y�l<CR�͠Q-�N�0#V�2��B�C��]E}�SM�����2B���=XZ��0wT�e��n�|��9726�s;�m�Q��]6��$�&u��Nq�c,�J��z�Ӹp�%N9]����-DH��6�b���wH8廱4��g�0\C��ޜ�F�9]z�e��O��8##�5����0��oLU�N-�O�շ��a��$L(�K8�{&�Z���\��co�
=�3�xbH��ZD�ka?2�e��������AR�G�X�N̽P����ZiVP�@L\�����s��bXW|'�"�V��	=�ǩI�"��X�����	�W�����lU�Ф�-������9h�AZcgbL;9�vI��KQ�?P��Ӊ,�Dz�6R
*dUp�:t��w5��yap�әD7O��!]�2���_�{���HPK���>r�:gЪh5iI'bg����ɡq�ʯ/s��k��;����ڌ�,	DG;��"@���*>��@!�]����<�ƚ�����M��{�����My��d\?/��_��]�UJ]�" ��ԋ��<=�-@�f¾�*^"i�Ёs�d�nOR��� >�(�g�ѕh��M��V^�P5�/����JK���⠅�8o�Ț<�Şl��QF�7�$ɲ����=�4�E�?)�~#� e�(��A�V6%��0�e��|	U�|��ȓ� V�U���X)�Nk�w�FD��-$�r��)��#�0�"���LY0��!��a����1��
r�R�b�\#��8���y�E#K�(ֳ�sKU�~P�$ژ&,�5�`4�3�G��߭f��R/�V�G}���P���h�1|$��ܗ-N�㙕��@���<2�u��`'��r7�U��k��C�8�g:��§�!8T�0(��	*��a�_1f���'W��h�%�<@=i�/�:U>���w2����͑�7�m ;U}�B���1#x���';�54I��,��	��OU�5m�Bb��^#V�`eU�r�!����Q,[�
o�1#����^R�*n�nX�k��d�|$���,r-"�l��b��%G�u��=�[~ .dVsW!�h��'J�)��$�eb*K�.���d�����,��+^D�4si���gӬ��_&�q����^��*��"i4��K2yD�^Ϟ�65N3� R\�]4v-��� �޴�}*N�Ǯ ��!����"f!�w�Du�%� L"������5��iɬ=����[�[�x��\M��ǎ�Z�/�.�R���㜫ɥ�����*�yT��u�X��u��/×������يv�d�1���N�\	�� �"��5^5��%`���:�ބjG��**�c���_��Ε��[�њ�����'��,R�f.���7��ð�zBw���[�f��D�Ue�0�ܞRF)i��+��c�P\8�T�n}.*��ԭ��pW����{'$fv�IA�C�@]Gd�qOs��>h��y��Us�Ι�c����q��ds6�����~�AhRa."ܦ�n���N49|�W�*ZV(Ե�b��J�z�]�.��6�INz�H�1�4K�C�c��*�� f����A�a�UG��{��.�����ԫ�Ɗ�
Ȑ�EIP��f������cf��z!�{&�ܘ'y�(�d���Gk�]\'��H�H���x+@�g�� �=��m�#^��9�s<�a�������E�K�T�R���6�Щn�K�j*�l����ҦiP�N_��(��{���)Sۧ���fB�(�N�5%��"� ���~*O�.g�Fy�i%�j|����W0���Io�#���Ѫ]h���}