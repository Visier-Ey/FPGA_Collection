-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
--pragma protect begin_protected
--pragma protect encrypt_agent="NCPROTECT"
--pragma protect encrypt_agent_info="Encrypted using API"
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
--pragma protect key_method=RSA
--pragma protect key_block
U+lbJ/eJSHMIKK+m8AY6uMyoy4umlri4Jr5H0957GghVLHEnmM5w0pNKkj/2WeVa
h3Awez+1wNIuIr4o/EVYq8q4bxhjEg8RecWewS7RZoGU0yX39Eh6jA0PmpiZ72d4
t5fcU/jsy/TEZmbKR/r0fjE2PflWRoY/Q2ycqSOUcsiuJDwm8ZgIvcIsWpf539Qc
N7REnpySzfpF14DWmKSLWj08VFWNLof3ATAanRm5KZeyB2INb1NMPByo8Lu3Wmue
P+XLzgAGW7TGulen3ZLSRzSo1nGaUbagPvx/ayojCS6E5j766UYjfnieuW47yLIP
NBHQ66sGnGDXMV0eH8pz0w==
--pragma protect end_key_block
--pragma protect digest_block
vNRwN7PR07nIuGRMRXMX9EgJbIM=
--pragma protect end_digest_block
--pragma protect data_block
ZIobVGJo1zyL9fY82dB4qPVWuhqPZh6nkJRBZixztoJ+fgi0KUvi+7chEdu/amlR
UTrKjQoHgCzXciMUx8n7qWRjg5BdOUUwZfJl8M8xNPklHbACpsaMD2ZY2mnt62ji
knsn4hBFovtKLgNVAIY3cky/DA/IJnbanyMpMuV0rkSQF6GOv6OB0bVnjIryP7dU
F/UEu29MFE0k+rPSkbCgI6hhSr9y0NtVcHEWj1lEupbWZfFRg82YOhwOG5zcjFfA
k/4J+8Cp15Cv0sLDuUULXg9NXkv9vzGGnIP3DhERoXPcnFOrcyvwOrZqgSIo60g7
caeHWHBcxEQAuD9l6TgyYtgJYQQPEiE4rhOhhdcwo1L1PCukvHor3RcIuUAE6X3o
SSBbjAmKoNN2nirJGdHlu3dj3Qhb9jUcYbeF/AlQhjI6UQJgCOgeGDJeHC1WkNzr
7iHflq9DEYF2OQhy/qFzPKUIAjUiIYiKT9pJEyAA00/ccNQREtXrRvip+rB6a6DD
8q0InzdQPLLRdaz/82tZfQRXvFeIEkc/jr9hyCrKWzV65qeAgjLGT2wycL1eltci
ZWM5p/yj6pBPETe+pzqZiM9YJkMITuYixJP4wo9it0SJjAhLlfJrwIgHIvLeu0G7
CXZbAT+W1/GFnM3uOkTQgg4ex/4WMUqIQBX8CDrbh19vUNsT2FjVTI65gGx0tUw8
D6XAaPwqk3Y/TSXRZ+T/dgq9K9KZyhrEV0X2whrQVoyJLstcAl34+UMzOqa7+9wb
+HWOU/vaUAsKPg1zHHu3rTJGYj9U9Bl5+WYAvCaJh71DUMZIbooHxok1IF2wc+jp
aiDY9ZHeBxs6/zyIAEG8aRbWq0mq1ltIcbJijnyR0YmEOeq3GOT7FJ+yAmYdmBDR
SUkpHTg0ZBbJhugPyF93P+/6dhjirPcMdvYTmEms+Cmr+69T26lBVL6ShHzz7H/k
62iAkTaLp3yUUkt90X4aPrERG+geJcr5p358ZCNcy5jYX6gsLa4q9H+IwPfkpQ9i
bF6N7g3uVJ092CltiO2xyKNG0S2CCvJTpJAnA3h7Tlw1+6pgiNdXYRVj+iZ/uooV
ttN3kAnPHzcvQA/+dLH4kot01ub7vh05ZSxUE5dbh4p+8MynCGv6VMC1Seml2New
QMBKts1VgRvYBs8SV1X5ZzTsp5oZs1SK7tKa0r8nt5d1zHR2dpkxejHnxWxStVly
tl8BA/GXwMhpYytRwdn4mhK+Um1RY55pMKaxGkSfJ1mx5tT6KrwqBLP7t4y/7epc
XAhMWereZy38jFOE4c30CHKBpOs9mhUns3A6PRO6cMI4ZB/Ib3Blme5KeJbMgis6
QCHMNKrxhusK5Ac7muNA47KcSIOy5GNyTbUtJIPYknJwSAbtnJMxskFxYF7XZSxo
ADxq9s/KY7qZCU5qnpWDi33y5alxD/9SgI9IDiVOTFooFEa8OYlSbNvMl0++F9TK
OxQz7JglBRegA8ODGbNMdSp5nF2XUL01yojQKfLcyXPZM2aU0d6dg/0tYONv257X
8BQ/cyXuAufXCosOWVcZ+B5GjBIXFUSRJI/2hlZrW5hY0GqQm+l7PTKKYydv68Iy
YsB7EiiTcrm48YknRgms+zMXZfsQP2YUlB398Q2S3PvkdQ/nDEDPoG4ETlzkQb3m
MB71srT2oXgcSfdHYsW7TUvN+32nbz9rijK7NKYaIsQrMJ2aF36jPkckOPGQV6i8
CqGtJsoHOBlmjGh1iPpLHrUbwSZXQ5oXdHC/CCeT1IOupvWGtwjbdeCoryH/Y9QY
QzF1i8JLJAMHYjvz6T4JXywjP7HsTC6XHgtF5apcePUp32+f1FRKxdCPvGyP+hWb
I0XKMQSUXeu6iYRTnzwIBQuLwF/xa/yqsN134CD1MV0RgMPQ2h2Vy/g5hpEPWNhQ
jRcq/XGvFeKu5ECzrQ0EQ7t2b2wOYScULcKs21J5gEZXr6hY8yL9WMUFCBSzX+qt
SZBppthZrM0wJcZBMaF6s5z0IJFfXnjuKahjKlAMsX8V7PGu55Zv/ds5kELbKZym
CogmRPasM2OFpfYBc8OkyyXF7Lbta6nd1TjCnUYvbMSzv83yccZxBQ3UIYnUaVox
54ZratSaSzJTk4ubrDGDkXbNJR+G+Lwkb+XyNVipVz0TV4+eJ/gjekxhPAkOx67d
B5WWWET3l03BpS/wcqanqxkz8PkOjAF6GB9puNznEI0hn8RnBBuTwUfzK1MN3Ggz
5yxrAKBApenEeWl32WYcqpOd4AwvLS83pZOqLvK/4MgbAUMFYyDgwJO63av5joVT
ngu0se5hfS8O/1hVSdsCiCOidmyx79FPmi3rSMGFzoj1xXTvQiqIVP/w/GcSp+mC
okOsbAtGgR+132i7DDEy8SVomGmjiHDghLRxQZavxShmWuJ3SWGO03maoRVBEzYp
t3balHr06MwJkAirqaCnzZGjwvl3KvUZ3UomCcmajBjkXL4BPTzzdYEikDC9PB7n
6UZ2DIVQnxzggs/F0mXM5GDYjye5/ZV4ztwL2AHbYEfnm1ZcKi14OC0qOyF24aRM
fPquE9rNeRTjXca/C5Bndx/Lk85r+wumWAtUil5AICm08h6cWzYG1DT7VMY8Pkzt
3wAFeYM2y9oLCX7V7QHvRMR8oYONAGZ5kuLXkVdTVpNrSvZoPpxyfFvBTPARWtma
ax4THtqr1s0LHM6755TcocQsxrzdwI0VlDVVeCSjy5+26GGbHaKIjZvI7NIecA2+
SVrYGdHzDU3aUY9WIxddMlBuJpUDzkFzB4zUV01e+BGaRq/BbyzU/eTxifyPU03o
5jzYJc7IITJy7KWvPOt5QlKOwYRPjFrBJQv38BD5xKt8TZRPvxLr7izsWlRiQDBV
x14yeJZOdMbQzVGkqR5Aq5ByCD2T47iIuHNC/oi/Vbw3/PgD1sv5WUSXQg7bBvhU
JeJM8X2LNdmzqqfl2/Y3ttjMG2aswX9sZpzJnRgXnQSnEa6yhbaJ6MtGS29VSNRo
fbwYZUymQmCyF39hnNo/erSYouPMOZ6Jem/TGS/s4SucFJP2ygYcJvvT0hw3ZH2d
T60Ke0xkCxTgQ6iQUvAvXCsmZ/CoO8SohlwF9F673KAiEvZDf1bl/jxp2tVm+Gbj
NvooIUS0vUWToGNEWkmnJz+Kcd1x4d6+E9sZH+zkERlOFAXETWrBZ8KfRqE1/dnA
Zma5dpuPijsbmEDV+/hpO0PX8LbM0KMk1h/V+HhFNz/vI0g9FR1ws6SoefeKrU8i
8lyCGfBVK5BoMu5ev154q5Jr0YKlAXtCY3HR8xTCWlFK0jOlB40E+G387Z5vLtCP
mRitY0NRAEgdmF9RO3g0vsigyiixC1l2TKaK3KfPVGjPuGDXwFgBpc2kkYIu7tmE
rdNvKYgfEqrAqEANNurUDbwN+w7SiBA5Kr4D6Ad+tqAlKRNyYVw+TA/4tQeHIXAi
HphJyTbwQqmysx0T7hFnGAHH2L60JWXAmIgWluGodPw0ctFPPgK+8V2K355Rr2Th
/2tZ8fARh0vA6kYBF+EAfVLNzR81AySjamjd17mHFAbTAZFfkOc2bc4jSXwhhR4M
8lUkawyFZTqNLQAtc9oIepmYdYjkDNUOCoAMlKvJfzin2ctxFhRUVX6fwvCSg+JV
s19I2NYSLhL4YbLSMcEdINX2A57qjisbatL2jLQNNrDl/jZpT7poHdkKSVx9SjNT
Yq21VrRmobLpZYdIDkJIiNh6vTtzlmD7qW0o1WO6TjE2tlB7fXo7i7+sEYymw6b6
i1+NlhZUm9lG0XT126MkPmAJjgAlb2YYR/kgohpzRMxyjdM5KvPGW/hEwf+Xv5TK
N1BQslfyp5fE29gMApM0jFuPNvHMcFD+55L4Qk1EADPKewEOE0dKxzm0Fv33SnxM
kQikxSGeTrnPIuC72XGacUCEAXXuVQRcWGg8FpOvQlVfeAVUDz/YZ+mMs3+yII//
LFFe+8gktsxa6VtLhGF2hKBhWonrswN5n8ArndLOzAhbbCmPuBfw62kcu/C3mUxT
LgWzjGXsCfEX38zZVe3N9Q27GhcwVpPY542K0hJ0YGg9MtRbTdFJC/BVRhf2k0eq
/DeqWNETWMoa1fl9nUNKNPjgD7SvwEuGD8h0cLRlz2FY3gYfeHu5nNzJkoOja3nB
mh8hHhLaFu05tuyIUvAncNt4jyzkZnOq7+YzB67WiStLgxLrPQUGgIiil43c127C
bvc8p9cOQDoCjzQLGRWIUG+3/2msSO0cPHmMKBxgi1egUHYZmDZ6EhGNDonPRqbw
xLSlv3ESDfNQcFwaS3nQ/Yk3Y0HiXpYKc01wWJkt0wguUMA/y84ULLYm1eMPCYCa
FdktTmmrfNU2jLxy4q9JvqE9qY0kmeHC792SUYFiI8vjCOjKpSHwwIOqDTtxaymj
c4eqIJpKeQ4/0lpbqI1FuJzYQRtnsu73WGcw+oMwqtdjWdNwpWmx65GDPATHears
mz1VXPH197lqIFKYrgd3WzEhlvOl8FshW9eDma3jDYn1PiH091LouBxCIk845toc
X3N6dGemWYJ7jiERh06b4bXlkmKzmPcdBT2VLB/xyVGN9haSNjEB0yHYhfxqXxro
8kogM8ByvEHzgr7G3Rs1ZnqeaeFUil4BIyCUFX9OUZTdKkW4H8Ua0OM7W6ENP4pm
up6fg021DFV1gVXrTYamvBOphZMjBd//zVjGWJP2VmO+f8+Ajms8PJheHmNs+Lfv
6hiJW7eat7zr7Np6Ar3zld+1PabkA6lx/cvzHzOUkw3KhA5N6CLgUbYtpx0J5ARd
cXatS/OhPDrI8zesqy7Jg6ms+MhdcODKcWPM29MaQuGMMKzn+nQNvb1Iion6OOoq
FaOcRHiNQAh9MkXT0OE/SjOybMZn1GkTaTLydu2mcK1o0KbM51VkYn43BcDuxDt5
seqryvRb5vI1i9q55CkjxIjfDO1J3Xa38B2Fj5HK6eJgE770/aGZUaNnUeM1tna3
lJzyBzd5gpI5fj5V1RTIXBiAyCo3HQLTlS3hYbmtG1vug1TV+iaY4XvEqRPl2jos
VWnYAMwfNEfQ9WhWR64F0GgrVcAxnfv/Z7nklZjG/n5EbPxv5SHFMLhfUONCHT6g
EL/+APo05saFuGoJ6D7zr8WUDAZd0FFjq8CExaAh2Q3w+ocms1z2nOsPk5EEyLiC
oQ+9peUrUMy9mW03wpSFlZpn0kDN4Yhz+nNsoo0zjhIVqdcCw0HR9JRytRzMdsEo
Wm8GW2GDbdQdYgatPtlIptIctCY+Pdp5/KKAzvfq1LqwuUXYyulwfyC0jDmjLJDU
xNjnd9vcY2FNrBO/+SJPgxNbp6wiuWH5p6bMH+6eCuYkAAT+XXtV783kJvmWMY7h
lZFJa1L8IDUQpHZgpnVTxLme8r85V0vIFfPe3krcb8Neq1mzr2ViZBHeL9ABWymk
LpN1equBOPZjRBjkPQRrjlwoOz4ZrDbJvm7LTkwmLrJ+HaYEZhRvISaEZ6JQy3xz
6UO4d96FKL2KOFOCtwOWD05DAWT1sizqPteD1c/K/7mYKQNINC8l9amL2pAOppjP
K6/5SQF0DU36+GRB5bt45A5+j0P5q+UYF/MXDTuldFioj2chl6bj2+zQZKNyk7Am
KHOCWA/fcYHBMD/zMJ9jdDIOddYz3ZIgub2VW2RogJpDgWsS3dkjGbzYk9TUk291
prFTshEJvnxUy+LydRBQeX9J20W+uVu/rTATkbA6Gx2csG2mwqN8cR8tJ6uKV74U
Ri5JKk1Ahf4MUQqQRfwVqaskuh3pm/QubtKS1ZTtkxRsKzw5hrfjYgsjGNIm0jhU
gWIfgay4L9S2BBbI5DvlxyJReFyjRkwbVokCSJpjNiulL+z0LcCOd8C120MfSQqZ
8UpafYxE+cAa5KU5zm4kK3TdZLr2ozxQqSn0bRqXTuQ1JWood3DXv+j3LHGeth+q
nEcns+Kej/QIia9JgOWlmjHK/f8HEBniUqgjcD8s/Z85P6kPfbctR91EeIW1Pkwu
DNJOwqpu5otNmQ3vPQfeG7wmA/LvM6WJU7zJd4bFoL5NHJYX6EUIQ1ixBrPMvNvB
qBjurCCrSadgz3eOV6fjylZSfhg78aCUkZqbTWs/3enAE6W1hVWLgQgcgFkt7wu9
MOt49+MMWzh3jAA609Do/xnmdh/UBXk/oV4nKrAMdZ38bXn6piPzdEwej0e/T4QE
2jCFCJes/fLk/z8+SPfxzXzM6WWON0+s6WKXFVD6kfF/72fhS7b9N04Vm4w7Kwfo
pRxc+QKnDKNmSfuYofLAZDmAPl8mPnUG6Fg5VuK2Plx7ZHUAnKrb9FMe0eRXL9FL
YoKw//Rag24cA2ByoAsuwzZcFVTnvjh3yjnLStEYmZ8+3G5dpKTb/u7ZxNnxlaB8
aDfhQOE7ectDabjGkjiVyggWmw5t9k5eOX0S3W8EKKCx4KJQeuILOFE7J3qhQ1pu
95oN37FmBqJfpqrm5AVUdxsVrYlJymad7yXjq/8Q7/crmOn+9YuSJ2AoCLBmZYD9
tyUyj6on4JUwQ5o7nZwK5XJBlEysSXgJiT+dlbtTMkYG2rguI0yS/yuLSH3iQWS4
/bZmIA2Md7MclDJaCMrs9Tm94RvGpO1rmQ+wcgNRlCchiwL29iI1b+Q0hwhFjRoc
VrvKEZwwSfWWoZE1kSMeMfu8d+S9VikHmla3rUtuXiKM4o1pjw1bHNYxQUrNcqW5
DQ+Goey77R0wVYH9RlMssxSwI9GpoUlibZ+exlDOl0DMQodqJDZDF0B0mX7Lk9s7
kapg57vaBwAdw9i43+lgou9V97tR2m3NPDmOIIexYJbv6c5P2mjux4Qj9AIack1J
gu8wytOmu/QZmdNkgRRaGbkfFLfo4FGJ1hCk8OilhIqDRXZFPd6/XwQ8m8UOqp2Y
874Ht1H7W+SVVI81Hd1R9nGrmI4XWauQyNDG5Ul9xviehnvaP0/Br8Q0Vu+9yKOh
BJ2kyg1unrtoy1r6bsn/9gTegtQjSLSjhlvimixxbGbEgHKTVTafRJq7WAYSCt3V
8oYl1ljaEmA+G2fB19F2cGuRqc4jXrGy2lUFaZsxM1AlHHwJXG7if2G60WvYk9F3
Zqsj3b2zaZd7oa1Z6oxwEqeStJEywytvznzA2/KKABHh8GE6CG+oegD2boNP0W6b
hxKyglKSryfAs2foY3AYpOBYYvvD1p8G+kdFJppmakaZVWGOglxxHqpEfDCCYTX1
KsmNyYERKMtp4Ox6FBxINixWa+zCA0xmwKi5UYqTa+OTkD+/84bASxLkFqAofDiI
V5BQNpQYOSSOizk07i9mlreoXBatkf1kIsrEGjLAwoS+36MfuDOxSnsAgCpO1jL7
Cp28DIqsPVLP2lypOwPCLdK6YJylT25hUebnKskHxFgYKmf8OUF2ijSnF1tJ3XkQ
nAXeCam/fvNW9IKzQ05SMhnmuJU1sBvAhdDCDaej1nz1Z4PR+cuFNwi9LqretQ45
tKSCB2B3dQbWu/6ICcWUT7K8ttLem0nd5t/OiP0pKXsZnA0KmV3PvBZ/cok3j9WE
L/qso2HmoLI0gu3CIkkibi8Qdyb8n9A6VzpXo0KwzsQiIg9ZjY3d5a2H8qNax3jI
xR4Zvlus/kbwsnrjrbVj49bbesDWzPQ0co+euA0/jJMm8HoUfAOmQc8PmcviYF3r
DVoIgJ3Gj+3T/3zuhea1RNhCH0Q3zhzw1Eh9Abw8c/ehevUWNcqcHWBn9AD1sFSP
fGl0A9EmxY+8TL110a9gBPvx82thmAUTgY6LVqfC8Al5WEa/jmYmmRnC9uxgQ96r
uYJbFRyaN1ayVKieVPIGwUqqBHKrn8UenqGWPUCZ/xvLlhsdDebWliFocyig4nZm
LCxWNtOSgonbi5bi4ONRq4zQ8qmY1QyCA1EHzu34Xzwpx+IrdSrD0sY9yI0WPP15
69IjR5DgsqnYtHaZrghQKGkkIcSr0XIOZA/FflsRIqkMFEMXnhMpbv9dIg0NddXj
oEOk71N6PiKxfdLPwTxepP0YGScnqBgGVAtNF+sViaTn8FMn8ctLozVctzpfvthN
r7wauL9AMmWP7jahZe97GeM7Fiexp/wR1Q3imOTdL479w6rgXTRaqaKESFNweA0H
3eAOpahhikaiFk/kFMhQ2sRQ/svyZ3cQva7xJKWQmbSjad3xR8WVjpCZsuh/eWje
Pe2+OIPmDKogY/FBfEZM1b0inHM3+sjPU2hEIsvnH/nyNDkr2k9O5mxEKMJISY6y
8Eq+VAIoE5RQ7BjzCmQXgtSd2xEWPnwLFrxq9v7zo2RV3ZJJqm4L0JllDODkGnsA
ooCM1lGcgL5D/XDLa/g1ebczEnErEAgT7XPAxYX43etu8TjnZ+xy6NxIwAZCKQYi
n5VfS++xRmv/umA1jOTGhX5fL5rnZey6WIWvds/eYwkXfXWNxCrq4dU5rXqPN1Hd
hdF6YH7jgFV1yPQp4zQ938EFhBZJCrU3DM6/6/+izl5JqDU/90aQNhHvbI4hhjCi
wh7fktunPd9QRtdPbmdx7SyHXx7XEXRktg+p8qjWWoIz8IcUTBqjkZ+DCdmOlsae
fY41hHcpmvYeeu5eSrcI7VYEKklcT5jJzLuqiyfoHEsYRcpNs6PTzNV2ietoZ8UO
Lb/GCyczdsR0fN5+72fRPasTL8YxxnjuOBxFItIUB3v8oo1wr41Z02vVfXpgMbvN
wjhynQ/glYqdN9Q9jjPISMgXm5uPnDmBdXhMsoTqhjd4Un0zSGf0jvM6Q+ez9LSC
Omb5ygqaXD/uLBfBY+nGnYH4x1G4Lw6onQh3mYooCVUQ5Qeb+XBMr0B4SCUgdGNT
I1dWCS0Ip/3U1TV6+enuxYkg+QkZNjRSCdBa8HJ+Q0dH17GSqJt0GakdSmnWJEc6
panNyH1+/suV0xjtoA1iFP4bV9vUfnzHlneeF9ECoSGaTm5z/1iBYBbuq5R36MyV
7gC9mQx4RrnBQy4PN9YnlUMypARab6bKYCt9GlAvJ1XqhV6Q0fnJtWFuD4uUd6P4
f+wtAxBd2TlDV1O+098Mg5/C4CoMeUHl26brIlPzYzNtc6/AId5P10gMgXrdGMbo
tna9iOAINCt8/sKzPJhekEdLnSpcixnBvvYnnZjpdXP4XePnLqQDTbfGEsKsMkib
o0XVPUzpYS3nGaeOAQC+g5Z6J6b95PFjXH1nXXJdyoPN64MffDN1oCKu/k1/wJyb
YOAgSuutPh4Xj7DAXW2LSGy3lvDcvgkgXW4Y+a2JrQnoVOrRILMzWdtOG3vchkqH
Nt91eA1T78QoMwNCPr7SB4iJLowWohNMpKNyMIEXW+4zFTytH90Sd0Qnx9xf/tS6
7q3KsszBGyRixWljXtgExLaHTq236s6kUZ/Q0msQ/p7wSjEybdhpw11ANjCHbPdV
khkdhdIJdYg2vFokj3itZhr9IE7XDhDW6DbBHinCuDTBM5VJLGDGFfazfKiyWMQR
EGet93vTvreduJc8bvsge0MFe+ICqygLk26QlgRebgIfskt1tfCVZlMkEBHtdEKA
jjoJHyBnlTbkCj4uT5A60BGQMB7oIIJiOU3RCg3Ay+OWryf2aAKij8BwuDElxfCk
6ZArFrYI+0QmRcTSe8r49PYcvO9sECUN0PBpxrCyzF4ExdJ9+sCDiWuLhy4DOb/F
pPhb70t1B9YCHdovj7mH3NEZ12IGb5siyXkGGVxrwRbAmlim0VAPJlga8VaEnPe2
SDAD195kNFSStAsaUmL5xRuUDLFJ385AdGIgtzg0cuvzX2eMG6e1xAwT1mmIiy9k
DBl5Rcg5ZYl22f/n3gd1DHEEl25rp8uX5oAf6GJVnz6im0e1x1YGBibOD8+0Icok
gu7zWmwXSdha8x1MFxw3FiCmh9vPWmGKGspxNp3E9MxU1mo8mH2lTBf+0J6UHMUz
E5XPMwwPnTPq7F/fT0ZMEsU2CG1kfHYRIfqRp16LogV9ujO26FzIKFCX3LqTRYPn
z24VyYJeeUptDOuTW35l3mN/fYs3iumM3SL6zFMgqBYds/H+9jiPSwWJHIOuxKZJ
/phfnTVsJuaoVR89cpD7uoubBUDckKhyeu/24f+77OwysYV/kCI6iZkwtTjKHki6
/dbtv/t5ldp48zJxJ+tiCqxI9xj06QYJ84a6n18PSnWFSa/4Ig7i2VFFfOTDEXY5
eyc3abWx5E+YFzySmqMkgAuhDDqJy3G4JsSAiAhXCZwAwpc/7IMy9REhrzT8KVrm
6TT/n6/9YSumplPbUqbCV2zSuLRLaodLtcWctks0FMqGZ4FTTEp91g6I4hJ0qfgF
M5hgG76elmXtkI/E37X74W0R4Ku86IS2gFjcCuDKvTzrHzR+mEYe+NvrJmiczuX1
qW9GkK16sueg17MHY7H1fj9c2CODtJRJNdPJLm1HAst7OXd0RooadQcq6y0S8Wyo
v/DTH0f8eDshb8pUelL9bIc1vFqvhgcXW2whc3TktUE5/hrTQPAv67K+Gy0VALmw
JfYDRMQ8odmRQSgt8aA9/8PwcI4YI9Gq/OFjqCWYG4nPtSuPWaSnP6ijTwcNz4xm
BhKACPnTodbu+9QDPXuNCABn/T5aQtPm1eiXG9+BsIZMTGBegEDYKPcaIHlxuweE
7P/7dHnitpVFAymuHypCuyNUQfGwCzTcHYox/H0COEV6ook18MXRSkG9H0MWOHkb
zGl3fm3DRf3nRPhp82mrDaegfT3Ym+MbfdRdAh8JBZbGfnFBuQLUV3zRUm2rWyov
eCUcpe5Y5ZZ14pFzubiz0ePSEDLkTPGNu2CqhVvPb0RGtM1TYGI+c+GFko48XZ8i
H7rJFuWhS20BX2m7GjzaIs9FTqp9lb64GtSTm0lU1+SRP98Sc5+L3yjI94OQ76Jw
COlBAdztpTCAwe/gqpwtsdwsJJj3x0+m31ugA6JXZisJ4GgOzU/Z8InZKz7oLG+v
NAIWOcDNBBxBqShsK37wF4HKnokriwzW0+pFFyWvPvxnRsBNUuxOPl9l7XI2cIZQ
lQGH95359IHtBObdK/AFJsh+mdh20IeOtVzWrh7onv07UcU/6rtarsJpGg6a9ayP
K5/L3LACFfgBZSn9wkyHugRMzvRVZxQqS6EOt9EF1D0E7SFOY6FVPL0Duip6w0GN
QjMidbkQp/pakhPjp1n1j1tg9njIU78xBZLcogqMDGgObrNlseZ0EUBFPt0Rbm6Y
ZsoWcgNIoO5hgLR8GRJo8LZ4kOm9ltCVYjOPPlNGLZDSR+MfStRgtwJkTXqwkqfL
4vVxRILt2qt73d/Wk0ieJfgMIWWGRwTQdp7RSKyxkYovBDneOKrtZ+l9AYuKI2sP
atPh+VOOkEEji8J2Hiw9jhRGTMXQWZM8OLgpN22rG5XlGF7hEMyIokcPAS1uLDNg
3ZZHWcQOlul1wAtCLyHZVBCZxL5B9C+7W8kDHmlQtMEpSwxqBQJLPOwre1tNofTD
nFaMSADt13g2OR4R2Tn/6O/XnNdRSMQsDtXrvbo/nAtaWpkLptT1rws2oy86T31h
DwfuKZEfSlUUyzJV9ubbe+18HQ+KKuCPBFxbZiim5WvbGauc/mn6UzgVEtN7Jn0A
GVbx5sMfehcL7BlAPWgzT+UKNsOPF2QeYLDHXr5XV9s7YzTlh02Gx/j3ZC2BLzyh
EjjBPeXkf1GG41WVb9uvbX3ZxO6jB5JVXogdsVMJuFa7nvrXYgqTeGls5/7FLueG
B3IpquLaVJnFK3IgdiSGNFa9d22jgCEf5AIPtlw6eVOqCv+iLOqWs36hb82nrNwT
PdJ84JIL6cMSVx3fDdu4YO+HtB7y9V2Y9kJYLIn/mmZf+LAdiG99MN+UDEpCoyyH
vdW50M0YtGOS43yxdbwdnXCyiUZb2eXndvMbd7TIdhfcsi/7BeTn7JQ6QSkug3HN
eXxMN6TFGOVoyMAclm6ssfX0ae1Vt1wFkvS0Jv7rI7u7fGolgdqBrFWlHDFIlZ8d
zlcfMzv+vOHBaoAOTEaDnfSvu3tGfnrKLVSvJNxYbJMyM2HepL/4B+bJ7q3Ti+wg
zJfuwSWSEd1HN2VGrsu1ViUJTWJhrOk+45wB9NI6zBdNqejtFTzdJk9OAV4+pJhD
AtkS5DWzzWyeZg3DD442j5k79GNvpjncRlD9gAmFLX2EAl70805EsB/PUhLsWU0F
aBskySPXakp0h80hyDPskwohiBvCiqYUR5XA8BBeqfIfyAHG/CeqOnFUTbxU7qkG
d7fFnQ2YoFUbNTtZ4DnrR1H2sSYKlJ4vCaRjxrPvhTCdsU5smpIpYh4DDe/8EQhx
TxxtdZ+jik496Ds3kvHBzSU5kqqbcxKqPWkmUELkhc7sUDMj5S/9UcutnCjat6hY
XiQz9rBRds7I307dFN1J5IwhG3Z1vs193yEg8h0M6BSU4QX0EzUq84gqsAkEh1q3
NK1mri1KUlk4qq7Sv/lQkHkhc31uPCZJIPYW6OXfm+CJQa8VKShsDJzzzufhZcEz
fNhNup2lx23Y87Mem1092c1+FD6EMIc2ezq86YOJeZwo+cLGGsIzbmi+JNuUT5Eo
uPCZAXFIFEFQZOHy2LLvx1e7ZffYUoJu0w7Gbz2PRmH1uExG1xX2KmDrrt9eRuf8
WLW6Hj6hNe1TrdaHJ6THkpiEafUmdlz1sMfhWG99oWAke5eLqArXDgr5stBh3VC8
lcNy8/K4MHfKo5W9vfcNi3YSmmTfCrjsFmTC5NbI5D1GH5lrphZuXZBxXpWIEfgp
hV4hy6ofSDD6zc7neU4wk/QII81T25/FgEfKx6HWH7ehBsBqldlZEn0YnNrnLnB6
nw8BOp3Fm2ZKRyPJojRXIACgnlL+8G5LdyMQYIIsYmlovKW6KHlxCZyH2LPIMrxB
/Dpvn2CIbyv7OgdaJa/zQiaJ7G8IAXHRuBCmhSxfCoTfDFJuZPYU+gbJaiAHUTLL
UKqf4xxHIzXfZjxz5iq6meZUYC4YnEWH0BfC9I0RMHRxZs0wesIy4IkqVAJLhtIY
pHsZxAYqBENJhRfmgo7IwpfnpWquxKRL3tjJoh6mPnutuedjeZ7pBbrRvAnpEYxl
rvIbXIxeqxiLoFUVlFQBSFgSQBlxUiqWI+C1MxQo/UsUGwEfibTQDR0/JJeVXy71
OSrk3ZBfFOAX7gcr9lk7e3p7R7yzaUVy67VggysldR3qPObVnm07L11csM+w7mum
xgKm28ht2AeGOmC1eaFORGQlTR7Bx+oCUvKSyOT8csc+R69QSHDY9JMANbzFumTi
TxjCsDd5ljUDGHN2byDRBEKsuVbuY/DjcovIz6NcZvoa4iFaHnGzNEF1UWvVhjhx
1FCfxfY40pVIJq4KwxDHPSWTtU0r8G/9HB0FOun6H1itRY4rrpRJwdbYIen0Ga2U
ZUhrBP1ZxTKIgb7/35Qw4HXeOUIOm59xGa3Mf/3JcWWEIr5UqPkjWyvxfYr3HqKf
MjaaAkH7stKULrPw4A8vJIQYhMlc3rBZ+JBnlOYueV4z4Qe9Y1Y4uwSifdfzgkDa
q4xgFLx9DJ1TqzimJc8BH2CMLdjSZ6p58r26m2kCFj5lmkGA9qgonxyEWRT6/Q3A
pm/xXB9gkzLu5ms7HekIUpnms3/zxS8pqOY+Fz8uw0mv+L+hCp17To6fQWYrYNqS
ryHFKTL18SzQZFX8rW+Yhce28RpaNojstGXqfSn1zyLou9SKfge9RhOwQh/RtEdn
K+kT/l0U+au6imZpKTVpq5xim+WPbW+Zgqo91utM+KhjlDNh7PJB+ucjV7EcKDzf
DlH8RW5tnLrqPYmpoYNFFwKpxorifKCPhFCPK0iBeJ2Zt/W2IhcxW7BixDZTwfYO
bDoq289b1PWjxyRpJgJkMufz4wGJhNGbaoJiBcm1XPZUolONmssPxpOopHaM1mGv
1WSJoGYAgAgWDfRryGTk8QiTZFJMQpsBU2Cdvvc1kjg85f3h648NypL5+ABKgss2
htIBWNn0GFUnoe03wgwZE4An0D0/CXUUr6YJosWNXpN1ttWdmhSwxQvOmI6c/AOV
5N8wkM0AKaMFb7Uc5vQWuP8Sg2447/RbgiUExPTqYzujgDGwkKD/6DYlXR9K3flx
IwKk6BfKpiHigLypz8C917R8aY/oXAPJ8t6FjNL330w9jcxTCRaklTHoAqI3Bco3
a/U8znMlgkQS3FfJ0vMSnwCJDFEi1g9SzBqCXXf3dt5gWvzs/D1ET9rDh2WGBMgp
TpuKW9qO3z+mGzJL3ixvopK4b48/8YHjgxEhbzH9jjFp1x2vPNQw1M4qB09ny6/+
BmolHiEVQuEFfNYRMHLYYzH0nfbREhe5E6BVNdvlVq64knvoqSLE5PCCyM0trawu
LY2UOHt66f55F2fe+Be6gq7hu01t1jop1eigQKjJHozko+6wK2D/c+P48Na2aEdJ
p98tOMyEoi/81UrXAT24d99dp0NAkSLnbFynOF+9LcEB4OtWL1o4k1x9xUjaavTS
Im/GK2AD+a8Ua4fTd8ZTMHlHDaRyWMJaWz/rYULoaoK6P4RCmn3bSDxomGdAil5Z
n6NJ0hhB6ShrDOnnFAh4/qN49m9yPKwQouM9DrK3tbLajPl6t5UZD09DCrl/cRxK
FVLxPaeT3i7HYL0kq+PyMwGZdmuKU/uETE8+NpsGziKSylRzFxfKFVfQk00x6QIL
cLOgFslocY5yoghsmo9f9h/vOvYMD7vrm1BPG0d8Hztxf6kjs5XwZj6Dpgq70vOd
fCaY2BeFXNmLbOOUnVCXOoUjFHpbGa08y4hIUYi3t4LPnRpPC1YaQG1BtyCB0u5l
ajDQaXKy9U+q0DuNQgheOG71Q4e/GIkb3JZS63TH1RarPx4jYnZoW1Zztqu37fnU
bGd+zKiA04idTJLC0N+L6ZGepr+cxyw3uwa9roqB3CSmXyA+gtxECm8TXBTz3goR
aHahdcHcULapkdbTjaZY/kSdwKGnq6hIvfyEHIe2rsG1wO7Gpb6/QjsHcv0m0z3f
4QK4gA19BDMROrOcYB+FB3UXCqxRucyQ8L8Pp+/dBjPStFKA69tlRyt47wac8pjj
bXGc/BqEgus34rbo4tlTjXKQic7AaybWbKYwpbpk/xep2lpOomS/SSy3xWV8BeE7
a9PLcMzCi/esYpLtAi1E8cZ7zqpw2r7O6eu6J1CfGzFu22ClncvEza0NWt6pdEov
ra8eq0IjXM5yAiSF2Dyk1Nio1A8ExBkpd82yLhgLmt4hoyR9jvxcNcHE/EEbrclq
FEzFg3UbRjshwdz8zksYDF32qxcG8uBsolsXUvzsqMfn/J5ExNhAnzlihx6/gggN
zOKMAoDr7XjB4lx5VdiEuU9Mon8TarQsp4WpIbufJfiTzCPCFNA4H7bN3L41psf4
Z7PebLD7SUdVhvKf7h833GlgulH5n/zgG1eRR7xGNmDgQSeYGa2q7NIQFkpvln4g
+HwTWvg+/7HQhBc7tw3IuTtx2zY8Omd2WIZPPqhfyIfwGagPT6OiHzY1xK0oJgqn
zOPuFe9QJMRhuMXiAzFZad46eOJ8gAtqlcFPi4VXl32lN25+JkSrOA7R4vXUGV+e
ahRZsLo/1lhOaI5k7av7HYc6UTke+WciiQ8swAG6lvQdz1CiHBhX0ADwmzfoJWdY
BB4XpJnMceq4L9hakPABcQLAKEUy3OTOsloi+8ed86UnNNvxUf6mNwD1XsNFxce8
kp9BEUiGIT2lJRw4DmFdRenf/0hMQ/XWneicl29NTGNt0SKjkcNXc6bBOi1CaDQx
8bBuACIsf7tyeP2SUx4fLc1U/Zy602NZUZtAEQEbAfVT5KCI7iyCVcuSIlHTLsmd
EPd5NuZwxZTjVy/KSQmU83tYTflDxISF9FHf3CRVqSbG8i5QC2d4RRCeMp5b2Aq3
C94KL+UNExKKfNcgZg57+ZlpqXDESVHCm4ODJa6VDewUOU7r1AevghVj29SHbHCy
QO+gQ6ogz6B+uWN1qJavCgKRnfEfdzICiHQCvM7aLRBlfbRJXGDmYGOn0F/Cfyi8
KtYLl0ojlHCcJDr+eYZzmjoUGZVaBczAkOrL0PqdRnK87Sygfanh88RXYn7HN66U
xJkfYRjeNrccMI+MRDkx7nKilot2JvglUVPYF3RC9hAY25HchY35PqGys6mKUu8q
3wCdVj8Td32Ves248il4i81igchTQInDowLdzR4g4eIKLXpQOk7I0GeL6aRGMaFu
ZIz6nkmSpzQNHBqN1Djmz1n97Bf8mu/Z+qd9Bog7eJhUSKkj8xCVrorUZuE/yVFS
R0v7tyrChkViLtiMOHMNWV86MWj7sHX5ZQg/zzjfjACrpBIggIBSLBbJnUtK4uSp
sbkkzLqiyYKeraEiSpiS5AGb47LNTcURapJgMjENmSmCFaJXmqmWivvIpZ/q4GUQ
4g7bigttB72k275DjNJ8QQrvY3qylU51s3DK5plgq+jdBlAD8qXg/1PROUiOVPTo
yPevS/GRWcj8g287x8ianqbE0qHv4bzLlz+pXUFBUc7Evj8fWnvYxkoG4To/fx42
4IVHz/uMNVgqCK0r2LCOFR/EYG+7QPIipUGEgH8rPenspjO/8e80UKIixXr7Jkzq
Vp0DwoDl5gR4gad4slT3+uq4Xo5wkfy8uE9zH3E7fGY+1gbsGRWTxdsxR/a+ABmD
IxHbDHddRT5fp3PoTWOfX07ZuJl0WAiZK708+LX5BEPSU2L3N95xnV/FWHve5r6s
uyfybrh/NKn5mU9T/8jG9IPrcKdEFKnKAK9uLsaG1Q2JuwthfZ4AUfnB4cKXo94h
Ih5m9oVdivZAP/neIvQoHH2e2tHAoQIzvGPV2PkcVocMZq2cktjHZrJ1XpTKhf0A
TvXDNFALopkWWXUCAaRxjwgbsbWUI0tZmGLsrXrCAqQO5uxK/SdOL3TFowhMMX2v
289HZsLgedOPOLBo5OJg4eFX0xExShpSDsqh1O/b9bFn7/pmfPRB7XPNDbZgZjel
5XY6XMrur9BENHEYfEVbWmyFMy6ZmZW+SStDsfrpwecKisVjn1JM2v8urTB1HQVD
+WqllWuxXgtAsqZIUP35pLF9u7ovKOup9hU4U75JqgE6LdRXtq2L6H9BLw3LXqgz
4Y6MMe+uq/4hhnt+cosAwT0twbpKzbNHT0Y3j0HAnxy+CpzYCTXQR/PYnEBTzHQd
nC4LA4DFBd0r0oKiuiBELT/JpUj1Pcl24KyoM8tWuBoATZO3h6S7FLsOAg1n4mwh
JZu3r9bKHZH0YooBWmwcrOIogNphZKSNsyfqfmWaVPxGWEbOUUX8JPIQjJ/TqQbX
fGIyoVxOcZfqDXGsHmwseDM98gyTTmH80dWx5UcMyGloRDv7U2VKPZslqL0bECEN
AxhmaZue3grLQ4qeCRTZwQkK+x0hgoW52wYBN6oNKZuKx10vWw7pfjF1U59fe7ZQ
7ZsFJ5mrRf79Y5i/kZQqwdDF3kdd6Gv53Z2P5BiFc9mw2Wamw8JAvvXWvK/Q2Gog
7EFErzubF93rS/fU+TylFvYv3r1eMcbMblo/KlZ6TV0tqz7NOID2mFiHo9Nuv9KO
GaQzLQJBOYFOk23TuiqQf3l8OotnKeaN9HF6hlS+ftl6ocNwTOQWpaH5xmx/8Unb
fLwkxbN/h9cUXAaiTYUpHDAodR0KGO8mgXehPrkFaYJex5wV+CpKgPI9BfvxTYR1
1Z5yxP+eYJMPW0rnjge/A+q2lQ4766/efbbET+LaxGWVsSj7G/j49ATThEvIC6UK
H695vunlDOu/RchaQ2v5IZjLb5cmVL2urlit7mnwgWBP872mBUWFpzvd0ZRRVeNf
y7aRPuWrklnYpZiKIexDmIf8usrMKBWTFSaCaKYdS3pLNGnOUlkigdbi+RogJ6L5
h7P6z8i7F2HDV+X3H7hRPwLLTOA3sJos2RJH2x61wAhUuw5r3Z8kJigmFCztoeT9
bQJvelxxzlHygtw8Nn8u2EtPSExWKdurQ8uUhADFg2Vfb2xfNcH8N6M1DrMxzVaK
T07WgcEGnLSUtsnP73TUNfEzX6Gk7AbCgxw4zOARUC/ddqTYKxa2b078iZZPtYDA
74pSbWr3icqE+t4xkCfazft/SUVCLunVxnjGJ3hKhtEQ7knJ6g8nfW14zObQuB1m
PlldKosatEW+F36vL1p8tj9f4hPfO5fsHNqXzVLGc+RCs24c/Kz910C908usfdCJ
zPykWDUhTCNs8cIgeboLI30YvKCZvk9ZktLeR1HzudIjYml/djN58JuwVTwFgg0Z
AtHz/0dQ+gyiddouy3QuhLLL4aIiHFBPn9RrVaYPO1jI1KKXlXjqqCh4PT5iLBk3
Ifjqh9WyMEW/R5bulLmopHumd9Ma6kzpJTh5FjA6iUhZBsD8yY6EfEvQFFLoFAmV
H0RenOcijdrgukTwPdmUda9r27VpP3SjZfi3e1sJnc7gYoZvGfY7ldCuatVIRbuF
wHZQZj+UzK8ghh01sPCYeFcU3OW14+DZ1NLh1UXZEtC7WNpCswtpz5y+xIBdSR37
3u7q1vcu+/Rfgnci+bv+IrXcR8mhP4/BrytiTSeC3598pYP0Uq96FskjYYR+2Wkq
oaYH4BMnCcgqaO8TdKMriH2CWfJmrBAzRGL9kvFqXU3qMUSaCOIAXY86UH/bVmD8
AW7u1wxB98qJGTWB6hRo77S65tb+Ql+Jmt2UoqNt6Ghgc+veYyaKdQ/r5F9XA9eV
QhBsOHkLFZEkKM7w/O9ZNyqNmqbNw8E8PYCegb0nU4YfNQhvzxS3PpI97oqhFAN3
sgNaq4Ary2x2Dn41Aa1tCsac+BpWGbR5W+CxNYRzvR7ZTcxrnQKzvqZTHC33vw8N
pXOQCd8E5vgE3Ms1LBC3aRBeHme4VBMum6/y0r0bXVg1eHwSJnswNJ9gUH+8Wr0w
OC+GbKmOE2eRIiUi3G888faMJLE/FT7E7Hv/KOIkk/zATEo5VGPqhFreZgHKcDQ9
mWPypapFKufFhL/Ru7xpMB8g7qgqNl9YB98mD2CE/0SZoLWvj19DVPX5DaDVF+I8
RYhfNx5kNNaLGaetJM05+apngmt1VQEMgBf7ckzHG3QKtn/VUoGlUjPFlmo1W8V0
cD16vU80YEH1OoAtxq2L78OvCzy2bU3MtWqzFn8vlGvmIQ0NNHA+GydutclU3ci1
N9PmlWOBWTvXilQFCvxusoJPk3uItUS0thXY5Ijm3J3VXfGmbi8goj6ID3ejfXUh
UFCdMw7ZQqu9jzAIBACjNi/P/qJkNXm9epVIF9ZonPnDy4Azi/WYCZfwSGF3/5oo
NvkLMe+Xt0RGAFZ2lvripPENYouvdwba56jXyV3fNsQBIphyODnNASDLrmPB+kiJ
msfT+1+Zzm1pRMC5BzG+a530q3VnF3VrdI0tsiKZwoBpg78INlJhXGeQjDjzWNR4
ScwO76fP6BQA9yQ5R5oOasCaVTTl1G7/fHtrRyapg84rmgBs4cqmy+o3Ze9eqUZi
Ter29CpzJ+i5J4tPxCM4hm40KnkGvRdn0xHBIFh3ty82hSSy47ztx28g0P/kCpuo
g6VruMZRYOWC2khVEw6TyuluIasqaNaXhx5hwQtzxGk3bnJotd+STc+uSp6evief
XLdw75On2Vokmt7hm2MoQ+/upPQeRhCTsayBe7tf/pt/oRpaFoW1/JGeXjhmdgVL
F10tNNQy71EwgCE8Whml43sy03L6JL79dVP3ohkunusvmpMUFaSdQWVCYwb0xhKJ
puRPHHmYUWB+Jhl2DOHOq1+rv79ubvmiDjsPg6MPNjQYHGYIw/7frUd0In4Wh7z1
EFgvfqtrDKgzrPJOJHkTlJGBAYvbeFMjhvwALFbSTM+3j5AsUP3pyrizq0froxSn
3sq/VsFr0Ca9sLNm5ozrrYc/0bCAXxzeHMlA4XmChCnyMY50Sibq6QUp/+yLovrm
sonLcJ2HerCrZG9rpXimd5zRuOKkeCwwp5FgbaqWXYxUFeK9i1d7HP3rwC9Xra2e
cWfwYbIBuXpYyHKq/0Qaw3Qqrotwf6Gw8P70FrB7aCLQ45UeIWGJdb+wDI+geZVW
PvXJVrc9dpsMQL7eqPhvuz68Jk3HcewI1a6puNFsiJDW/XuuPS1k+QE7iVxhRaBt
k2fzytuoLiv4yaaVCWRPH7lwoFzOWo9ARNICmUHb5GhwCLuXrAcdBLBHbQzpZFHM
u5WfkNNvICMci1ICJICUlgkXD4Y5NfKDHP63TIUFq2CLvsHFCnr+dYjrm0kWJnBJ
ZqqP0FYnaxMkJnHe4ySpp50iyEcNfaSuuwTMjbgY6GXkAAPZS9efkGTrEomfGJql
ved5NwL3i6JqR4yGVhT4FfcpvsP9tC9WMl9a6UF66wCV48wjbiTADHvubxczxC9L
GIcwdhg9rspBXyqjBlK6u83Q4H+/jn17TULai6FsULbP0ckgETXH7HpVjsTD5T+I
5nMtZZ5eyt/NVtJLANENB6nm5VYnT8xvaQRlYpZEzMzmkW+q59R3tYuaPAzWT0k1
i4b1m8hpzxozdnKvY/RpNhXNS9wtBmXtsEuk9IY3GRBwkBnzsGrAJbh+h8N8oWz3
JeBgbkK1H//YpuhvuXYFr+qKq/8XgeEQDvJCeZ5nuF6UPRg4TKGRLiiu+ed6YwJF
YlxnxdzdXY4bfyJhrqenBIYDKArGg1FBhHA1UaLMPLvf3u3ifndj6Itj+H/+yPZt
MeSJs33LCkBzZRCxgVb8OS3t0B9prtvsj1558L0rJrSVta5KlppSjk2qbRIJoO6+
JA0dEG6Z41TB+5LiNW1HmvejLHjKMlrv9x4IbwtBXKnLM7Er83o0/KE1AVw4C6gh
b/OPB1c7TTOQz7iHilBQVPKKmI3jexPnnziXlgVZsljxLO1zz240LknAnIt5Pyei
jVkhPMRg+7HhpKLuLsovL4AOx5ffGfNZ07PIwROHU4W4iqVU7zl6JJ/FUiH9iqR7
/pIg5oZ2EVgZ9p6IeVoBEu1QZWVDwUxCCuJ7Mijpr+oQ5RLeV/yWNG5C80oS73Dq
REuzXK2X+bXGAew8C3iC8p/0ekRalZ7bCN2MNw+sp0zOx55i+sPPN+Cq11Y1L7xe
az8SibzgXQZHRoY4BAK2/fAH7ExLtZsqD+GI4jVKSUOVP1QjxmpRjhnqtZwYlbPv
HedMOqhQ2Y1bJ7RaJW2APTbCN6ATf9Na8Ml+oawWj9yO10xHBIV1TY+F3Z1NoSBO
dSdisOuoB6I13blEQFFsHHrGQA5dDDPtJURaGqU4o+zcl+lfv/1bJr5hShIjc4Gv
HfRcXLsUh5JNNFBrDpRhlVpHrwH3fzRhKyde0GVpvvQZ4ynY8999Ky/mcK9x0cwy
nGheVJL+36JFBmDKs+uvrRd1YajfWCe6s1jItrcRPaqXdyv8AtWaeS/lyd6kw6dy
VDQjKzTGjqZq8bFsVf44eJf7z5LFgdSa0BOgm3nRH8Yxx+yHI1w1ExI07lgCh3rp
Hr/wEqOMTYsKzcv9HRIg+lBni57SmIN3wq6AD+8kTQqd3AKIcqjqRPzxpStiS/yi
y1ghY3OJDZGxNqP6UdFBCbpXrTXZYxb6vVt5K9+6cFFnzmOEuTQERzL3Tz85Z8ee
XJvrk55oORzWPm+zJa1cg2j5qN75+zDYuYAfi44iarc3CMAxkuGwNjwOhBzC+Atl
Ein+bZZIRdUdhQoVDkFTJz7MmFXKXhXw6EWBtl7E+CHz6lzIb+BErT1zEoM9zzmI
0N/IJ3npaW266gWEAN/aGKPRh10f+yFW2gOvLYONokNhMdpb3FKWUMNPK7uZ6rJX
KSyd5XotuHeeeaPN1OqIgHGVb7s+MC+0ymLwUz5wGUIKK4i75nZ2WsmKVvxmcea2
++ddg+AOBH0Y9/kL7Uvr9Bk4SogOlfwP3q5/t8t3soaZzP9UmDB3T/5+iESzBrIP
pKC3HpFzpKQdhGR/IvZTusHBCc+aMfk7QrnYJexgSx2/sOKCzPydM5IzreMLnum4
8/3oxb8RZIcjLEMrGkcAeuij92qZFdDu/VSqwByMd9ejGjriEnGmtLMrHiaPEW97
0d2DwZdrgxpTJ+3Vebi02GZ5QDLVgHF2muZZMlsp2cwFSGJQ55lHSG78122Pdxsb
hS0vdF2qG/mNIBwSX1dBfWSyKAjUQt/UlciLB1KBHQF4fLQ2laMCagEltgJfLBcS
2N6STYEgtxA2ic4lYp3ZJdl5rO6bSCqJWlxvoFtk5S5UavEB8oI9VFeb/DtH1o5B
tXE+mJpi8XGCXfjmktBv0h5MM8tgM6itnvnofOu9BzogWMDIvLh+r3ETUZ0t9sGo
IhfX7Qx5PX0KxbVV00ewrjYeqAFzUXrHJmAqd85aKcTsYKxw/BfTXoHg2yQi05YW
tmSy3HFE+4fdKJlf7yQv1SPUZpslSBnu/vcpmH+AW+JUqbf7CgMaR3LP61fxxcFq
tKyE/tD7bpBBd899DL+/z/XNmTTI0Y0KGwU+c94T6D4BV4Fy7jcw2tUOKaA+qlDI
BSeqVNonKN1OiR/cIy5gjrvwYbk+L2hy6eQXoR8W96Nv2KW9+a5lGsnQgd+UmKKs
V1CnZCXv6ZEZEamkfNBk8j5tq6xc1+6SldwNLZ8oAqtgSC5OGfmqmLK/fNwUH4JE
qxkhAfB6JRFqQEDkskQw7Bf6GexBBPiAN3+Z/gxNKrfDGDBEEfMwa3wjDG4Xo0xg
vIvdQp5n1w6tXholbnIi+saQQK+ogE2YXKkyFO3EsTiSi3QDKg70UNpwGcTekF8m
Msov8bUNADHRT415DTWYK/yfUIsiNdWghUzxfw7R6rUvxsnASptpPOJxX78aASPl
ZiEIyinGiZC6zbsq4ATewGgFk2sOqA1HJ63SeeRawRy9uemRhxU9Tj3ha+GDnirL
ju8cJ27PsV2XYxTncMMSiFo/juinO2inZBCJ9VdGpRf8jhTpsZOhnOnAR7CR4LXf
iVZHXpkcWquo0JxuaV8DqgwhVt2ktmjaKnzib8axr1YM6/nA1pMYBTeyeLoh8lC3
Y4GgcxaujOh4OMpct0kkKKtwlUnIyPRUPm0f2yzxMESNguUUd0NvdyRiDNXeHbIL
18w4QgGn1JgnLiVi7hyBeimcIWAjIOSaj5bZm1MTJuO618g76R1bkXui6JGDKbAd
n+OSUhfzHyc7tiVisJZcwsLSD3YNvuS9Ix8EF7pwZSVRw/B/gXosIlfv5QfiVGzd
cO9g4YWc1uFLcTQRpHLU6W7AoNNh5Qh6OZJan74e0GBUX+rq5Mm50xSx6MwQ//aT
XNWHvfs980RIU2nA2sHmGTrQucskANlXOoDsqr99jEA43esyIfcjPQKH2GCDk2lo
r6CWsA3wJ+W/oAEHOaAxlugo6OFG88gX42hdTnctBFAwMxyaP/Ws9EuIRznJ4vJv
P1I+SKfdOEsJ7Hjg+cTAgWp8/IRivVNna/lx1q68Llya9WJRP/bbJXdOufUXNk+M
gYRO7MsWUWuph8NCqtbhPw0Xl4vuCd3GX1wxAvpIZUn2AiZXJ9sEBzVBWhNJgrbm
xCvXlGO/WAvw22GS7LDr7woyEVG0GnoSKy+5J5Pzeks77A3IpIYH6e66P21b1xvO
+0g4iK5iPDDKMK8Esus18angq2a9TbPxiPwFpJk6vDqr8z8+xgPx8HGBXtk4ZK/9
gCQkBMrMY7QQNdXs6KfJxSAYN4h3KhxBtGUStAN/cvkB+TXkONu7uilEny2cbrUC
VhQ76KHzokM3FeaRN6yh1UdozShCP8KTjVRU/vV4p4NDzsSEvPZOZRzPW9rPAPF3
rArRl7V31qpokPOEAlgAoNJxjLUG8wI71352IR4mA8oSa5pJpRVxVt+DTBeLEAoZ
L+U3piaNs1iaf5Cpi4DHMKlkwV4AuPGFJpDgCt8QIelhpVdTXoAd0Pn+V6Lqg2h+
xcxBzuDV048A2WAhV54Np0sf+h9JT/Nqr5wonzxTA3YcpcpMt4bS/2y2pe+BFAq3
wgGByJLNjC7yVaLDXb66peGWMl5YKUYxtxMTTruV7kosOsZuW60AjZhOkIGqNgS3
A2S5d1PQwlPaKRi8927+lBtknQcL8EkHpeDQ5GsMP2VvXgRAyDmOHSQq/z6i0fcL
sCr0OtKWd4B9+C4nmdq7EqJJnrMnXsMaVycrR3sv0fXJ3BvkKiHy6PTooVyzWT9P
Th9akuIYI3qsM4yHeosHIMvt8UC2/b5NIPzADPag1NCUMBqN1o+hx4aR4XzNqXSM
tXDVtZzfe5gNLqxdztBA0IgtuNVtundBCagNljeLuAUyP9oPHXKaRloNt38bSXCy
aD1OHfzKOyYYvR/YCGFxCLV/6FHTNJyJHCHs/F5wsoIZbi2glmktP2gIpGDJrjBb
fvp6qawME5OJaesFHO0xPnBAGCjponJf4gHhSPBk8e3AUca7Evqvh4xEW1Pt37DU
tYWjuQ4BWn0ELapWCVT2Mewig2mDAWhtaUfdzHZDYpCA8Yl4V1MDWnd/IY6snJln
Tl2r43HZvBwKu97rPwq77jI+aeKn4CCPOtkHXd1RGZSRTfpgfAtjr8DO+UnLOawB
NqyPb2Qm2+b1x75CDpwJYAx0oQi9MSgjNQtcMaGCiC3HV172ARhDLB5Pt6YlkWqr
PETQT478MNRRhu1zIEG6GW0TT6r9Q7oiROrTjWu1sjFVJ0rsBRtDq5gwBesHPevD
nMxh+GOH2TkXaY1Be+eIfbgc0uN4dIkMmGhqGsG3OQZ1s6VXrvpJOBwuooSEFXVN
2qOOa96EbXoSsKER5WJn8cnJYZ6kj5p6jYMQUr6pXlzdigWI5S+XcLo/OY9+DM14
3XqSZmunN+mlxaXLzfxG+D9I9ESRKylv+1w8o9F1fJyDsYo0Aj03FouuHdTu8xfw
KhNrkMC435shy/AlfNdRFIKS7ehd8ktnE+dm4k6MO90tAs8uPZIuisO9UfSxrrc7
reHTf5IggLF8H7/AqjBoWpMZvEV13R9GoE+53m0bDSps6K2yd1CDlwZFO6Ku7qfE
KQBp1xKuBnlEVYedMgjuT+PzEYCdvl6BIWIFJrPVVk0lGPCwY+SWCgzVMjAE6a4m
xMZg3Idn5QKr2iHMRO6QfwbL6Zexm1Zj8phjvIrDU8Qhf0Ms/+2NQS3rDJkVp24P
N6rPQBAnYSjBpjILMbDqJW+1FX7QeN4xe5SU0n5j3kpsMFrg86QXDWs8XickQ5sZ
hSqE1XfDFINuJ5z9dMpIrBDs5D8PzzPaXNGUTzRPQmkWgW1G7vGL6PDJ/HtXTHZc
6+NjgK3PTIjtPCfopeHoGRxEMT0mLiT96mibdnIJre/Z5Nq0GutoR2mMK2QN0A0a
fcbLVA2mumZOWWR45WCj02HwrN0pSlPJVb04wYIiTD7FWCIPqXATlLFwvZFZ7OUq
C4Tq5/Vzc7we3IOGcCI9LJ1R0C5eTijUdqmYhTDjt5QuvJHxQB5p8pUiDw0IUgPS
kUsE0+EhfvQHL6k5uqBFyXR440nC+FIGwH3FaevO0V7aAOmp7Y52bY6H9MR05rtF
wkWh85qjiadUlSNQnx8R/gJ1ajiVDfIifLPLnTp3pnTpgCDFqD4hmfdcPuUM490a
BIrRPY2lsppCUIJ7bKRhWcNyEYzl8Yjx2Rmd3+mEis7nKQTAOKWSq0cL3ZOiT9Pn
Xc9NRX41+on1v2WTsOemapPWqKqFb8Bv7lG8d76rV9LoJjWmd2Nubhxo8uobquvz
mVBWwlhHc7HJqYyfTfYmMTK7/mR4LwJuSjgv+mWl3rySdV9xZu1Lwz94QNVvSB8b
FrPp46VEhtY/EBwxn9NPHumHvAjP4Y/nW5uH5vzsPwEEhwjaX6IGX6yYRPb04I80
P+/eK/tYXhv6h2gtNithiUjvZkKlS16CMX2+OdG+v7NAYFpreG4CKzOSAlAtBDc1
Hj9vcvwspff42eRi1staUCa1tjJKYQhi2BQueouS9mI9wNR45QHfP8+0S/SxMHUF
rCR5mWb4ioPtaR7vpwWIlmfFSOkGvcho8mfmwGH/jQLAPeMK8yfCM9yPeRFgN7nH
/NR6ogBA5OJbOg51eUat/1kNUiUXmpVn8oXM7EXYraK3paOtrDb5lUexGkMjeY/o
k+4zmQHwPRZ/1IJdE20V+nDk3D2p4r+TxPVSFK+QDar9nNv19yAJGK4b8P51mvL7
69ATsxEnDSjgkc90qth16Eto9BWfjoXHUeieESpeHVWyer/qWbsHGNCKDSlnz2zN
4ZNxlYO9z48Stzm2tVgeOEaeflrEA4OApwPP+eRTPUsKZfV+Fta60MuAFhl40ykf
QD+lhiX8nUNLs9tY6+Fvm/knAsoLrVgMIz2ckpT2osU+kcKGgIfaLyBKJi+Wwzfy
Fkjeyd8gSyOsUd0jk/iInrDYA5Wk4gGtZKFA+R/2lB0Y9y0B+q3T7JoZdDAIn3n+
/osXLduqmXY2InbIMWK47UkieM6fc6SMRUSUH6i6FMNv9iywC2wqBfrwRqImfZeK
/TBUWU2l1aCAgSFQhji2BwmjLgRdLnJYeSpVhE3NNK6dhb87Z1DBzNZsQdYrvt+m
U3EKsO3TwfR7rUkrHwXFmlpIq+G04Tlmv4z6DsqBGsmLew7Cnd0KMJGGloVlloI2
q3kmF1RGEhMUamwAv3YvW0QKkZMPL8IjidgFfPFG76BW9BR0HyQ428EH/34VpcL4
WHJkRlh+oEwWmB9GEp7x36wqLwoaHVWpE5fdrAo0DG9smL8f8Ej5LfeJHYqvrgSp
mBBf1gd1eDdwmlsn/LIAzAl/DXD2vP2vssVYNBaTrsSIcGbQWd0zC7csuRrfNPtd
fFT4OYG0ryGLNf8Ozog6yVuOnQNotOOHdB9+bU1V1rBZNaEWDEWBUwQwZIApX+3Q
vKnUKPTVCW7NRoxgKpSUC0/sVuvj8K1IKVBK/zODN7rqaNt5trzhHdUzDD5S34hM
6IngokhnglMLvTTdWxQsYfjF1M24TVDC3pL1vxcbGf7LJnTY+anWd7wYplmqppoR
uAfVQLIfYyMpCYY17x/oNI/qIgEDCoG9w0p6fctY+mDjeXcGXwlS44RFW5/Na2/a
4twHQkWkKr9e8VmBRv+RAtA/07q2nJ6w+T3KzSRu1ZmYhfvAScBdFvJ5w5rWkc+N
BDoedOcgplC/Q8lDVuP8taawMOqIHxmwCtVSDplDYennYg82ihTyZXq5h0dgHV3Q
0Igmph9P/x0QPBejXMQVvaBCzxl/7qgDCzjdkzDCji09/boUuQ5tE6566ZUnn4ZB
F8uA6gJA90/aGpEjWzLrBQM0cvBSPYJ/WX2F9S/YIRoKyvCwX8TiGSeaxtPYw2+j
ldAgyENUjZDN1x+pX6I8ImMuLHbvw53r7eYRCskYJU4pe/xliDtuI1HmUeTm2hAc
4I8XhENib2y0tNKlH8Y8goF8NkAmh2fcW3ttm0T4PAQP/fVBvhMEh06uHmpIno7L
bHEHYB6zD1Asp6u/lRhTAmtd2MjpMtyulljX0vj1J7kwyGgICmWn02QnHxTK8e2s
GW6K3QjTK9vQR55Qfb44FA068vYb/6izh6+VRCNjca4qjMJY5L2RTJvHgt6j7tDo
JvcUOG8y9iJL/PbQRHpmUZpVs89P9jcgj2MOjsKN+3CDXyqBA+PY3GIiBbvRMHe8
3JOgZ8UqN9d5kqraDpyhUDo0Zt1m7z2zfqFtffVZ+i+K8mlcFgalM75paJYigi35
mRlbArnThYEjFTYAc7MGQsTVrviAoQrDqnjgYhqMhRdSnNgmoriHE3NbFc5sEEnM
ovCKX1DQOR9bNjeNvRAmfOMo1zi3XUl2V50OAxreVWsGygzRGo8l4X8CZP602owy
akDThchPvi1e8C7tE8bd8qMxwMPuXcgnG4gSJU7yL2dj8bfa0QVyB6mkynV5GSDf
WnmZdftscsDPO5ul/9Eqq0AixCCircMFWFf8zOThHXhps1E9p/OkD0FHeZAwHFrI
cKgBJ0pdUIxzaUdsZ96par3C8Ub0DzQsIOBTnN1YUfUw9Akt+iiav1XFOcnADNLh
R0IzQvoaUMV3OZ31dwAEX0JouRbPBLKKxFJIEacJwnS8qwEhH/H7qWzeHmTMHoVO
zDhAPmHqGnyfh5Cvnt+favp9MKqn9vpX+T6t3K6oMCu2Y2Rb6Ztvpor8uaebGGNQ
Im+eazuMUbSRFfcHy37VHy/bHmm1C3aTQwdIdXb6p+BTJEZS6ZGzmiYAR6xIziZS
ZqnxU3Xdh+y9TzV0ci2drpHIgWp3JZF4Ta80jyHPtLJBcvBYbE04CaRfURrxXX2o
zQxBm2PponVHGjsiegDURIR6MbDUOZ3zMcmxEsECmw7RMF6Ets/3pnOA5OjJ0t00
GzUQoyY4pDrDXFvomqhn8kR58CcNOrBsQ3FXPV1KD37TjPEOnhxaTY2V3O0nBV5a
bn0pCdYamZiby0kUzg/suCqfgwiDhE57D0tdZd8ryReBk/E+5SvpNsc0cgBLwfUw
w+7uv6H23+d0/yULj1q4ncxNaVmp+TD115ectOSM7lzEIU3TZwkf9I7x5IMU8vpJ
LHI8qRUySwbfL/sVH3fNOWI1SPhvw/SJrt2eRl8GBnnhOzdR+ZnLtmh04n8Rq2TW
K8mQ8a5Rdsi7OtVChEXx7QQ8wRtEjWpt6bGgdH+K+ybg0Qt9wqOgmh8NRPrqeFJb
d1WfFKwe6u7XOBPqPsc9r9iHFVuDH9Tr91YAkj/h7Td7fZ4MFOBSLwfRj5z75YGI
cpCz3z/VPDPjvM2A4CPGPR9U0xXpaXqZEpWSPDJTiOhe3OlEk4JsoKOqGs+hI/++
jL12zgFxq9rblMvMSsinu6ryU/23XbI5/83iZuvjfobLen0/A2Lua3QiFUC65O3M
gPXteNZ/pvgOwQhKcbge21eZbMG0J7eYI3LTcvMvrDtmebJsIm7tIEPpVSOd72fX
lT7yx3zKEPkGLz/R6sLydmJcb4IQE4u/UZhOZIQYyLfDqI+5LbRxIKCczeLDNz6M
UanFExDg/zewD1OHfLEGSsOjTJ1xvbCbMwf6jn584t1aAQGvfH5nRDmUGTp0UoDz
DKQsw2w8LCnVc8wwceq9KWSRRedACBYigt/sMKp5hSZ0gmamhCoddTyP1VIRsthF
vQkT3hCvu5LYiDED533gcg1BItTPJqCXInVgdbbf+xHROyETx6A2hkVGQoPDUw6i
h/AlzP7Zdqh3xDrHjnE9IjYdNAeo15RwpKiNmUcz+muxgnJbj8UHSOwCFTxJYPFd
LRDSV7z8e6RpnPqhoyHMfcYG+EIYji1uJFWXrKVyYGq5v0qeHujR9ti902tyuaM7
xllutLeR4xKbP4bL2UhmiK8OP/mC+welRdvNRodiKsBaAW8GMrIt4j1Pn8wYUOZo
MNDz2Nmw5/R8Gjq8o5vPgLbX6UHUeJJKj1bsaEp1XBku0fpNxWnXahYkT/NtRiV3
WCCGpzgIDX18eulB4cuE8vJQGf/7EngAYecAarM5E+tSGXRzAOYLJtGbUaTialMU
wxF+0a/5hQS867wJ1Jl9/4QvvLkjZ/5w0zAn+t9HO3Q1YUhqndXpEyS8dQrWSflv
K50hEAOgqKL1VRJ04ibWQybO+m3DWJJAQZ3ixsmBHnZwHujeCGqDqdo6OQNMxOLl
sduJzE3BDBXhuQeo30qtzvInth+TLYUsy84pFcvdtMM9op+L04cCYlbsdMMEfxY/
Geb95QYRyZU6GgZIfOzBZG71dsXd36+hNAcItAD3uYpLZuzR73/MhfpcWIC5O9ar
hi84hLsS2XjH4s39LyaSM2C9OZew1++MnlGXMqwVTrgwHy2pxmsUZL3AcYHm3r9l
+Z2BLAiRYVgV9YZdsbEGdVqC1zbO11I/vmg3TZkD5v2agvDLyyzKiGkLcLXItQgz
/9iaDz1i05cAkux6c/tDV6KJHQIm+9N5/yG0lq9nH/zpRdNkAhL1ymTI59W5Lw/p
QPJ7ikP1yE0fWM4J8B0wqrdeCjsyuq9lXkC566q4ni5r0q9AYTkpzKoW+3ywOZAX
Q6zer5TPdH+sn95nqRs31kO8ENFRLuu/taL34JZRyyihwBH/Kr9PMiPWYbRKPiF5
ccPAzwBZkfTBFcijFVGcHZLIUNwHirgHlyGRmT9WVcvDi/7zs4sI0dMMWs3NBsOi
JKEigplC02o7DQdtkO2WkqvsRw6w4wWQu16sckogt7Vk9y/h7NwZXv52BOwarUVl
OyFA6vqXye/sSTudL5AAox/dhW2vD4CF6KzruQXdS8oDb8wgpvyOe6ghpfyn3onH
75eoeOXN5Tjf5oz7x44IXISYaEyyqJ+ccPsbTH6erknpSz6eY25ndhqpz00TYfdp
gbGNigqc6wQyY+ak63eHcid/cInkhAMSu7etCCNPo26l5Ik4siczPUzJ+5YPr/av
eCoxIYYAgRVODnvqVN36ZY9wPA63py9KuSB+6vABtLLz15tYXYW9iqwmt6ykHYWA
GN0j9wIXHX0COXhP7htzExPNYa2f15EJF9Mj6Ps5qyGel+50mkjsyBYRtBF8Y/6d
CmpJshxvklgNexVohEt0bsJ99L8r3ztD0rm7I6AYRhry3TKy/2ri/ilMPODD5nOF
hCMBSyWfLUb8qKEhdVmMPG1ZcenkOAIWEFNn8epvX/ZwGECDrMSNW10iZXjtVOCs
HIDMehqPQ0JH8tdgwzBWOerE/X3BIEUwK5EvCu8YLUFb5TGTSAZ1cjgvM+6VgaA4
voqLrrH0q9AAR0xsumeSt1Euix22q+rLt1hHT0nEBVxjjvXSAwalQ10pvdwaPZQh
9/2qtk1dvDwfCPt0il4PQemy4XP2SO7gAKnveH+e5qs0R4ztuW1/kkhgAdPKdLII
jg3hHhhOPwM2YiOCy+zU70q2NWDLqbU4vBWtkJU/OoA7kyz+lwvSDx6fnmuC1dQh
sFAWB4uF7/EfYs4rU2B0dAf9+SyR3wRMdq9rpNB80rsx+YlYG2nIS8FKpa1/MhB/
rzs/186pixHgu23Aiw5z5DtXpg3Fs+5Ng9pPUJ/VKQWX2qtzv+7l2KJpcNDIvdoq
vjroWMqcyRt0LzFqGpXUrSkvP0YIpbeVQicua0kbrB9Apk/OzrjMuL8rTmBSA8KZ
Cof6Dfh0hs6JqmPzDopwhgUxGRCsvIOdNNSAHrPng6E+nkeJvis3h1xXDb3CNHyK
YyIf84vywAB9drZrxIlTtfRSNzmWg96R5n51q6ymPHRhVMVJ7YxY0AQuoTKsJOwi
5U9siwMbTnmp2QwxMhgQf5pNGTy7ob49Uq9y81LjXbASyL0Aj/HJS68sp5kPRqnK
6hlHrcJUsTdARiToQYJLWu/xF7cDkWUV7FFBFeamrpRKUFmH+9wMEe/f/nZgXR+/
ly97RI27FLU7UHO6A13dvvkYHB3X+nJtCXs1786BPyDlrte1H2zOclHSdxBvfBBg
c2mlpC4drxWb4mf2AGlLyUFdn3frg1JWu7tUsilegpmvazwgxjy0axe9ID23+5J2
GiPNS/8Ww+7Xba0QrILwSb8Mzwh2z8M6kPGOK/VAWXPW9fJNBuHJ0VOSCTL0eCXz
zP5+WfzMlZjLMKSsk+pwdPZ3eG7Xny5my/vSy6DnE1/lYpkqXOMX+hSbalKVrO8i
MQfpJVhmmbP0Jhn6sf2+GkykWl884uzwtXMyeCFkoZ4OOfNANwhntqnqB7osVEG1
wiKmXOLBcQpHA7A9JDqcT2PWTo5j5ZU0DA5omSO/s8dQlElhLh4IGunq/v7qw5FP
8hY9O3OiKBaT7mh24fQZeaCVA7cCWzKV7qq6rLGhOLLljxOr4ikyLP3GBKIyT6XX
htRLqkWHlP8/jWhonJZRta5sg81KhMCK27t4kBQY7XgU0cJIKaqQOTmJm9Wz4sSs
I7VJ1KdZ4oEVcs1hXQM6uXcxqOJPcZQLToIeptcEfomZpb5fcM+ijXUj+qZN4HdI
fw45jBt4OvRFE4ChSIGYTuEHefKQADNbCFjEv/Xso97/sBsOeYFnxv+pQyP+kd3O
oS3kiWL1b5WqcuJqSgrwlOthAV/mVeap8kYcFwe9Is7OULDD7SdySGVLup+pvVwv
sGVS7XC3f5L1y5zhVMQ62uz3EW6AUaNvn2roAfLozcRZh8mikLRr80C0NgS2BYrV
mBRS71pZ/6LiBd7Hj5FuYUBSa6md8EJ9bErEvXh33p+rwZ7Hsv5xvCvgB2nf9Zph
wP9b/gUDB5Xwc65EhDttoUwM9G88d0p0/WQOCYmmG4IPyXdiOnsdnFWhj8/uqRt8
bfqGdVuplce/3AYuuIX70k431rCu5MJP4K26BQWBSBaB3ToSfDLPgcveWNYQulAy
u0xGvpSox1vUWqzyq+07pbhSqKVEqc7L3l4ITLgVG0fKrYdLOPG1NXsBJw5tQfXw
9v6S4m95GvHTztq3KQ2vaQSHXejjaMv6YAFCTLBy3iewWk4+IJIGlWsCaOV1FHC0
X69lUe1Gk3FNWj6s6jnVGi4YOcU/63fApHWU3aAztObi8ewtF7nAf2BE5dQJFcGY
bDWL2O38wiHSxaMJvjCBLyCaCnEUWF6yakQJuATKcpPKMdbxYotx/yx/UiujOFnC
EnJa/B25SL5LGON/0cwE1UCTjr4a18jrxrh3SAMuz/631QV0yLZfHzQ055duEw7K
P3SI29NQSyk1oslRcCEt93VSyC91+It96+xoFlGwBpO0MAlqECD528xdqI94qCTi
R/l5VmDD2S0aSa5mLL9Z0uTvrEAVcLxAJU8/9ijn2iScWfZQfB4Y5sK0koUuz0dR
qRM7XmmBRMX306XmMfMXcvK7YX6KH1oB2vLrO3DDb6Mw+gUlnUKkWN0ABlAn4171
dfCb5w+0uHzH0wSQrAaJ+2vCe6XpSJaTNHX3uu92beNWb7MbJMxELWfRvNyvCu8h
TUQpra4CGxEmUA0UIwqqvYLWvEXXWMeumP+4r4ulpYek4RTf3wPlTHpO7Z+964sW
eH9cUJ+6ZKApDOpqZTFpnBvivpAqTewLRe2eRbSOELIdjtGFJCv56gpxvD1caEZH
7JoZ+M5rSFfi8Kg1d8YUvFIxvZ+IwvcEd/lN/Hw6KSHtZ/y3KwQqhTupQe/2DhXz
ByICyjhZPIpHQOrf1hDBirlR2RvgklPoXirOSI0yYWdZCdeVDkP/B9wLH4GgzWdT
hdU+RDQqh2mrgiGmPrgxn2aK7Rxuyaw3N3pHsMWFsY5R4L4UNK01HfiVdaVkBN9e
5rpvYdvsMGEe4VhRgoIFcw69j//GFaimEGuFzdfUIfUxT6Fb4PpJThmx6g0UA3Xr
ur0KKDTlZ0xq1UFckamQJKw51kTkiTnijKdLR04tI+EuVS5zO5EbSPtPC/0Me4Bd
4onJLf5C1zLIOpYJMsznRPfO7sC1ZLLbu3LMjFmGUBK51XipNDYDMI+UB7kDfDqY
9+1ArAirMoRUSLw2D8yVKT1Jt4tvnBnpJna+u9ZviUGU4JqOaHmqKSxa8kRiTe8z
uvrPoyz3Se9+k8a92V8RmKDfJq6k74Mea6xevDn2H4t4XuSeKtP3H3cu5t22PRkw
yqmVI3Tf/RwjqIiA3f3LzFox5JBWrNuVT8/vFm9jBHOFuSUH/OnM3jU6+cKnMKGP
xNxJz15liDeAXoAPw1aJkj+9kVbjA88gFubHIeS+wpAJVx6JKCqDbHVz/F1a7Q84
q0RGXuKHdSisYcnwllB4P2+l8f3erA2FcDp+5iM3KfWBZX0fYFsBlfZLyBy2OzAr
PPvYlsX5PnvqaZUH7WyxrvGt0/0euAao/PAlU/6t5/dSI5qYje4wHgFq3XZu/iZ3
mDrFfzSUV3nXrnGCOjR+WQ1wihtELmPxwm6xkTPS285EMU49tK3RGwGtaJNtjZ+W
tKyeGROq+Ne0J9vrPH9sb5eqcVSkEyLx8Ds2NVCGr2Jd+DEfISk8UlEMisdhhda4
4BS2aJ46L09h2ApcJCfdJGZBXp6mZ5Y5Vryxew06Msxojq6hpHmQO3CAhJ7XJNS8
Fzj5u4cZY64kgckz6ZxhW104DMj1DF5RY3XOa5jASjc0Vs0tXZWoEt2PYsVpTjc0
WnTLyyjVv4IMHZjAcap9FSIkOJzPiCSMc4yBJ8nzHRecgs81QpqEU8Dlg6adRYAe
d2tLyvuqoVrCaon7XS0iPa5HnGFpqyS2hJQ5dqhxDsF5EuS9V8wVoLRja88EJaLs
MlprHVZ4wiEnZYxhgHrFDFPLsxYGEzGnaPISUJrK83fIEYC3RnUibqaRAxv1/BnC
dYjGsQYoYQ230ai8Mff+qqk8rze2IN2CpfpW4g1sXZXdUy/QFpZBG24c85vvMpeo
oWA4CIvH/dQJUVWjO+JG466jEkDoqbu3Kowfwn+MLY/ybL9YEOOijtMd5Gedi8+G
rfc71ccrhbn+yOzXdLGouR0rI0lx9+iKr/zWAhngDLMNJ2lUk6US5Zf7uEXX3bMe
bobyJOclwLTAbhj/RExs0G1I5KDKiAxUEvTwX2GUlXNWqdRXc5En69cHjkWrUxdN
KumrfpTVppIEEGbKLI6wwD+cxT9DBwJwg25i6/UQU9Okv7qrS3sYsO0ehZdQMja+
FonQvGclC7TW9hLkK/VmuPMoXDhtyOKRlCuN+KF6qcb3K3mz+niELDRRrMUjkRo5
7hj0k6D0V4JnfecEzAATRbodw4/YdtMRImDrGJFQfevJkpNfRETwNQYJ6jftiSbd
lT5pS8EqrgeeleKWldgbGeWzJHAFfySlcicEcBdxLBx4JOaSnvLz6njtYLvvn5K5
ffv1kIXock3h/nvPdSL2UN/w5Ere0dijf2qATFPwxonbOICrWXxbYWrHgQaGQU5E
mo1DnuZ6/xvGaqJMCgqOs3A0a2w2Ca9Hu4/+dJ6olhLeKc5sfxF1HRQqzBPkDXUc
TqOPD1/1rgYCw/ZhgTWVC3PxUv8ixwL2OOUu41IJS9HK6yXDHs/sepMj0UQ9D7Xf
2HvRZkfyArq3GYZTsCSogf3182/1PkMp7B1TykwWvMU0a9GOpKLBrBKFVnQTSFOp
ONocEVvDBrBjhF5KtrkvYYGdkY0oZIDidcBAY7iJ1mV8mhXsc6bxNT5Mio8PkTdZ
DYK/cK+UPanOkE9pJZk1I7NH8zukjnFlOPjQMu4DH/94rpJ2J+MM8kG87d1T3on/
FC0+HutyiPZn1NOcJe9LtbvtOZGNOFet/R7vKoZeh6UfuSfB1hFG53PpMzOqS07R
qICAHon5J4JgnEk6wZwjKoqIvRnIhsSif8gCxPtttWoxNd8hyoTMZsPXofSuLGSU
31fEP7A4Nkl0qyScmLQDkZ4f3rnGv5cXDdFY7eYDuPvbpmHuo1g44RvEg+UvnJYW
JtirPE2q3MI8GT8hIbyDZ9EZvO1Sp2cE6mNGTCbEanzVv23D8qvR+EdgLwoBMkKO
AUM4Wy16Nhcn6FQW61AgsgaRpM/m/pDQ2uA7lq5QFpzToHYGoPbnsUcVjWe9AlMu
VtBvuiqo+p9HXH00cL/4aHlRuj49fR41ski9xgX2nznGFsbHSFwEBFv9AVSjRjEk
Kd03otjAcjO3R6VplsrjPelCsrNxa19CpRKHwxpST3vTI1czM+jxbJk6iU3Sso95
+U1TYPyxhanI+ss5g+ix2QAtvl1qT4PQf5BZBNz3bN5lH9Ub8Jt/UgMeRVwKs4Ty
GXr1nCWXrUsQa90wG9cc49DAuZO6ny2rH9fAswB7hY6etxE2X4YaE3YUn+41huyp
wUAsXuDw8yZpQg/gpy+Vcujsi2GJRdaj1A2VA9UKAZq18gkMN8DMvKGGabHKiLTw
qGQNmWCe5YXk9EYubTyCy1q03p3VVIwSuc8UOFUc/m8QjK5424Gi2h0nK3i+escn
bN2QREeqd/ntyP1muNnAyz03jIC4DOETY3R41H6b3L7F43sbfqL2HZDzswqGvnzF
RoWM7BlxboXlr7gS/QB8X4LuAxPbpQ6sLQ0SwSTku2iqn7nhGeXxbac85i8totqd
vCk5VzqzIOxBPh4+uveFgUidoe99djAaXS8AQrJhEvAHzbvZf3zM1KS6cYsKOkUz
w8bs0i4J3y92Nyt+/UoSV3kxpgYhkZ3fX7a3Zfbjp+8JdZM084LbyUvQMg0WMSq1
K590+c3Aac+wrSVS6SFhlhKRmgc68cznpqmV0aiQ3+6VIjNgdHKTfXCmi/fsYaDQ
np8/eIe19XEby7RY0LVRSnjeQrXb3/1skxFzciEDJqOLY+tbF7mMxjI2TxaMqCA+
ZtE4OmMxAR8t+Y/daQbij+DBoRYD61L4gCxLamdcY2NFQD2mEIbyFa08t69wMANJ
tDLtPIYZzu0GchnOFnnDU5GoNZn7JInoeFCJ9arOSutAEJQMNwCsl+ti+Gol9GHW
uuHJigsg+QkIpMbHTLzny2ItGUw0qCjx06hVjQ+QH1cjbn4oj7PjPwmkXPzMluE1
ORF0b02JhQPRA9dvlQNkjOk2WTdm6irVgO0BmX5BbVaC1yrFVSTmHBroynQD4wHe
apS0HGDdLZZ2wKqEiEu+91A2TejnfshhVq50Y7NAyLcx9ziKXgiE9Rz5toxpntjh
v7ubpvcsuciT1GlcCjBuVOCaOPS0lK4biNwBoPw1ccUmKy3UI5GzmplU4sNuobYy
X1Ch0NZ33FjqFDuziw9x2cZUYvnS29+KsAcp5UJTsqbhZ/guuqUCt09ddDCixgG9
ih+viIl/YWqXaOlXPTvS6veOcCPpScGvTNHE4zO9kXX0yEWfCUTqwvIhasZXM+ck
e616m0yyEPWNLgJv3xzVTtv3E8QLxoAm7M6QI0NsRGWqT4GWtycDkjaMoFxXrTrm
CYgoBkGMnSo5Ar2npyQQbC8FWj6HDUhamGsnFO9GJCOwMyuI7vYnxhpwzOebRBJq
Z+zbuwpnSTG++StKlu9eIInX4OzqabjU4fny4BAz+l3w2usWud/J4I4OdwNOHRNS
DlcV6agV1VVsvxEpG83R9nehQXfJOQ4mN4CUij1EZzhG2ETMo4uBFf9OuBIa2wQg
SRhAeGKuCXUhPRZAM5mrqf0DYtXlgVSnGjsPDMpZJ6eKo0vlXCV1go4PAKJ/VS9b
RkLptlyoo2I0/+V7Z4kdUd2hMgP8uI7XMJBYFtjb/sJO+rlAzcn3UpBZJe9kJkGL
Mah0RIFKIQ4iegqNcJil5+3XNboMiEToLx35Vi1Rn6LVkIvfQBRzTCewEaZUJwXE
IZrk/PBKnTAqChO38SYEaPvVU8VJMWKOnErOZZr6OD4w6GixwWfMrdLrFQYRgHP9
HV9GnuNh/hCMH8FROyq35RFc+h3+Fb8pHi30u4cO5HdnvjcFdvkyX26aViqv6xvH
tRpvYZYTQjgd4lLLeYbzz14G3+qTNkf4hKOpHUsADgCfFl3IW0abaPP+b8LH7bsn
Onyn2veP2q0CUhZTsptm1XDfnIMmHApkWVimwOLhpyacI2r9PiguvKuFx+t89Pyo
owjRnzhLKr0W/lMubXmqp8VcUIqTwkD8abAV159zJTeJzmF/ynhQlOD2mPEWFTPW
dZwhdvf0GVzPrmpRBLAjI3z/KDyt/gNDOkMzWgrZ5igAQVgT/c/Cz9hWeKzZEQk2
NHa9+iuqyCslf2Dqfe/ByWQDnQevCDcyjU18lsUulSHN1E0gITtN4cySReK2kRP0
z+4n3IHdwMrFK3x+Y2EvmrCQBvxoD8pNiJFxp5SRJfQOkOkViI5qRwYAfIUe7c7r
u22HpylJBSD+4FeGw7WZA9X5Jm41YjKYE9D4LvHjJd5CxFdw39FDTNmFZqLpaH6P
uAIoidkRVnQ0sLvzor5d4mEuZ4aYMwAksMeqpMbDsx/DAJ2G90NgreLm0fZclP3Z
ycwvQQaKQIYKp0RVkSfReruP42gsaYUl2vDHm+DEy7rLufniKnwIwxTO4+ieB1A9
7euEIb6ZV5tA6ZVBCq5RQuaH/PC4ygb4inilzYDL00VD5W9vZNfy7UujYPQwuag0
hLwW5znP3wLo/2qihYTZWceUMebu0PvJpaozDucVHgOHQi9wYE51lEsHEcvQutY3
V9W0V633i39YqV8ipIP07ItDTlnzbS044qwX4okCq4zj5FbKgY+AD3rT0QTOnmvQ
MGvEwJ4ydO4ku6xFzxblX2Aw28xD0yGIvXAgvw6ZMqfpFJVUJillzmizlPPSfDXI
dqqYMSRaqF2TjxA0I+7fbb5tUKeVrYp7t6wdPI1/eTAX3igmSIC/FEsL42R6QbN+
2o0WbrmHtlzsxgEvCCt1j+U7+HSI/P1vs3pTEbjqY+60Jyn6KA0UzX5EV0YsZdX5
OPLTOi9xoqggoDS7Up/+CxKsfhNKqQ0P07NqM8M6BenhtCmBJop7SmTbXte9T9H4
n5O/r5ZKPMSivFNX6spizWfNQ6lYLI4J92mTDHgNgAPgVaj54sqk1Q4mZnSoZ3so
SSCoNoYL/vXv0obCe88hlQSvojKVjp2GGDkJLUOaxacjQIGuxmmpOQPEPo85XAlZ
aKNvJALA7GC2jadOvWvYECM62MVfcLHKEw4YRHhL02ny5f85jpmTogpZkLs00C14
OLMbOXdxCkUgSVulD4p37EaGd/gEwj+P+yHclOBup5LYjd87nWcyi2CNtF3oA/cz
x3eq+CwmG9jrPduirarS54Vf/XHqLzKltrnZJZKm921N/07qqdSliE33kbEO2jTj
v3jVobtek51c1eevyvvWMyVZmAQ0saUyAYvzYXhCY9xUuKZHgVRYiSr+bu2RMvSh
TXKc+X3YJva6GUWWVole0ydEofHSB8Ofkwdcro5FRrO8MUuYL8N5+A/9lTlkYp9h
489lMeFxIjojMZ2rdY2eoIalYPBdU8nhy+ZWvgU4HozPSg6Dg5iaS8VPMT5qb+O3
DR10sjLKaHV6fwFp77uKp0ovyXkiXuuvLPHsglgK64SJlCMp9hGk9jK+lcXulDWD
mMUIQxTyyMqYzEOZ1knsIai3G9sF+CFNOrjrNkE18nIfqG7ynRD7kDW6CpmWQ2DM
T/LQ+8LCFCq8FKBd5XCWPjbkDkhzKl71MNCsS/qWKKOqC2rHkeDJThhmYJEinO57
N4nQoTtO32CrVwcnvv+w4VbmLHoX5yniWMm99CBcafHvi6fHNpN1RqkxV/QJ19o/
Ja/tke4xMG53PyJogfyxV09sb4CMbGYO4UFystpVWOzbVwYw5IlPLlnjq3oivrhx
gxskD5Rm4puJx08BprAQ/0DnE4+lUGX6WDtdNpeuUBqmbvjFbciioE/RuMCKOxrr
2A80tpJJelRD/GQgIe9Z/kpgc1YdALbcJe+bnnhx+QMDBGsFwvxh+61He+w+yMtl
WlTMwZ09Z6hIyfg0FQ1nA8OBzcYwUJQ3ugUpO3GnbPZ5sAQQNIJgVtkoaSSerkjr
4oMaSEn37/tD8rHmF7YfXuV5hKzQE5ddA7PH5VqWXd5hLM7wcPkMLLyW00gYuN6k
pjfO6ZBh3XBvRIZ8xNy4tHxb7sSgOpZMJBza1y5eyDhV6k+6+DmEm7nWsvBCTZbK
k2LiH7CAniwcLUqOHWB/ggAOyrS7N0+vX/O7kXb7tBfGrJ46rjS3h6zE/WbzeCmX
P1EMRoxPKkn8S/1hOiyGSKVyC+JxzLtKS5JmrnU2yOIlMFCIeMl+ND/W66Sn3UuO
1lgKmjyc4qKocZh4S/gOwTdWbTqug84D5LCU3a+flqVx+miOkQdhsJhROUJQZXmA
evfdJchK0tkEEzhYp6jK18sDIbToxmsPCW9K+2FCMSP8tAIGanYnD8beqtQT+G7z
SIfutiVNGaBP3b4yLxquPFnIgi2K0zlIqXVOHodVlUGP6Fy2JGQGcWeJC6guDnom
bSE0wQtHomKjOsR5+ftvv9ih/fPKoeybbR4vjXOI0B/oSr9KK7gsek19KEWKAz2l
5ChyAcSdNXedZ8c5RfWLUdVxJt5C68pL+3Jhha/P6V83WxIQT4op8Ugnq2rFsL2x
or3fFD8phWaw8Sx48l0neQJeJXmxeu1zu+NfnlF5TKsFs/Tzi6kevzWnN0mmTsuA
FPJt4F7fsiQHR3x1BJjk4XcGLWu83++s3inGffBE9+6CIRfQDT0Acbop2GKqJQ68
VB3Sgh+q21sUslgawln90c+zTAGG0NoFaDbrJVpefF3NKDwH6lkJR26Wj0m+cd1/
ASqnc5RfMrjb5ha13zttCcd5oJ4euZgN/kf5BWSbPTMAFZSkHDlb89kxJfda76qV
VF30d1HM1g6+ZXwCMar4Byq+2esTwPvyHRv20C5qsQ3/82dnRggAJpFOmPExTzI2
T7QbI7G0qeduGXA4i66U0T/6JGnuHN+KVyehQi6Lvpk6+3WCK/UCaQ3PYgah8ebI
JB58ymXTA4i/6JBxaT8FVVm1IzV7IZHj6IHGx6FgeV+i6qO6DJidQcVlo/81O1SG
DaJFhnJoKleGewIHPPW8yJm0nYZx4OlkzHWNpulmbQYfOzZyOo1DdDlmTnPcwZVx
h1rebMYvFN5lUzTcEYn/BW5lb/RPr3x11aCzBrmXcaAIJ1nAN8jwfmmm98wkQRpP
DvCX2WXoM9boVXwDHEbUjvxWJSqMfr0eulc3eQahvjhT05GyKbSyxElv5VUX2HUw
oTjJV582iWYfNw3BiUN+DAplAWT9hBTzeVfpr+NHZUhV7TtkxhzIWzDzrEq+lS8l
+/VjNpycfCbToOe0VdlGaZUJqDcfN3laTe+dKPMZmonKe8hK+aR5HLJ1ah8Uo4qT
aL16HCMcP5GqpUueJW4jmR/hwDzHohYkxCW1Ao+jdGAjKzMVS2NdZQCwFUVWMPX2
JD+FkUFtZT8s3we2u/gMrntmqoBBdRsmHKd6SoGK3T6Sie7o0oH4ZgEtBP2gcFr1
mnk1xDd7WetS2fzlh+7NYuiULCCMF9JQe3DhAMb9VxUmDqKZA6GBH/WaQWIyjyw+
gUOVWOsxR9t0m5ELsOzqfNvUgbrFtizblZhoGr9TJK65TFJqkxdguG0GhhM6b7bZ
ryYRPO96l1JSDMTHceH2FSPLD1MXudOFTrtbx50fUC3LWE/utgF/RihQnUxExCRk
5skLyGju6OJmpR66WQYuJmp3bn8KM6PC7lUCDpX/3ZMlP7IYzvaNqGO1AZcRb5v0
4ZVq8EXmhz5qVHUFgZqcT/QJ2/OvZTKZV9tS4Fi1Z6Eo8qycSQNoyNMh+vJECK18
ep7aE2dLy4FMiU8TrUZPnOqooldwiila+TYU9jkXrA0J6Z7Psod47b7T9un3i3hm
ti4+TZrDNOPFEuvTsHJLksPUOJ+n4+K7WOoxKxzQ5pjL8fkwzBOtF5Z7mIiliWhf
g15d0u+MKhGqoDM44lYjEmcWRRJu2UR1uTy0VA/iaDBO+1vqiNOocWiSLtlzXOeE
b5K43IGQBvDwqJnEFa+dF0VKnGYKeWClLIRgjfwpnCjQQsTqhzK7mVQSFNIqj4y/
6BMJYhpKEyUG/TaplDeMdiTD2ne45fxS6JQY4f2Nxrpo7h38dGXGJAz8dWJHsrc0
wanG8dW6dmY9ocoHlXJhrI+cP0mczcOSfSLylyNUU99Vg/ur7Xvx9HR6s5DG2VJf
CF/JcjSmevu+xrEMJ+x1yx4Ux+trNZTnIi7hKqPM+eCba7+KIQD/CHqP5Jhq4WN5
q3K5bI4OYdC5quNxnKgxRzjTOeWkPIOYoVFxYnTw95cQ6rdl4wKFL2z142dI0zVh
PgrSOMc4s/InnB9/uyAEuNm7Icpq0HUrKmPhEBw1dOeY4JTif6iajR5oK+oqfPFh
BRTuiUXkXfS6+3YjR378t4IUWlGSySfCH5YwgjFogAD/87ojphyYAAG+Dq9B4I7N
eGL621/Y23CDBlDZZwWJ5p6rPmICo3vB6g6p11DUbxeNaF/N0iP5CdAmPvW8yR+/
8T3XxEd5NM0jVj9qYFT27Cq6hIbeb7YV1b+W+pYa0rSw2Tuy3yJ8gImTiygFI74J
ecXsZWdHgS5fWzz12z4uYBWZQzvtIcohWFMS6xzjHFYRSRvRmulu+JtCh3mlThFZ
J04ZWmRnN5lGmavGuyNJJo1HWuRLUaMJjcy0D48aQJcAnHqJaR/oxFFM0bIE1UJB
2GnZm+eCXpFA1sb21E7KFy2pTdmLxrNTM2+jhIaSjxpfUyY0dvk4u9Tu7wXpWjba
W4r0V5X5rpSQ5zL7c5QDoD8FeTo9kzHF0vmLL8/EAjhdzmjj6udueQZpsBZrL0j8
IfIJ7+O+5fP9EYD/SIMbapBjeIINcdzeeWAyvK/mmSmzDSzsix4IWVj2Cdg7CIBR
wXzcuYcyVuzTtmvnst+ZMXejooQxomByHsdLj2iQZNMJnI1+lLQqJBp2L24iCxsr
pg8CUmg1ctOHQYymh07XK3qbVf63N0vBQXCaR9rCXSaphCi7VJC4VO2rA3kZO+9u
FSxx0QUqpCrhZAofz0xN/xjK7J9zXNFmZsKfO6t9C325xrhwQqhzLal9XtxIIGN7
qMO4Ox2D12vkfaqaEyAJ4M7knSRlKhCLLJA5neRZ1Wvn8qfmD01sCkaq6pDasBLt
cHo4kFozFWZYCHgnWHPNPV1FE/TzFjrFKHDebWT0tCLyrUYSokRUdWpTxOk0S4pq
gEIFC/g2XzDB8dNwas/yJ2dLEKO2oTW/hrsfj+SNidHJhl0h/Q0PrcvrC0yEOjjl
xQi/qg5MqqCkQYLmL0e9wtRvZnyeBuTMAK0Vcy4DQtTUB4zWOuXLm5M9RH/BTADu
wtaWODC3QRp5Rq5neEYsiIxRRAzHnECRtUkmwqXqt8NjiCeQxZqEvP+6Z4hpp5x8
gisr6u6/kZTy5SXCg1z7qagffq/FSUXhoYdvGBP0KoubdYFbNpZjkRiYzAGFp5ia
8dhmq8kWB+k4o2N6NkLG2GqXaDyG1fFmXolv9aL3sWH5GE9MipzX9DTm44QN6SEU
+6Nxnk2TIzUB2UM67CPJFnucF6i0PUrBmbyyClx83MzXhKddACrHtQeFr242twm5
xXkSlwbKnQTs8+zHyJ54WTMyr3i5gDJ074IkXz/QZ3sIEEKLYVlAm5lVJQ+jQ0Fa
sSNezrbULoBWBc74m/TCfHXJtnQs95ytKxWUaiQljxBrVP0BMmZfTaLBmVntGxFF
sx8lmeUMz32Ub56J3LyYt0ZooTJHfoXAztl1tXz1U2OVcj1RUw32xyP1j9OKln57
wFFzuzk3vc97XKsZlkxWNnF+DH1it8uGu/pwXfODam78gevtjiRuxvh46xKG2pfJ
CHdexheAF9UYSF8SDpkB66D4zaETV/q8Rax7GD+rnAXfvcS3MRDoX9lOyzXtL1f1
Mko/yAL+CNOuNCZ8ZmOkqYxM+8W/5d3+53zVp0r/z3I5gtn47yuWDX6zSBJvNNPT
YcPpghGRdaPxJTDa35CnWz/n43Ffc15hP32OAGbnj+SmMNsEeZYEvI10nzFRw73I
QL0Yf8z9pOG4D1JOeDKsfvYHpkYjUacHWRekrX4BMSSWUGVSX5TH9uBDJ1wLUa1x
Q3KrN2ohmQu0mDy5kl61unc5I3L12VsLyYPw23h4qfO+N/DccmNpJkASphaqZK4e
7kFYxFtHVcex9UZ8pnfwmDXO0cCY4IONi2ab3sa3fmHJvakjYUnt2vdUijatMRHO
HTpQZVTJxsDHwZB6Z6uJH9QXChdtggvYOaL9n7U8RQ8HqO3kIG7nPB5EUcFVThny
wHmM6FoylNY6tHZzDmflMsJA9HbVShvxnpaoMu0adv2vQm8m31/LT7Dau1BOAVHY
l3L3EB0fT3VZT/0vg4j88+nqp6hkQMCVTPOtQHQRASe4pFWhxaoPIHFzYGrCFYOV
jdZflT9wh4W3fs3leYClOrhC468TXczVN3qdLeu4+HnOvyEdQJL1mx6s8U4lEuBr
pnL/MYCZLHcgXP3uWOVBcGNDi2c8OQT6oWt53jK5QUzfS3hSBqcI8xXfDYgGNUE/
ov37G765jj7hJat1Fs9x+auCd/UM9OIdr2Ywk0KxzyCvEp2ccV87Q24Sry/P1QMR
0SdIYXAqJ3dYGMDQqcXvjr9Iq4NZuBY7AzW28ZL2EAq6pI4QvHmHmmkGIAPIKG2Q
V5JDlMKo6eGvG6qfwnZpzvXboVdAxs1YNps1vezhd2cbXwq19voyisRCHEikwrXe
U8UF96rLywtkioOq2R3GZ9euMY6ZsluPwxYmO92i69HgzYdpsiJ4JESy4UQGpHtH
vXACl4M3Iv9Y0MDmTj2GQ6hfB0iFD5o9K6mOkKHrbIAC6NDpYQDLf4ZJQeaQ7vk9
9yNDid7VdOFgn3jHVZpjD+MifQW8OV8TO1oRgXUtmRV7RBSekuYUKIaP4nFgkSaJ
rp50/Yqb5YKsCGKawbT/+9QyvUeAoJY5puPtEa/QVZ+uO57519MGrFeKuFvl+PQ1
F8qHZxfHLqGvMNzO2zFurzVP3b94c5P54f87xe9joHBJ5pHJ9tXtliKxgL3JvPNi
1KuKIOuxRHZXHyMEC0/8kOG/kNwNhVWt0cXDf93ei7IjIU/piftqTvLQG0CrjkUF
XvaTZ7P3YJau/Q6gDwJoxeUES+ggr+OYdMxUfw7863T+Ye2iBQuPT3oFQUp+vp1i
wnX+mm07ETQckMlkycCdT703n1toc6h8mPIGB43XoIyMSK24nxApU6QzKwgZzk+C
ReAjOIQLNC0VaZeNE7B8G85cp7iuDwxeEA4jesraBRVfNE+l/2xbppxVyLR1al5Q
ZcYBfOCn9mgS+w+82/2VAejaj6lAXutxdmmCmbuaxAsgfDsegECS+07r99JCpT0D
MZU4iglpLK4mlF9QinqHtAPvk4RLaiFHL3iyVKVJL7dCGjOwXtDLfWq8Eq3CpQXy
nPJkiA8W2EWT3rVxEtRuabDUpzSOFIyxxraupotiDIkaTyhlKiUw2rJ6UFNT3/Vo
um7O4N7uGsn3vlrClRRCRDVTNBON9mBlV21lAg+b8SfyhpvmtaYdv2h1CRnkME6h
ytT/6l/ZQZFMnsms/T1zh7qvPKLa6iMcY246MWU23utqyd22yEzriV+8XXXi2Odu
Dd3+Sk2ST8j7bMuYYRAL13QC+abXuCeTBjXPVKyxlTm63aDWJUwQ0U1TGgpPkoyq
mLX5RHKnf9I5sJjpW+hGnpMpFGx5v+MU2K4TkrYRcoWlvydw13baBpLxlIkqO3q+
dPg240b+I9eAgYXYAUN1xmqD4IDRAaNzJ3pKDis65eSFsXgUkXuVkAA+GNIcqFK9
nCQOGFD81sg7Gn2dbn9DU/2PJ7KUlaTNAMHlXdCZJp9YjO3p1/r6wR4Rcfz9DeQ/
fYKC00iMoi1H5D9fgAMv3bWx9phqv6xOJjTAlQnTXYEp1qznW4pliWp+bFFmU/Yc
Pw9zfEc1UIEkYm95pXGbGn8pLotFaa3VPSQPAues8D1KX+m6+DlHLA3bNEmna3sJ
9bpxsJ/QeT+bTsMXmydP8IADHYbPRR8pAaIGHu15V9tAvDM7h3FVxBRgaxP+1sQC
Xf0CnE6vl9hAm8DRKWcKESI7h6ng/bDlPv6fKaCUBCrBr19rGsWron3OrkY76gPu
QGgJGBr9+M34+mXYp0UNC4NyTAKNbAe0ZVuHmnYL4NVRi7VfwEda5WjvjJOkVaIc
VN37QT1ZOM0bFpHxamz/ROhH+hCpr/QMG4T5xMlHItfpA1mS8KW1aeAh1L3WarPB
y1+bpvE9K9op2oKOeicXxzs1+0EG4IKcFEUzPcEI6obssP7fqaGE+IEn+wZn5RRN
6/3q9YZE7hi0VYkE8DtXBf2RtywRNtk2+eh8xyrPYfL1RcG8GsadfF4lTBdfJmv7
Wq40JX8EZI2gxGZStzzTIGoj+tW/NN7H6coSJcXKOO4lnRXWBnRGfpn3Fm4wxevK
U8Lad6YQritD7TovS9iftnxNlIZMQ/ctWvfO9UG8if52uYycR0yb7Dln91m7P5HH
cjXz5IYNFZhRvr5nyfFiqmSQsTweK2glDfUCe9JhOgeBVJB0voWFK0XYZ+vjAxWQ
l1uEdwl8COQYd+w09QcOTGl9Y30LwCf1N3vi/k1Rf7t3lUIIDSH0x1KzcF+idMPB
ijAOs45fwPveXN/H7S1Ggt/cYnb+SFFo8/Ehm8fC9BHPQdJqKp57xexPmFCPV4WW
sPAwIrDYmsTRjCh08WkecVL7UMMqn0KtX/In9HjZdsEXg0wDtZaegoT55Ln/dXZp
KI0WqayR4n9cFZCmY8t+D7PEVlsWB9SZBGB36PFmLVXpDrJbA5ptIpjhn/RoFuvd
yIuzkxm9kn1dWB2coC08JanzD6iy4zMGW0y3vLP6ZuqBxRGhd1LlhNjYIxF59WHj
UVJ9oOnj/QQ4xuAL3uQyazEna6r6FVfU95vWNhm8TUTqSoDa0Uco+VVt0EvgWBZR
ahsNtGgCGC54apISsGo7lTfLSyd2viFBGQ5QU8y/vDBFkvlr50163Obrry6RqGEw
AiFd+v5xKkdJWGHz2o5BnHm6mEWqPpbyuDdKhWRtQlJL+SBGf2R1LMIMnnGAftUV
DGDNkyGp1u4hL5lz58uEiQ9odcU25fdsxno/zo7q+5WMf+dik8IbUHCMlb48TvQ8
UguA0H5JtcfYswU9/b3Qx0AV7nimOjTiMIRHR533sNcSasjtnGEMW9zyz64oKcCz
67AEn3+kAF85Brz4vieT6fUaGnWY/NY0xbJb6NBUmux+w/Z721Ktal7TL13iAHc1
--pragma protect end_data_block
--pragma protect digest_block
V+DA0PbEi+SnQ3y2FttfD1LHIAM=
--pragma protect end_digest_block
--pragma protect end_protected
