-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
--pragma protect begin_protected
--pragma protect encrypt_agent="NCPROTECT"
--pragma protect encrypt_agent_info="Encrypted using API"
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
--pragma protect key_method=RSA
--pragma protect key_block
f1ST++bS1VCI7pvYdT0/vsOCIiPTIMo/RE+X77DqxAgBJ5GhMbb0IG8MIioyBXfA
9q9iaO2fmoXFenVds9czA4K5Li3GEZx8e24E1DGpm9YMHbkbCz2iYHxFKm/LbWMy
OT8x4HwmqxiS9yQYum161PXCSoDBwPm253Sr/BJ+YhNANJCpr8m2V5k/Gh31Sy3V
r1zLMvusFprMYnTLGYwAyMuNUKREq2ypdmGMWwCinJvrUPSbHuNtAR7k7Dte5uBi
d0r5hkJ7RQgnr31OA3tiRA3QuKvAMZt9bk/DZvSvq5DJsyGoy+RQdep3zJwdzoGO
Z2V4MCOyUHpPqMn94/9zHw==
--pragma protect end_key_block
--pragma protect digest_block
H0MGrVZ9t9pZVSSbVlqmcu0iatg=
--pragma protect end_digest_block
--pragma protect data_block
rc9MXrunYRLEnFn0ref38Xmvzq4bWv6leVsqEsaom5oHvjjTXEPhje9W6lYTcroR
nl6mxQ0k4dxuIQwfXRreAo7p5IRDWIhRtIkOezUP5/12jYSjiwZ92jfRDY9pnU8X
tyNQB15/Z48u9j8iYXwVw3d1X2AOCeIjP+nZzI3MGtdYmRXitublyyRFNyG6xlDl
Lo8um5NClpr1l9gV0w3T105BRGz1EziiII1ydZnfbeEJ1RRqlIHL+7lS0uZWKjWn
wvu+cIbLBAaz96xlEwSMh1Fje9YRuuSk75aRmiZ8/hueFrv4A+hX7SA454JUjWlX
wWsfgQOuqOOa5+wPTIV8CRBHhbApJOi5TBCpPDOBZW2+MWljpibW8QkeflhAJdUb
8H4cCXf+4avWodgGtMsbvbNaOXeIFvgSuU8HiE1u4evXwLltyh5DQ52vrURpvUTl
7YIQ6air2+H6Qh5P3XyBIbv7XK98WfHhj6MbEUvcLxyscC+reqaUhTfpjwWV0poD
UJjmKx8X5rFgBRJ/aAuPNOO8fW4kKeSCHc8pgmNiP9QYp5rxxRj9Up8IqeCKanag
t3NAWBNXcDjqtTqJPE9XRjnOyAPwWHHLfoLkQuIoCDMnDO5OC+9YnjYpAzyKzcez
iw6Zq+Kutj5LcuFt5AodbZwOtWcMBB+zG8rgxndhSBAwBpEnBDlk5ASNk736GctX
4If5EW9fDth3QTG38lkBFnSKL06pSJjIxnIqTxz5CBdDnMco3J0LsDgTVhyY4aey
0X1zIhS/e6Fj8k1oJY23LNqU6M8rQaNMoOouBbxQY7k8dfCoNAC2CObjD+07yXzk
762xBRtHXJLa8V5VIxhboRu+4aGLFtP8GmJrBrNg/8smPOdpCVEFnMgoQ+ITt/jM
h+4QaGE5KOU5GUmCi4zuLfwANHM5b+z6+NvkzAmHqgotgpJzFKPiKXblhVxX6gti
Ntb4OqdKu9Ea1Ct5KEICLsfkUAEs+gbwGZKyVxZuQi+R3bIGrSfC/vY/kMazqjvC
oxJqJ3divXwmv58/UmkNYZmoamZSAjl4IIm1eNgIDJtnK7I/sIhKJgJtkWQrj+rS
IMePG0qs+OQXPxrdw8OfJNb+gLSJN2JzWmxXuBuDvbQoJHVzUHY9BMAnNv9bqq2V
F5Ej+v9yqnSNnFpdAI579+CagW3OrDQDgZRQqRmq0066Cx7pfPkTyxX5HUmOCo4F
2zacMpw/vicJlGdpk+LLGgLPyMdNp/JF2kEoTtMaxXQfWt8O57OzbaqnGmuq9pGh
I/3q5VNWNardQiGP8mJP7vDdov5bDuflAc78z3G7ap5O+j1AX8aYUh+FNdkuWGJi
WUQ8Aty5E9yw2mRAVN2Hb2IqRU8lZOyhElqW3W9WJJagFrROcE30Kf0DcqgM1llM
88GU1x6BtpI/H0f0TKkb8fmaACtNnG/UBbnJeoDsAKT/3boxuhzbw1XWVAHhMILX
eEYpnwRNztY/ghoo8woRnVBxvsMT3hq0WygoTXSh0cQa/8On+/+TEhgpaO2Gtv0z
vrGkx+d1jdjj+4GK0gpKgG2wwRb+0PQVRMW69qbd9rQjVZL1dEb72SiFIPTGZKeV
bDYKiYVYPDqtsAZ+FYjauQ+dWV7BhMUYrTpSmIpe1RfgIQq8e4BuwDGFGrFx/yA2
YB+MhmRhd7SDeZw3Xh/8SsHTH4gT5+kBxPIAqlYQZDMwZhPekJ+k9TxoHv7bf1O/
vqle0GCrxTexR24ABhcbPi8Nu0hWAsjUIajofUhr/QsuhGFyMs0VzJxsL5LdkdN+
oIWrPIa6mO620/beCKGoPVtjnq4DCng4SUJf69YppuTjsViKC3a4zhQ8kFbVAuA5
v+lgJ5SOvMS5adnId5ArgP/FjEB8fKh542YUSCbXH7V0JdVCVyaqYJWqCWJtgcL6
LHpnELKL+ILEvFPYLUWrcigRNQSFXkJ1gB+SOzLFIeIKAcgBUPN/OZFYw4LVbAuS
K5NxNgMuO87A1lV1gr9ubP10sqMbR7dbOUYWTz0xh7G6r6+P7fYvuNaSf+RWysWW
QrwSERbZzhHdKtx8RxTvWMCBjOs80s4s2O/+dkon+qk/x/tl6qH2xY79lWJbk8ym
fZ/xzguB4ICiBLVByE2ORN3uUbTK2FVm1E066BtmPYJQyEwxrx3N0vsBqeqe/cTf
Re2FRhRNWJG0/JvEQ8cc1eC9LrXUYgmnCHxZBJyE6yC+Pb7aAVyiz5QqrJfMIFmI
d+2ur3bXBtTgujh0ZA9tHmhPjFm5iQ58EPoCJ8NRI06Z49Lzy1FWqe37v2yxV+Ua
BgDrWYSrIVf6q+xHDkaVesD3VXEBX4B5X8xm6RRcqfBUd7wkqiAfjufuNvKOlU9g
xUKYnVLc1UKAlqVfGwluzu0EPjPa+MWcuFBjxHtYlVi1pjvTZ0psS4TMT8psgdo7
xs24nu3jOtpWJQlPuWNVBWuGrZkm4nNBlHd0l+uZ0z9qCx3TCuz0Jyf5y5B/RlKZ
2sV5Y06VrReFoPFw6zUVrCYopOU2oPVhRWC2HHVmiWtYtiVT7LZ/5QZNCq/k9ryt
w0ZwSMiFAn4YywNimrfVqq/mBKBQLGnzGdDpqtZ5p9Fc2yLbcGk654DVryiA93c9
wVIvJ5nbC34KF6ky1ivOApMOqWdBTSktVP/bpcTvD6CKdzJrlHBdFyN2puhxpfGi
VXSTgov1DV/Uz6dvDfYZWTxiVBfi6OpiVZ1frsu8beacVjTbuqnmY6LkiNZsPxdt
3+mcVV3Pa7uFbIDr9LV+fWDPJnMLGnRCHNfesUDg/Nstfs2ORakx4puJPC5D81HP
QuZwAIy/oFO+JGP81MSKwYiSDCtOIXLUDHXJiJfaLV3o8J67nTEFiHI5OzJJ1KfP
QVM8UOdj0oxQ+ASyS4cgEyJsY90OXRw8Q0fACATKvdDcy0CNTDJwwZRXm8lDOIe9
3Kmqlt8g6iPBJ7VMi71kpxuFTKb9N+mqYotRoE5b+5kb/FWrxhXq8O+JvRftUt+H
NlFkqMXunuO/4hkEewOizcuZd68kwED5kGSFmbs1EFQhL9cti34fEl6dalWa3SuV
Uiqr20oAhQW1i4fPawT7CNK2mOOMU+rEvq7uFnf7Ip7iPSQUy/5/q8JCHgGWphDc
rrK7G/qgYon9/ez0h6wRPLZHA0wM634cTzj0nIKwfIBmpYalSsXSfTrd1NpiUYkP
ShNTto2jmBEiX0yEW3Mi9FhmDB3N2+AkDMX+V+KFgn5MyMiUaTc49x7sS9dA4koo
YHOd5zuiLFkAIvRL9cDkHbywVybelRFPvI29CJlaA5QK7JxFcAijIReb8Iw68c6H
oKOk4A3w7TshZfVGjFagBomUGMJVRkCwdXXspBrpmHCNSDYcCGhWvvwHTrbDutiD
Y6Wrr/q4Z8r4BOhj/e2EfokaxCMB571F8YqXzj55/mEW9sicyEN6ZQD2xySXAsuA
C3Q6W3eCcceiHhDfxDruc+bvU1WHxZ4mg/Oy3DGxIn2/0jjSKSWD+GXC3xbSYSdd
DzoMC+S+zaO4QOxFntdgl6ISGlmUrUZJ2T2CS6C5AxDEdSu5U6cxZx6CmGwL1Jcm
T2xNlafc5AaqawOwnr1F2JSnKtjW3RPZqiLtM2AuQMZTca2wsc2LpcRAgIlWHjx5
fPRrpnACsyZHQDn4BJgV6CVTeIsmZOQgR7lRQTEvyA+ZSFXP6kU0qyV+SR/MMGZ4
fnDysaCmmkZAR+NDj2pjgG4gpqid1/TdHQpEedvvtpnW+2YqwhlIzt+DC/QYdCkD
rt4VnJrIh0Whx0j2sMRNi149ejt+ZSHRabSJczSJFk5htjPX8XeP8KaZDqFCou0M
h5x7pxy5YY6iSWMsGSPour4mtYi3VjYtmoBUnSrWZZ3YFDmDwItnD0JRJZv4TnkP
mGnE4hZDrPmwpcCvSDRmpmvHXgeSz+qwNGmmi7Yw+8js3y7ZXmivsgy+bSl9tobT
mxC64U3XdSD+43UCjkIPhb8XSAcLf8Pi3WkrnRJC13hjv8VUffq1VhP4Lb7yRJap
gWGLi2vdo0d0t2SrjeyEm+DHlsEsfgGp5khapxWM56MkJbfZydUikjVQoBRs2zqL
u3UrTG1E6b7IJDMiFob+OVi4ViNTcC7CZ29NBFqmAxbyAC2Z6+YpGgCYPNqviX1V
UXjVoA7KCI2ZhxL6UiZGq+h7TUud7F00nQEP4baVcTEa60Oiq4M9ZYmoEOUsxlZr
vOQrIX+3CUBdDJd2d6q611zqdEOqozYz7JjTS11Ad0sX56BEaJ2gaIqOds3sqvT3
AsCwloJlGg19GCrVn3+Y7ONeXwzRJxirswEr+xrxos6JnaE3sYg/T/JxsgxvutYC
5yKXBmXeCFn1nav/HgqbU7Gn9Il42PVEBuagPyYSvlwG5wJx8m0/X1P7yJZjJLR/
VeUaiGEXJCYLv3+LLp4/hggMFt6C2Y3BnVjH9pqizfO+ymwAwVr9uTLyZDTFL3XM
j0nwhuiJGeKiaIFM6+TCFyh3y6eWtVW5KCHuGXY6+rpPtz5PEOGfTn6eF+ivY1pK
idDaoP8eo5UYHq9WKor5SArCm6nDR7xuER3aUvB6UA/AgQV+rE14DelEf0e9bjEM
OUr0OS6R7wkIHzdvfwsCPSkNmRWz4+fcGA2PeTnpSZ75T8yHjGkZyJBKOc0+qXW1
h2qanWj0aneISZIuqrFMKupee5NGNt4v87sUJSNAet0d85UrZS8pjnvZR9ln5Q63
qk+LRAl67xsi5tfwNnCuin/Jn+1zdjT6FLnR+RAiP1gV4R1qZJaWBGk638UjShKD
9W11wkRPfS6FLH4MS4iKaNmaT3qnRcyO+nn2kBQLNd8m3XArWaeHmk+/biqHLE0g
Pb9eKCzuSYDVR/Zdg4EqO9xyNRYbNUb+ta58EAIgvNJoLvo6PDMGFMWU9SECGbE5
rP1pa4Ce4ciQFwffCcIpB+ThsWgJiCKZ5cz6eSXma/ovUWRUpHIjljwGslPWKvcz
KUh84/77SZFhXBl/pA2B0Q0r/ny7hqhyet9vJCB0aqFbbKXDUv1cbK6lSkD7x9KG
1+u/1goOF6GTzUDu9iK+qcImH9M379pEPqfRk1AXFRS8mQkSHXcTofyNKUILRIj/
+G9FOhf+ZYjC0MRKD6rrQlOf6As0lkC7hiUqBqUn1pi/fc2rppbkFlaTPJlS30Lp
fOhDnC4mDHAtLrUIKYf81QTl0LzLc/3PGHkuBsGixPvPFQ5pD9AkNZNKTGtFtCjt
p+j70ISGc97ZV4vCpOicsIE0+r4EGuxDS3eElLyR/7L0Fg0ryMygt2GTe0AU2Fer
s3H9ZXLo5XfWUG8VTePQ3uAdi7s4YDVMlgNg2DEvivoV0VCyVGTRFz8F7k525Bdj
da6v0959Q9gqh1anJCU8z+R2xn9MU+tuZ5C/0l8hfFRobE9Bx4Xmt9fSNTrtvCT8
OKXORUEOxCt0NkWS01hhL49TR6YU0o3H32rnZWH9fLegpzmGkbM51oRQ4Fv01lY4
iVdzGJCd/5sIUefDyBgL+vNC2kVCDNAU/QmAfhx9V457AcF3a9+qAcC/eueSJcN2
gIPulfUSAxDyHNavSkeuOFptX2Cu+GdS+IPieVrxA1YsjMgPZ0RGXqPd+7/kZZ8y
I5OcR3+UHc0dhNxWxcuMqNuH5LD9CapR9YXOuE4WxqGF3fYxdACbAzl3SNeeXrxB
xudattr2iWRLmEvmSrEB7PMK6lhU4Wh0o6wbxKwb2Ua0T+N59kjHG5z6vnTTw/H4
+Ms9YdLceOUmyTxgw6pnqZNIfhJ7KXLytmavJ3qQYNw8O3H/TtU8WEG4wUNP1YVX
kvWGA6W7I9P/fM5BCWheKCs+nwr1fP+cD/mvAlBix8ezYfR7wOL6HdP9OGirAQsd
n3EZwXwWshFJjxRXu5arygHkH11szBBKI9WzjMni7FmEaSg5rxTG8JvT8gCOqWkU
NqtsR0n8BVAAy8ZxO/xtace2Xtg/d/jViEonbPuBly7M2wyPfmdoMF4kqcAuQ6e3
2LF24nJlKkydayW0XCXv45UTo0q4MG+9vrj2oJaQ2uxtJkYjSL8QVakJ5QJVVDpL
t5aUEDZBLcmsdjiQwJf4XYh7WjBWm+8YZUWHYCAYYRaAzTa88liHEhuJrX9LaGs5
t4h2LDzwpvAIro+29VK0lXDom04ZJX5RDAacXK65rDcjDgjP07lHYheey6rr2q2W
/MZCMuSTtPkFWFarmTs27UgQJKIXKKdmrCF2MoWuUlOU4jLm6mr8wJrYpjrGvWZ9
sdbgxoNHC5iFdgftyIJgzVjTOJAghZrsa+Brl2DwAQvmCtKmIHg0jSVuTxUlJ7F2
MMYBKAqNHNizVfwEa4+NRtjUdEOqiUSmii+t4+73BjezhAl9FbHXapf6zFwCTsCu
CLMFVfFXQ+u9KY5URhzEJVL5Gk/iyHeY7p3URKksZFi3LyL0PqaIgS0Bho90NCcC
6jeu9p6tP+O+0r75t3l9p7JVz+VRmv2WZa/rWY5jYIsEdIrC8D4YfZ/DBQXP1Vri
pL1Q8CZmJMFRr1/jzkqyTA==
--pragma protect end_data_block
--pragma protect digest_block
b4oImmgODRjaSTTQAj2PTUzLhlA=
--pragma protect end_digest_block
--pragma protect end_protected
