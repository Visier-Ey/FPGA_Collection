-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "N-2017.12-SP2-4 -- Oct 23, 2018"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
ShcCT6b+AmyFx2+Lf1DTU/CpUvJA4rYXHZQCzEoANMpbthRkmNDLmZ25h4gesb2V
bdHY2vDDtBY3Sar/itUByhQCFwQDP5qDVhxIo0wnM7s9a2uKrhPB/mB1XiObU4iq
yVMEfED3jRuGzVcKPBnwYfHDo3VPc1Ix36evTpkHwW4=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 9440)
`protect data_block
b1ZY9zbWiv0WocOyJvDSt2VMG/QQ1muxNCKEGVhzbIuwMIhDwuAftZxL09CjS8mm
zv8hSaQI0IQs6BKj4fzALYSg0tQu1/wCy24IBQTMZ6j5fG3tlY5T/BJ/5wqYwntW
q3pPBcnav1b6nRPzl3GojztQKjtBHEDVJk4e6ZsH7euny3cS7kuOFbJqfGetz5wE
04fdm9SQJMVyuySlAUKa3dgEg6aAjJjYcK7C1T3altW4g2oH7S3fgy9gNovtv/54
nV01Q7p8pqvqcDNdgoVdT5xJwU9W0Ox0y64D0s/xCyPCQBDlunAO/NvsmlsqJg91
UHk1NkJ1LRNmBHzXye6q3XOoYgoUGC710VIJ1rIelQori7yrxm8TXp4/ShmfqqCz
tG5I77oVwtO3r9EpoB6/d2Z2PvrcVnRJbSS8WWwB0RS1JSIkpqbMLZ+4+K8HaZdE
kdo79NcPMsYbIi8oQ8zJYw0+PqfdYjD5r9fp1pyjTzyfV2++ZJTuMuksGvJdu2Lb
ljfFnujoWCYhYxACoACmq1pVxcu6OBoLOk3LmehAWFdbCRYEM8kkNo5c9lW+AU9h
O6WDoqnc2rLGULEkrBlCqBUByojHYWM8QWMF0CIO/DzYCrrzwejjhmOSc3OwBQHp
jaEom2fT91DoHv8sIq63dQvEuYSV+ASqJoTsQwpMpXni+K00jt2H4zVHUMrWrPYa
VyOhAc0LdZEoQgFIc5kpN+e9eMBeVrNRltnlv4098b+pVjBPPMsxF3XHgJQ2505T
zxE14G/SLgvmxDYRZxpM8DsMyZHImLAkysdP7uKNxmCG7n6DlAWanwyhqEVkK04/
PAQZfrnhTfLXC+/QUMoc/KO54aJBKPzc2Rl9DyFdSMCPzcMVi9zBJrHKxJNJKg/P
VTYXlP6cKwEchtnFnManX4m/W6TebScaxFgXAPi1DwCSuTG+Cv8Adhx4pCuXEUl+
GWfFTQfHzlzzHvxbmsZZP4sbNrjxi8cyNJGLQ0Uq2XHvEBmViA0qr0vpKONTTIkB
1UzumwZt2F2hunZNd+3s3f8/aiBvU4nqkuIRIE7H7W1UvBAqXdbpugEd87TGqwJp
me1jqFrymJZhC8ELWSibIXLLPnO0EPZtTLKqHqZLy6JvyRQIZRwmBYH1fHOBoRZl
vcb2aiou34orAd+6XBuR4B7k+pxO8Ac0r9shvWEA2WJ0Xw4HT2g/sjdXWH8QLHd0
cWwPfWmnjIYjGIy/+XrSl7nSGIpSwEM3+aN05uIIWcqL+swfmmfXMQHbxVREHEDR
gRWyuX5OEH8vdRoHGYWNHriYCpzm0JbOWBk3K3t0/FSv8XvlD8x8RWn62zfQgDTC
5lA0y3hkchXpFY8JtdsEBT7HnyV5aFLMXwZ1C7okU2Vp+XVjH0zIEa8/EPQs7yFK
galdqeaE51quT4mzW8C6fDVdDXbD2DRuoV5HvfEdP4zZG/1JojDVWsshpkUYmKE9
y1bIycoR09QdmWhnJw21PXRNCrd8KDIAqrseruPlIre6ND9xvx+aopkBHG5QQ7oR
kAOWm9Qg8pRTcH4eu4lQTF9Als7rzwyDN7wmigQ0dpUDF7J2XRJCh7Qi18XA+8Ux
NIe/c+0e4HDCifj5nxbvmDG9Vs0KqF6zC9SKSyW4Fip38n6N7VRpsxEyyTmtlMAA
HJSi7hufWvgZrCAMd76d/zPtEWvg5Jvnmbsxa41nq5Cd9nOF3gsc1SSI+Ckqdu3l
mVMOEuc2EopQHmNS+8dPU78qXP6/1HuqnzEuvzu1IRS5e2ED8LLKWH2btHjA7OCF
SMit8HnIp4fRnq6mYZ9ZU02HW6ApFV5LdQ4I7zpsl+3BIuALu10vPmz1aGVuNiox
xBLr4ajjjIn8kmbcbXkV6tZEick3rLVrW/oOxHDcu3XfdKGRqQ15BBQGIdEYhEQN
vq8gnKWe6q7XSyI+IRp2piVkjqBdkys61YSKc6TaMTfc43yaMETz3k2cjSm3c8rJ
KQHGoYEQouIFVuIniPt7KasU4CFObb9Mli6BhgbFFqoATqdhLAqhbrcYxCwe2rBD
/hsgQcSf7oaIZC29UfMkuC30DqyM9QlA7M7FAK5vlJ4n3GZB5DCd1jqbRIitI5At
gDMYclPoyxkhUphsqKWxpV1swJBqFcydtlyQ+tIpW9GEwpVHRoxv/9eMsHjf65sm
GUt1LjR4ycXIlm5kK+8ld5IzLEa4uRRmLOP4zJ4TcMO2mPd1nNm1qknriq/VsYkq
fxnVbL1xEu9EOkSwBBGsoX/XDiGDB2HNe5+5GmEv9jpLurhh1k56KO4L2lWTk5H4
+ONVyDdNc/xR2qk6LXDfK4wPl5eoqBeRtnPflPumTUBx1P9fN63aGQFlLWUztVVK
F8C22DwLLaHZjWOZYrO6fzHOWnca0mpkKxN+nn5yOf/cTzHiqM2fjFzr+fgx/mwx
rhrknJl8uUhOp+16N2/4m9hG8hSo1l98eQnv13XKt4MTxwy7OnK5eWwE/JSaJUep
6i72FRnI8N2ZBoKJ44endnrUf5TviAslgms9wY19Y/kHpoHuEdWWHERCKXRGCX1u
B02XMTlp2REOxOkhQSK4Kohfr9y6s6ZEtWF4mAAqsfNbpGhUICJAg9/MYbKld/SU
m7Z/c8aXBcFINMOgupvy691MBEl69K5xmWXp90sNA4eflsi8PxVbeUNgUd7Yjy3M
Bj/sLoO9WO86ltk3eGCMZ1XWt21Gz+Ou8LRTx+YOmIEm8/pGogKOBQtPDPVZU+uN
nW3tWL8h9fJ7Tdy2/ylzn85BfI+db8rDImPyEGmsRNKzRbeqNFa26Pyzmw+Vy4Gt
bTde8K3s4NmJmWWHf+Fn8497GvqWIoQ2ZIQfKXqOXG+0mkOKKYtOW+Rb1Q3Lhi2a
Ut8Y3ZHh7n8NzIIZKrdOrmRg8zhYGfIkNc8wqJWNoKZ5fsQA+joC/YI4N9SuCKh2
KqmKoz21s+kslK+iL684sEnxOyjDqtKCVecCsi++s49o6hvXC+hH4lN1ksSTyyle
wD7pZt2TEjjlxDLXPMggHVFvTBBMrriUQQgbi5Mp8R6nIJjYD+SbEclZIZBEbyOc
r5EW3ecQOKex2UJb/Z+fy86aUGKJndSViVQfEDWgKsZtqC0ctxb3V8B4GTkPZqKq
ZUY1C4UQGfhicZwNlBWdCp7qgonXO0g3CSgQHvtBiS6FBteq9oS/8t0lBd6dbly6
eQftu8J7R0tJtpW9ZvI8J4OvBpjKadgvOCYUuLULZU1OmnljUi/93HgMnD0Y69XE
xWUDFOq9rhYPu/jPeo6bdAKvPapfAR4yc/cFGlUM0dZhyZGpeqxw537SAhrVjSNh
Sir2Hz13/0y1W3+YRTRDYJIxfIvGHfi32zTBGBtgQC7RLvPADjN4yBbO6qhorCLz
r6IZ/DvNb5na7scu4mKDO+A8blQdUQGyuf61E0tFAR2DDP7pMm6euS1sAqnW3tvE
02BbztfnfPlDos9rXhFPH5WygydTGkco7QvRqTgJHmeX/ErjcEdubs9cRrrTa5nx
FtZNOZKLCMaGx9QPOoKTlZh7MPfFdPQgprdo3OUsBJdoqmtZyNVVWgRDPYNp6/AZ
PYOqth2BAnP281R0T1NK17Ay3uXvk7ZnhL4hzIWmSpkThi/YYcY/eGREsVPK4GXq
n9cibR93qr2FNwESuzZ2M73Uuzf33AiBmM3VjtbadP8UpitPwYEdcH7pw/s9NQEE
eXiLLtlxApjFVP0bEorL++lAWba0SjZfKJNhFXoBKwOFzj7X7/nVqpUItmmAxIco
jF/UJHW2j9wn5W1ACWQtSYejad2vUAGZ5vRdtr3BCDpj/tLTw0Vi6Wfrz60i/kXk
oH8N06pcWLsbmfrLbAQ5UkKRqf7i01tgjyIxy0WfM1BIc7U5eSHC+lERffKC8FbQ
x+kE9oJDsTVwVbow6chGpBpY5UBwiQr7iTXb+aJPqW5N6NEAIJsuaMvzZnp6vTjr
xtSt7TGAfEzW1OH6TZ9T25AB2mhfFqiWYSag5wQk8DHvHad9sLsJBtSyu/+BYQ6F
aAa+zaQ950Ai+pULQwEQgqHOn8EXz4kTO4uAZ56h7X4oCb5cBqMnUSe2/RFgRLrl
W9uDft/E8lJZJg8pkPU3MluxWfqhZmoIN78IIOSM/TKF5dUXQ9k6vxQjgYvw3Mvd
E2lUjHxLjYGkzaiznL7Mmi2QtSElpJI15xC5Yg1SdwFfenGXuL7kdF38kqCwsUWK
pJp6xwPidUE4Jej3tLM/OA3RCac+Uxt9lPqgeeLqjhTdZVsNYKfzuKKPTJ9ehQ6F
z5h1v8lFDp35S/Pdv82ITwHP8EGxDtnH78Xug2Mz9QYL8XwTIL7HP7IdFzI6jUun
gldeblAtqCi3zdrzqUebnakHxleS1aF1NOrK33LoiHcSX+PP3F4O0WT1mljHGMKm
kKa5zVL/DBrt7vlaBVlZH8P+8OecOIU3ZH2CxHrOmZub5gLGB34cFpNvUa2kQQdg
J3XDh+yGHXQf1sTIiEW4cdgVb91FmnscOzqV9hFdjItDC7shtQHUQYbNZhlO5mD0
waehKSWEp2j7Q0s1/kviMvRN0OGVQG7raE5I9Si2zpK3WKxaa+YkT+5qyE7d6vif
8fXrNDuwMmnydoSQlofRu5BWHSWCwuqs0s2uLc0Uzf+gmZiWxh7juATp0cSsn+Tv
pMHeJrszoNL1V9MP4moAmlyNOm7V7nD+ZBUHhpCD0wnMirILydWqAcri/x8QVmry
Quj/rsSkbrqfHguA+mWhEjtetgL0bdcweWKXWccdsUSuEK0gYuyMGWUOunEh2Pj9
FMxESOqMQrCFW0lrTeHCTQsW/QitGzagTQrvSjnfOzLkvCEcJ7SsV/8IX1vecesn
IAjdIp/ok+GNrJPPq4rAqF8AsMmugG0IdE4T7pWtUhQR0GCInnHHi/zkkD0lsag0
B1LTrFYfXvOzhK4TOMa1m3BPEAVU6eO724IyjS3pFmow+sro1muUsh15b3esoEIw
TKRE71Gohfzre4tsU3qVp8Svj+aC3nYPhfpGZ/rJhZwrS4ecrBWeiWC1YA56fPrx
nGnS7S2a0J0ULV0Lf7IXawWoGeH3lhQf2krbdxFs1WAY490vZjVVNWiuKVlj7ERO
xoEgU8KQZaQbJvg0+GNB/NDP5MFKnO+xuiJ+eWkM+k/DeObsFqqMqNgqyM1bKLpO
gtA+xU46Jj44aBxAdpwpemXzQO0u5tzNK3orOi5bD0Fdtbozt5iT4LjUSQXq/RMF
h1Whb6hW20KOIBpRIIZY6BViUhdmtSRvxLF2asVxQ2yGsyaRqXMAYkyblHV+f75I
V422LFIjMJSIKaMw9cvb/Fu4UPmvyeyTqLxmkHj7oLfenHsqHzrGqQrKxyRQspK7
IlJC0mpm6p/OsH+Yz5qRxdT2/nCvuDoZYGsPa0uezDe0vWXd70DjgN8EaVipLIHE
BUqsz6xo+qlHsFuyfpLenAfDZ3rQHAawjDpY3w0uL7pnf7rbOS8XPl2WY1aZ4HkW
1QKnPCnwrCYFMhTGniSaiIo6D/2knxUC200P6rfybX1gNZix5Kh+lMu9YkJgVeyZ
pHgJqJ5y7s3rf+T8o7NmpvXX8lfeUsQTFntgQTd7UV0bIpBOFfHxjfd8CqA+9t6Q
YdscwOPh+4EDxZek8FQe8P4+CX6xHRvGqVgll7LRA4fwF8xn7V6ylz/FfvhaI2WP
kTbNTxXM/TxcoDr/seS2oUJpnvaqEXzN/pGovKyVKHYUqmv1o0fIzLvThrN1QFN4
CafAhnWjL/l6lGrjArpH0ezC4XgpJlhGCnVJkoZsRZW+G4jrZGPyfFhsIJFxglF9
848A28mdXles0ATgjpYqp4X0P+Q9wteFBb2+FG6Dxoc3aJ6rbEo4LsQtWB4slGQF
PVYtDz6gwT1Lj4ufaPwJqZEkIfzJrtQa4vdS/NHvzmpWQilqikoZZwRLwVr9ZucY
NUx7Grr/OUrdsJwbTInaeEPnOB6zWmJVo7ZsxPwjIaPr2ItkyfqWUnmIY4EUBS2F
yTEnDRGImlDoG9he93SYlpA5IUCBD+I0JCAcmcZnUYZatTrE6KrE350CcWa9oqxO
xHW4FG79JHX75TQytq883U91GjfSO2lwD3hbhjVBdVAI2aTNoSsI+DD9LIGKjtIh
4TIDr3LxYqFAz3gU2+mAXfNKwiKO59B3xZWxY8PZDKt8ETaotYfEogqEw5Ctj/Yn
/sIPknpoLTK3Rh/LNjRkNpFVWMttqRobHNg4Buv/HrH9VfG/IKfFqG23pwHF2ux9
pG0XMruqffej0WRvmyKoe7NHbKaDgWlDa3f8oHl45o6ExQ/FiSHETPLteWMLKAlj
M+A3f/YzDV9DUfI0s5YRKbX3xtMWi54zZJuqTrPjHOTzn4ZVVu6vtWsB/66OhHWq
wyINpB8wilCPcgaRsvabRQg9XILYRMyVhM151ue1y8Xikh2kpaEbjgeMuH4uBr8j
9xudVO/G/ixTcoYl3Ae2kqsMnqRFExYxngxJ0hkXp7+AzFwG7ZuFWTmZpcS6BFwr
we7ybT4zs07gZrCkNmyo5hH+XspWZ7MXsJQPNHdZDGsbwJykYiajnofjmW7MJI07
TwmrEI28j83gCY78uD1jyAZVIe8YZAKyW7adBroBaz72LEMLJ3IckGl0jNJ3BzW0
M3iSUIAmS9nTmv4/h9g4StMJaJORF2sGEW82veFx+F45ULZiceWCPDUOBe7n3jBB
3Kv04i70MnI4EIg/B2b8A7YBXivEBWeIyNaMOATsBCYDmzc6OM5RHevFVAxUanv4
CS/j03boGFfQCGbPU2xV1Vs0ktl53sRjcfPOi6PlWdJYnPaB65+Ls99fahiCct7k
MZjkJ7HNCnlTUrkAbR716iUiZmmFpJU0RqBiGpVB6IpCtZ8V22uk3B2spVi8A+PC
2YpFNJlhOitz5EmYOs93xxdaGT4i4SsulFJnUIvOqdJloH5lwr8DaHzYRhkc9MSl
qrwEjUuVDcyk4ZnbPf1t4WvU8FWrxq+iEWb9BluKCkqLHbUjnuDgHsPh5ARTS52b
UHeMLrPVp36gB9u7MPeGY6pbaKI58RJJqqnfxjDVWAVRrntQOSeGZmzeiSqel6tt
3iuODyP6yt7LFuIGRfsNMog1ul8xw+2bl39ZcUXFNzjZJR2DLWqD3MdmsXj+y6nY
TFadRJIZ97rFIJhA8e/M0PnPoa3oPwDB6I/It9fFUJb3GFBViAQqD51E8WmnZm3d
8ylPbqEq6C32vcyn8z24doWzAZagto+D/PKqm5TLrPjRliQycscTkZpdPPO3+s9k
bZloaKxSEqwKga03fASWr1YW9KTX7xbgVH0SjO354vazmtYIX/6xVJL9IkfSlDe+
J8GUGuugLNs/WiAK6wX3dyXIPMAmCuhYTV9Tz1ifwEY8cCbbVKbOx/SltgLtVMnT
OsauUoa5wzz1ETDrms4Yhhq76D0+gHGFrnp1YaeuhPHjodox4yjNl1dJ0YXzmKxj
o6i5sQtqhUGBXHGRf+eWEDfF8bwNHKhvSFl9ZUxNbYDFPUye1REssweqLH+ap+lU
rwhV5ASY+5Gs6WAIynuPoN6J+lW8iCwRvjINwHp3Z7iUsYBrwPdTCRQWmB6tPEua
kpHz0MjeGeSRaMy15W7PFO8bzFgSO0w9R2ihoIhxAng2K3LvRAZ0UKdqWlm092tH
9QncLfWg4GJzK+vg0g0lZz4DICj+Sket4/EW9l54wrtnzxH0eNUVMcu9nf76nY5b
UW3XYEO9sntW2sDbj8aCp1ewLxicZjkI4V6T2+K8U9cB8yaaCrr3bHQUGjCDZ4+A
gxuvlqlbQxltp0/lTIUIHrN01J9kZKdYBVSHXR0dSPEoyNfBHS4YgllcFu0XnXzx
VrzvZe676P8Ok24om8Z9c/CPxAVdBoAQl72iAPMoPmsrci5d5+WDwxR2ajXMVDfI
CmFGmkb4WZaZ9R4jIrxr+PmjdxkTgGJ//ufH8aC09mmjGQ0mD0ZkOcrRKDxmByrF
ynFVuPdZrS/iK1QVslinbnphxr9/c13/5i1Qsc5ftNUcBBOaxndVhuHA0uDkCOqv
/6R15l/opeHYu3UYFFP9b3JokwIuXXvWl11mEIGbsC/sDxqEUTVwps2Wf+2BFaDV
JWi3Iy/9TODyzfjj1DD/gBsHe8FEZuZ6Ggv7DTLZn5Jirp4hkXhoMem+lqx9BrR/
5knfzVt1oGIeenmGuvEg+Z6Xnse13cXxQdiO+6J8iL6VM3IcOGzo4Xbdj9kkHGTo
WGK3d4kk25K7zUaS2GqaYazTGyXuGSYTG7OnnD+yvwaYsHaIVXy/nZ0ot7bLna7p
m+fLAXFku/7z+lejNAXJJM2+n+HBMdK65eeItrPDOL2P6LAjWtrFQgXcmiI1Txzd
fIA/tSDTdkVWCH/nAkh+ZL8Yn8JsjiEgQZnTH4TldsQ2BidXXxMQ3sIMPebh3/PL
xd7ejOUntVZ/H9xi8Q9tOiYTCdra9ajYfWIdULjtzCiK6UyYv9BtKIckX1HuQ0GR
NWnM2jJV4Ri0xTVSuEeSVM2hAGo0wIBjd4Izy+6f+FAQliXmtQfQ/3yHWQwuILva
P90WUdAJlaiAd/HBCED9dCmI6ZcRE5Eztc21yZxWUuMW2iIVtzLRT7gL010ioGnK
NxfpAulGEOeFpCCjgrVnjbvtbHM82NiqKiPsN17SetrcFfhOksCAT1abUXwoSozp
1uMLV3ILu/ePTNLaCfwB9pCXfWL1q9FO1UPoyQlu2Zq7fULlKfeLlQGiQiUObP6z
HNzd/kaoIaUIFnxMxUSWgnjPOoKCeb2pSDoACVH3o70BRM2s7gidXWOJvOzGPaWD
BKqMVR2HJ/gjtgjmIeuwqlPrW4vrh+89FrtxhsQAxiItSJK7+ShJscEM/Afs4RE6
5sHRn+pitNgEyM1VSnxyQyOjg5F0OXjTJfRt+pA1EKweXUrdSkswnlUUlVILJsl2
GTT7uGJfeZMc4d58qd4y4BkyIn3LpY6v8B0KryAC25/j8DzyJfuZye2xF8DiPTHw
75pRgipnY/dMd/TYq1oqvrklmraAYppK+sz9vGCWHzlh+O51lOgSQkxaZsx6JrUI
FVQWQoXCuOi+ldugrVpSOl3cHH2X9+2LyuBTnbgs5rtT6aBEzPzRymAYfftWfLXS
g+YBzNJ+hgtY32hXZ7E0hZcWN54JrnUZY5iL2Um/sLZZHEoMXhWOKsz+3oDRVTGA
5TNiAEHTu/cL7WPG+MfA+050qvqYZ/Z0iz+9+leC9djC70WTsdAiOxkw8aNw6mHl
TF6/qqffDMhqhcCPkQ4VRWOdnKR0NtaV1PW6VnBSuRXRyQ3Fj9F6ldd9/EiWEKVl
h8lv/6AtY+FyuAnfA0jF84W+/xAd41GdP2IBErDDfcb8FQRNxTUVfYxNtNNvDbIM
kRvzhyo1VKWjBL0dhcpsn0j7sSegSEOdIEoP8LpsC/71kjA+4AlWQXydrHrf2MAk
Qtt3SF94gxngz4Da+qSk2nvxZ7MpRffon4P1MoRDXw8NRTdvfDFYDJJtrUtYwT03
XmJDeXOH6eS4gduuzmgt1XxB8rxAksZVssww6k+qH9OA87QsyqdI4BI1NIZlBxpr
1B6ysleV+m2z4imFRXazDbzuX9qqtI5ncddRBwASX4PQYCwE+6z+kuayuRL5e5fH
MorPafBsEnvGgtmtmRofbdsh3R4mo0NI1RrkkLAHBzw+xASOat0HSLrrNfBvPfob
ta1CjCwV4LDCZo0jN3SasLFRYDEa2NG2j+j3YNvm2akvAGcmndfLiwNis9tJO12U
VcARIZU2IgZx5QNbjpsYjlXJKj9WHSHX2xTfXxzRKPcwnVcTIOzSAoXsUiIqQpyd
5ZTNEw6SaIPa2rHuAlb6/vyozcDJLVdVdunUpU5VFC2VC08+8wWZqemrUwxUF5BS
MlVQB+bXI3LgdsdaayYaeQ48l+qZIt7X6FOCoMDogpzsUrgMF6y+38EbxESpbktS
dJrN7+jhz3YFzxGkomtmj0joUNtXJUN1QVz1MO25lcTeqS7WaCWuCce+w8ia5wRM
gAeJ8GGdYAJ6UwqxTLS8JoB3ga6P1+QmcdyF0SnyHbGTE9OT8nycWc3dqsfjd7SV
NbNXzoasYaUKoY/O/xtNAApg/VjH7GWrKUEEHLI4V9GP8XmMMPVJt1y1wv7+h/ch
dz2rw/HMoLLXQwT1H2L2PUj/l39soL9xz1jqvbuG+1vTOU+rt+0/HqoQ5S0x3lNE
uKQFQPupr3S7Dm8tg4yPL7WLIjhqO+qFnKUBku6mNHNLTcsNiOglzHykzSPc/126
UL56MWwnMxnWzrCBdCTIfoHRRU9vFm4O000kSazxYvidJXcmG1sT3wmaYGMu8GXu
ldWbTLW/sV2z06SKp33BLeXKcehGVrJuIqaDNEPif3omQw2GGGFV3TBGIHx0MeuV
RdBOt6yRgpcu8O75CFeMMbYk8wRvcQ7pjyfmdYE0ehKenatfC4PwHQzKhwtl9ag8
aJYGI5xVIe4O+YFj3mF9zadKQp64Z/X89IUfIOro/FPAI4LYx/5ydzIMa2IUFDjU
DOGLxzNOocCIgySrRdAhqIkIfXKDA1CvHumUW1kpB4UnqrJQlT+gzanJ51txQQzi
RYaE+TmMe1nqEOrvYUIe4S6nX9lshJ8D8sbAhyXovCwEv6VcVbuARRv+VKswjJPu
19cCA3oO+8Z6DKbwpfFI8cNsuCs2eym/8756CIkecNWOsNS/WwUWiRHZTch1UnGm
wv8N/9g3DHkjLZrebGk01+RtHh0nr+zyC1IJrGBwWxQJyIe3lnh6XGc2L5FCGPVG
C47ebKQ9DG13iR/aF0yRGaXUdOKx1jhd/i43dPNFoaqKIGiNZy3lqaYhwB5hjQ5s
SsYqw/+8tf106Ye+CbuJyRp0uRN1AG6V3zwdQiBy3uZrpSXvgkbb7WnzjWsJamM8
4DM6BR0WjR9cujPntGTLnqXI5259CfLzFUJ4YqL9jsWeUHOlEjf6u+jgEDP66sJV
mNJY0J8qJ7U8A4GG4ZtWmIHFwCK5WHFjjv/lkPjd9wuCssICalo/d+FruwBqUcIs
kVgFNIsJUbxEpJnt/d6JLvY8IjMEX6NmIDhSEldXal2f/XEkFopMDjPnZPHWI4bm
lXT/K9l6C7iCxk21QguVe0YZZsJ+cYeLcsE43aOQ7uL6xzGlQoFQQ87vzdqEgzlS
aIv+04qk4pZU4Z+GzdQVvBQZ15F4XdD1VBQNf8u5sTRqFI2YntY/SLuL60yqM4+H
BVeD6iGh185qJlYKjJNUIovdikcTXoW7JsJqnGVwhFcOIqfQy5wY3I6F7Y/eOGk9
oRWvKdD8q3TqH0fYw1N3gMDZuMcvL5bdyYOBD9mutAaTd4b/5MV/JR49QRKjgUrI
dXGLSLwP7tNc3yyDwYjQUZ3hdNcaolNBeThXyioO82YwnX0GFKgAKrbaWC8zn3/e
0pMvPylSJg5aTDwtFhLvvz+ibyytCul9t7EmNlS4VuZFy4ASnTQW6iHgNsUVfinl
AlUs87bL2WqYqTfjTA8TbACz35SoBTrh3a1yFeXF47xV2qwOl2L458UxZCuFE6aR
ZhqS+W/gUphca2W0SQyUbhB9sAsYFN68+KpTlDL0r4OvkTtNp42MTVxL0gskcGvS
5N1luftXl8KGb3XoxGKs07y0ygXah6sgcLBG34DJGNzQeh5Je4xlxH30535V0FBY
rsUjJikGpzjD0AattWtNyYasQVW4r97KzwZl9R0upboSzBaDBLpEGBr+OTOfbi1x
wzbsLlA4akJ2sS1oJjMdF095n647X0rUZBhAqWJE0aboDUn/RbbHAhqsSxqQ7Aa3
qSDvbR9oCJb8yZyQnsK0Wpy+i9B/85bbpi8rfRa9z+zEf3zlfp7gFvayznWFXEYV
KtPtxC3Ol6znOV/lVPhhJaYYDe6qTfrkcfxCgd1XQBcnbeSAOSp5+AI65IBjmSx3
+5Xn6wdjcaNnP48Sr1dTbsAuGQD+2UIEZ9O1jy18uDT1dX/g2YDrz9ViyU5gKV9n
ZKjTWTjL5OxuysIpGYk5Ym/HBFE79OX7SQGEBQJbGywdNC1F4ztl3Ehue/rnUtpy
XDWfhHw5/qatazAtfoDeeWXaSTsZ2xgT/GrW85bNjwp9IjEovMDmDS0iEBxZLoc+
TeB3tRfgpNkAnwROXwg47VY9Se1WxlvcwkPQhWf3DWLqCzdOsumr0rl7alRejIjj
ZG/FVgagYswkXyp90MF6QESilK1ol30t1cj8iQYLP3d1KdyUpKAXamV3g11orGle
K43BdheUjLmEssT/NqI5Ibopj0AI65kn9H3ngARhoXkxXdDwZ7OinuUk2kieVOc2
xEwbCthLpXMB46B1lZfc7nsnsIpTm66VKrC9To36BfT9nZHFCIBrp+1M9BlebE/5
Cy5VpT8Mj+i2ouqUMi1VbwMu41LuvWXQX/xHLC5nCn5lf84fWwXRaObXHYTk7C4s
HNBTTJ6ED83W6JyqWl4z3fp0jM06+i2Cv0snQ7OckItp6NPVpGIyLai5CaOqRdOo
7ryyKwgLCkw5w5G9EDq/5pQxUD4NG4ue6CP8yw+XAuU=
`protect end_protected
