��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���J�l����9C���%[@ ���vK�G%H5��ۙB3aԯ�g�!�
�:��JN�>k� t3�[r|������D�����P����gbY:��6��57aj8������!�	2{�/�x0X��C�p�=왒$:{�wF�i�^�@!$Z�I�|"���<.*�� �<4B}��n�)!��aLb���nj�������cd='^�^�1������.�D�K������h0�leKܡi��#j�~�g��nzJo�i�����^�"�/���Y���5H;���{�:du�2�{��ż2
R`$9�1O�g�~�2�T���a?���8�W!ɻ�1sq��^���J�ܺ L��r�����^p�R�h���S���g���#r��l�<wp;�hݼ/d�,{l�u�,�l�JT��R4-«��Ӳ�'�պ����`��f�����[�?a�+�0�C*��a,+2��Yd�Y��|�l7�L.ߺB��+cO�0-A�r��f!fXQ|X�P����#��0�K����\��]�A����B�}��J���ln��(�� �N�a�I� ^5(��+������斁!��9��z��ؘ��$>AR���,Wt���oK�O����-�A2��j��̦��O�ؔ�7q��*�+M���zjU�|z�T����} `��H�MN�����Xb-@ѽ��O��N�7�09���Q�F�voɻ�P�ar�KIڠ+/�K�	��D(NQr�܇��쳍��1�̜�O�q[̨z�J��� ����]H���d��3�!wil},^y����L6l��f�ڥ��_���wQ��a��%�h��5tT*=��V��@mt�َ�Ƭp����������s�d-�����0����A�I&F�Y�q��P:�?������@�Q�r�}u�Nu��&����z��)�M�o����0ws&�}n鑲j~��@�d�}��/'���A��E�z���Z�%�gs��Y���s�䳴�O�o}�����Pt��q��2z�P�[u98�6�`���W�^�<�O�?�r5UXjXb��QPj��Ѿ5e�F��ۤ���}�1�'�%Q+Lx��*�i?��&�����Ӳ�B\�����1��t��X>����V+�g�~;�����n�,
,�����V>���4�0�q>�W�9,��|��M͜��f�
S3G��1:��z�u�hI�)S�mDDk�w]�m�.f�$��'c��r:?�=7{�w#E�D��OI\׍pwO�΁�V����-qE������?�=��VX�I�xfͭ�ۀ�p��:��������m���v��kЀ�T��~Xɓd�U�) 2�U�g�]@5΀���)�T���
*�c7��"��4�a7���!O�4=2�.�g����A9|t5uߤJ-��Z�B��<�}eAw�R�^i�xAj����k��6�yc���ˀ�v�T�{Q
|�9�*��~���>��X��|�5?�ӥxv7�&�n�%+-��/�p�|�!������o��J+h���1���*Ź���QL��(Ġ��(�ĳQ�e�˃T�/ڴ^�;CU!�#d�8*g����,^�u�"CwR}B���ϴ�@�%~�%:�8��!j�!O:���*���b؀��,��=�`��mE���B:Rl��C���h���ʥv�f����:x���C�]T#���1�ʡ�1L8h1�D
	�򸐤��g�4S�^�Ü�;�\P�0�"t(��s���K� j�yI3�!.�e����`&+����]�]T�%��Fi5�x.�h�I���j|�~��a��t'��\(m�ƌ� ����:c�ػP�4��򍂞,��/d�S��8A����%"�0k�^b���+en��=~��q���7Sq�F�z<����M)��h+Y����3 O���G�gu��m��U̠�5��]#技��F��)ΑV6�:gaY��'��Rz����ty�m����s�s��̾g�`p`�.K��,��^L�kP[�w�Ng�l����6/r�K�>�ѵM�8#�!�� �|B��ږ����6�Q����Gj&��{�G�s���*����� �10�����q��w�Oc��wU:�C���Jިiew���S޿9����Uf���	,!Kjq�O��n S_�H�����Z���eW��(lP�>�a^��f��a?��Ǹ>(b���+�u�	��*>zyb���Kd/���`�w�7�C�!&�'(&I�ۨ���1T�f�4vֿ`�|������|CJ����Gk
��>^(y�� �C�&�(�El�v�2�t«��'r�u^�[�@���?h��^��s1����*��5w�2��	��ә\�E%s��D��_ϋ`�TM���׈f_թ�M����7G���clm�;K&�BVL����hU.I`,�*�7U=3�az��F@rm�(�r�_�|$gp�jK@�e��b��j���ܤʬ�)�T��,4��*i�x��q���1_�P���� �}���3[e(�5����{�m�� ��)y��s���&���N��A��P 8o��;B �;sB
�Y�91��z7���*NF��f_��/Ћ�.Kp�F��ow�YR���XJ��v�߂L����?�X��]��N&��ct�$a�.<n��r%�L6�'�\���\c�?p��tȅ���c��֍�^�.��QU�$#,���AK���䠆����3Z�[ȃ\{�;46��n�e����ݒ�RI�G�ʳdp
�;;͹��^����$E��J�R3y��t^���u.{���T{�,g^��!��� Jfm�O�y��%e�V���	d2�����Ǔ@��>%y�?Sp�\d�O�S���͛&�Yɑ&���:�&`����GX����G��L%�6��6l4��E���\$�����2�%��wǯ���3�Ym&&etY.�?�S�����gv4i<8Z*9��1��<��q��Aт��NK�B��K3:3!�e�*�骚r��o��m���!nn�;�ݻ�P�ڑ�9nq�l'_����r�ӌh%5���x��W]h��u�w�Ç�"���X,9�+S�6
�ʪ����p���8�	G�����A�`x�?���
��xaD۵��n���Ld��E�~�p�:����44+��-�Ͽ^�˶�- ��k���䉻��������є����g1���V����f����q�}p�GWZg�l!����o�� *L���F�*e�|)������P�����fe�Ll)���#|�˖�Oʚy�q)�����a��p���'�:u��Z ����V>����K�ֲ�o��<�ո;P�&�H蔆a�zV4Z(��j��V�i����z��~*��yX�ٙ�}���Y�|/����#�w���o���n-�o�A�p�ZyeOG��;V���C��b�pQ�Ub��qT�JRE/��r��*��ؿ�1�܄��^������(�|���N>����"A̸�p�~�������2�[N��07���7�>�~H(&<%�XYO���0�/�r>�=�G~���*�Ƙ����L1뻚��a�;0���S�}=����� ����~?�އ�m�H��#��|�I��P������+RS��6`�h�K�BR^<��b�����Zs(�m@�?;^
c�fg�F�n�6�֨���vĢ��O�xDt�X��@Z*W���*�A�9���u)I� �N�}��	1=_�Tҽݜ�}��R$�/ۺc�Z�䕅s,ME���h?��:�9Lfۍ�1���׽0Vj�RAYP��%�vP��<����=^�t�Nĕ;���M�s�Zބ�u&����g�T@�p%>��a�5i�5�x��dL���V���8H�Ii.Ԃ"C�SM�F��᪚�)I��A��hU���k���0K�iO}��-��i��?wq��v3#e�������+��ˠ@�|$#�#:L�$؍x/*�%[����y��(��A���.(���I�1��h2^�d��*ފuL3S��w�,f@�.�lV�5p\��]���Y
��߷�����j�u�
�P�b��eJ�bb���]SA�kp_h�B��_�4�M��\�P�/Ɇ�d��D /}2X0��w�#o�j_{��)0l�9$z�����װK��ИZTfha@����b�Tɕ�(LQ�S�4C��
I�kg��!G����be�c���Ͳ��� =��s��{ڋ�WW�`��BX�zc#Zb��o�1�k��9UB`���/��!s�ͤI��1,7Bw)Y��Q͟\��}�}���lh�>��_cW#�qwL��*uGjCN	��_c[y�M����\0�u��H��$܏i]yD�g�&boA�N�o��")���]�wd��-2Kvu�p)E���LTJ��E����qD�W�.$�xeރ��ƒ��	$�2h�ǔ4�7pW\uZF��w�\1��ލ���,{á��1���Q6n*�4)�߻sB��(���ļ�|���ք�G#���'�B�~*1U�c^�U�W���a�!D!� �(����!W���3�D�ŊH�zAyS5�!ܜ�%�>�J�K���|���R�������C�OQ�&.;�_޴ 	��X0tr�⵨.�c����6�:ܭ�x�l��xR�ڍ�I�^�s�nF��+��Q����r6��L��KU'�����}�>y�@�긾��|�T�q���ep9S�T������{4���AJ1qgdF�cFw�4B0��{�v:W��)jҐ��= M���Vu��b[�ʸ�7��w����2LUc�m|�j�9��U��ťZ�,���h8UzӦ�T��Y�Tf���yA�?���́�F3����=Qhp��HNQ���3��[��ϬL��G2�
��)��B�`����+���W(�bq��,�Om*@�C#���_�k8�����0Ű��x����ú�_دW�;Z'c��8�Qs��K�#�oW+�[y��vh:�t.�Q���O@�6���!� �_�(�ٔ�;e� �55|��E����I���@�ܷK�G�+צ�d���3ʃE�L���/��8�ԃ�ꜬZf\
�'����-��],\qz�	�UÍ�����79B���8"1K䎡��W)�vmo�V뼆{�]�O�oY0uW�Wf��T�𫜓]=)RY��n��bAZ5
a�	�j�1bVC���C�o,6t6�[t��'��yӋi�����>��<��d[�@���=0j�L|�g5��Ӣ�:5LуE�T�8�x��(�J:2�h�������zܽhC����8�2��~�k�X�ֵ�p�\L�jd\#�v�P�@Kmip�!!he#˽e윲��(��'P8(�Ń����e�� ���S�O�q�f\^{i�w2tArdh��Y���^5 ��'�sb���)"v��a�?bg����
f慘�?��d'�ϩϚ����S���4��`��f���_͎����ӻ���r���T�]�{�ä�É��J2�Hc�4��;}��
���nJ�І�7�=5�n�+74��,z�UgD��Q�!K��u��nU�ĸ��査}�$^?�k�Ū����1ޡ&�̊�Rm븝U�B�䏸cܓ�Q_���!��d�Aj-h@���Bi�7c��
� EĿq*� �LX'�x$�������e�(���B�N�C8u2��v>1K���LQ���j�4����[p���r^O����� �ٯ$Um�� ���5��C�m�:����K���=^ʷ�����ىۣ^tܷY��.f�Hd�����ʁ�����=�j Jg�561����"��/f�W�'K�E��Y!�T�\��Š�<^B�^�I��Xb.\W��6o���j�E��+�/ۊ�y.�@�xj���.��_�WHW����c�6������{DG��M"�1�����w���R�&��Ř�WԗB����-���[�EB+ ����_�>D��~��G&��%��xT��U��{CW6�O�k&��;�p�[1uIp��zg}o����{�{��W�Ԣ�4�i��n�J�D>� *�����kp��NZ)����s���Tػf�<��*˕��p_ۚmeu�>�j,���u� �q*��Ҏ���n&��T�1��t�acHd=	"��\�28�ߡn'��@pJ���ی�S�rҦ�L�2�I6��j��ޟJ*D�=x��~Ay; !:�x��(�.��g��;g�i�m��@G�����.�j���GGa�%a��*L:}���q�s!HJT@X��<N�׋��i+11P�6]�����X�C�ey=�ӨZ��}t}�
�|Ӊdf��`��ٕ0[��c��	�C��M"�Y��M-HP\�?s�0`6	���;`����.@���&��I�'KG��&��������:a�}2�����p��.��Ϟϑ��_x)/�^C�<dĵ��J*J�:8������ H�'@�鋝��w��J�	d�g](Al��2�H(�lG ���P��x�����)�(úW��� iг�|Id�������in������U��]n�#����;����4ɊT])�QMN��e�}�^ �"��c����A��������R�gl���LV4ͬ4)/�<uRG�x@�hVJ6U2��IM��:��U��z1w�Wp	ު�"��Π�\ӕ�M(&O���}����j�D�C-�!�����/�(�r���:���;�Wu?��1E�#uz��z���Í�ė��f���]n�o-�K�-��<����,mp�$/O��e㏃�^̩�᪄1KPRY��1:��N Ze#;���NP<�"�4��̒�.�\Z�w_��Fvn�8�7�r��@b��x�Pu9uw��[���`�@�Yd;�?�k��_�+�7HU%U�z)@�~��_oz�:�L�6��37��%�Hk����5����C�z� ��s�[���7\%\rek�# Z�JZ>H��&+�+ys��+����+�Z`���t�{��*�Cj�;ά�iL^�xR���IY%'Z\�彌�
b�%�4W����:x���z�^��|߾�/8�<.���(D�'��O��r�f�q�bq������
}5��3�%�ȴt��0%N���d��<�p?3D��i��T4ishj��o債8F���5C���J�]h��~ئnGz�dQ��G~�Մ�Z�3x��Qf������1j A֣E�o����-?n���Mb�K`;�7�����3�f|�H}H9���E�o��`Ǣ� n^Q�<֥����(?������ƃ�*؝��~L2����cEn�����P��&#�t�r��e3 �5���76G����u�nܑ��
zQC��j���z�7Ebg�G\]���3����=�^s~�"��G �kf�C��/�����1�P�ġ�J��K'6=���i�KcŬ�Nŏ8<�`���f����F���b�X]�k�jVP�a1A��"�+�R}��/[w��r��N�g�����`9�F���Γ3�ܸKe�-k���x͠�1�7:R^	�����b�Wh�N��ᔦ@-�?s�x{#���P{����������iLe�/t3@�=ok&��m�?#k/x/��x�uP���������:��"����Um,�s�qv,8���՝{�%g���Å;�	e�� p��#��ͩ�o�ʣ/�����6�(<]a��]4�y��V�X�I��u	�0+s�)V/��A�.^/�G��d��ޅ��(�2#e8�:�+*/Y?�G/�ߍ�<n�!��pt�{(�o{'�������?��j��D�����!X�������=�uOZf����	\KQ��;%�*+]f8�@z�>*�rS4x�')Z���2V�:��_��c��2OƓ��R�~�#ȡM��MnS�9�.��^�� �O�BV=�<��k'�J���g�q0��"
p�Qgp~��w�!d!�c�z��2ܴ2őx�~X�'|�R��O
z�*T��v��T�m�S����BͭcT���9|/��B��+.�]m�;���H*��fB�2��k�)�
��~�k��*ü��,篔�"\ogY�U^����û�N �ek��;e�D�������,?`��ca��O5ײ X:P��3�c�w�g(����L� �X q⠦J�Ĳ/t<ePL;G��B�!E�U��'�#�n�}�_Q]M���E�0��-���T�x�G5z���y?�L�N�xf�g��Ȍ�#�+r���,I!ʮ�Yn��T Ma���bUg� 8�@����b�7;i���:d:]�g)_�Z!�CfXE�8�c��<Ԗ5ye�Te��H[�	�n�A�r�28������
�)�c8GH	j!��wS̅��ˡ�O ճwpAj����Ws���,��	�vS$G�Z(a�-`�}N�[���&m�,����V�P�~Jp	`t�m�pc�=��%�	�Ҏ�/��<U:��,u���L
�W��!tq������T~�Tw�cϦ	@��vttb2%�B�/VL�1J���[?�3�/�r��`�,.H?�p��n��c��?iő߬z8��7�@�9���͆S���H)y{�t��]b��2W�Bz�,�g�IZ��)mǬ� 4I*��h%nB����� �2f���V�������]ƿG��p��O_}�~F��
 "]�>ψ���c��;�Im�C�˘�����_K�(�ZJ"���5%�{�B{�FX�:fT�S$�����!�燿�Z������I"Aގټ(�K��)"�G����r�R�4�w�(V1*`_ƞ��9UX��Q�Q[���樵鬸���9�~���D�ʤ��c�쭠3faz����R11^(&z��9�u�����x����7�x�g?a��1P'M���Ig�����:8�S̯u.�A�[�}z9+� Z�k�E)e�Y�t�����s{��\�
�v�~���%��$C�_in�ʭV}`�����7խ�_c�&c�s�E�]lŶـ�$X��v�����1�� ���,z��J��%#�D��)�I>],�\G��#�A�D��+���>�4�s8�{�{�l	�p99�t��U�1���I,�]����q)�4kR�|��Դ@�m���֘]��<�p�_��CHw��Ɯ-X9��K
���j�`vH�í�!�}4Y^��ib4c�8�c8_(�'䈂}�=��W'[F���eG�AS�x�:P]�Sb���[�l��ù"/�J"޼,�L��!9$��֥�]��!����B-�};)S�L���VY2Hu7U�n����G���{d[��/�K�2���R}M��VDהɺ�/_A�@=5�����(^��O�-SWYvMx�!r��Z�CԢ�ᙵ.i�Z�*��V�5"���#��XZi���*mf��	�A�l��k���9�����$SL����r�_����<\�|�}�󰑝��S��Ofލ��u��1�t5���#
�i��x���$
0ڀz�J��*��K�<P�J���Z���!��x�T;��7㐌��aY��꾃����.b-���H�f���!�4þ�Ԁ�iy����(�Om���`FCyL��7�(��ǚ���~ �I����'}��ΣB��Z���p<�Z-��"��M�ݗ�޼6��W̨q�r^�d�S9�i��ѠS~����茼�5�h�!3����5[�&Bu@�Ҽ�(�iz�4����N ���)��;$\������`�I��ӫ��S�x޺��d���t��9��)U\��Kߧ�i��/7��u�=^[sfa9���߼��cQ��ϙ*u=��{|yS�,s���A����7�g�+��3�H]�m.<����Q11��B�K�_��vZ��H�a�&q<��z��Q⒃玕D�Xӈ ���y/��B�5#�_���ʌ��蠳�n>
|M�?w(OH
�x�,g�S��Ȣq?�������=f�WàK�UJ�³o��J���˜P~��Ѹ�Gg�D�E��I�{U����9��cf|�X��V*�v�
��<KY|a#�L��H�-�3(��e�uS�a�l�V��� ��C?���7��iO�����Z���PS4(I��C9�-	4V��`HS�V;�]ʑ�]��B� ����T�.�����x�	�ɣC[X�)-k�fËQ�n���B����ߕ��?{*ܫZ����]Es③�ž�����j��]YF'�h��
�'΃%{7�ߎ���W<np�ص�p.��k5 ��x�:��*���.͎����� (���'���n�,j	�Z�u�2TV�i�x��(���%��x�X�#fN&�%�����i�����6t#t���ŗ7wa1����8�|#
~���.��߽;����.l@��:��j�`���`����i�@S.������Η�>��8?C�q�� � �ũ	�@��\��H�V '!h�4�R �4qϑ�� �	�R~�P��޽�Rxo�H���k��}4>ㅏL��kV�l[�7χ)��m�$l9c�#����Z��:��N��r�ҩ�t���&��v=��#5,J��sC��gF��>a����v`���l|@v��AiHf�a�nOp,WT'�D��Yfy_�4�WXj�	�W�@���*�Ӿ���"����%t��Z�x�C �`~����G�tX=uv�N��f} �����b޿�TYgʦ�C��n� 4��f%:�_C�>���Y��LQ� =��MM�Sl�p&E�j�X�:8����ƈ.��Yè�i[k�C%\D,�n�A&ntw�:�-Y
p�7�_�;�;�?U��N9ο;�p�S��*�dQPq�B���_r��|��l��YMf��&Ѵ��� �!�zV�h~�^Q����6�KU_%��ś<#d9_����ݕ���j�8 �<��`�������Jf`�R� �E3�|?�v������\����Ԕ�\��{
��k߰=��aV�p�xz��T��kR� ��i�+
�C��H(��E���(�6;�dh*;�&�9���+mg-����A�i�&�*��
���53D��{ʃ̍z�x�[��F�����)̟��7�?DH3iF(�*��h<�NZb׳�A<E �4gb���k����[m�,Lj��ܙ9�1l;�J޾�NH�4��y5�qIC���V��26�������qRD��qZ�Bᥭ�r��A�G�B�,�%]�hc�m��Ҹ�\��z�GN#�M�o�O#��X
V{��(��:�,��T�-o�c�/j0\��|ߑ���`���?��?�n��u�js'|�y'�����ϕ�����`,�;v[�	�*I"�{�&�y)�rG�C����QX6�tg�p'�?��KP��-mp�ܰ�l�^�j)e��]���R�i�Q�Y��_\y<��}O��3A� ����"J��8q�E���d�_Ga�$ }7����0���F��ʒҖJ�Q�G�eHshU7�>�/�a].�C(K{A~�C�w]�����0D'_R��osa.@z0�._��<���Sd����Ӌ��m%+x'�ԑ_ko��U(8�;�8܍�	��#��
Z���,��*�@XA !���0�'���	�Ć}�>� _���#!�l����Q|�O��gUou��WKT�/r��<�0�C���:ĉ��E�3!LƦa@B56E!N�(�[zu���j\G�����6����]�����V^ɗ��TĨ�a@·��E�dxA��!P�\�-�_r,vd��+	{ Μ����N<��������f�������kgn���V�A����|t����w����VS���T��!���(��3���[j�\e(w`B�6M�XM,���7%�
��5��䊅7z��/��* ӺLvRt��ã�P?��[���V�y�H��>�U�a�X=O���!�"Y0X��S,۫�w/L+)=����o��MU�^�� �S���cD3ԥ-�Y�;ɥX�