-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "N-2017.12-SP2-4 -- Oct 23, 2018"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
sGVU57MmTPhHovckIdtWIAL6rnKTU8CcnoSm6chJFBX6NSYJb5YnXVbfKLR579gX
elehc3Qt5xw36Ar5KxGZWgyUC+6y3YLe8xA52E7/VwMcuHIFaGezEwD2Fp6WEHjR
cljOdlB1HFh+ldNVeXvMO0MkC6A/avwIPIHxePth02M=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 5584)
`protect data_block
mW+XPNB6uTTjuDtF/K1Dq/5mXkwuk3yr+KD1O/OBeMQpNFlU8v5OEqJCBnbdFnba
TTnbbINo+RHKxIAGnHBokjt8WWzI7jA95w80wRSyOikb9nsrw75c+23AIZMjnwaH
iGxvL1ilnpntRWe1lMtLjeOPAwsMfR+OKYJaAKJaOBDyjAous8lLRwWTVZs243qp
41F8dzHEqM+OquvZmPbIsm0QTg6bXNEb8WzNXvsJ0FEi5d9dtpllh+oC256/dcHv
xyvk/GB5TUZSVyf5ohtmZ1lMUKa7NtCHFHGVBSNe7fzSBrLBPJu6HymlKWk3VJUI
N+186oVWEU0era4SJY/PktyuG1v8oB3gDHGBBIc+/EaTtujmtbrdMg8rNuSPJkS0
8H93edLXAMQndCjGc75vmLW9fpG+RtgaP4I7XRfLR0BdObBcItoXWXmc/5867Hfw
Fgr7nZBs5MuQx4DLdFTZ5PCgq2PGf8hwk90ZpXS1Q4iCHwD7aAmZ2ucRq1K18Kut
x7M/13PjccpEgMgprbEKNl0ZlbmKGqbc9oAG1njdxq9pxfz1DNFlfpCm5tEarI64
ykKg2h9A/sM2squxWhXGihPJ4BcnkFQ5sQOenR/rGQ6KjIKZa9nIhhxh7ueeCoQ+
luz1TgUJcmsgZB92RYSXwMAathcg1AUVFKEVujZLBEDXV+EnzNF35YZIfgHT6zmm
mV0Vhp9JPNfg6qvgdxy31orHI7JdVT06jsFpK+xWyOf/OXcxmhxjuWpIMGYnY10+
Ogt7jtBa20KB4wYC8RbqY1A2UHB12ioMWQix/4XF+TX2Wh4Q5qp28bkXVsV5U8ke
WQX415WLtZHa8VNO7/Rf3UVLzYU/Sjp92atGZZpVUKaUArcpEEnm5dTh1RmJyMkL
gpzjRfu5Uvax9c3KhiEYXfIb516FiBbzE8aFkeyofSnYEUgymS5jKziFkyTDSlE7
OCoe0jaoqZpDte2pRLqDPfTobLMEvZAfbxM8VGyfvY1KShnuEs7nfmp1o3eFJqxJ
nxJsmIumszvS9aLN5OZB12LFKtf7HokD/mzo5FiPbPe2lhhi46y0gE4e3bmdbjIl
0jekcMi2deMfeaPDzj9iGCMA/wxtZuiCjH/5BzyZIUdWECnZH7A/C4B8Dr+CegIp
pY2bnc4JDHg4VS3QYrYa8Z92eoRcDXaTJWyOkVtIQnNmmiZh6WdwEJOK9LNbmC2l
3OzVMLaoSBR5LiuSPekKCb+E+4UuO4v0Bje1h9fMPFHuzOLA0xw3eS2QTWX1WGAs
Xh//dhrCWJIaGgGsFFj4yGffVtvp9dkt9M+OEngMYmCDR1HF1hsFMhdSW9hWYkZt
IgNnsXQkl8oVBvHeHnllPle8HT9UsOfBuG1atVAfyGui4S5KhlzOC3pQ1B7MCVdx
4TlRkQGljAslzWIKAwowYDxxUIJGu3sW+38jFdsryf1o02SqjiR4F0q9QKzPpMZQ
lqiVMaHBiK5gw18D5jDkNYfwWfbNrTJCxF1lyxmjasfq0+xXuGNFld44OnY+eRa7
vVGyfZKnfHrPvJ6EZ/MG5pwkrX9DKwz6kYGujDSlAWlUYsn9KRZTIFrgnBUHD9z1
t3nIxjhKF/ZKQEnsCsOCB5YuIustoRMcyFLGFUv1lvZgx3HtgsmcMHrP1o3hkoLq
0cIdDeom93nzvijt+kes9s3CEHexjU/ypvSGU1myA+EA9jBDbVRkxMqDxxidf8dz
40Icrw9XIT1T02CEQcqBwXa0geqzM2ikotLuTd0Q5MJE/UwqJ1y8MYgotCey1tIB
t3/JH1/qttnLmlbD/O4lx8yWFNdJY2h++V9XgKKp/pkxgZ37wG+HjL/81NRxpGc+
ARnn22L6sNqvmvZVO3g/G4Yh/uQwvTLerJNXd5WFbhBMp8wOvwja8N5itBDz01bv
Irkumu1H6MWebVluEBRuH2x22q8AekHqBFlSfF1lkflg1TDW0xaCgEh4lS+FqEUZ
29qTsK3atNA8MBo406jlxgBd9mMXCjVd1crh1TJNpPQ0CdxmXl+u17ohxTBDgam8
Qkm2JXeCOHE3JjwK9JwHLRcgjRhzObygwpl6/HEZFl0YnijsFligPwQuE/Jo9u2G
kWcQlaPoKKCpovTXYbrQh6v3cqyd+3VZDQJhQ9VJYFzXo0DkOEdcO3LSGJ96qgsA
XtqAP/JcjT1J6lyVaVcCFnx0lqlSOSmX3S6Gx6xN7ZWIbRvdHpzwZ+HdYijit4+H
htCROTrZlve41Bk8kevQvmSolrS4a3DPho0oIbKkAi0cQvjubmyhFEQZk+LeKnF1
+VelOEK7DSL+26IS3Hb6wVfN9NK4TWV8jB12inQdMWsg5VPvuLx46q1PAO1hLQW2
yDjSZVIBcrARRDsrUReqdZA0O3tsn8aYwtrXHChszYYvugERWJGgEw5f2hCJiQB0
3VEsF+hDfLAHgNn6YRu+pXaM5H5OGMS5uMREcBklDU76H6LEmOhQP3eTddiqb8CX
wdLIsicDOz0fRllVzNK4a+YP76o6TsS8RXry7Fer4QBYm4vEPZpjnDqeeu6mE1h3
/SnnW0MFWlVEi3q9G8VnyiQKwtBeoxXNuaWeDS3unl+jTMEaV6CZAEjjVx/hHfys
25J16U2bKlfQ9L72oM/Qsp54Q3oDVLLFhArI61ke4J4LqTuLs5jlKDGYeT1iSnkC
GeuX5LcKQjxCuOlaetf5RxO2MxKC8ZfKEEkIinvkVJBRlkE+zfsqqNjXrCuELdrr
fgALYUg0PFd5M7jGFyow7VZZSrV6vjxNLUpJxoFMrRQF9AZJ8ipbUH0juJTeEqPh
O3ugdughZEbSHYsekurYksra6YeoeS/JCLpcyxp7W+N4gcukIN+ffYuyucEGkvKj
Sb5K3F/3KScC5zvboDXLwJm5akYNKCu/yOjoBX0O6NbXIbetVR0ONBfAWu4P7lxL
fMHf405TPyfFYtZQrhqEcde8f/DqxplD+lUDLV5mQ31t7Egt7k/Jdxl5bf4bGK4I
Cg17knisLzws4bh9MX+Az/ulqfA7qvGfktYhZSVJ3SM/Dd3lT5e0kMAHn4gh2fkP
Wl9T9SbL9TexOPCkLCOd/sYN+g9Az/5BFO5wyk3mGdDfuP88QjfC6ZtNfRRisr9j
mCmXORj6ThcXb5DE4gDMFO3Q0qM7ngXj0swFMH6cqNqu9TJF0IApSAlkpvC4NrbH
jC5L5LGpjniy9CnKlK5d2XpooIMQt9SDulWZ1soP8HVopR0zpLkjlhA79TbjqcRw
kZc6KklELYiiywZ6SkFYghk5rIEkQ6IVDdNCDB2UIPyCeMoNECizmMES5cGwVDYb
fwMBPTkRG+HvXsjbIK3ZMvw19F3mNHnA0bzy6kFxJFctYJqH7lCi16qt2LPWqMGn
n4QCM2/XIp2Y3VRnjY3kmRdsXzAtQ5aj+5rtBv4R2lfTs2+gAV+FQqVjUcSWgiSc
NdVkkExoxPYKwCA3KXXjHnwyPRRR/qD0TI56N2AQ+XZVrpo3ouXsHIe8mdBVReUr
BvgtZHSAb/gp/IQ3VmeibqGSUGwkAMKGXrewhII/ruK6/OwbPjRPZTfg+r9XWqol
s23KCHwSpHbIqbBGndAlWNDnmZYHPQjCnS5df1VfHntL8RsvUsQSqKnlUzcLCat+
4WtPm2PuI5IhpSKpCtWTVLhdgTKEQ2/qlzD96DNFmO0W+823tNv45tcC3+qIfFmu
0i78hnPaZJLry1vVeU7fo9PHqG5aTjyemy0W0b1LXQpDQDLUSGi19K1Xd6OLPDkj
2XI7vF+h2s5ZZ4i/sT06+SKq5WZAzikw3RLee+ohKctG1niElcHmpDzzHcBzmANG
CV0VOI4C0GwKRp74X5xkEYhWH0qZOreuY1RoITPGH9SRpSawCzpoN9I4p+Q0bmp8
lYozb9BmS3/clUyrkSJdULMIwqHsIj4dAZ689WUneMMy1jxmm3W2TqR/V4JbPiqs
vyA+QMLbH3omMEI1sZ0VR1qJ1KVCOUeAZTSRVmRPbhylvmWOMAQ5W61G8vGGt0dy
MHGwCrjvf/6hF1lc3Bk5w3SLAq7yNQZoCkypTQlh+dImjeFoe/TmhTMv2V4U2R6A
UX2Lnck1ehI9+IhShGrfTelIqje/5dzNOZrdEeSV1Z7ll6N7KuAPNfGjjLRkY6ac
VMYORNoksQ+4Pf9ZkJrrff7N1cjvEcdnc9LMxIQEIwAh4/QuETBWYxgT6tOY/UkO
FM2W/iC1S/+9JT/oXBNG4jl6xXgqUZ9wq2qBqJRJV4DW/nKHQvje9b9365Hx0Sy9
k883hRgjrYVcJADLh9LWx8S0ehttHboh4PROTrIezd8rV5Tkcgm9HeUgq1qIejTF
LCOTDtPWWO75G1mPYSg/ObpakTob5bn2pVimwtOEbjKroGZ04tOD7379c3fQ9jlw
x6u0VSEEGIqxOnFnFx/7uGwlzsKkeOMiKdiEXUj+SZNT9QrD3NiB/VMNrpPWcqTo
kwPH10W/ImZkx25Q3kMCeIzLvrXC4GJICL6CDTD2uZaW9AD7rGeWOpYc7ATZX/m7
69A/9PO0GTleoGWqK47bHP9nH6bVynqZ6CKWRiAGA6TkU3Fwcv17yXifzAB00Ctx
VkkHvU8ZxG57z1AwWIFEeQNjwoagxe6m8dMmogvkHBMzl9EktogKYAedlYahYHW4
glb6aDcrl1PxJAENNRAR3QSH/lJpjXxcJESKG51k58cU6FyOzYbsI5Z1VM0+Nv03
QT5fhm0PU8V8PJ1trSYM2Ucz22zYAHw0YlpKxIZQl/xGeCv3xVN4SU40nVa7PO9F
eY22GYxr06Lj5RlAkr1DuBFVFODUk0qSaTLKT84UNr4iLoS8j4P6PWHdmVZjUAj7
18LfGmKgeyL9nZdl8hhyDS4F39OePdP8wrgHXPc0i1h7OUViETXMR+XUk5YjKhi0
fnzs9nsXjDkFNFVxc6hRTAkBobfs3KUDO2U4cpsCBWn3QbipgH/iCxIih8hSYJsc
2LYCbRhHAZ0C9elP27HmtsiKM34Jz93TiutOBZSmCuuobKfVRwTWoiSRxjaSaaEi
3tU/gvsw9XI+/xdGc7Wbgpwa0CnrBBMIYa7yHxhRyeGudiYzbez3koLERg5Lz/+c
PPI5N1HTD/u9JxhoFP9s7ugds9f0NB9vFNhO1RSfn237zf4XorYAPdyVdnI3EZiH
u/gh6Q1/Fl2dnj8TDWXtGNK9rr2m3Aw/c0tONie9KRV1cK4RVbIuCYhqLgR81H25
5h8r8TKBYfZ5Zv+Wv2odo5tGui2dDHNmGoYSbiIIjd94gy62TgOXHQ0f6chEdv7s
/K9lFlo1ZXDWjBO0KjSzD9DP6HP5iEmR1Rwtc0ZMVucigup+5Bgo1SlxP2i79BCW
J41SlWujwMdiwUz1MXTSb52OMBREPdj2P5e1Hav86kvnI6lVWfhk5m/kbSAY2W0+
/UiavApZ/Gzq0o9Wd7Rr2GOItKsUXDjcZMpS1FE31B7gUGDyxRo3zwaA/Ki7xtFR
Ynkm9frfRpm+dlpkKwc4I85CTL+3wdHv8GMMPALPYyTOwl+WH48YBcyJ1nerYs6t
L7bWkb7Pl72qKiRFLBh2wqxQ2QNXjLGJauoY0HZOrHR3lFBEWX7R7NeCnhMLadPo
RxIpSgfNo6t2WCjGr+qLhZ0Y8Wvfk4YTAN2Dz8v/SJgIcDgGCmRjAZZbOid8E+FN
Y5MTG0PmtZ6RJ76y/eNCNsH+feVagQkF7lGwqRG9apEJ2WBbcRs+X7elBzSgZ+d3
ERLr73vFM/n8NMEeC5tF1s5+UtMzCdEzUQ1x2HbKagfLP4c4T35/hLmodMHpww70
C8IdxQ+VXsIAbHbr1P5aPb+FwBCJqHfduK9kCFBPzVCBSeNd32uGnlImfbINQuJ7
U7ry4a3scEOZkI73doLk8JLpJ3ncxfs1EcJE2pZq+B98Wc38SuIuHCzwAJlR2VPJ
FQ7T0l880H3PrkQis8LdUpU1V6UqOO0a2Uh3EtrMPdNjury15vsGSWrHTZv/IW3L
Hij/kxDcPgvlAVfwSOqSBRm1CsV28Z3hbzQDLYENAxYw9oY29qDp9Pi1v+xPWQTK
gDRaOkYcgxai7GIqDPNm4aQObL3ym/eI+1ux7QNIqAkoae1fD8Q0mgFgSnZnRe7c
wunAx2lEptwuNOLF0pYfpHXdvELC4ufRXA1RA+BibnbeQ8yww7S/n1Og5qZFcwRj
B2RJvJTFGuyZnSkBZyssQYyFlQ7BJRJw5cEbrGI+zxNy9XyJQRQ5M93/AXFXbWGV
cYLQG1L6pK2GkhrAMm654gvHQ6qAJP9wiRYNb2x4ayW8apRTQYXTmzZIZ8e2Uitz
nRL480iXKMhyx64HgLO1aZcfUbefNr7p5qROFXXcWwVcl94769g23ZRsuffKpJIe
6CyjphrUTp855gjWYhVQgZl0a//UAQep91LvXqxWkliT0zTd13AfIzerXiq0JJAs
IO36VsTSvdrXhBGSgDDf3XqEVRZz806A1EbS6FB3otSEIiHweqEZ0AkIUJMOJ5sw
L6hoUYAiPH2aLR5kxVesxYhzEd3lQFCJjw8hCv+5+az5fz/5zBTHJJszVWk2nH1x
uieYTiDHwzEaXypPsNjUIfvmflIVPJpAZChxMLFBLIx6aTqYchNe1imwoJYXnOyr
uMQHDU/zuhSrzcm3Vf/SEiw4JCZP6Opbm224rQ38rGKShp2WOSdFsHSwE9IkzmGf
M9xEvTl12Yr/zAwAN/8RU39nN4RkxF5mq5ekiZtD+TptA+kO1uyIK4tHZQAbdM4z
lK2VLd16xbIjBAXSk5PdJNSwNkDu6g1SmEcDrkg7l7iy+ti0l7x+xY+MEMPk7m0X
KLVj5Tsbia+tPMaI02nzFL57HWN87pCjQ0EWXk9xFR2Jdk6e/lw8AaihUMyQyUtJ
Am4YE7uIw+G3oVUajQCtzx8LS/nhz0necslqUwYHtdGKC97TJyepLU16RUg1FLSF
hb2gOzsQTK889eRq5bf/F49ikNP/c6pX9iwuIcVfNd3qkkKKQiY7lsKA2onGBlz0
bRIRFMbIg3shjp7XiwUv0T676r/+nNWSrEM02GLnDyCqHO4PFCCI98SFi2rhAwy6
ri2wCV8rAJEtoL3mxUWVfKcS2xj4LbE7BtS5ZSqUhnDo3PDLfjoeDpxxsTAgV7lP
wh2hqI6+hEGVJNnifcBaOLNdy/TGkoB6yPc6imR0eTDPwFla3mTBJbQN+x5NDHLb
i7Kcd64K0VLKRDQz5Apel3pyCgZJ2KsoExqr/nYruoGIUkQqL18QuVqUNf4LPSEd
N+j5uUqGqlFbjUCV9rU2vqvLat8cwzcKUf3nabXSArBE4r6lc+bvxvn/SwZqCdmn
pbCugbAC8DWy9LnQ8lYHOsdMfIKTufUxfmFY2fJuiIC8yxxzJjOUaFgDbZLbsB7u
l9q43Jlk1Yxb0sW8psuTFA==
`protect end_protected
