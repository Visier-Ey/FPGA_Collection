-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
wRQzu/Fiy7UZBw1H4kCNJYVzGE5a7Nc0ujWSV8sT0ymjiVjqQs3EGZfjfp8uKizn4XSrL2sECE/G
7tkZ6z703l74RCrnVE8JyAVs5MqxqelOWV5Y454kn2cxYbM8H/MGs6OkNuKS9fCor6/FoeH9pVWe
89iV2fuZDaUmWpFMlOdeqw5OHP3TZXlVFbIlHYQpJeT+GvfvF1n4gGcBlRimn7c0DPE8LoXbmWib
S6GjvX8gFAafjcOoD8PWEi5EmoBCHr0j8rzpOt4VChLJTsBAhH3jQkc972BOJmE6eEjzLnzR/fO9
4SZd14Pbk+WTMH1+mfCAh021eD91b6dfaNHKxQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7712)
`protect data_block
RHlON9/2Ryc60adlJT1gZvSCA24Fih2v1FBQ9TBP8u2YwIGq3LIPPw7+pHTRtLTNT7pJ5BNSsf5u
doGdMBPXYIzdkl/pkImyxevFN6eObPp71Bw84EyxUc74TNcyJgI2do8092uNiNAWXDW1EN5g2btZ
5BRJKGKx+LgKUEt75xJ5sQjh/G8s2SQ3H7WrvIPi3bE8QHyNs+c38JnBO1QeiYZfenFNx435YJp9
61LhtdQu7B2Zrd5Yn75kFj5ZZ7/2sRsCHfxITRIdLlL09/kEKb0B4WVrtVqK/UmCyYK4INltvBDK
rrf7HYmg9vgc15cm0ijniDtYXCw4h8XBrvObzBUhFs6JML1L2dQlTbFjOSy3L/xw1zFcwZmmqJUQ
lYzXcbWw5UCYNzbHktB2xGclaEDAb0JCsgcyMl6we9sO7SDnrzWzu7wBAKX7tknpCPWP3qzhZWE7
KJOJxZ+jVYqxa/nBh7pnVSW39kx30kW2i+MZ9I/AvjlwGy05qJQcxz0gIP+i3jjcMY2SZ1JZG8pf
IhNx505ulVZJNWkcqUZKsNkgJAkC2XqB6S7IBgysAhvlhj248HagatSVWcVajawzKKw2vlS5mZh/
1mRRJ1wWOgc+jF9xStaOwWvdIdWJopfY4a22/FYdEd1/7XG8mRBwZHi7q1FxvGU94eMRugjhZ/eN
7Y0Stmv8ewAITQ89g2ka0yBCDzwoCay45z/fi68I6Ew0Mln7GX/0/KtD4JRnjydLL1WrTEq6Ce3W
ZDHdQDa6kBs6NCUCrnEWoDQP3jD459npY9KpETE4zss4HCBIif9r4tz7xn35sf6UEDi02wZUvZg1
xfjkhaDswTYPcpXlTyfAG4Z5Y33iFtcdoacfgi4TLtRvAQT/Beb5qg3MdvR8TYqFf+pBgcHC8/Io
NCFGX5+rZ8z1dZbHYfavFK3MV6XAwixFzouRjSLpHaqsitVG1C+MSpjQzk7VA+kec1VHuV8mHOJD
1IVUBjvyHibyBK6hCApbxf/IkK04aSIvI5AEMuyWAUocNKLuape1OeouV+YSlMeA10H1Mpx7fYQt
ykzm4uOmmw3VtVnBQCnyGWChfUtQgFBgzCjrnyhrO1R2o/Z+p2o1tb4aOAYw/4ShTwzsF/+i3/jb
Ll75fqxF6ytVjmFvCRq+yi+acIfTkVTGQDtd3Ou767ogl/lOLdPvZDl31XLZOXxkokcWqJWMQSXx
2YSV2Z62Hw7FKWDM8yozIJIYQTkg/9+LUBVGoQUNJHrtmGfkHvg5wuW1Ahj8yaPEIUs/QkbZ26jz
/IThlIWIJK2TJksyjW0Zv8NhQf5C67n07lRaUHRRXJTc/iDXpUBIHjG3nQhMxq/IKEnp2tYNyrfd
CG4iNO1Tk9VfUdcBARtYPm7hYrBRv4KWD/oH6E9dKVtkVZc+wIWa5CDOG2WdFGp/ZSC3/N9ji3Rm
3oDouSw3JeZaK7dbvGhrwe8jYGgmuY0u7gHYwNv5P+cp4q2We+DLqox+PVsEyj6YY82IoYQQk/Pw
Zrjo/uYy1cKofIftkZpXgiUhzgtZjDPF0n9yRlGRzLi4IcnnKYOIsp7lTA3iM2OESUBZenIGdyMS
S7qXpg+Mf8TpVnF0MTf42XsDTnSS1aXVpbQd2UKjSy2xeKSye2qdhaOQdsrKk24wA/tPXDoeR3NT
HMIhNqW4LBHJa7ISkF37/UFVIMi1udXr1lUGiOb+e02anNG5krIFkFqBcHtVwF4pSa6ko+TKpDXv
lliKgg4E9RN08XYkebtt0Ur/f0HGzxf6GLEFm6jsL0VN2PX3pNWXsYTB983oPUHXYaZJJETZVSQn
c8UuybsjSbP61F4SafX5hWVhTjgmorSPOwehQHhuzEToAQecUZrGGClsq/kxMTHEUrhkk4qCtQzW
ZRUTsC3oLuWBRlx4ZazJ7ckRMdxZXLWvEOB33ZKpwSBel/kPazY5+2zntcHU9zUln0JRmUG8Ut09
prZmu6fY1ZjT+AYeDKCMOc58kvU+hZmJzNfzzCMRB/jJ4yqSciheOivTzSy4RMvE9kiUY9gn8lUj
RkWLOWDK+iKRfj3mHcI/Lm+oR1NTbqJdfcgXUi5OGwxDauDUJkxJmCxuxdO1srZPyfDrbDBOfdtB
Tln/ZrR+wj1GmvkG6s52c2xoKgkgiYA6CisL+kTD2G6mLhHQ9KRVTV/9jrlsbZKpU6NG4+Qo+Suq
yPDftUInDvlyp9gFSgxecRiApnnGLMr0PIpU8o6WzKXAJ9TjkDZ+Ca4AXqJ7BaKMLb+TtAh3I2fg
iL6d4xQdjBkAcnF8xm7XRZ2Yd7dCLvElPM150tC01Svl1Oxb1uz3UZw5ojb2iPR1fQ3eGL1LeaUd
lt/8mMO0k2lznCW/r+L196ub+g6BemcBD8MtE3+QnYTGnyFB8Q/jADQMPBoDEiMUOvyj9iQj6vDv
qKArA2AUjDvN7TpsLrjkSu2iaBFEfMCbMRteBkZwIj9IxpUtAgJHSZ548IfOGWkS8ZFoHwrG+mXq
fSyoU8Yp6HNUGIuVxDXDGUpse68XJX5umYxfWm3wAekweBhfm/Cq37afgBgIrRFgGPd0OrYocOHB
NxJomIE04ywHV3Dxb525nD+gLb35PJWJ87yxSFYg5FnN0a/RkXeLc04AlgRUaN+JKroRdotxm1CV
ev/LWRqrUx/KLrKfvUfS3Y0s0B6wiK4VWSfbm63N6IMC2OLRsUi88pffMA9DNHCQZ7hfH5oDNbvt
qS2W7qWrtvPL2P7VUzEcE/Z6/n4UvFgMir8Ky0QraFqBDzQVPAq7HYsEfPvShTsPVoGnoqmihsQl
c2fVE2DvXXw9ob1lRO18ZKf2Up/M3MiKdKnr8QBeDhrgkIOcqaNrub8K2QbOzmY+FWG0BB8Dwfja
DBmsRz7J9s8dR7+AVI27Dj5NYXVmOBA53QNOMd2B2sRcBhr28xd1zhwsijKKLyrUrTmdz1JQ3Ajn
AIWIbNgDBUAzeYTHGzqmYMbl7ySuafcoRPQajvzfGkdXnlOEwFUkGHVRhJitwtdrnZ7fBMX/GFhO
wp3DfZkFNb3qR4ZPvSRwUpVJijnSj1+aIYbzPgFazvZat0bgpY1ICJX0uYXqwcS3Tm3GeNDskxeK
BSvuwzr3EHRnjR+gtf/tpnL50GkXYnVVD1ShBJPWffEVY173voRIUzQMVi4fynbY3rqXyx8s2n9T
WKFduOKboR6zOerY8jy/ShEckAQkZtUs6uBEFEGzbUIU+UHOdDuPKN2EgHEgGgbeagy2xbZ6pzJK
qLRn9cRoaHz3aYfr/mlwu2ga1O7l9Qir563BQQBHA31+OShLy++ZD1Mw/kbfjKAzL3D4GbqsICpv
Ugnzr2KodJakKdCAbO8xmWH1W0RTT+Nve/qTbtHYqNThiWCPQqW/TkL+jKYP+WfBdWWjikGAceud
V8OJk+hbgMk/RTVrKA6KigjOWARae1dUiKwRTPGa+62VwKdjCRJbqQ4LtV6v6JWbYakOINjP+7ax
4KJt5cwmIS0DJCIW8EW4bLpfkpa6Sra7NPIwlQpkwdUa5on0/9gwYTbArMbLH0IZzQQR3gbZIqUQ
mF1tyhs+I9Bd1BZhaTD0C6pnlUsgbMpWv5lWVcuMKwoHsLK5NjgU+vIMEOe6mduYXKMhNwIRxuH4
uXvwPn28ZaHFIrA8F7T/g1zlfNdXP2u6RIET2iaSfAiN5IZmRJlOX/cL44Vlf2jtt1cqIe6mkxzp
sTNQ1sUq7diR95txp0/hA2guLsPqOfn15SpVw1KVmb+eQhZpC4taz2ASGn+gTyxupwo4BzZ3Nkgv
6m6jP/47bqLNh02ifgtst8MboRKD9KW123yv6+ib/l0QVZ6Cycl0iXQah7Q9G90KBCEMYBnJUx9A
9qZsd5lcRH3grXz0bGbPLgBMyxqEQch8lVFkBD5r9AS+deyz0Y/n4ekI0jQ7s//R6thvWwYxJSg7
Sj0kAGnGkYS1hVdbji6kPYgx7rP8xy9LDK6w6uRiBGnLD7XqwEEJaXgg0wOnlVJH80iM4kOAu94W
ZO1dsxlYb5WZwNLEyp5BONbiQXyXmjf4IaHxc/f+ZGOOJxG26F+dTdSrkaImCcGQZU7FqKHpVnaU
GHJqdqR60q8PHA076gnhNT8mpeFUrie2HZWlp8RWAuK31hPKvFW1GiJ0JLVYUpFBbkUhIqIMLcPD
TlqXV5m9M9lVA7kAAPdH8BMh7cMAsVPr5z1yEfw4Xcfolo5SSBo+zwgkpod82hSgwLHQYTDFI0I8
1If6qqi9pWDC0Z5FSxyDdJoPU/2HBrGulJlpFcfFWRcnFOBPrwhh4R7I7YOvqHaMQOUrdLOr8kjD
oyshxbwzCLvtIfPM+gs6y5m5HDVFDGUj68mkiXbXiv6pe4iSXQ2eXrCBLr4y3LeGQbN3IMXEVQ5y
HjAW1Z1mO9u0jonmC4yvNFs7dyoeO1vorqQWHyEJ1e165+b6bKfqsREi4rePJPx/YGbUKmoj4kJB
NUYiwZsFT9QMOE8hFrRX5JymlbEIbiiPx6xNJvWuFci874GhXQQyV8YyiXwk7y+ddE+bZF+4r6dI
kMCciG/1RS8Jit1HkxlAi0HfcOqS1mTzk0peMcR/Fnh7Pt5DN7HP8XKfu5qkLCIZp4e00BIuAOaP
g5PQkD7ZDh4LsL8pNREMuqv8oGtW42ktAYyCuZNst1+Xp5nIlFhzEtu2fv44OtTxk9nD2XbCE/Rt
rb67NCgxv463QCKKuP7MXME/IkrILVCDFv/NUzbJ7DA27qwM1IULn+9npyx0tEUZDPCKqPCxgQO3
s63fl2dzPts9itbSNeu36p3LUeiuKJvHUyCpwhhCZkwasrVAeIguOslcTALyi5s8Eb+PgpVhcyOv
/Ua3dRdAkTjoyUopGJyN9DfSRhS1SkOQJgaUbdbrokMw8OG9152xU4xgiybfYb5Mzc8+UGWVP1q/
/2su7YlEFgEAiyj5goZ+j+wQuFI+cH0rkjYokUO7q1gLpjcyI6lZYZZdNTh1vH8EK/VlcrRFCtwk
QoNaJ2i3DQ/hqGYtbBhziHX7e19PQ21CqK9W6CaNPLIDD4wDv4mEPqwpu1Govykxj8tObEU1YWEV
cd7fMv119/Ba92/DPdpZOrB5uK1pPekEu6TuEkr2nGDNk3I21SCYHjB9sbHGhHNWxN0FbuN2g7iC
FRFbo68OeoxpY5BHgOHkPm4JK2l14RFMy7VNH7nuJaaTJF0wtwmAUR7fV4WtraXmS71Tb5Qigs9L
uhTyw0yizCEq95SAzBadv49tKN1gsNECy3nEKjPXYNoHNAZGCgn8d+s7Dt4Cg3YarBLoOBJeHFuQ
+g8MLmI5nY7XeAjbo8+pA9M/F+V1MfbblWy6bChrI1+nwnw9Vs7tDW2TaH7qcEqnVV0BYMshNyI9
0qEf1LXEhBlzFBD5mei6GOfcyAyCsqVxY2E7tUbQCk7ynyRwE/EME3XQ/lCQ7RQNAO+J/JfE6nEn
LoXdotcnEcOK+BRFWffxiNYyi1gXPCOE6xdL3AuOoCZbxxspNnX6FFyz379C2mIppXH04Es+4U+j
lDvYcm8UUsVRGEaeywXYE215MXu+Ajakc0G6xNIPHWQNTTWRAjzhhh4+NePHuKWnAUQ/PaMNgClk
luI+Tks0a98trvNA2KhvMUDsXMVD+iO0IULq45vVgJGTyig0YEy+p3nLYNBEn2BEOOxgvsk82pXa
5jgJzu33NkqnoiPRmJyDkdzki2B6hZ9zYyZzVbJru5POE0JKcg7IjOv0f7DhwwJnN7r/l/67350Y
vzboGorCMZEdD//Z3N5Lwy23wQBI31VYgtGqKAxTRsdeP54Sw+CvcZ9uNM6J0lgZuK058GDt60Cx
Cof7x9bdcF6pghz/H8CxksFlxWN6gM4GfUCfrAHH5rJR6XaFmHepADmCBhXKOYJJx0KJh7oDDWaZ
G2GnAt6+KYgE+6JjF7nSOQKf7pucR/PKRhSJPZ1+8ikvZXg6iYgu4lRqXQSupKbMlvrh0OHtp+yq
ptUeMCNJhJAxjAoAy36skDsDtyZeT/o+jCC43uzJbmPMemRFcpWDU5xM0Ln56EFsdv7MP/WcPJCD
wAJvV+TcPEWZ2vIR7sz/Os5dhjEWJIiwbmbwicv3oGwWXj8AqXPuVKJGrIsrMBUsr3m1lkl8CVle
JTET3iy7QQjcnS+nTrxNkqKHdV0uQr4cV9b9nCvO+UyFYHF6Itzg0EKZhKRvsXLEd67/1C9Jnksa
S6g9M+kGaWc+Pd4a3t5t9Rd++Qo7boeMhUZCjZwLGZJOgPC44PNNaz6pMWv6C4VdcuD20AmykkSN
0GLuV5At/g2Um4SQysyg6nop84XNo8xV0agthwnI2Wuj6umxQblZBwsTtmlaMK0fEb9kyrx0+TnG
CC+nU9TZFrtWNcgBc6mmHKwV/D4LjDq3oI5d1/fcXKLSxsaedm3Me/KkupF2DwjWRRMLTdrR4EYN
nQLA3TFZUjaKyPSfIZMGA/Yj2slWvv2KbuaVxSoDsutMulOroV/2XAzwFr5fpc7WMVnHpxOeKBT4
nnrQcRrw9S6X1/QtMQ7S5uGXVy32zw/uri35wTiW1Px6DebfZo+ShhwvVKm4vN4Pbr99rHhpgVql
QYU3erpNKkXaIB4muxH3jqe1YwomwgnHIKw5RprNywySGNpCGnXvEO2YBKFsbW9qKkRyFH66LX/H
cLqK4AfaNMGMzCSklrUNcl5v743MQVViG7fsRPcqCsn/7elCczZ8G6mSs7BQXXJ3wLMLXLXUeZHH
PtxcmQkQfQWZB2bgN1pXggmQ1YPpoK7+JZJc6p/dDWl0HMjLMgINDI7w21COLtaxABLN5hYDcyc4
VZDLoHKCBODXCVtMgPkdO1vJ3GWkbVDvWN6qax7CHbs5VzB/PE0CdNk2PBsTA0yfjBzEUlaTavH5
f2eOOOUsgDPWNWw2N8dXIkvlAGWHiSVRdiabqa6fVNWdbuApVoUQcKB5PhOr+/ssXvEuIT31yYAF
t+BP155cj1Jpdfjn2poUt5Ur5mJT+1E7BpF4A+eb/rpip1HaqobA7DSWjkaEkjWxre+OG6tEXvXJ
K3h2bn9Ecvre6AzySMsID6D/W7izMokXBDixMyzCZ4k66ir2GQ4qFQnDvaeSrcJIpcU3+90vjQmE
HkqDNKkBDU7DrmIyxPBqelSA1CgABwL21VjK3LFFZUF0OqSixjhkSKNMKo86zpIGCCGAcbUNpbx6
DBacAtb1B9WBYZ3V6rEGEEjm/SbhgMvwxpUY1wlc8DOt5MTJzJ7N+r1Q/asmE+u1yTSZqxBbQX1W
qnCmxH5rQlK/CqCbxBPnGgF+sKrG5iUt02B3NWpA3n1IQeSmhaJ8Leap5zlIOH7n0QpIs57DIZyT
iPCR1QXJ/0sGw0i00ljggZ2PSbCt+uRyyLUsQrSkXDIZ2W6fHjD9Cm6JXjJDQMLXfAce+7cTptQx
FLPA1MOf2waQtiVpAXOyVjnybBgvsaW/Fa3Iv84TqzqjgUC4h0dw3+j0s+IpAYRAkYGweM3CEVaF
Ma/JPBZT0us86hKntT0VQ08hOgk4JJ3qJA/YdVXF7HQyrqzfnEpPXtDNUAQIuc/Mg10N9D1Wihst
6hVR5h0c2gg8BmxBM/Btvs2mgYr79JK7gtoicTGrkTwr235bkiJRo3xB3KDtL6DMz6rUQaf5xPTG
qdC4TxCxVMyDSYA0WDcMgk9n7ZoIOP+LZTkypyUFFmDTGKpGNzi949Wqy5CYr53y3X/JSfoaNwAv
M8YGBi10ccSkz/KMfS7vgMYS9GtDHUZs6QnZzaL0qewN+TZBgHpPr9U/bOXjI8+mNlaf2VdpVuwE
r02muqKcVGXrBAukh5GhubB/6nbkMiJwsqnpnooHV/i7lAO6GnV2d9GBrtnqAKe/HLxCAqDmrNGL
oLVJo9jRh113kZjDR2+H70xADXtOFhYTda0KoUny6CCL0a5jwYpZr70vXNynScsqo1gs0wYQ6POR
wiTCWe/B4jkYFQ7HM2omLkF7B0DBDSXOIJeUnRiBugVu9q7i44moLfhzNHMvJr0+Tz+t9wPXO1ZI
xxd3zJozdDR5chg3F8a6M2gWq2sa3PPXpo8qY29term2ryuvBSyMAQ2uoRLywKdliCQPwgebWuw4
ksgTC4g4DhUx5kDajBfqwUEUVWl5wTda6MUm7xH0aDmnQm45WmxcpELT3z6NbmTVdpQbmFABXez/
6d7LyR8X1k5Hahx74m7gloGFaB/I89Y2JGvcZNo6l7MY9yOycA+9fSrdwWqQxtM2ied9KGhGbplm
hHHEM8X3JfaAsSBhTbG61ZP8NHTDzTzAtuVS20YvCgXoCQ3Vk6hkNk+uyWx6kGTizz7ev80f+0ZU
IOI6qjLZsmiQOa8gVmnokn2jP19CJsErAqbhQAj9G/Zado8YniZ9mu+k+CDeGisSoClg9EfFtn83
0T9UgJdA0acbZgxoKIUdlX/S8JfGDaw/Gp7jMA5djwyZNP0jQlJy+WFXXy38GH7lUW/e39JgjQV9
o6MO1DFy0YPdWuboSeuy9wUvDHi1Es8ZBVfIpLHfkdWEi6Wjhtp+U+60rv079VXZn7p+OZGnWOct
XsPW9Dd0foJCJpGOMAXuet+vGq4nxKlmty2deTNQKkuoKyHnnfsWmR0QRprjeyVupwG29NARGfmN
HE44tSYEwODBnNoo1mcesouUTve0pexu+GCt4tqo+I3qh+COFKMp9FfnH0EATE8+mD5tX/wUhuiD
Zh88bSIj3yXxs1uoeXGhKl5gyITfRsgF/xcL3v3JTpHrUpK+hwEdNu3GPd7j639jFfF84Q2qfQBR
bPt2nBcmQzruljRHdwiOt8/h8jeGrhx4wHlC4TWh2nptgHc/ss7inz7AmdlBvUME4GuwUhZv1Dzt
yHNxrgXFhmIagmBSzxBtxYXV2qn52o/FocLWPhlpvwONyEmowxep/vuonsj2seN91nhDsb8ej/ba
ha4Bv3cayj+CqcQF4n0bjopeID8Zkm2Uno8xm8Fo2MtOQ08o6t+weqvX6N+M+RExNJ18devPsPz3
LazqXh4jqNSw+4vCdUdYn18AtP/ct+BceYDMxXHkmCXhfMvZ3nJaCvc7FB+XCnkb1DdeMQiAJHV0
ILdhR3CyC8rZGiAMlcBAV2XL0mf5Hhdo9uPZ/ZUWZk52G+eaw6t6TnJs1kCFzfKMdxDZ1p9Qroym
lzfVfq4BxTL2Q4oGZ9eeo5AOgU1XQoIQpMp9qROytJ/RjTbVGoMMzr9dfBdt9ZLTV4HTFmnoJsKZ
XCbqFhsq97GNEXW/ealv+TPwPwaLwAlUZa5fsR8rolgeLBdW7Koogz9mkccPnepNO2StqcjQrGHm
B7GET9/Prkad4WVorYoEVlbTGP1dOFZW7KnZ3XPm0AdIGsL8tiNMtJqNAXWdBHQtwPjtS/LYarJw
PaCltJ/nfLgiMeSMZxuvYFK9zIyytyRkUwCsaiwxgPeJgYflGh1XAu0CpZxGNpLh72iqMudhhL/+
WR45VtlhxjYOelGDXG8m9qo3SBKLH3n/lzzl1/atFfM/RornzAZDlTvY2Vb2tHA9kbdK4IImcMY4
Jgs6udbrENY8mbR8Jo15OVMhkw9EJVuX1gCrockdsbn9ueG5HKkIOhVvNDzTOJH/AMRSKIynhj41
eLbXYdLHjSDwzvr5WpSET0CPh+dCEDw/gYAC54TQx4ZkU3LQTkmkFFpaKkwlfK0ipzf8TOYDU6pr
9zeTaZjTSWOPxq91PTlJjvDRzBnSoGSUkkVHOpS0PdgoMO+scQO2k5UhuEatC2O4STVSr3Gu68i/
Ubiyz7I5pCDWK9Zv7/656ll0g2lJBNvmlkCjJI65dYE4SAEpHnyT6DOlqq/RhnaRxE1vae5PVEd2
WWNeDFtfYMhSah4FWi2Xh8RQoNthICT7zvKmwCXTQn30cDY29st03SKLWnhRgWX6lfi8vRyMDir9
9N6f6wjkfeBzwsC5J1OLdOxZgwkqf7f8n7EYX3u9Iph7dUjTeHavmkE9tnbTM3dt8GJzl/vSbxHi
s6jXzO3oAjRvovkodKAtiH617e5pClPqcDSNOf4bbhaoR3041skROTHjJzmv6T1ezJwNZYFI8+R3
jOGa4fQvCD54acfWQmDV/SbKaG55MEcLNmJ0VCV1/x0ZIIIZgwY2xTOBtrM0qNCjIRGHgHaa6bPJ
AuKikT4fDI/keK86/L0W2afZfjjW9VBqL/jtXAFxvBQMA2cNzHbtn0UNzaw2S1/rOCJ17E2lcPWV
A0Ju3dmmAYqZrY1xjDQsngo=
`protect end_protected
