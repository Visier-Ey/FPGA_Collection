-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "N-2017.12-SP2-4 -- Oct 23, 2018"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
2Xyw+Yr807elJ0bG508jLr7NcCl2B1aRT6ngEiZ41dQOVUYwCWItJbFEJWp45eNZ
NczI6OIhpKPn3yzbWG47kkYJNBHq8QvPx4++NmXWa+cqeUVR5X8NQH/sTQA1gM+/
7orgZCkc7Y0JoSyu0yTJ+KFq+BcR8TvdtX7cvZS/WOM=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 13056)
`protect data_block
dcq/1x9qBCV5CqwyK+o9DW8s25ZbutI/02kWA3chIHx7L+VnCleOIRqROu+Bkd3u
7kyE3dcNc6duvnqQCeJebBsNeaAiXFOnj6Yil64ZgvIzGERobvvT6MxQZrXBC9UT
b0zIHihxoXqJDa/ifG2rkNay0wlZzDdKYAhwHWx9uLpqRBIzEOZSNU6tvWNNOYec
ABuNbairV6/Y1FIlBH6bSa7FFQ5kQUVVuksvUSqOs9y6SxlzvVI0aBEidhNjVi8b
n6/63JwSq0+bbo8nO9BKJNakmLex6vhWREO/fbgAIw8Vd5rHnPCqrfXfGDAJygCc
Pmhfe5P2DpoXFbG9YSZvlKUEA0zOlTWGulNml1SJKw794s44hWkBgedqbkG/Ej6q
7ajgDsbVuJnxfM0vUWnT+0c1vGr8zDJhMIg7hg8fokvrKMB1V9mv7M7cHxyCG9zp
djv2qvHIjfWVyxCEuSrJuE8VYOUV3Rq0gQAc6okA9XIy9e6evDMcfb6VHKIzeJCE
KmyG8V+TchrHhxax+wqsJro9bclwvIb+nBQEIumn6s4MRmgHuWC+CYAekkKyVZN7
PFm7/4ok2aZQxZZnPBF8+CGYnXS5br862uzzBmZh3Fc4fa5P9hm+U7CnF4+gOXBc
mycpcS5KzDFnvbrGqs0m9HK7CnhUhZrG5KzMrJdcUlOLKHOvdH3it69Z51GKFFgM
otZx+g/r8zkf7QGplSY4Q408HCj3Vn4Lj1fT9ZrjBnQfhiChSxpLNCYSQd3ryCFS
vRshPc++2miOFSVZP1MCNbGdPvrk6BVbnid91rkAe58GEHZtau/NRS+EMLWuc/Ob
XV343kn108SeyQ/4yx+L5Bir2kzHM4bXAW2A6UQtP8aTbU84w0ETad1BDTxXJkNo
gpVsO7TIX/Xf9hnt6SrdCZR8CfmcBY8b1k8skR6NixkjCF5E2B63pj5ebNb8s+Q3
A3ysXpHDz+W7L4oNUucqPIfM7+QEZj16AsbyAPBfzTmOOJ6REIZMA8AuQ/y6Ia4h
cCZlzx7Q6Acm5w1fwNyKfLSQLT5oFL/upErN7GA5O4Za/XxZn/jdWzAnyq4Q6L5I
I160S64sil+vu+ONzXwXQuxYw8bCmJfaI8R2wGLupaKGTyeaPnBW4M4eHs8cj6zQ
h5eW+lqIN/yiHGU/3Hp1IpNW4Q+Lnr9TXg29qoRAJBKgAczuUjpH4Av0MlOfWuNf
u8Crs+FBVOYca7RDQ7l8Z/SJmovbDZLPufPj5/voSuQssYcbMitwxHUyoAlurifw
YqUuJv0LTwuPYMzFPXdpcsu99OmxWV64tqP7oUm4iHEdfC61AR5sTqsequLrbcLE
kInxhXxu1jmiatc9cwqz3csCCDeZ3+sqi3etCt3AY4EHorisAUzZt0NTm0DLOwEt
SynQIqUB6k/PtTwp6BHi1eBuveH6V41cuGdBW2SPaa1fWqpuHogG2gM4obwUfQiK
tFCVreX8l399ghmNUS/PTUNVQuVaJTkDd0Gg87BVP0piI3Pxlny6v9rrz0p/lS5d
FTHAylMBKun3yMqjtqXblCIWh3WHcweRKiqcu4wMWzMgubZ98+/eBZjNReNv+qcH
pjnEMwL6gbXlTMYVmj6iRLKYS601vYpzSnF5Tv6nWHZYIDWadckYpfPr2gGngWvO
x+pfTQIy6ZIMm9svmQ9g4X8vPVAA3Q/89lcMHF2QpMVZnjw3ihcejyO/iPgIZ98C
cLFoZrUkotB2iVq/Uapv0klmU+krDMLdR7NL6DJgHRZRSu7eXJlqw6xxRrqxqsNX
q5nMejz3akM02MxazceAFjGCIpgLYVisqdzREKOKPxV4shtTZwQZn67VTd4jh+dE
rgkb4bdPufQA82l58IT1/brQdR0eWgafBfa4RS6BpcQIS/KSGozMP+j7oPnWcsib
iURpHnpUoBG2PFuht23TmmdwAiXY22os2gBCkmiKYu2G+Am4ccYj3BcoYUIVnNMb
lV9Vwd4k2v/LvGrIYqebzM9jUbWmDT+J1wgUywxvR2Chdau8nqoUnX491VD1s4mz
ZsAqm568jUl7hOqeJ6YsS3RIQgme/0o7U04QBDAWfBKKelgrKhu0AjScjKZyPZDq
/TxURjUpVOHE/XScQEGDGGuEfTaLQ8BZcJLq88URt43kiO+nWLvb5E/8ybVC+b/V
oCIixp+Cl8Y+KSoHhIMfdPM7sTXq07PUNe/PVeEArcq88bAiMPqGelGt6fezW6GE
quZcCPSuX21ZXdTTZSyIwxKy9UvUEaskRwyJgiVi5xYA3dSiwIvUxvUaJRP8CBRX
x3i+0WORO+852ZvTQ2a8x9hmXT2Khsb8pCaZAJFiW4y7kCZxSFT3A4Bb2xul94kW
WCwpYLAJPFnsv+BLympGJfxkLSxey4qIUqzfvRAYnj/WoCe/FnNl4EArvtCA9LcT
HIuJzAWNV9LU5YPhpLEmiDwvc+sJPLBrz0R9GO37Fn4/f1taR97iaFulc9fMx/jH
87qKfogITStsCc+QW6imZcnNU8xSbxOYpZMAMU+Z+ETJ959XEmyKYi//U4Kn0LrF
N7fe9rn5YNc7DriLEdfGu8W6d4E+syoutZEtxKKrF6537yc96WUNXYJHBlAuOWF6
eQRihv4VJhT+/qoppNSGo0ZhFtGSOm/6tBpascOBr3/aGMe1NAZ1BGMwMWIlN2sD
cYhpNAFBpEmbiBEb23yJYCcJ/GuYVju8zEaKx51Lxl4Bb9blslmYB6jFrR00nNYM
1U7e4+itbKqX+V6SNe6+8tN/G2hR8tkjY/oYn6Pi6ftnoOHbt3alPpC3lErJFxHx
ro36t178EfLVn7RM92Z/vUjGcMY2p6MqYhqc6T9xduMdUMzrGDnAY6tgbsFiGmG5
tIvDCsGXs6Y8Mky96Ec8hqIU/bQR65xqz8ssmqli4Tgijw1lXgk3uqJEUyE7CZI4
NNQxWNOHE6t5pN/VsB2mL309WDbk8KW7IpQ4Eu5slHiNS16l+RQ6TyJQoDI5e9Ex
r/ysH54ngt6/PfYjjKLW9io83r3N/gsALx6jaETh91DIrSi29W2vVwzEl34Mhh2B
sweW84LQHVDav9KGOoH54QKWZXpqNYU6iXdfpmrhdLXa2u1PoAUQSiNz5+CB8tDL
OjPar7SUxhdOgZQtpvLOTiL0xEk4XJ1dcDiJtZUpWMC6oOu0SFJbYACHohd4PstL
v7cdqE+Xz+j1oKEuMQKRqDGXfQfI+uXNjy7LaCYExQaCLztGeeRKHHifxZf66cAN
ix5Ijh6Oe5y4aUUEc9d8+ERWu0iV4eiwG4DuNiEqXicTRnhIaF2U3DKFaiHoOmXW
CiuNT4aqb/DlOyXNadrGeC/RZ3BiBsjJkCeakFUZ1iMTuPoPIAbYncn7gfLF/NcS
lkaVt70VZrhAgGsgHrXS2iwYygtRAGZjQCG08VVu2Jq8MXvCTnJAxmbfhh4zlqv8
0WQXnws8HsSRtaaHCmHEjOpKkqLDxQQ2msgWW4Wo9CbdpCWF3HXNQo2kzVRxb3MN
CC26YBqkeisoT6asyNnCLu7oHmqpQoxkO6V4r1uSHARDV7ztLXTLCw7uT7sJjmPA
NFrxGE54TVc81dylrSnhRAyAz3FqvSu393UcO9ih90Dn9fZnGO2G1rh2+pXorf1p
7qgGpQgnKtZWU9mInjiQrIHnhUiNv97aHA21uyyTpC+MUntJu8YJAGHRtSB+XqSC
sPEhFMEG0JmCz5vjZO0jUc9wEugzOEKmixsXpJ+Or4epb+mbyLkKt5hc+zTQe7Ko
5ZylLv74wBhUyvcC1BttShEena87miLwYdRzpg7x5q/9MtC5aK4KxTJfzufj0lXB
+7QZdorMgeZEVv10lbpPK7dFHAmkfcFswikfb154w4tsxEz+ZVujh9F3bmemdZ5A
5glD9Swq9t26pmN4QDHt86WKdwBZroNGmcQ6m7Tgsn/aEOVEAaKvKdNX0SWzQXmh
WX6hMiZK6/hZpM99Cuyqk/omDj2sNYWYhbMv2cPZF8T7HeOp/mE5n8Ad8Wu2aQ7T
aL9AW/oZktO3B27JHob7usQte6s68CIBsBbVz87DNQuQRZ0utGHbptXQe5R9qjRz
5sDaP+BR5aQmC5uBj/D99r1NmNubhhqtas0cc76r4YOp/VlPzTGKUAEhLtLl2Y42
uUyBb/Ec22MASt8nVURReQE+a8ogqbo4GHpqnFAVBGkjoArPsflY1e3qinUfGgl1
6Y4nRbwZIMZX1LtrzNNYl7sLlo/Lidkzcqv9CnrtkXfIV2MIsqnF6hyVBU40i3J4
b5KQCbrPJ0KY1vtgxQDWXhV8aIIJA7Tusj6GZ9rQZ2MZIvigW0jDYpR7BvNn7dfI
IOE7ZsMyJ/x+XX7IvbuN4OtHZoxVysh+jfLUUWOYHPZ8s6WkpmShE5Cb0emW9Eny
1aEyowsIw9zucJP1hzwJSRadY3o3aXnJi7yokK14mL+++OC7P/tWhDJxcaNWPGzB
rwM0kdoHroc5Yn3SFi7GbQkTCMF4yPjr3z/smdYAeuysWCaog/C+mNX/Rn8qrpdv
K8eHZu5DEKu3XlyuK1edn1JaSZ0XLduiVxI7UXJcV6O1oovq0tFwddoHM6Eeun9y
0kiR/e2Fn1QHa07HHR88pMMk/B0bB7xYJ0wX4SU4Xo9jocb2V73/TqBfFOkpEKIg
73VJkt9I2cTz/MikArHwaDtWYDr3oMmhp0dAXVR4X1qNxeEIkdvr78VLjKCEB/d+
ckEYRMCDTrH+hWlQpsvr0F+DvgV15oXpejX8NDMJp4i0e2RaIzFQuZe58igmRF/x
lNtGtgE/XaQBOW6m8336zut33tvczJspFcEXWs4ZGcL+hfWpY0mUn4Jj5EpkRMl3
/eMNeSYIokV1rGmQZLOWeLeSEjAaIYV1kWde/OxUyR6AJ762iLId2Ie4M3SERVoE
7vQZCZ4p9CxuaAoQBJ49e6zEi2AtMfmNJno2UF6AKa/81g5l4aqWGck+T3b2w+ZV
mUcjntXFWCrwbc+P1iwBWbFoRecUKbswd3VD5WOT13nblD7pflL+Q9jP4YvC+d67
L/lDyBkPTWc8lsKfHCVJA9Q4Dy0fFRrE7aGrgi6yrFmSsWG7FwZlp3+qM5jUINnu
keqQuW+xhoUtRvUOpotf2pSW1iVMuo+iSgxFcXreHrIkv9jfgxihcrBNO7Q6ZdmJ
ex8cjHN+vIivzrZyGLiVQr1oHN8jyxE4Xsh2H9ducyTUNb5C35HhEG+lS1MOK7dD
JJOdYYxmMakcW4p3AQUjSYcTSr6G14MskJjhuGNY2+Vy7JUbKwFM9Pa8qDxv0JVz
F73nRwxm5G8PpWjlnabJQzQs8/C5gbSBnuml7hM6JeJkCm04J5kS/d8fpiXTCYrl
HIiqeseXD/gyVsIu4p2lWsG8Z9WqIfNwIhIcY7QMo/1gS//suAV+N5illfCP5rIW
iFcku7JZUUWch/6v29Eq6PvIKYBt8Pq9Su2rHD2YWZSXEYlcnCExA03kOCYVwK66
3MfE6G0iLbZooAIA9f9GRSBf6ac5FoNz6pXYn1mL5+b6hRR5NN43HpLKBiIydSTx
0XS9PcB8C2dPYA6K++XK+llbWcsZCKIrObhVzfpNot/GwYrHACUYdfO8Clf5r7ws
VpxrBsSPYeyZeTUKKcljYZPYQaQ9neO0fDOxYWocgZYgDhw7Gvafg+FC5Q3TNdki
Z2b9CElTTRYfZKduXOfrVjZYRPhseKFlp0wUD5A6Wyy2TTjaJchWEq8SDjExvJqo
I2wLHvlNBG/Az3TpUpm8EhzVfu2P457agJkXtWtXoM28fdryjgDcmCqsXiyQ5YdC
JJoIMJrYXz5sgkcCkQK5py9Fkxi9cVELGW/DmnUXFznshvojuNlxnvGExJIpbcUV
/Ey5go0WGK7T8wR9dVZzVgO8SYV+3NkgMv3pK5p/4cD4XsnXYhFShqNl+Pasl/P5
IzoOCeg/hfx0J2xDXppFHmasSriPbsT8iFPwV7iG0UJx9ngfsQT0l/JvMTWo2spP
417b06qX7GHBoV7KtVkWAOIvsifQbqosyJUUn9VqjTODuLDeeRoIl0y/cj0pp/KL
4bPdAOiPGObMNew7uKMs8EgYSTfYr4OcX8etOVrCi6CHITCi1zQw/Q6ykFYtjpbe
On+XRNrVBLlvblpEpBdhRhyCCuq4EDVb7vkRjz17i3qVeUODcts9ZA0qfmVgQu6o
s0TY6BZiBOp48H74JFT6PNvKnHJddIghX2feevsLSZ3rJ+aBdRqWdYd2MBkwhhZ1
prRt2StjjYVsFReF0XJwZidTgZAlrbaQDoGCxJP9RdOM10vuMz6sNBmjL+hkpDg0
xWSMU4qatbpk7q+2FvW19hKzruSlgyhCWcrjzA5WQlJtQ4yt8fbkCibdPuyvqX+r
tsJlrSvsICs/HffHiBI4jOxW3zJcQTRlgszfSTt6/eRmnzInOpOJzwENf5VTRV6H
J5oPqLHhvWa6S86we9INz2ChyeLOOnFjXSlqCpwZXxgZEeMwpTu5PvWuHbjyDRge
zLyLkPK3H8FhJtgtUEdQ110Ylk551tifCc8XgDoctU2iGVZT5ONO7Nz0IuMl3YGe
xxcbhiORyK/83INmLfVFdONJASJC58B4IF//9k9JP5ZzFjykGiOeP1Ey//MnQ7ou
E8+ntDWf2rpn5WP5V6eGhM2hi8Z4wWOCX4ctODvjXa+FmAo1E1SrcFDmcZUeFELd
yyKr4Fmsyc/I22t7OfG+gfiXHoUTFP5+uZ7vIPjVmgxQIFvBeh1FpoiR01VzMyxi
47LAxdQf82E+sYbYA1h7u/nuvFFzDoXobl4IB1Fie+hnoA0sAfDm4Kt4SdKEYJs0
k3PfNrNXhfzCz9yDVGJ4IHxfrT2sd/qYZoegT7qAK3ASmGj7RIcwlFqGn8jrcb+m
BykI8CmtRqvmVcsASxxRFma4frKGFOWvkOeAjqz+Bfu6b2eIL5AT7d1ECUb+Q+Yq
v7wYZA4mFHrtqOAbjnUTVGW+hds2B1bGfEx54c+DlF9Zcphx5z5RwmcDrJIVfvoh
wtIMwlD8FF8AC9iACjdO/stWB/kFxwi278d6JARQWY8ZVnbAhJ4pNCFGe0t6gCKq
UHd4q9dC0H2Grwjl8XqunZNsPaxsUOazDzT3p6XVrxNlwrXB8R3XtBhA9bWj/sxs
ZFJlDXAmlrY93+u6EYhIVbVebe/RHnfRi3RnjC9a5OMmR14gOevvztvFRRJ9o86i
H9NNR6ihrZeF2UvhI4To1HESiytXCXczTWuuVRFE6wSzLaNGrTeteEeJgNoU2FbQ
LZI0aJaPk7RmP+ef5NCXbLRd9d8WnYNpW+/Nhc2WaqJS2MpNZiaMNcnUBK5wZt5g
nL9M4Zqiy6ZkLq1UG8ttV0FczVfyR+6w5B5O0iQIokHDfJS5cLuY3ezUxqY7RN4b
fZSJ1LlH7jlczTyoSIiOAug7YXOoEyoiYhnvAlP5tnPxZ9mMsaeJsBxE2z/geYLa
8UHIuo5evVFNnN3/YWtg3Tu1PbWbunZxGkH350JUnSmZA4vcZBy+8z74tAtiDYW5
xpUDrNX0gDtRKmL/YftpUfAC7MKMZ4vrGKWZh2IBqyZj9Fb8CknwaE80cu2S0F0w
gWj69TigmcqUM7z+qaya3ef0KHBN5KRE7rNiFxQkVmUAjAV4L4vt/J3T/DlmiOnD
cXlFNYBbqn0Yu8DCCglt+6NDCcEFZMMwOTsuOwWx7K0VlO3E8GW0NOXAjD6/c1Wt
oaIoBXDQM43qvBzrntDWdzNXXQVAzgNBislcZQfX+9M48flGWIx1nTKFqBjEAHon
wrYATqWGS1NHHptPHLJDDKCDkCZKhUTHw5tgVZcCDnc4VFKBygCwf7cH9cYt0eFn
PDefN9s+XCgHZi8DOmomXj9Z3o89JuckRIQCyIp/GIZU4GOxX59hJWdK7ItzgqFx
YRYSt/Kb/lL7DhIaEDUp4p5u9hr3MA8aIeiZfbKfc748Fr1jV6BA9yTIFIY+mltt
GcEAyP8IEpGajarfkeq096DC2mPgvPAFyuL41n7tIW0UizrlVHCJFFz5VhELx8y9
EF9OvblYmzND2hU96/VI7oSslzjaXqbzwtIQnZEBCc1XuSFmZfWseHyePtWGKFAv
we/Rz64LbTCjjbs79FcWZYRWjOaRQMVR5L4E+6+aQWxdw8zrFO06XyNu0+Jyv9j5
9JvZ93vWz8xXq0APFM3vObczgf/u/jjJsj0P+Zdwy20mmmluVsbEYtL5PyLI5QNS
ZYYOcLy9BNIOEQ+F1v5RgbbyTaa+96x7J0rDDyYZJ016HvXOBbzCSy4sq+0U03zK
3DSN+eHx9Wx0ZGMziau9aLZ1z1LLk9WCYgUZsk/fyR0qU/ME4gQ/y/jOHnO0HuRj
pmll+QXSme9KCYPu28oMgUFi720N9UAqXZI9gupuXaprum4sfwxh1Hp2+S8CpObm
iOAeGoTHMJJXesqzTp3FQZwa5/ZfRcnpgSNRCEZ2zryzZ/65MotvCGWGowuTYO6l
uyrBpREKRkxAf7T1eRw1YpD2W6BU7FJ9zWcAWdUEjw7VOeXag8M5vQopeltrJRDF
KahsWwva3R3EsSksMs0MIwRUZcQWA1Srw1WJbIX4jxE0PNf0osDPtXyZpLhr+u7P
zdlghC7eMMFcYMsutnzWA7yzmpcesAuDpO22W3ZxcXchZdz2/CvkNr2Obmifp7qb
V+SfRipMKN46d1PegOnWALLdoHQjtKvoB5ciHE5B5Slynt46p3zs89UbmR7JuDiR
wFIB8xnEhkIzpko1MKVk/9zB5rYKpArwROs25Katy/qIfg7sWJEbS6mg7pXMyrjA
3MXlVlWbnHp/CHSKC9RuPWsJ49cFXiZNCKjVN8df3AKn/cpTygxc3Pu+nOj8h+S3
nXd8tLrBerMURrALLY3LhfIzFWsaWElEjhiW3jUnsCxanWkxxEL1KQfdlukihtRz
azUC3rWzUgQVVKzbBfbUy6uOYXIfUtg9EeUn/PRR2rZ0TdwFjIDvVpW5YGkyDszY
swn7U5UMo3eobAVTjrKYsoOdcNugkbj4qy9uqD1CCoRxO0Gh5UNvL3vVi15iLfQP
k+kVv3z/uLyhUA7uYIifs1JqwFCsHe77LiRbAA/TkvML5OokUsv1lgQEviFAg0aU
C3wQjqCD+bCTks2L6vE9KSd7Aosl8/OgU2b+2eNhb7X+KtEz8oasE1eq3gbUxAd7
k4bikkPhc/4h3LZGJxBwuW4blq+dt/SfvyziAYM8UNAKeGDedxNhTAeD5xY4EWLL
AiL3tqVGpwrKZ1MLhGXmYerXIuMkQDAOKkW02TJxvoTtUF/aKT54CfjO3NtqLjwW
eE5fsGUjXq5adgo4MRYAKchrGM6P1Tf0RLrDy7/irCWA16+5tKtTg1WYABIZjhcO
qHWLhwT9bikaXqarsVfNm8hR4OTz5buml11bXXAbgJ8GB5Lenskc64rOHK9EUJOM
PlQNALAa/tcrfcS7ZGfL8wb/Z0TsQXLjDsKlcrKSwORof619VePrAIfAa3/PViXX
52hOUfvbtMvTZxNRtRzW8nbTDHbzg1+w/EC+LKwH88Adxm4L47+3bqodjgMIaP58
US9vp0slxZWPr/8Z+baTZRMzAfokRp/4ed7OFicbkBfTP4KHxi7ldU2v5l5azhol
blAXzGQYkJVZBSvuHc/pR89Bw2i80e6uVlfAmp6bPDhuuB3edaJGy+ATAXOGA2gp
xE7wJaJN6n/qfanzkrHA/E5Ry2uH0sRh7IErG5yWKNJ+AenKC0qeG1ISD/bXQW+N
D+1QK4Ja8QE96kMOv7Tvqu1aeKL3358OulkjI6TwcDRhLRSlZRcm5srAoA+zytfo
CrA8mHFaS8qWo5g32AyC/LUdeGWylQ5Q0wh0PtH6LuJfhgTrMVzf7fJxO3j2YKGS
MkL+6E+LMaaBi92S3Kc9eChdeLct2XbP8jS2j6GIo75HfsqrWjw48SWAMo19Sj8e
/HEWMHo1Z7R1W4D1My4MtzHRLQiVNHVmq95AhHLLH+xAiJO1vHgYq1M56YZA99yt
4YTuSMv3Z6eWmOMxzP2n3ii/gTRRYONXqBP4aH4aM9A81HRDDlGqHdruag959JPr
8a2ev+3qdEJ+jsj8RKJJ2//pDF0dxMjjHCGhx2hYspACxZiXeDIYR/hJGoClBtDT
j3Kuk4tk7FhFYLhaN3w7Fl5L7OwMaj//2cO5AO3z9X/mQQgF0PB059g/v5P1uUZm
HiZ/DztyH7M5htjsURC08ufhxfNvmLjSL0FNknyI9xt+I4Nekpr5szhsVazoJRMz
lg9pyHCae9/NBzuPJrZeAenWLpC1bssmLjN0606EWscY7NF1ClChY5cSRb02IKSh
aBBrzZJLYg35lDjHQj7eNE4vWeVZgiObjwQJ8rlEczQhJx1NwFwwkvptLZKtID2P
W9Eo6SDyjICr81Nzp8QjvP5yEXHGkxn6dKXuhM7qRjS7ZKhYva4DAxN9b3Bna15Q
PzXML4FHtZtuyfDygx/CT7Am20FH/ExqKxLNF7EUTSnLi0+Kjjhw4XnlOO64yD7M
/0ktCmB02kklxDJZVQyQjjU9rXg2rNXH2IiOSXDqpu2u61+mh5OukY6deRAEiMzl
QvYMGDFfVGV1XvAUF0ymvjGaTU0m9b/DAl6rY4YIWxLXNo7hhClVzmScED+swRif
4Uo6GOrDRWMG3eQHhvi+McIOLXnWRDnvRIaEgrIue9pv8t7pOBWg4KvaoyqlMI9x
PA5Q9sLNJE1y7ojT8G5OanWHTAzKhPkRKOIcIBPZ3crIvGSWngl9iM3oW0LBZyhR
9g4jMfEh2IV4dkweAcNxPPH51/8HSGE6a+90mYkn1xIBNADEHa+GKSClL7CT+gGs
t6yO7VQsUTaX0S3kp/1gDkFjjbmGiatyleQrq82IwwJ2jIU3CanKJJ3W9sg/cWG/
p5wEvWwAXJYLK8RTDE8mXVuMEVNZUaka3i4S7OtlVC+Y0rwhcTtTWkdgtxladYfy
Z8tbJ5MYCazUaSBtw7sT3XM5+otiNQwpo8nx9GKSNICCWAltO1M0u/HQCuyiG4Ub
cVfzPCb9kADPlo7Y1yNaeMzqI8T21bKAC7vsAwTTHLIYcCktAairGGOvFAcVCabs
ewYt3XsrXB++Dm6xmRKWGgb+twms5A6XfKLIw+tNZNGL/mrsyYn9XpyBhCoJ/9Z3
jVFTU2z4ZRlj4zik8akhYxVlNHW8hLS7Vvoeg2DJpHjx3jkfbnCKQdbBSdvysK2O
EvLl5rA7m9INGOIe6YfzIsdw8J5Z1XOf64I2p9OqlTL6kyPcBuIpbZL8WocPmm0A
PEP3D2f8xVKhNtuG6FlnSv2JRrL9wzH5rmI5lUdbINIHjBoQ45vk1tI5ihBl9K+3
OrsM22QcVuLQTaHxEUiMWfxJR2YD20WCrCR3m/8WL0qVNYU/C7gqmii+GmzxISl4
AcUtuRardYvuzFyGaGQSqqk2Ho5e+w71j/5/x01ivIr7LazCTR05ci8GLQqPild6
vayk0jwIJQeXJi7873Rhag7Vml9O3n+xPFOHtFzijScJXFA+xK9tZe6RkX2ZxtpK
0ks2+odqW6pkQPCtR6u9P5YBA+3qC2kKKD3VfXa5aqhmEsKGe19ASGrExmrazGl6
y1wCVhGLx7b398sX8QjkYS7Ws3SEG/pWLYgVDXnrtQ+xrsI+ye428irg5YrDKnV6
d14O7pl4acJr4AoV3SfsV7nIHVskF484hvtg7S4G2LWKWG1nn782RAFz86Yy8qdR
X4Zx57zbiyfyBfNoH4wZm28NosqAPS8K7xw0J5+vwUMqMQ+oHxntZ4xULbBbCWb4
zx6ZNKRvNocJygbTp/cP0FvF96pnAs/n0HKLFBIUGJmFpjCyh6fJhmWr1ZnS9fRt
8DHuj6v28I020QPrSms/YaIJT57uVwUKZ6OJBgeTrKChN4BFsO1xfwtiDWvS3ClH
vOp6Y5dA7K+vEU8JesO3eoezyDvWdPaZf35yHvpKxcsaws3KEhP8zbjy01gdx0B3
dEQ7Z3iwMrt7GAkda3QPIYgZmwvi36DFdnwjwjV2HC4psS3Qx5iWnyVfU5L6j/Da
sG+vHVplCIMWnzQZKl9K8QcYCkuHN9ePiLO3JSv6O3zCqbNhYXOI8tjFta14k2GS
Xq/Jdi8Gnc4GoLpuKBDHIJ0pqlTm+htw7jFaqRk+OvYvO1aL7zQjgE2tEwdHfdnu
+1iEc8O42cK0ibK80EbnNhV1fTHtk84Q4HIL+zRfEXRginCcgb9/bsyrnLZmx4ZN
GlMRfhTkjQ1gq3dt2E7wkrdACzHqev3DRgrYawpC5Qd9epYGrt36jswfe9n1MirR
YA5f1G0YMZSI0Ze6jj6B05vYjepClQm0h5FQ1aU9BHHXf2oekJ0Bxm6+FPSksoy9
+rfeaMaOUgEYw+C/J2/3VBhHi8Joq2y8xyEkMQjtEIt62b9kXbd/mTw7xxUrSZAV
1iyFFEd0uAAS5c5HQgEanYjgc3u+yGvky3x753jZKAMN1oREtDrCC457Z+LRoHV3
0WZUthpT/aXsaB1EWI3WKOiFxQxAesi4aAoYbuOEPxr1srYxTHgoqi7d8vbIWCGk
gE0DRcU7fPp7ble//s1V4f4l2nkU7cmNFaQeQzPZsrTlX3uWTClM7aF1Pdh7xHVM
Jg+i/Qfwj9rjuX9cZR48C0o4CYjJHxpLvJwONpqjP5miVvnFd9LZH8Y60INwBovI
gYFIuPR8ziqMV0boT296oZyS9jYjJy+MuBh8UR+qY26JBYmgOUzof/7ZZ0rsJ6F9
OWKvDRpowdTrX8HOeerogwTaX0YQnkR/UUox8j3m4v0ZnYBc1JfNzzgfXJ7lye2b
ZYMfWIQBY+WR+KwEU8aN0jV5Q00Bp9FFIRKzAtJtaWDnDlqFq6vt5nRZdFW32Crh
bU5QS2FMmyd4zTjxoBZYbPcGtQnhyxEdwVJN219M5fLyZII3HOglfd/gYrfGc9ir
z9rpW+Dxb435rQUXVic/B59g+a3Q2Fs+Smt18ZnA2elrSOR87UAJZHFVQ8tZySTU
z57Rsn0SH1VJYt2gBmxQFLveLmKo4TcBK1HBpN5SxWL4nggKNu6eTbQEInp7A9BB
UPqvOcgBVly0rnm8U1LxwjDBgmF6vStWvkxMcJT+XtXijqgiq5mDXyJk+Kp1KQXB
bHIJOMepPPpsWxgaPY6VHMRFVL9kyqYWZdZ+q+cPSIvePb3RSPYlzxFGmEHm8+00
09AWIGDtjEdRsX7Wf9DkFSaSmVyNlWLoVyPTh5strwhgjYcSqL1qb8FexljMsM5A
JX9ImS81P3Wyr32xLuCFg2n+hPv5u+wGWOZho3HIF41+5gNrVOFif2hTDdZZPfWY
LVFmyQnKDOBlwxaxXR64j5Nn5mgdXNIZol+qm5EnGjvu5wzeYs6RGLVHGyg06xdu
cU38O8NqXH5qGvmmbqU3cNLIscsXrSYiVcFGNVP7bjUvhqqOrg4Yv+MffOKpzxBe
rBrdkoQvxWgNajQOlEEl80/9SBbp8swHtww+WplYOMfQ5sXa8XbER770fEO5QU9w
1v23iCQ/bGFWUAa4VzrcrtrMmQVHeZT2L2sWetN5zggaI5m2gL9WhVHDAqXyp37c
azd+swCrgF4iK1Ne2AoAYNTD/tGZ61z8cvu8cjalFFUATD8YfwPvm8q63aH/16qM
aOJ0EGjrngD1x+81aYJNITFYEMDaOubgyXLNja5DT3wwKwk13zdBQx/tYo8+E8YZ
XjnKBYQXs42KjuNnF6tYS2D/H3jLFH2s8EGgtNoNfBgvauhPVldG9LWs/RcfWFNv
aaL2I+YoiUUZQiU+ag0414+EcnUFCEszXHJVln3J90zq3ZoaN13U6oizoGhpEJki
AJO+vn6yxqJU0HqsN/ELEQAbtHErGyYk3SuRuRGNLyVhEEU8enCEUU72oOoFJfSl
MgvGaVZIZj4wW6kbEk02o1dovO4yh5ihGa23gWizpbka4ceGg6Cn2x46uNc1XV93
wYtUWewNhfOouY+4kG9tke152r4c9ZDeKSUaqXwpsXi7dFDupYATzMEF0jKX2G/p
reCX3FqjaQpLtEZ3buf+Frb0AjawOUpqeFIwtN1DICdGPiFNI4neF5+3GtUMqe4a
S9BsLAM5tmYjfZxM2vTv9CPDkDwkOZWcsG6oHk5pGVl9aAoBg20Vn/5BSlnbL1BU
bn7eaUj/HUfLnVY0TxM/ECmf1s27lEC1JXGCekEp7rai0YwC798h/LMY9lXBRJIG
Bvf6RE0zsqh8PN6KE0yMNeX70E2Sk//FkgqmGxnAzTyJQUfyNuSmpv4yzUfb9wns
DKpvbEX5FxmYgoIz1sXp3m2IrnGs9DUeXS/4GQ1z4kiRQCwCK+kludze5OPdV2as
pKmnns/y0ovE2iiNN/M64OZe2zbuoFr3kWNJpcY4QxLtw2JfXQmqTqcmYmpSZOFh
HT20GcyjHknZElDdmKpcwzHWufk+2CAr64bX1NmmCgzeeo5pq38tGj5rhxN8lqX4
KvDYOwDqNcf7xX3qnzxXI02ZMunYDs7zZrEH7nUmoMwaPSYnGpEL75MSGB8sdm9Y
NpPNBDtOJ3huW1yQz96rixeKUGv4/KpIVD+ssTu1CI2Fowh5yq0nSwRSKnAoFaVR
L9N+fZ3au2jfHvKKmRJikoZJGWAucqW5SbBHceA2Rqmd/ksPpvLUrZuHijTifwy6
nB7cQ/skBy7sDkwB5qIOsQHECnCWSzFvSDCHGLLPOJa2pgWxUW2lLjxnQ+JkasKv
NR2syPGOx/onKqjdJXG+SwXjxtTnlmbiatuUXzi6NL5SvH5AN5MXDLPSxN2JS82B
AnMU83WQCNJVypOQaGPJFodevw0ZNSta4NSRlV6L9hKiVmZwle59z0/UWtevI/hW
kEybuK6RKnl6wwO/OlRgCwnNp0mLuHwCF0+LA00E2zETyRgwjPOqP2NE7nbDTD0E
HoxMFGnL66M2TZogJcJ6+2rfyFSUo9g/0dUDgxh85A+ELFHMIKHjs5Jy0qTYGFK3
PVTBEg2kJCu/oy7qDAMjEJLR+XLklgjiEIXHd9Y4Cxwvs8Au7L+DpBbTMcwl6WIR
S8xq/2FwtQZYsaWxBVXOZdtPvrzIsNEyEr1Lc89rQBnlop8fFn33N8FO80g5MMZ9
gu1EOz3lEfELAsTf5TlGz9UtGiEHm9z5KVPa2HP04YQ+maPalWQ8Xo92uF4H7Mwe
9ZmELn+4b36BQ335Z1nra9O0EL70vrB/Un0QwugX/E6pKGGkYw4naoFYOHTw0ldY
0ObCMNpR0C7yBu4/vwkLgP8jdFEDS9c73Aa48eQaPs/zgTfIkoZCqXRLsGrY76j8
wu17rMlhtHAZL+bI0p1mmg5Blgch/JbynwXKjYy7PxkAEeLvtsNgZLBMNuyrx/G2
xMN9tCRvdQPXKqfP/G4vxjJY12WQQ9oF9Yp3AJbX1P3X2JyOnXVDLWw1VgUmqiBc
8Vct9X6QMX88c4uyvaDj3D46zXsyKGMskAteUBs5RcA6UOZ+JeLp9eyeUwAxsMDh
ElAYtSDGv1pr+Hh4n8lgws7sMuELkQrlHviaa6xgOAMVK99dxfBGFwZw4vzhWoeU
MIP7nbzAt9QhpErjGbrykC2RXzblcnSihRgMq5afRWGsi85tCiDa3FAcM78YwYdT
phssHIy9nHcXsa3E2jnWb0cNguH13BHm9xGkB8L8ki7Eu/kegNbt0v7/blTQlG5v
NnoFP5OvN+7C5Pt5Gw6No3jI3MDH+1y9OWqXKmjueLjqJQW4KoPMlfuHi+jCxsFv
1Rr82l5H1O+u36q3eWSh1YDk4IdMJTTg1w4wv8bkmaSRSudJUe0p4YGBEFPDSYzY
Qj2I5534g+qtBHZcBPwe4fkHow5+hhmxBDj8JV6RbeOC0DZK6JiPHcKHMFEo04Y6
aB9XgkauZj3ZWgWrW9lelOXABBqDVH3bn42z7MWlVaixuXkFaoKdFSjb8R40zm3w
01QrntKRr2jSsoPAGRAObONHzh7aM9yiaycbp0PRf+25RjzAaK2pq4E85j7Bpg0g
T0RTOyvoquGMhKGy6tFBwdcNDqlW0CC+ib//cED39gPUShLM61/d1EegK8m+Orno
A5wC19SmolV+NZDkMNWI+3hUIUNGd8ooHzK6X+nbJLGV8OZRxL3Id7mEArTRu/V+
PG8dn5QyhXmdqIzxZ1hgAPIkzZMwoNDsOkaXnOQd0kLXDtz7sUUehAGSzJzXwex1
QQAm1UU5q2+YrMiz3q20cmxHkhJxUWu/dJLHQ2m+ijaLhcqILwrqXdOREcC7OfJD
6u117oLMY1/8gG6W7aofJ91bD2AQfpenjrHuBfK4yA1LA4fsVo++CWAFwXAzWWjr
/SE/E6zQtwEOeNtM+X3xpIQJkY+Vxh28DIQGwP0O4OtYa3pkMf6i8GBad7jXM2j7
8RKOBWWAsLyaOl3XqzEMbke9RMDDT+7bYZKUagrCxcwgqnyBddGvAuYgodz3SmJk
nY7aRJ3g7t7YUY7zkdJOH3+gqP+7m2a7y0fLbyMuGvruybv87hBJG3uV9Pse+4gh
o51h6ZZ0HKaW8/MvK+cB45MqnQnewKfi0rZhG8UWsmjXnvO1BZlSDYAJL3C/Q5YE
0HKVVBCEDmrtH3unYnUO+C+RlcdcSExTD7Kk2Cv5YnW03ixj05vMgqmabhxBKa2/
7jGcmPIugPU0Kg2FdlBPheXNKGCrxV/J0YAFPiS8hJ+IQbtTXVThqFiqTpa8kr3s
M8yeGjvIrnhYXNf99TBWSSKPv63RdMFjCwVIQzjm7z4F2SL8H7ptPxtyV63H55zz
GQwyQov0ApxAkknJxIB+cENlYT+z02/o4kx3ZieJelGBn50iv/3j2tJ7Fba10oD3
STk55uI02YdD10tbOZbzuqERh0BELNKnTHv0U3Hl99dAjit/wn3QrflEiQ4ZZBJO
NUgOsALNRKeWxcC/Bqb7NQ/8pfZbWUw2KgwQVE04nZuz8lVq8Sk2OeiU7lq//PjZ
YvWCkB1sW+yacw3mLEvf7M0x3c3OxPPshpyo8PaSAYbUhF2r1MiBjIA6D4qXblL+
P7MgVUldbocZqSGXfWaIW9I2+cLXUQRV3rCokL8HZEXHQVf37eauT9mKHZ88GqfW
HwQbyAodVJukoW+uM+INJxBHCriEtEbbwDgBC3Fn1rl/YdGXgLb3SPL1fiX7FxMU
YnNY6LhHi/RvpzQxm/xq5ssIzLLF848t7swx8Zw3fSMBsTIqB/cV6O8QbWMkzt8P
A1YkU0vAnHt1FTSuxDw8iXZOH+bpNYiANm2QfiVbJFMihlcG0nxbfQUssIJHYT0j
AFKM+9cbYpUayiNMoXzHHkpSIMbpQHJkLfa/3GJSTKXYC79w2cmFybRHMTYedltD
`protect end_protected
