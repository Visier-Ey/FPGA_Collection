-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "N-2017.12-SP2-4 -- Oct 23, 2018"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
MIODzXUXbBjgVLiAHUU+TKH92Dqa2bRE8APMNG9m+z8PTqQHX9Fc0wYVzodkT4HR
Op3xKpuYBUOmjTmg/OlKi6UKIFTG8zrwCa+ST2R3vNbrLxUWSzZ+8Ae9Q4mKs4we
L29XA5XAOMJDKvXbtobqYGsHc5pFAJgbEccQPv5tlkY=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 34720)
`protect data_block
jydBcD2bDXNd6z1CoqJ9e30kCcnXekT8OGYFKRGr+i/zskx7ecFeUbxczf4I7LAC
2WLTXrNCskwmmfn0FhtDXhWRRw5wMQp1quIvabJLHDdxp8Szd1a9Y56VbCXVg+he
PjScbm53pvSzEmwHZLs6+e5PY4MWHwWIIS77Fdre5k0dyHG+j6z+swCAzNXwq25j
qVsqCvj+cmKAi5SwRfmKxfVZPNieqL2mTfJysCuqKs24NOEcIUAjlpnDr4e9qBQQ
feT8BwlCizGJ1KnlGo8bNa0OuOOEoCWBHQyUTw+uygUgJExIHwBLDiyI+yfwDJQO
dTsghLUZjRVEVLLYoEStP4+CEiveanVJlxyrtcs/5knwDfY7RysH50uEXhQq9Oc2
oxgyWiuwfm/UsIvVMWHAj6O9PMNbmkvxTuyhOG3g8j5VComkDLI0MgV7rVTAu/5y
ySVEDhruE17Kysc/xqZi4jTJrnauu19No6lcZbSPRsRoatjLxKoesVkmwC6OEwRT
sXvjMXk9dWAWTskPMMk2Wn/4lTpvC3h4YkBsJZjMwZkW68NTLcu0An8ftqpaL4L1
PTHWiVS7BoAavC1Bs2l63jtqexb8tlzJWcSVYo0m2YUjMA2ijldk0bw44AkXFuZK
OiNETcjW6ai3VHsuPOC3EpzZmxsj0ffTAnqmfuSxFadZOmFmQuyTS7WQwA5FCIC1
KeNPZsvzsf7ap+8ybROxbv9aP/OnPdXASsEmzf5GuiyHfFUF1OCVTWO71D09StXN
PXiov/qH3dJLJ/TGAeRizqPNR8UcB3/ZptOhUf+eyuVMUd176tbgW8aWbCCPUc/r
FK0c4zC8eFBepPPz6B/zWOW2/vtHDdkpJga6WWeHMBGlWaBaRva6/W2t8UWxqvMf
8lQ+YA6zI/D3bBw9QgxSb2YshK5uc0QcHTGJLBo+CNnMnrSjFTEqS+C8o95Zju7G
STvY8wf2UhEQ06ADsgHwRpjxZ6M5PpvN8MTQjRt53V5+i3WslcsYw/IbY2A6zJ5Q
Gn3jhbodGDSHLvT0cbcvyVELvyMt/1fbGTXh1zTmBvQTNTDTLvZCxRCZ2dLcT4CA
W+jLx4kSgsKChUqHa8LT0wNn7mz3tzed01nmxLJWbkjjLeG3XU9WdVZ9IaEnQw7a
JEuwVBFdZmg1VhJPm6DhRD6sKE6pkwdbwXGGMrQe5evr7whnMQC7emzTDMLDxO5O
D/AMzMU0VOOCcn1+sIO9XDodwCha/hyleqsX5ts4dDLxlwHIOHDDswZ+V2WZksEZ
6W9iznM7DMQ0ARVWvdxxRDkU82ooBmPMY+T8UjxYno99RBSMau3z+Lm+2nNLHD5V
4LHMcb1CaP9QqSt3I0vXBDwE+8mQM9DMLiq/tRiAuFddqpcjVXsWXJ1b4hYxuYkN
3YWH656pZknNOUF1/UOhgmo4mjqbenxQywdlU1E34CxkSSOfb3eTpt5mdmwfgVJs
OZf4fOvCZ+XK7dGJHks9DblzpWhIlhBHGv6o9Nz7r2edmJgikz6YXSgZ8Lc8s6c2
NMB1Pg0KTcNAqCgGGaCjG2QZa7QfLHeqOfPISbo1yQTkBVxpxAgy4Zl++TcJEsUH
Uv+cBL2Pr8H1DT7nEiTALIXb+zdTLLfiieKKPXJEmMAgus8lyU3Ra3HorNl/UMXZ
Ki5CVkQkKdntepMv8Uyrqe5b+zgNxC0GyAF9SSmKsFp76HMHQLOPJbpRqPpbWrnt
jjztoBg4NwtKnPhil1sev8FBsBzGIOH2Au84mcyoZydrY+o7qf6eaa4KzbWcVymq
lkNgSm1XS0/4GSJosS1fg8bG8RZ0bOjW+kTDnDkShLihnaWk5Eev7GVy2ZnniJ2u
tqqMXKq1ETO41XoMjQOOLZHz7Kr1k2kKaluqO9eKZVNt8fVZCug/TMSxe4fyt4V3
WtA+rDqjzYVsWD0XuG23ikt33ZC1Av+GRc5Rlelqdc0r2AE8f0f8pgVP8KnUC74r
3PmPtEEkLvWhwY7YkVOULs8biEty+8xDPrEuL3Px5wnMMXKT+U7qABrGxA59Y3Ay
CijQoBQ7kESP0oRm368OZG02RDfCcdtLoJoNjgw2/DIdFHU2C/SGP6dE0fTtgTCM
ec079zUTDPhkjENV3kFlJvvjd+0J1jr+y/SM9jxzUVXDFZPwJQ2MEgmyOg8agspZ
v7C+oA4UJjEZR1vr0/IwDSTma0AwLvxqLuJoDmTT39G0lFmI39TRXFecU1RAtUD8
Tg/RIRbneaJNJ5f4j+9v1yW7MtEFxT+a/er6YH1Z3/IaxSCPfCmrnL6p1jhvxd5m
zsjf9eWp7PYRabgFQTrt178dP+xsHk3MUhqz1fIu6aOz/8IB4an6mMB2beU9s0uv
/c71cK2XNiwI/SXAA9bl1U5yN/F8yPlJUEkxrQLw+gY2HEhpPT2V0LNTNa1J5dDT
qTfQUe6nZ3Q3tgtblrZwzPtuIb6yO1mvxNRHMy4I8rUZbrP9j7h+wt/SIsMXaHsS
PprrfhCf9ejh58zvCWUHuF7Qj0EkZajjqMKcfAMVhG2MrnX+cv5dq+wOdFwL9Sm4
SIgeRkQ9na6zhWVdMauvGIPOTT/KATOvEKAGJfBY2Ne7KhdUByWjZ6M8OzneJ+B5
lcYJjjlmetL7/umptYiFWcHl1k0Lnv1zDw9d9Go67zdjg7HARfvK6CZyyMpEYT5c
+kn6ral5hLh6ZjTSuNAKRzbUeFSvbFG0/oVs720CrNX/R3vk52xPWO/jeyY9k/86
j1ugXJiuXljcGOSM4ms4Z7JTVJFh9Fz+q2MK1bXMIQtzyGUi34NjEQCJF74Ta44T
p8KS1O1Q2Jjw7pcc7DlDQHdDLfg0wDC1mb1cKjoxs8GaweBEMzFgH5j9g67tHarc
79Jm2RdCP6kRRplDS0uIReWEfdIksnMAQGgJYDxLjL0q+xGYHPZBRBEOcx9wqfDt
0ZEwF2A+1wYuvKGSVbbRoasFrLxvvK4SRPu91wqlhXuXmJEDxYFYDr73VNTfGpQv
McV/5cs6pl/TKDz4Glmgon9GbUqfa4rCvdVVAnqpKk6YKim+kYBu0Zm/9hw+PYu0
DmXp35gNAtEu1SO6+cwz1efWtrwZncXXQKRvW2tbx/83nQEIn6TirvAoMbzAWnI1
Kj3XdOQKWtBij8pYXFzxr6iwDte/FzK6DFX3SwsSjTn5AtI6kzO3g55xbX01Q2+j
RBfsMexqHlEDIdCneTsyeRCCQQCEI3CTKYG7zmBFXQnX8aEgA9Xd4ScRRLhuVQx8
0HcGyOfO6Wxwxssv3njiOui43x/VIzIinDwkXPhF5MkfdTxKvlQ+JUV61LGBOXqU
IWQVhI8hk3Z2lcegDw2GDyT32vBI9DN4UExlu8urOLI15dGOZsjrVrPri4i6sKST
tC0Tb1zelAwEF9VcYfD5wG46tlO2Cp3TzOoFbDSS9YdM3p2Qon5ZXF8zraMkU3D/
uqwqUfP6BqxZboiScU47msP2CVApCGFpXbg3r9KiJR3jlbbpcFps+/dn54JfXREe
6G3Y9ekF9FSeB2U/qQmVsIpu2AISnF69gczLP89mVaLBMrHEiAGEehtMUX2iprJ8
rkIjO4Z08W3/HBttxIz0ukuVHlJbVcIx8rYw/KCwmLerSYur+HRRSmu61v3BRfE/
3gcFk5q+w8YRFDcJFLNK5Q98eW3WOG59r/eh2KjeLzgrSTiJ5/EBPtrGlL0uhyto
21J5fhMJOaOOa+hARFJmbTH6Mr/znytjeAEK37bDLzARPaVwyzKZpBwOx6LgGz07
s/tTghgKnL2UFw8uRl844U+VvBVB6zIwWTfIOGkS1HuhfJwdCuu5tbYhkL6xo7Be
XuC1PJDFaPYMLyGhqiy/FQV5RZ8evsuMMRQTDJgL5h3o/mqmqFkc2qAeINz2GaXY
E/Mra/DgYhA8Vcy+SGG/LS9E1ZA2sTM5lOtcVF6O297DDCgvlpy2tUFI+W6fCW8C
NagQp/nuQLATMpDrdAJny54FJAGuTvJ5LG6UbGtBrGlhtk98BdqmEL3+NuWuh8Dm
KvqBJBDLPQKe65TwmkdbJ1y8DKOGoMZiKv2qkpFzgJTYdAmaSwqEsegsdFoLV/HP
PVS2ojByikC3v45H0qEtCeBYV/QS4byT6BN9CZ3nZWOtk36pviR4N3Utp8XYxO4/
YcGlAAmdXqA87v65SctuL4D7qxjfot3EUjZGwJztmzaPMJGoSlqnp4Xzp+vYeyBV
lMVF8oK7Abor5+TCQZxO6F0896oTk8/RllTocBMkW4wqsST2R4RItaOLsOQ66myf
jtcsauMg9SRNLL6uxKOr/T1g/PEfC+j6Riw9Kx2b080Cj2uUotHaT8JuVGVwLV8G
WwFBY72pMz+2qb66dp3pO7I2HZhYfUtr7P5piryu7URZ/hxNiB6WSSW9uX1KzpS8
tS0UAeszsChU88GzPN2gkdlZi5jt9e/nI4dFAEzo1BPxLRMBpBShrU1wdoKBSRpX
29wZxPUll8KHEuBE3O/1+BkCK0OcxNp9wU9Dl8o8QsCTryDhkL5WM5SiUzQ13zSS
dtfAtfMEaTTy5GeEIEGuxJ+Ug1zpsmhAfD0sn4ZOQZvvB87ixczSqy8ySwYg27AE
9fagkP0iurCTUL1CJjM0CPzLmw2LgHmd9fxBWrXP1IPlGScNiWGj+xkdidlrxSiD
ro3GeVOj/AxrYk82hwrqGaa1TpUpuM9bjcCM0PMhpmflEUcZVgtLJyOP5rqYQAGc
gohyGQSv5m6i/dpauKuVtAG0awRBZPW9UaYm50mLixwzgnsXRRVBbzaiaoHSFqkl
zNnhg8GzggKnqpUCi6U4ze0aPEnvysa1Ah3mO2fb3felutt9Xceh/rBP5fC51C1F
eSH+/S04k/dVIqLwd1vAj2X4jkZQuQI22veF9G/cBqtnoS0XT7gmHkhPCvIUiZmN
fbnG/BtSSDb7PqpfDviJsmTAFAP/AK1hAjiZkgGJ6MwWweorxFSwF6ZjEbVgURXC
kvDkMizO61bQOsjuYSK17y4KikRTOsSBiULOGioNlG3QNv0lDst28z+pNprrjdE2
HGOYNJFnpa/ar6wXM/tHsBU/D650GYILcdSGMDfNpO2xdgHluo1UTZ1aN+vUmWW9
T5a7S+8LGHS9GvfL7AUwyaI5c7SmiboV9J7h8S7mmEivn6aPAbyPzwtuxHjv5PHP
jLaN8V/zudI4GMfdB+hPPkBRbxONPS6f1GyOZUfstuzFSnXdj0AV9OdPWVATs00r
beKkFCeamUbm5K76DRdeGB89WOzOP2Zb4322pxXX3neXOKey60kAeDIG/3B8FREJ
aBaShWk4vSyEA0JjXdQd/BxHrWfZ4uvlbH7BeLjwxqlA/oW/eJ1SvaRtVJ1azlOR
R54AWffSy5NTvHf5I3BOyE0h2IKsyQcFA8hBeVmIpGf/JqREJQ8LVOt7n59ntuTm
j07OVydqZynA49IhNJTeZq+KQV64bg0dDr7IoxBOiZNzyNK+R8Rt0LKMOzxOE80P
ufe/OUnK1DIoVDJTtcosMqlCLN+kJ4O7ks/Z4SAoDDxXyY3A5gRNobHU/8hj6VVa
h6pIZT4BAfHE8xpOqZSa161bcoJkyG8qADywVfikHXGGammpS2yF1Ela+GOHQv0F
3rNn8BDs/PHq63VO6tfvhX2WpkcgQ5b7rrD0ssmBG4do+rp2QgqjoLywbn//iDqh
+T10qiC2TYQ9i1HPzy9hwYNtjxekf9fyIi3qUOOihdf0/2Mvnk9DAmODfYzpNhMS
73lB37/UB8Ti2fM8FYVJFuedxB8hWR49Le9Ki4ndPsaUuCdVIn1Vo4ULv6HT7KmD
Btq5KtPZfzqAkhn8NppEJObU9yHSquUSDqMn2iKFjspSIkaxPltPlo6NBspY8llY
Zr2R/7WwVWPOkPnQZfko6/xwRMMUAnK+YARamV3DWi4nYnM1MN14rgAArsR/GylZ
oDaHBUAsjk8cBhxCnibBaBcgTAMKy8ZR+iOK5ss7pUbAtFY/1xf7FlmOM1fxabUa
up25ZRl510RZODtRQ7CDt0hi3HESCH8NOtUx79Cyg7AbNDsYwgOcnT6JUvllP8oF
bpt27zTs99SyG1tLcay64pry2k571nDX4kx56gT77Nrpap0VQ4RWPcXRxvO/V7wD
HOKXpl7NqTTAr7XV57Kjhii4WmRNhITgrY9BPqIai4ftYY2N2mx6trwlfdGG2/5f
q1kEDkqz/3/5kV/vVLl7gqLA+P7rldsp4KvOPvFPycSJKrXIqwTa7f9gFmLaG2Pf
/gliFuNb01YH12Xhkwyk7jfwRiIvqEdSpip5euetthOJtnmUpwWoq2Bujvbq/ZYN
dUGgP4KWcsjwsJTKKKzNZKnbSPpVLgIaNgyKCS83SHakLIPtTkidK1c4BnMm3aBY
1fBx/+w8b9WKxMZ0krsyjvUEBToEgxwTQNMTiO8/KvnDXIrZ/fiy33jTQeQk2GA9
8ZuVSznGICmodk25o/gwaWJg6DZaCSsCuWrARnyViZBCMxGnxCa5oKbTrald+vEZ
yV+MGze8n78FOh0nndtIOIF88YVgKAT5h+8wQGg3XNbzPl8b4EIdSm4agP6O+WM6
pnFXGF5FENxysiXDR7tmmSxGMpMSqGnR55KDXTQh1NN54HShGlsq3+PgU3bMLKWU
72YLQbMwmknG8swNAvl4AVQTQQ/JgK93zxiIKG5pPCDvHHJBLcJI/oTYzoCki8Df
rNlcyIx4PIitBe9t3739Z6FM7zK3uHK354KSo+S4mMe252jn5lGqYO+ytbOqbJxi
INNJajAKHkQ63f4M28IDFD+c5fEU66GcDEQQEqxD1+2Qi76jrpS0g5RrJJW4nOCb
HxIcSAnHDeLNf64vfUHbbEAjsY77hX7XRI8Lf2wkkSaHzfsuv9pyt7HAl39+BvpF
8hKMOQI0mjegwiwIiiu0edUJj1A77Ow8wMk6Ks1SJjKyHmQ6G88wrhLNWDn11nCS
aiC/xByyYJPQT2Cmhq/hzzdv6ro66rnUVdRj/UgsmZvMU2DbCUn7ubVE10jKfn/V
f5qCvuLtBQGNZu4pQEsdsFfh+51/ASPVbx16kAdjOzJTeMTb9w0LFchFVbBFZgpp
SWQ1R/CBwmi53jBMIZYmZZHq5R5ec/KBmumSgFHrIhcMJWcOKuDkkJOMMP6YOGeP
3Vc+lhl1AdjviK2X788IPFUPdMdCK6jW6Cey11weQ6Qub1ZrinUsXAt1FptwDgwv
Oo08J1iDEOZ2pZ5+kqK4AYRnQXEDlS7jsfn0qsKgmqGEXNT+3eUCdvbUEntyV1Wi
bPBZiQSdUnP/B45j69TofxMWxh7534ghYbcnVO0HbgVVaYgEMzkDxel2Ws158UmN
IsBpnI/MjrhI1/Q51O6uGiMSzN/PwTRupU4G7sgAiqYxK1IKQeSTpOxWvo9zWRX8
n4n4d06fqnnQuPV43mWDXmUGOiUQW/tTdDY3cR/IMeIY6Wt0Avf09N9ubvfUE1e6
bDUA+MvMGpWRHL5kYOaCG765O06E0kPiO37fQPAyGExlI5Rf9hd4Uqs5aRNsKt+i
qJmbf5j6GSHgz1n7Zd1sNiIvdLI3ezWNpp5bCdeikBy1lYMCpjl6azOo7yGxCb28
Z4PctZj6iLXpA70qJVUj68YP8VQpUY28dShpNcz9ETopqFl2VvEAoZMlP4UJPD9L
BvxlqgeU3OCGUwKaUn5nAo8DkbCDK1iH79aPpWlVVjOVmhx7suL9321C6i4wnSkN
YDSf8MUTm9Vaa0RlkxIuVni63yNSzi8m7Bzg6pafqNMcpEwLNgkJpVM1XPFGSFek
33meZQnE7SWjiv6a4RM11WlNSkTg3Ez80piBx8tx0SztbNHot4tbuQToAe/1Wssy
gnf65oy1QvL9C/pPRr945nfELTwywaUsCJ3IoJn2d0W6+Yuz9CJLEtsXG2Kqfc+B
TE15znJ2iqBrj+VkyHA51QMJQGLcwnhSBMRWFwoJG/LXm7f6ZciV7XY0U3dv0X7O
v5Rp26svFTpX6RYrVlCK2nom+jECLjnnNpzGwTWn/Q6ObjKQGYPbl9zLOpgw8McB
ghF+MZbbMbveYDSOHyKq966qxbnw2n2VWaC/1OMryo4EohCmCienjQRiekDcOCEz
EcrfZhnaccC+BcT92ZOhcWZMMGIeqLcLqqZesB/zcAg7AXSGtOL0SSjywc+xsPxv
jtSW9vTQy+6jqS5FJ9LKOiJqhLT5pmtIDh/gtM+bo/4NGdp9LtDpuca3Alxcp4p4
bmgYHcxVAcAUL6+nK3tXW5nzbhPcytEccaRnv69nwlXRxr+5pbEyRfZM0jtR63nB
yOSf3hPGDoBUI7hHmXBE1QWmul7INgYgge6XVKs6HSiA+B1Wn3LoVB8UR+zk+jsc
NmbNmjqqWzXSElmMb8bYjl0lmBZMjG6NOR/1k6et9T50m1Dl8ncfC/M6Zy89GWZS
1lpwnpDz8xdJdV1KDd8tTYecEwRto298OpmdWZ/VaPlWBzX9q+oXMm079OiM2d61
1RxPQF879okuvHgvQhC98ifbTD6Smv9OXP2dltGtvEsxVxxFM+QGhFJC/c1m1iNJ
0G13twh4iCYaER62bEC4kDxnLvh4xR1vi0ZTTZXTX8qPVumZpKA9m6ShANhx1rT6
mlG/GHUufcLgfmG8dr6IzAnwdzZLDkOodWPS0SKlknNF60aLCKcaQZq4UPOA7Oa+
Gbg+c+QnYzfvbNli+bA2La2zLVspAk149ztsOkZYz08EdaNpZy6pA4yPqSb6G8qt
Ee/L1XxeS9H4kI5iBi7lqsIj4pcEfXLs7D2XPqWFORSmc2Vkerfr7/Gd5Oo2od0K
y6CwD7EkZ96YWgsH2HKtamNz2INCmgPbm1DtUDeYRi4na1WBVs5b1AsuKMN+ivYC
EEUObJDaP9QywT6dmHDPJDR/xp98ENgm5SBf18ykvr2HGM65DAmglNbZriXHqHnd
cu29/4jwxHWAC9tlwW/RRKmiPbzQi/gQcOGDXB2wLm62MzupBRNntJxuCZbJIVPo
Pjugf5O+A6nplLcDUhfjCipHRMPSOJCke0FGHeqJqfgGrUT+hLvs/yPgu4515BI4
/bQIWab6Gqd9WtqeGfZOv44u49y71YNdbIFfgnO3imbtamebiXl/iwRoHmLIEuMA
OL9QKP2hJKIdj1s/v4IgvF4GceFmGbQMuR/4+5ALXtE1U1moytbJjSdno30He30W
HBAIWaSnJV3/MGHTESv5nJdNq4g9afus4Z9wEXkYn4UQXNJKzAqARJi6v2yiZOLS
0wOvBQGxZLy7xqn8Oig8H/SJl38+0CIgEums4/7Im49Xt8gZWVH5iNqSeyIhOnC5
wXUWOYYKZ1JfVNepVHTMu64buqCW/tEsWDJ158B1mMJAdaq/jeufw0uXSzdiZIUr
TjMdjNMetRGGlKejPZXKndjiRZArU86OJzLVKlq2LJoOjuON9O5fvbH+jeroUIzj
XlsgdPXCZJTfiv/YjtcUEJAazgGRW+x+opwhqIGOoD6jeT/3WdenQPw0k99vX78N
sulh9/EUrArLBdpO+m3OZOSz9EcCZLwn2HQVo78MLfQDcsgD1Lpjh+x8c1/pSqH9
tdyI6RXMdFxryUskd/a4/Tr2wJGAgHsj4RYtJkviboZbwW6eOb7bRDtJ1mmEcsiq
vOktRZtFLdYKxCcdjNcdiIkjSNKkMYX/rpHYVBcCCcoYmLAnAnriPtIePU2KQPoP
Q7UsQy962CLUxMTQ4tOWz1yr/7zCnMw9alYgBccfIZVT16LKE7wrWgQPud0Nst7/
tDfVgtZ4gkBy9WxBsWyNlvSWlEroJSfdBvi7UQH9QkCwtCMFSi7JT9m0rU0cBpZ1
XfMVCUYBM1s+0cfv5aXY3zzzPmSIuBa3kE9NMTU1RAWmVfVr8cxksVwvOodthabZ
djqsff4dYMgH/ud9b6PVhLIgOsMdxHVNtf/uwbNGUCOdYudAmgKz+XCPsJ/69MAg
recDvdsXasZLmG/yITxplLGALScVuD9oJkxojU2xZdxvZdLhFfzFEnlxG3S17/+w
Z0nQzQF3V1oGcFHMlrx8qWlDDWwMsUK66dn370FzONhRYpBU84neSt10DK29JVNV
qOqfLYIycO1/VSZkVKzV33vazHwtrj9XfCCxRQvxElgEDXmIXXLR+7B1S+njgwjS
k+xFyuIHx41V5nZv+XenDPntAQTyBpJOqYRgthKfM4vl21MVAAGEfNZLnxdS7oUE
vVyPr8N3TKTOlKgJtk1N1EbRQ/5JXNaXITLTvKxbr5HZMPvnVBV7yvAStvNvpfJ9
apfBJFhGFo24YZypyG+SolZYWUH5j9PS4bQxcaL3x0zVG9UKc0ACf53/003Ttizd
MDCZtbLo/hxEtcqPUUrcoQeZp5e0XGUn28oTfq+op8WoGebBkLm/XCFaTiwDn+0q
pjAMp3S7H6o2T1LJWN8Hz2mf2pOYozvBRS8M58RPSql+4AlNX6zaVln2u9s6yi22
w4YWZDhEZ9peCxUufezwvkAj6AdtAoXnwH0Gv9Dz/hBCBIYeN/RtV1kJc4ekd+6K
GdgOU7A+/vdxyOzfzhWtG9tKBztS24YKcmstB/rbiu7Iwt9ZCsYSmBQnmOojSkxc
S50Y3BzvAPvwotknv58vZub2IB+uMA4VDAnspZXSVnQ8dMSW8KumzRhCO+4m6hg7
1G71YPBZt+prYDfZGw+Y/KhUKOrpyi2BWMpD2Bs26uQQmoiY5/+KdfqKIsCWozy2
ryBounHCYF5N/dvZielK1XluDdBXw7xbzYy9H+VUX0VJo2gQlie2UnhmJSHmDrgj
9D/sGagyYDwRmmtuJ4i/lVBVWmutpvIvOyn6hOwSFKlBdLik7UFznmF9VVztm0bX
uIjZXkJsx/J/SGn4CulDwi3N6xpZhFVIoRPrygUlyKmMFF7Yu+RLK2Oxqyk6x0/W
YU4TuM7VlBWPWCmpMfPWj1aEgoKTMh/Wcg1/7z9+5kOyji7+jDTwOKVji1VSiJC+
35eCdd+PW8pxIVlvBhm1U52gOGLwetRms1+mgeqVs9fQPm68l98GkAx2T1ek52Fz
CbAoYuxyCPHJMbUD2FyPYFwFtfgLGVVnAnqXqzORFFAwD4BC8WpwfW7oa+4rFhxr
IdDUwgVKWSaZ2ehczVjfF/9480rYFcCNkf/HiN3CteW1cIkBiaigkx4dgUKMPCcm
tb2suFmhP7YcTTEcNCbGtf9OScB8jWhlrjI5N7rBy3J3eVaS3vvUtYps7pmSGG+Q
pveEfGE8F7f09bFn6tx7Fyw7gUPkh/H01PWhaQ6OT2GBtZ1H87HTcHF6FdUVBFC6
A6rYd53ycj34nk391o4CTvAhjBHIt4fPIW45Kg3qp+OVM9BnWslGTfj4mVCv6l4x
SbgWXhno+MoxZcqyhd10hzkQMl752b04jmtzFWvEDgD8B4KfZdS3mzAqJM7INEn/
R7qnjBdWQZi9DrL+6YQQKVgEle2ihX0HqR0YddYSj+tulwd2OionKhyfRbRZOYP/
OfYnwh86y/y0OnY3VGCtTGX8mmqrgWr5d7gkCrDAMbZdSzWBNy/bzS5TUtCrMKMz
QMhRgoSTvjjsfrCWeiCJEzVX5WGlUpIlWBXfAUr98SD0NAIvv3KC1yTjWex6TUkn
A2sm9GJQ6MSEk5z85Z9LMiaq/jplQ8srx3McFgNTN2WeXCQfjdb+89R47om9MtF2
HeorfufzoMF5SJApRhpX/WTorN40eW67IpOt/sRtHlH72fAm/v2rcD1L4JEpdct1
qn8pu+Gq730OKDF2uvRsZamAtMPF07vDQX5bLdBvzA67byV0cw194rNfMB4BF9BB
aPdtcNv60AVZXCf09qNDlBlS4eJqUGXpXld0iOoNZlS4KGSh99GHyxwOZkwMiWv6
0FngL/JI0OrMOjAaR/Hz+dC9A8uwhiESXe+3lsH7nW5U4HYSXI/bNlvDnwCbwzhj
jUNCu8pQ0jyAuIstVD5TvM/OZRZToI9JUDBtWiaCw7GXJqqx0MQIQxWAzm3Y1ohp
Z9QXh8HD741C3KDX78Y+00716/DPsDwYjuIdgFl7bbMzrxZxMlH1PaVmuCOpCOFx
Iux4zjD/fGkkU7Ce9NZ41dNXoKoMw3WxmiqwqdwVxgYXWEn0mn7RVWqC6VHjS2iO
GIWPD/6Wj0TkSV9nSp03KC/GuOGWD4Viq8eVoINJXXhhyYnSSJWXnuI4cmUEqkpI
DIGdd7wcuHdwsK6RdkFTmCfmGXLeNsqafs0ukhntgzZUoB3WHGYBl58/xIuJXfx8
eQXBQW1kdaGUeYtz7XYZbmRZIM0WUlS3lnbICjTg+jxQB52Dui3V6YqeuQ/h0iDQ
wF9CLOwaRNcAa9RHC7XMqeex/iguJUuochGIOjjt23fQp4mnHFW2J0JKrN6x81Tc
+ALT5QldlFkIOFK2tDal5TUumPbZ8NkiVl1TdIRuFBrg6RUCyt6MBvCCqfRZDWq/
f6Sygi72myITUu4jtbJWSMtNPi82yKJ0B7TASIpvcJwk6abWjll2e3OEbLRtsC8H
IMD7bnN/hwq/C+9cMzFaH4GP3gknGAdG50/s2xKGQmja4dvI0mztp9TjPEK++kC2
XGSwPc26XF7H4pDn4K5Aazho9tOK3aY3JWBfaS2E+TvQkXTklL/8/5DbqPZObu7y
jZa+KRZxeqrhZvG+4qpUueKVy/8hX3X1py3sSbWToY1SO8R4vUvysUvQdBHtFpP/
QkMgq84dQm9mALjWbPnclnJnx7OXHK6BFkTXCqZrPT5JP5B1YpfMfJ+Oxi949BZR
PPV63lshBftHWIub5HFqsz3BzvAqCkxVnpJsXB8B936kKpSqpabgnsmY3m1el1cG
362JZtYSurPKXI2K/WT01izBY+RBHNExWS4/hCjHXwBt8oE9AQjs4R8rglwjU0aM
0f+zddGBrLQE6IGC5PnBssooC4qdnVvXflW5XVORHoKvQaYShDPhZuwCvNLcA7m4
DzhkrWbTzAOa1lSpTNImeddGAOS/YmS2DZNbqJDrRqerq+/M04VVE05WfAXwDpG8
qlgG0WmK26cntmy+FAbUq+tU5UsvtClYeV7yb99GXRYPKmrWnhOo/XryJlTXr7gR
oN+dDbFndK4gL8RcUsQZQ3DLTveCH/Nle/Z+u5OblrCbUePBRHuWagO6o9V12LVr
3WgzQH2O+xTqfb0i6k9+Z63jLE3Q9LagnKdcQzeq+sF4YEVI/2wCu4iyfTmoOjj3
T79kdtNI1k/GJLRm1a/uvFLMtqha1WqPxQvWqZ13SI4NNG3t81eDVQdTTBOte26n
8IPUdEbGbnxP/L4rqvzKmflU7J/um601Pt60dghiuu8551ME1uahgOKcDRKqNGtT
gW7j4X5IApJylacmpeOWwU8zM9gfXIBRCTSnzHi9fTFFwRavtpXH1WRDbOgxYqfp
HTkGA+IJse5km223DmbwO4MAzHNa02o4twtK3uWIg/rM3ehF9mHQ99WAfVqdMjOx
2dOINwkwxWAb7kQ6yPDfBo/Cmxikx48UDdsMwucIW05eD67vN4YNLenukRlmJjDu
K8q+g5ILvkvDq8BkJeUhD0YKwcstO4235p6Y+wP7DHRtQ4zQwLnxNpA++n3dmhYr
FGtSpz9stbTDeqxxeeXNkF0X724DlM4wLJteu8T0wQr+6j9UvIfSuCU2l0rBSIZE
BS08Shi03NmzdIAZokQafrjl+TWUxKedig7zaKJYsak+XUR4lB1fDZf5B1mhB++o
Yelinfo2PSRq2pVj2ETvEmMSVPIZ3LsIcfnrFtZzQ4a43ayNb94VpXlKGe2lmT9y
hRzZbIBMnTVNXBOEc9cWzplkqh5QQVi11w0Bs1qaRBUANy2BOFSmJ4B6V9iDSNZT
hWhe3Gg2a5kklZicEkYbNqit/gpiPSvL3SWTevsWvTjOS5bUFMk7v0N66krSpDgi
EwU/gSjKCUykY6+VklEV9S5AczCZ+eIY1BuJFQldAh6uCsELvqZaB46OJceGhJVb
DLhXLiSTHQedoUe3CMRqmRkCB7pPvqr6zm6J/R2BQrWCdVtlZoYUHWlWT72yKj07
OtmPIlGlfT+F1VEk6EHJw/fYenBzRNsPy1jdL3YzfWfq8kTpJXX83TiIJljODPSb
2DF6IwfrQJFL19TdCJnuBpPtrb0uMr17DF6wEiOdr15wI3GNFKQzD+JwVXhR/qEf
cTV2rNKW4+2LfKZNX6dEfeVBu++AFbwDqCgNbjeeQEPTswEFQxk2zAG+LR0EtDqq
eJ1zaKjd0akosUndoU+GBv9xDB5TLgN936LFE3hTTfwNMx6KRT4PxUgZBmXX95xx
GkE63KRP7zRA3Nofka253Vwjld0Skkk8HbptuDzEZYY3OwuaNRAi2RL5FsEOZdIJ
AluhEEHf2liNCYmG8cSW7Noi2Ow68bFSL8ZIr78i6PmtwKfyt/mdJ371VhXPo2gN
Y2mLe7/NPopcUqqPR28hF+aDaIEWdyetJD5c6BmeTkg8X6e6txuJaydlsKC+VhIg
Dk4sKpN3FOeGYz9BROJVP/Ov3O0gQqsuYMjoiaepYKZVNlSFV6byEaw7mTyoa+Ht
NHiObT+auFFz/elaS13HZsEmu9760ezsssXmXQbzqUwI3UtaRVute5pxdD7Haiwu
8q7EfKFoPwXKHaOMRnSqUbpiR6mbbjfXqjSmHy8qL3ahK/4S4cuvHmYMVSzdgCNk
8eRZVZUZxLaTvRifuM10hFUc29hSsuaV8fbyWB66Dh0FTKY504RLUNfnr/+YQdDX
c/yZ24oq/wVJ8hx8f3NtS6XHeE/wvR999jlRJDygo0JIuH9zl6351b+FwzIUADLy
0fJyKhzhDUtlI2Smbm8GCuphg97sMFcTN+P0uF86YDjq24qAIkJJQZPtK9hivllQ
z4uvMpz+AnWcn4mlqCltOrsc6/lBlbndwLMdNVy4nssYcfFf744pHCyo6Wn+ts8S
bEu/0x2KZVcgnD5TbjjdKwOuxSnhUeZTunKsd1GkkMVXy3uS18UlbPWWmfUoPClW
IzKxV9xGm4gbEq9kpIUfRSF/g/TRstbYwAYERND/BZZRDSelSvL/GIsLQd9x65RT
nVbxbb2oSp5JEGOI5OgJRU6TH/yzuF0nJnN/jFPfDnau1kifaqqSsmfmtJXyYlTM
2gEZG9JKI1XuY2okcgHvq0NnZhT628mE82m57aE0hp2K5Cz8gb3QwxdhjuqBUO37
w7uxzPSbjapSMRMzzbejAtCum8H1D37aQ9++gjh7J8IjOg98Jio3LD8TXiW3RRmw
HiLuPQ8ZOYsqrvkhMUUqF8ZVtKlfCPPJGWcMWbzuX5gUmHFh8qx7+9uMh/PU5p6J
4ueRi7sWsxLdVJedSnPDkf6J/fpBmj7rbpDEFOZAGhHJUA1pCuy1VLYaS9w5ijlg
npZKN/dJXHwVcPGCJEcAXx0dY8at/pdUCXbtwsvq5yOh2bfticsJo0+Qeh7T7GAu
tnEXeREkCXAZ7cTP5oZtnZLrg6URnxAe3X6tOgnLD/dwLdKDBDTqdVHONRSkdLwg
H36Zl0GEc+JaO6+dVUILd6E6G49a8Z/aXRj0fKX0oP0pkPtbw9yvg0wyoDWt/Tma
iHPGYrf0ZUI68czSTuIRwlRF4BBjMMeSO3JpyECz1f5QuIwPWqqhVMhoCr27dwbX
7Q9roFUJNJIYJl37Xm33AwEFxMQfiKr4poDwjfPAVLqdYkizgyEC+Dk38qPKjh9Y
/vG3FTVUPSUMv5ELOJVl1aV9phGqJ9M5KuYswXDsX1n2ejBTfCbPlba9OMaYlmyc
z0Ibff/yfvVoGUwohMkglrJZq9Fu4UvBlANhoCF/uzbzhYlBOJ2pl5ZsMMOWx5W8
Wd/NddHgmXWlyD2ezRDr8xGwlq+How1d3iO6QVK1fJPnYNZpLFxCqJedrv3AFgAv
87htJr36shrufj/wsgVbrboJSCiWdUfxHWJIiFrYx3INVgaz8VSJs8YpGMtngIBX
qiinVEFzbGNmAoDyGsJGOmPgIxjjFOK6le4Iy2kf9AXX24kDb5Ih7dbaYqFeYOZ+
LjSDP4LxIhGm8oVxyRHL9KvHMKKDBQtDWdPC594vvy9QA2tx1fsCqjS4JxVmBWi9
j6JQD166U7GKoZhvNW37E4EOpcGFR9CK3g9BFryOb3tEXeSfTlCX1/lGBPgexcfO
kEoS8NGdRqKM6o49huFeA/MOnyTaY2JTIN/Je1U7jsD6zLPn8Crb2m9GgBsK8Jpq
0m0zbrpxhV52HGQGL0K1BhIH8tL71nw2uHIsT29TVS8J7/o3MycoZe7gJMaGC0y0
aTkxi8yjyoPBwJ6KGQ8Vmli6jQ1FzizVMGd3gXzE+z2wjTDT834zdq7olCM5frmi
t8O3JOg5VtwN6JY73oYRR+lcLqr2o6PdhUXLtcOVF5TJO2FkfQZbvnIKrlwNWD0W
oy7ko+YCIQmzywyF3xAQZyprSUTo9XGDYkxP7eab3PyIPvmN51paT+Op+77BP0a1
ImuNSWMzpEAxEch0QZ7SY2VgTzXbw5aqAl2MZnCs/9df1QcmfaIDAO9Qe/4tAoNw
sqweYyUxjNwgAANENCIrbvLxz/c/nQ1YDJkobj8X4KmTV2yDjMMtQyoB6BGs8gJw
u5NJyxEGCWylTXlt8NXEdrhwlJcDOvNWaBvdVoU+9bBh4qiYmRlTelnqo6Mqkqc7
21PNI6qtQXd9TuYrwFeH50ORfDdjaH+I3fzQL4Z4q2XdLscWxJyrxToIuBrOOmBY
LxpKLP1/faXjA3CVMaTeZ7YD64L6xxwG3UpeoF6Os4LWJ0b83MukoDZZKYNi/QqF
sa5WQXqYoIU1NBbLs+WCtl5LgwIL8flVimvuPsgFE6tR041ksu7+2BVcPvePTBUl
Gzq4FErOTYNhusUsC5nfhZvXT1fAq+bTWZca6/Z37twcGDWolikKCC2PppKvjKP9
9Ak4uxKIEsRnwA10RFXLAzGGJs1bbGLlQ5WF5vxWpvvPacclKpEoTZxTWCoRFVft
+FoNiiOrhQYVMRJONn3qI5iWB1z8BHFPbxQCWISgqI1vEvan4yQVWqTlubI8Ty69
Z7QuRC1VmbrZL/icno4RwDuPwhPcm0rH1QlJnGLMPUZGm+t2/tDMOhW8f3tlwe4Y
fbzeGeS0KEORFZmd5zIw1F3xOmt6VzQyOYXwD1FKFToXnlsApGQqoDdJltIsdQ9n
XI5BSo1lf1zf4Nz96KmPdWRJAgLgVXNwebbEVpPkcPEDHbF5vXIFycIBrFWBxnWf
kMpC7+BFrYkV1ary8EMqKiYhJtvwIWAwhtkqIaQdVzJFnl1WzbcrFxtXWmNWo4wi
5eGudENKdBiRQyR5VFuscgO8cDLAxHeoItqEU3D2l89l7kpHbAX1HJdZ5ZAK7GHm
NFf18gH0uLzigqqw+eDm1vkWAuVV+pu2+wcLenWAMDrEKkvJNGeNpQDrHGdZHZ89
FXIcYQkpaNZO5sWyP8h8X6hTMxuyg1rqsiJyOD4Z3k9yxvFOf0GEJz29ev9RpsIh
AaXcZ3rSDUpPYcTYD+nMniCJYIKssxSCNjDx46gOZ+37wwmBKy5fmFk5j5xMBkev
w86lV9ZG6QFiOADvIxf354L8qvlLvMYPk6UhAMBYAWBzk2/FPgSW9QNVLW3/dsB3
bq87yvzY+TY4MtEHUzhbAzr1KiGgAylgs32VgxjAvLNKzdje0IouVOo5l2+izIIg
YBoMlCc/ustO+9hPrPP+jFmmiS0U+hXkzD15AEUNQYb8awNtxOlfUVzgWufPbdt6
1AStJG3VvUYLHeK3IszozJ+LHpJ3Tvr5AS3pVIdRWlRN4/QpXwQ67DKv7PgRLNAP
MJPFF9wv1jXVd7y1HNczOad5QqjupK8udRYEPlSwiioEBMC4iewZuW3QqtBPKrc9
mCc/yznq0y0vEF14ocOeyzK/hPauS1mBDtEdebEVbnfyjfIXNFZHjO/IckDPaYwi
V+12/4Op0OdrfhDTPC00K+JLG9LocCjeM0tytZi06T9gs9Cd8TybxEpIkWSCwLIv
GYcIK/dtcMgUtSUBk2sT4iK02WtiCdJHyIVQKTzLqiM0Ez+osF/waC7mFdz6uvCW
pnTYEblSl31rAQMf1vXQsYR69YR0Q3kL7hxg99TlhpfLIj02e+9QethyMKDMKXIl
OXMCoemKkcQzS5kBtGtbvxO7kqI9qx45M9CZ3XSTn5n8Nx6FDTtlDOUII9shmWV3
tqD5Lw2ocqUettfztPYGqtJCqR/j4YsinwXlTTorjNvRbLeEufXPDzv0nkezKOjV
zqZAFxsFgvcoaCIqXBgM9lKaRKlDPrjl2R0c0uxNEC59Kv+4lcJMCHdTRNTzQCRe
PBqI1cSQzyyzldqz5P0scMYGbE8df9RzdEPOrZgrp/Prwe4jF82UydlmHVibFdgF
4Ezo5TNOY3oMrO0giswWPiu4NlPAGMKgji8qKFJKITZCj7suwUYsfj9jyhicOtU3
jGaK1KYs2zbzoxNRWVAejOw+0sWqrOCgKN7SUSMJmXV0RfELwyZW4/+zgkVMdCuw
3kIB/pRQLzzIQ7Y3C7k+ZU3RPLMB0bd9oVvAjl3wk6CcTlbyLaNH/Bia3zKuBqZK
4QMc1y3RYVZ3P2SMaAfDW+cGxfWk8sxtsYQ46ShWzZf6Ef6rLfvhuq/fE3JPzHbl
ZkbSAtb+Al67hf9NWsnua/3KEuxoZt5Ak0pld9XdZ9NOS9A6OUwCzsYqnIu3dgap
uWIKrxGAZwJK0s8wQNvIauFedH+SmNhVpnyuK2k0hhswVElK1mlRVDNymoTLoHC0
NYXHydbhXd4n14/aroQ31//kf5bpFeVbH1z8pm6KX52zmCQQ/0UairrLhBLTuJVW
Rk1ZjiPUAsNLUWNOOaFkWZt903xHYsl8lZkkzc8XSL4M/veGQlA2ll1LG0H6QPX1
kbdziuv5mqYa09jwyYuGtFU/pZsHmjOTMoKhHiurVrwt7KAgOeyMBu3gEMC850jP
YfWIOgFMS3vurT3vkNG/K29xd0nvN59dCcb8fQzIfQIxamuFejgOg8xFlCDZ9wD7
7nJDrIqOBsVVnbw7Zyh6BEe2fFCsrntncOv6S5oCyrzXGF9IqXXhCY6jaJcSMwpA
KmwlVqzu/OFJmeq5A9NsrA4myWx0DZzH8f55jOWKE/mDevVQr3eU906yHa/VL4Te
5gRZWAJhImXJ/JIKPToelz6jpS//REk1PuRxMm0j2LlLAqjjahHVrCVKgHNUaGEi
N32nRKszQ4OZnwt5WQbTilhg71vFRtjx1rEuCpmW9Xiybca/GL371blkQ9NL8j7H
oGqWuORJEFiV4sERtFnAI3d5wDM8EJLH1XjoR1DyDnwPMRCQUk+nH1B2bS0KRUjY
NnOWdLtdlXsQdS6j+gyKI/k8Fy6uitz0zuTGjy17ulewviy/utq70q7pkysYRi3I
N6a548IvpBVEUbYcosnpcgxtWCYR/2VjoDqFHY3KMt4CUrQCYAQLLpSoZPvC5+se
+YfZmxodTAj7u/mzeurM+WCpLSabY1R8zdVJ4yL3Y25lf0owU0QpQXR8AR4Ne6KQ
F94S9kpqFJ+butTKG4B1vjrmdJObkQGbPnVbIo6gpEsBjqnwyycIffOiyrUGWQxi
Jv/cYWeEi84QT9BrpZo8Auik4LVpbDJQ70B1s7tX7XZowrLXd5az2eiZt80InP3R
cYgpq8Llgtt9+VJrDip3rU+G/jbg/DyFQ7hA+eAi2y1mBbGPSNA+t5ohhac7IkMm
hjTbRgLDcWYN8dJNnOywfjaxnpDOy1efG9WOkUoBhRCSpp8kv3uwTFfj53QTOMXn
XMvCtNtzFMSpGRkmHL9YjEVbqCdlQlbSXeal5qUhecD2GVrIm4NnNJoSelNo1FNX
gJF86weFNG23kFT4jxCoZwIe9XmW9RkQlTNDHpL91aeOOCVDlKeSW9esC8rrMFOf
mkoiN0NQdjN94KU36LNMpipiOC+ZivgtXDNZdgtbG5gC2hboz3AIhfJXKOQrPWWP
32WWq4aAa+m0mK2T3WtYgAXj7IUIBOioN4qpBaOHpYWXUPvjezIy8aUqbph9buUp
jir9lsfG1mOH7ydCA1Nl5YY4F7nSgaRWSHfaJV08u/P3KhKUbng7jWz3PI3RyLWe
UKkNJBVPm28cAhS2lf/giCYd/aBX1sGBeETXZ1SZyfwE1IEJ4lJtY2XlYezRl9Wx
RCdo0GUiRTxwR9OgPR9VZyjE66zDZyVlxJ08rXX0j3ObTmVckDxsxOGf3HIX3YEm
Y5KivF0ySt6vsgIbBrAwiA2w5USREcgA/DQYIViC6fAvg0DustrVde19jlFJCjxk
KsAZwGBBU5CZ17JjjeeI3GV5YCmY2x2aRwZbOV+wVwdiu5dIaKl/Sf14qzHtXbhC
ShbQ0bECLGIBCnidwzLqRNafcCPCsf0tsyYGPCCxWHm4FhCtNY75mlw9bDc97nx/
TS7y29H6vSHoPUmde/ICWssVbIA+3+Sjuhz0iN1eKinAE//ZPLvEwt8kCausRYay
sLqGTdjYFi4xXQKOsN7Jg7JPv/Oc1wzI1KCcK1pw3tDchK+NDcKtm/UitCYk8KPC
lq0joLff1osrXfs4JnP+nGepG8mt7MyoNH8iB9iHXpW8cxQKYfzHMb42r/EKvoD7
Lj1my2G00v2oHLC3ac2Oz0AblJaUmLTIcTkxoktSVKvDjFnKfOe328D16bCa3N1+
YiKKp0wVxfcaG9cv9bnerkhNHrB5YnQB2f3Fo6rFAUaEbNPnfZQGbeZ7KnnxdTfv
pwzMXNv0F9CSHg25q+e16QPmCFRmASAqOsxbAxq2pvRA4oP7bxyp0pinCEtIJffc
wGdAPbGF9aa99UoQp7pHeXmVfepzLTbKAV2fPUDAYJUEkmnbk3csT4oL7FwuY69G
FqeOAeam/TEMTKVHjjHX2z5UjfhH0Iq+Zd+bJAiNkDQ+Uq0djaKHbqRQw92EKIQj
cgPPUh94H0SxakxYIaIOE2J5cy1uhZnG1IiAElVwgASgY6rlQFaBTv3wXM8GRIFZ
YWFIIy/CqapEpOo/Vo/GOnUhD8kqeIKuB2QhcH+LlD7g0KIXyd4ClolPjaCMtZxr
yBOcWVfzOjVVG599HVV4gyQmcj6u80jmscUFxeTnQ8pIxm9LMuyK90Xen64w+mj5
vS5kHmQ23zhxONpddKSCWt7kJCRj6rtIbBwxfTiGiT6hBwR7Aq4vPUY4s8jmzvsU
oC2tpYBzX7fpZilpbwy92WqE/vZAu6FkJCvU4MODzn5J5Gk/5XqlKdb2AISHeFfc
AqrtgFlllaskwNUQ7KLnUGwwzk8TzWb/CNlgtHtJ0K06SHNoPaRbAs6dWKJBtABo
lr2TW/HLQM+uWBCpXk/5buZMXIoYIxnQ25NY/ih0Z5ei77B9kHirR1BgzsquF2gv
AxzKZ+DGKFy6LKsmCoy2FBbaGKnnYimrjW67so0+F88sCm2NBpQdAZhkPI/NMXtY
aUoN9NQ0lcT/b0KFRgcBERMFkLaNUrz4YzF8IzLkyGkdy9e1PoTlMBrPcDv0l5Pj
3rwWu8LHokJSjoxF4J1rZgAa0OlXjM1l4lATvpXanvBbzjTdhnsMh1ygPd2cIwW7
8jYuaWFpY9JOOZkpN0evI52SFKXfk5X/swd6J8c4dE49qLPd3Gy0GGMRL7MZ757D
kkotkzNk6W/tsrZKXzaedfsXFTRwM67OLMCPwRaDOhFhBEZGzBoPJHgTAoXMhRne
qQsI2STk4tXrnwt7Fo5xFjCO9fcfRUP7n4tkmvFH+ZwJqdyEMA16ErJ9dOG8f6T2
WeFUcJpx9WKatqUwmcDww+YSgnTmFKOYPFe9jiWy7c58zYs2mbgljbk8x8QM+AYm
BZV+ZNqozh/CRli0GI2gAuJoG7CWNdAJGGf5mcXQEPCNGiv1dsrj8mBYoyUybq8A
TLmD52Y03BxHPP643I+OHSZ5EORl16KvP2paNAwYrL3yP7WvNbsmTpHROWkJfs7P
JUUeq6BkrInyAhlWFs+dFvLUR0LGtU+x+tKb+A6AdP+JWBWZeS3qcIwaq5IOvwD7
6BqIG+2uMhb8Yj+tJI4I5MUojwCY5Jl1YHoy8BQ4Oaplz8RZA24XoB0j6fskCAFq
UwnQvfv5hVXnUi7DSCd9oUBYsii4Gg8AKA5HHHBK5TDwFpWg5hv6T2WL/WJuGXi6
cczP7U0z0kP1SraRkqrwBZ1T8opmg5VT7lBZVgdsTIhQgUwDgYvD8mLHvWrcsBT0
IgoRV3cHZdMWA422+yLhBSWwqNWTFTB+d1Y6OBE/xDly/11F7DYkN9e12Y+ZMX0m
jm6+ZAGXNA2sh5lwJC4l590ZgqPJRZWpJvu5RKJ57RaXl3/VaGaRiXPVz/X49PiW
7Dd9JgeMS4mr/9itqcfcuqrhhAVK+caP8X0aZcobOkDGcjOnHf76QI6xLrQyXhxi
+U0G1tq9gki/eGIwi7ryiBw1P7W81l8BtLiuDJIyFFKhkJR90syyH7Js40Q4KWpV
9P5uGCWYvfydsqO0EgdSnolnsDrwk0C2/K8itjR2UAV/xZ/KPQn+f0pgSZeWWLnc
kZhDBfkgLksWU9idREiCeU81J1vvr3IrPbZgvLSDSkqPBQTNMY93zXlqmddFKYvD
wqhIF/Uc6tH+T1EHs/87tvb2jIacTjknYG2570NbaX4IU7Xtu/Bp3U2lvzNELew1
hF3EtPHINBKChHrQW/Y/OMCBhz7vL8OW+N3wHJp1mawznyu0VoftpDS15bKVNbLb
OvOgqOaZu8Y1U5kCpDxhIVjailWi9zgyq44W10KnCBcfzZ5eaNubKH+PT0QxAPrS
jRFQRj7m2viF9byMUUSL6nk0IJTF3rHfJZmwm1Y40yZOgwGsycix50peKYnAA1G7
4CO7ABLmHYGItdszK6l5StePWNC39waG9D73y901YvoSd/lmdSc7TE+xZGvgadM2
+Kb7RNb62LOD1plLGpqbATrcaqITXa0JXcOWm5PyRX9+ZqB384ASJjh8pMMj+ddL
cBtUhNnTUDFrCSVwEVTsCJ7L4BThcuKZSCjdmTnNtQP70tz6/MVZJdJXjOWOKL+4
RtxUDXRLKEp0zHsv0h6zaiKpQT3TFUd7iCfv1K8KiwZtZBDYR5mTV/rDsm5vevlf
BSOUndqlETITV9feG03oeDgkTVb9IH/n6lP/lBWsCMtnY+4DVKHB4J+9Sbk5pdW7
zTNzoGvSWNt8lkMy8Bv3+ztj2MiaTcPRWpdpsyvj89jN86RqBlOKJ3Fln2voFQwd
pRdiEA6N6+aYkVugVQl6YGnDrntYGlK/OH8HxhjSVpn/6J68TTBc7FgRRq+I4xtm
XWnF74OwQZlfFFsbs2V69uMGz3JL1aD3BDCFIfZ/n52LipzU29jWNHp1MUrAEAH5
cd5GIEP5YhjBddywceRPsFl+4sxuI71KmdTlHeywfltV09YIixHguX8WlnVHdfX4
WDn9hJsOOPsAcpN2yNPbEqj23sUea1Qp4X6/VZ1idMNglJ6KCn03V1j06nIOvik2
pYjAcFeZbA+h0SPx2QYF/aPFve2u+clzsdq+GXoRoduHXCCGZQ0dEdmxLlnpTCQi
EjmiGfgJj4ON8a1XHBjDJwfCplwxKDc/q1W5hpGoQUvRlQRq2Y7jnzSutDGY5veG
FAHiSNu34CQrCKEWVk9tYtZOCLr/1MH7LzIyyIlW4PNhbMbvFd8o0YWAxoqBqS32
VjDkatPNwc/chhvqfAYi1dZgcTd2U5R7iF8tMRnEqsBISxnIheXC/B4D1GXJury1
TO4zqj9b6N5CTEv7nGV+jgU/4Opbpy/+RCEnYVQBb2VXn+GpBEqhWzx2EAyCvkI5
cvgUe0rsFp9jGr8eASswK+ZfVp4Q9BbcdGQi9aLNnAdPxTJ4wIsjiAtrAELHC6KV
5ffwDq5xQTFc8Ys9+7xfs4qQg9YI+QcpvLCJyisX36S+qpPyVZsR4Ia/ukpUSm00
oFhYYOOhpJshkkkBiGrg8qnqBZLXzBktPNaqBhKHjq+XLTRjgiP4MEik0klDiBhP
UG3jnrj0K6CWwTau5sml7uXoi4C7hA4Abif4zuj7OohV+kjr8ofKmGG1MCBbIBf5
Pc4Rx1b1a2WHEY37ZMLjiUNK7xcgcW93lL2kVtm7RoCbwjPI0Ltc0LIW3JkZJl9e
3h8MMly1CrUzZaLQoigJ5dJGK9SJ/pRDBTxCLl0FYM1waEJqSp6AJXNBdRnJYHt9
Cy8q00f+SNBetFXRPlUE4P2WMXsmTXUGessHPmfcXKuUeyV0OCASJJ+MgroNgUfI
42DlMcmEVJRFR0aie0TqWtTTUl3ralgt5m0i4E6ZhJFSmOC8qOj6M/G4sOJR5N5w
P192LGvS+fMc+yxtbmDbMRUc4IduRsWbPq2AZaYe874AOdS3Nx12V1+6Jka//vB0
8XHCpdfc+HR9WFd+I1NIpdMzQjE5VdBBtBKdxoTj9j8OzLHxuzL5qRwZYQV2eunP
aFMbbMTn8RRLh/rHEJHi0L0fgbOOlZq+ke23csbBURqR0cUjewaJxxzWI2pWA1XN
nkDNrlqC3fAt7ksX8ha2Ku45P+74QsowoMUXvERQbM/HC3c408Rj6cXHcOl9aatE
MFO+lOCDO53Cfye55LrVPaqg1UC6MuNqMUwJQWTW4TtjbmjnsGCZw9kdyH5B6csq
thuW88LnW80BJflGeyi8NV7pJb8h1z8nAAbu0DUtD+MglOhBov6+sMbtAHrgxi7g
BKny29Zq/xr45AFEtCUvWDSFdkTB4+I9yBhRvIoX2E7DOhFk2+ekwc19nKI2ZQnK
J44jRdFV48VRG7eBAxS1ra28uIILK/Uo43574xLFNBXCFuyQNizcUehQ5MYJXIay
VGEw04Oc6PPF8A3FbrE0QDnYbD/tm0wwa8irwYvrtICZ3qZFA14I+uwLCqep+n24
3HtWMIvCADkzyVErbXjSI6FIN8lXM4WA6yShh6MZcz4Gf8EZITmBiBpBVsrSj0XL
DcatbLqE/JhT+hzaIx2qL1nllT7UPfS/0lJ4zsdilKccbtCbfc81mKcpviX8HlBE
MxPfS3sibu83EyCJrflqFVY2pwhC6GsiWLCIHjGdaRv1DOYa168g1XWxFUppfGzA
i7+94eTbFhzuW2lG1QGWA/0px/NMG1WSGb+tqObakuZxnowzICCA0Is4b0/55C6z
q1BqGg1EW1Nd4bTC4l5eEh+JIeC6YXXKosrVxUUJsYt1yE83BZ3UqM0WhjpmIyFQ
8nBj8G6gA9aKKFEDV05BLKEj+GNciX6bgb2fYsZD8Hb0KDrp0T1gHpvwvLIf2W0x
U4Jp0xy/SP2WkRIXmUuVDdt9riaPd/6qk6gkbSaQNEjtd0BosgXKa60XKCMfN7IT
EcVAnagXQCLCVJfdpsvZCXxgc3bQyicQciMllvwMvMH0uuajeObmMrlj9KeuNGus
3aFvsJqaG9jdMwh5xei6/tQWNgqh0tjw8RRKuBGQO9lzNw2rOuOeFYmxAJZBr5yZ
BHXSvzRJ+Geeyrz/YRmOVVw3a8gZgUHumj9h7KVyJ2xb44wJAw6P07zkn/lzVrEA
3SWtAcf5OXKCf5noK48rWVbjvpyGiqfjuPZFAgvtQi7xg/kVcKjmiDwW3o/rev++
lA1sFAymBi5s2DgfLfCin/fPqqnpvzTe8O8cn7EComoCmzxGu5ZUUfpLxiBZ5BMd
8+lJsTL8NRwhgfUTLW9Z3NSkNKmI43p2KF1j4DAAUIKMcItn91l/XFtl740Xf+br
EpLwkljU4pxu/Ogf+q6UtbzPV1Qo8Gq4+GFk6ktELio8llXl1d3I/9fqJv2QO4Vd
hSdYtq+GzqI2pBIIf+vlxr5loO9FZsIDtXUwF/xn7ez6uA83NEExIrYP866NTDSf
79Z1PxyJCwWNzYkO0UNLQwdwtF24OLBy+o/LspVuPiBqgtX24+7OV71Jho8iG+10
HVat7ID334v0sUk/mUA2fC/J+rv7Wi1cD/whFjtmzfmsIalFocL7UnZ2vzL0tU7C
UHZ3qxxf0a1AQa9kkwUB0Tz7x1sKVoX7N+/0llcORHT92lJfYhwLpFsiB09MWNKg
YVXPhTAW4AnHLa8TGk3gFDRZZQP/lEunJooGPmr9SQWNXM52O5eFX/xZ9e0XaTzt
sNyLDJK5aSnQ3ZZsWt1fsvW8ZPNFIqS9eaktbZugEDCbDid9Qf3w35iRL+TgS732
aaYqXyTquQCQP4I+hbHj/N1n+Fh9i43rnpgIMOake1WJJ/VVNOmD0lHSnN8wW0TR
bmKyKbURSa1VtE5WhY/pGAkoKdE30ojw2S12+3bOpkMQ8pUmQOqeW4HzIJHPd059
DKcsBfuX01UMmuSaXDmSEnoqAD45jyBa1IqiiT1ZO3VuRTieBUnN2KtQLr6AiMje
XMvAkpOYiDGIPKqz1sW8h5LGuMB7Tae532ACrm+iHw8tRe9t9+hSg4KtQ7fdMHzb
93FKEUlWgyHwQ+caZzbJSIsM2ONcfcC8BXmy6rKQ5tbiqoSbD8Q6ERVW0bl/kRwF
ZrbVkUBw4/j4qVzAIzO8namPP3gHjUtFRVRKANgAH5HEvTB0KEyJnjRntW5kCpeT
jxKuELulRxU+wJVO8ZuQnPKXRkOMI4aY4MZlua7UZnmHn+FMfOljecdpg1kYCGeG
fIK0wD7wGGVLujZ7tRjbB0MSZW+D09feLhcBuy2yZYbx/CByRkOmRlsPO4+7LMLr
RBySHOblhTsE9BOXF5Bokplz3ecki6SFLXg8pfLlF+L8Sq1glou3E5fujME5c0Dt
MkI+SnaEZSEw+LC3lxuzayPTObouf/NGGjSj+hbch/36Z5QaanQ3lMWlgsR+rD+0
TCh1Ms/5flqxOIy8Jj5d4GH24Yn8eFVrsevnyqE8g4BmjixU7rV75XJKxHUD9RSr
u01K0zKtpS7Dd2p9igUB8dHoegWtQu6aYqNFoURxghZl8d7H9q0NZGfAv4oO1zcN
iEq4moFriWEPR23DILGRdLOJhyegOQzMTF19k6R0bFeRHZSU4WbcQJSVZAU9ZHtg
Y2tZbCsRWhSqJ7u5D1Oe6EJmFc7mCUdzPUZ34m6hGeSbMB7rpiEccvNptVqEJ3Vo
YhbrH2vn/zYGpP9YyBmYCPEKOefM+4KP2PNZ/yReYbPhnMVOZdH9lN4bsCD4pLBs
K7w+LNQNlvlmdNF+gzlzdf35h3OjY5kUmM2es5UX5xRx7sJHchi8HYOGFS/v8pSg
bv4ahJcDf2Z0G6B/Ci4jIoAzsCw0ZqpPu83hrDWsRpOIOHgMeJ6uunzin84uqiJb
appP/85uiugKUXTXBJXtoqbYVhi/DTaydTo3LslzEgDb4cJ7VtTJWUkJehpdHkHM
YJLC+9dJ/OybDAU/ZlbxTbASDchi3Mh9mk19TXuecuiDkommpnzWNHK+LtCIovJM
ESMYfN0vqpcBFxmXqaSuumjw/wpTWhRoMug4/8CTJ7E0Os9y/tyN8ZMBnIjWfDgE
wPa5atfEwPi0oy5eHvz297wfZXgv6Pdm4HCp+63DAryl0oHGRuusqagwPWiMa9H9
n2Vs5gdsbmONIDlIeYFxYb2hlhT633vclGA7LZ/G1R86XOUE5SWDFNsAmpJrS1jn
FUeDVLpeuLjzslta9M+M3/jLbz8h9kmmslsPpBB9wtmVL4tRvgmhWCVYDizCCZIO
oPlOVx7Haz8o4B/HXxUJDpIMHZA9Uhxkwiyva6rA1qRU6kzcqtkDbETQb3Qr4vfF
mxnc+QaUEFYvyoUKhohXqV6WqNfM2HMGp7m7UDsJvNXFCn/gpfge/s6cp2e/krEI
QnTtgDv4som72PGL2V9XKq5eM2/QqYuGe1bbM5oB3OeStepkno0TXT1GmKVQOqh4
ojPdP19kDn53k5UV6Y3HQeeNTm0mRFPnWzG/6jT8ZPTOR69eFjK+YcsdKCVEzud3
MBmuAnmF+MrSco+11JfXAZjM1ZQkvs3QKcRGPKrAciuP9GZU3QODegv8VwvbJC9v
hlyQvVJroxYhPs+FK7B9u/EU3drMnMTuV1Je1S3ws8b89JKFAEaTF4VI808hXjAT
ts/Aq4ZZG+zKpuSXetBEA5SY7clnBhzD/GP4JMINEnEnGBL4pAQc5ZKtIXmqEavp
EXR5JFSBQd+8m2jmdMBEBfQ9BDR3JvIbIuUzOHZYHp16xq9bA8IJVcIoVtvrYVC3
aHtTYcx5wpV0KoTjJmfqVjqEBWZNMS9GP7fxT3/v6qpGOTGLyhkEAEEPHbY8aP5F
dnEqJARZDDe4lHpuvYj7oKO2y9deqzI5bWGIjtv9+9WehxEK3+uR2YVFwY+BJVw1
v5D3Rhkd7Fqji9+bnB6jf3eG/RRn7fOhe8T9v/q3KdRpzK7TK0wEQ2a3oUl5dXLj
ttMlY7XcddWEynRhfMkuSFQ2e6i27aVBOSzupaeo5Jsu17CABimacB+LFNlvzNah
KM2UYa+wsksb0LiAZPUbnbs4IsHNeEKyBzB79xSbMTVKc0w/xCSm88z0PzICCrWx
aPis6hLHqfM3OGc6SN8wAmWR4XTFz/AiEMbJ274RV8c+w6h0r3hypBj8MBlEGxhE
xeNnj/tqfonICM6urU3sCmePHKwOS58MuL4D6O3YvRFePrGn50f9yURZR1Fttu7L
8LJVhz709wlMlkrIaamIl66+SF/iMrrO+dG5wcRzNFozd22GONPSMSGC3KbPT6lE
egUC5YQ1Ttyzr6B2cYXABT+32JJTNGV6KONk/8lDM97DXzIi8b6SOCXr5P0W9lSx
LQqmY0OuMGNbujZyolHDdMd0fFKl2QoxGnHSPz/QWKpYgMNX5jLpq5/MUb642Ce9
TuqSSWRCwWON7q5P7Dp5E6IH2YexogdD//67MOAr29GHXberkzTDcE1x5mO6leQl
buUL2fueRavYf5Uo6DME0RJqmLZkg48f9hlfpUjgQi+UaiUVbV6fGrv1NJ2bWlKg
hxnkLUC8UMLOYTzdlxKVoN5/QfHzHHAJE3foLq3F5Z2QSIPG5OK+ADgUp0Fd1pBQ
NEX8JYQ4djYUOe/Zy+N6uWmLeVRdDG5nzYvzjFFL2wnX0slG32D6k7ikrh3TPDmu
caResvPFa6MbyS9pk7WrWVgVd5SM2bihQH+vdiiuI++4O+vetqgVvVXlydM0w4KN
qVDxvttdkA6GFI+80dJAZjARbMhrc/jHQBWYnpKRVhM6QO/nC6/Wp3Jz3fsYunWt
INmgOa8RnhZmshiywUli1UWEB5zLtyoMF+TdP24drnBf6QfHyN2uInWf0tptzbEl
WmKGBEf2JDXWD3EViuGnrAeZj6TcGe0bAm2nfmmiLysg0bxI7nd/NUolQq3AXV+O
Lrx+gz/XC8xdkIIHpCP3Uv1uMTkY4g2UOnjM/ZXP9V0dme2GWF/KDS0K+NMicG+j
IKVRF63vz2kXcwttN+WNIf1DsL+Th+zee3NrnPdr8s/tcAajsKZTtAJRgNctA2uc
+BWlt+B+Aoks4eSgAd8h/UFnebljghdsP4SAuC1KYbACj1Ohox6lKngZ4cdChff2
Mig+XUSSZpKqIB9YhUqnMmlcmvucbzxLHjD/8u9lwUEZBqUprBSrSYRTFh8GqvCn
UqdeuRsmqy2SeFbFCrHjJ0b3RBTACPJHTHMQpMT8QV/3Wgyjwesb46VhFw8ZfSWI
23YwMwUuRT+ouruKGyROjKwQCbIrpobw3gha01/EGXvs1DjMxrKPG2RZ2aBfZPnP
GXFjQ6YA4V2n8IsEYgi/FveyI1P2HAD6e+sAkb7Q7m0AzbNhTXMLWuUPFzPZ4Qp2
rdaA0gQwZ/ovsbSVfgNT+Pos/U6FdWbyV5UWwifsWAWhsPMBAzjOChmtz+xhQWS2
vzxvrnzcZKaN2EGO0YWNTBwvjvsg3kpaCqf5C43xGv6n3bqQpOZ53L8Dxoat9cmg
NWUt5xvPaPVOZEckYcFk8rsV/U1IC8t05Pf32eEcfC1aritTzgvw7pbOK2+9Pw36
O6r43g7uZgK3lPhJpoA+e6BN/bK9OWBrn5DvrG6zlFx7hgdO+tj7IcNjnZEYBlRh
VbMjWGde/al8ffI8SXqOWKAcUPopJrqaubCFl5pHY+dwHweX/QhUqADD9SHA2EGc
LWFvrBX24FccmZYLUBgXM011TF5oi8IGaR3f7DTgqHCQMhgSKRCNS/ncAbDwq5p/
zU1TileXuCdh+1WS5zvxzK55DSx0UbUzutOkCZTEUFtjlLP0yEp0VEWKeK99JriD
HgaltK7Kdi9fYFJd9YYhxYAXIGvndqyskQqP8FTYbxSzoTuqJK9G3k2V/a9C1aui
0gNAv2u/NUZe6AHbY41+mDql80zmi5dwsE0iPYFNc0xuAtAP1JJ3tqEp54yqSsLP
A7nrPljHp6M+qqCQprqheihAiisT105yFPgDMTT+p7eKqUEt29KSGPmup7yaOrFd
fiMfSg70fSyf8lk0QB4KH+yzmX4CuSNQvrZf0kjLaA7f5BNDHXym5STuDU2cQ/BS
NK7JTPtp0B6uJ0W32H5u8aq+4pptN2W22a10cAkUiuVp36PVRr2YH3em2aszCFjf
fLUTroJIo7bJMVoYZStaPtYmcCF14iY0BEOhnfso5K9Fy4qR2bUSQd9kh4FDxr9w
Ri6W2fwCxs7CDwaDFAnYz6s7F1h/zt/m3MXA696SN6zPP5CBTdSTKJV9+F1EJ1Nh
M5Ree4ypqcEhi/IoaSIV1y1oxVE5eBhaRx/JRanZo7cguQPyidhuVcCtcntLgz0P
lkpDbp2Qg1T5LhfVXvgNNq+9JB/PNCtChCT3FKXsl3YlpGa5Y0ZZvbnXwV4TcJXh
+CqZaTTd2RcfTatLIdD2ERKgTyJZkD13ZF6b0JkFWLysn8LbHu4EuGMLWTw9MGio
zHP0ud05oh7D6CkQPVYZ/E1v6mzSuJmQr06uPrFMAUuqaRFtij0lez1HkposaM7c
QsjfEFo23wieF4n3hRKoK+4UNeYLR+wuikGtjUp9T0S0kJJBHFfJQoAyHLXwv6hu
ceOk4NiqUT7Sq0+uxeeRkTE916FCEFtajTtcHjBKYdY09g6+erjUMfzM7VS+lYdw
47MbATvjRT8CCG2I3hkF6cpFkzSlohXJ4Tmwz1ABBgK1G4oZ3nqc2bPk6k/ayKJe
KDZKbOVo+inWXKgXYZIhD6duyC7o7lu7osmD7dbH8a6SViDWhmSaIwcm9nBfPSGt
j6pBJLRRJhiuyMfooagqvMrBLRePvLCWQdpgyaDoGp+Qh5cwF3s7fEG5JlzmqYzD
BdeJo0BBRXcftUiIXBPMntXw2nxZBGPYXVKdwCflqTnF18rxKb6K/1xkMQIxxpeQ
3+5u0YcSbw7LlRQ5GkbOviY92SOmXwpWti+YQ2f/dXtCgztD3s6EwEeFwjO0Sl38
EqmEapjbPZi93klFP/HL8c3aydUeo/6lEkwjOPDv51nfTWQQ7BmLcbue5MEnBnjG
yfMQU1cqWw0JCogpGwUgNBEe3udj2JCVl1cusofrYTX/kaBiqZLsWbIuleMYd+jK
S/FHjLNpE/4t+wVU0d3RmGCajGjRwLmghnRRQTH02R5JSbtyMv+aDN4wBQkykW9p
E6ReTdXINnRJWDj0uwc1RnCzl0YxbeUIYwj8g6eUIE5sz3bPTqFo7yC6JPjJyuAO
IYoXOG9JmR56XUDw4f5JwYVhkEGv5rlEJIc/v5/YE22qmxY1voch02Zmu6N1vx7q
d9oAyCTvQrJpWd1FrHjxKX8AsXftt91oDEXD22M23p0Dg1BSeZGQnAoqqe9b/JJC
+zHBZSzIdUyI+QZoLIZhHTtWK/SdXqbtwfIS1Q7OQk2jADTBSTfvYL+2dxht1AMK
tE91cTxU7lT5rt/HE00+zg45zIH2OA0BTesYwtSMbzGPWv7C5LRSaqoN0hsteuFS
0E46BtrfIG0RXHboXqKlFrZr68nn0dv4R8LctOhsae/y8zG7pX77tPSrNYSw7igV
TpNOeNS9cBV0NMoB9Lu9Qa5Y6+r7dOM3U9u/LD4ELn6WDHzFTGkNTDS1ext+Loky
VjfN1QsMpgpbYvCTOqeSyiYoQ61Q30yZerpqNjqjB6MGTmj0TeFJ5snVGQzydNRR
G8TL7EQelegyj+fSfi2oBaoGRVy4g09e6oMrfWJQO6jWjrVKQ4faCX/DXb3OxcA9
R/W/e/L5MX6dvYUs9cXQiTIqKpx76JUUOH3AwjKKVau2q+3v7f4PKPIpkKyBMFTL
4PHHva836Fffegm6IiZYVAy9lMqwYHxNBluk3BqUb/8k7sjmP7+8TCqCONTGEzzB
T2Yolsh5yEKnamYT3tl0ztudwg6dR1z0y3wVIMSwtpOOE49h0gVGocE5qEqksMal
PrbKUBhYAhO62aol/gQgOAXLURmMjmAZxQeYXXt2FzKokEOb8EecnwqHfXhOsWob
Kvz8YLFj55MtA9GLEtdX0qy4HnHu68Q8GJmNx9Z+GBOY9Xlz7+z78IpJiRs5eMOO
SQ6d24nrj28/7n7hyQuwmHoskfuy5uV5H8N3I78nPwEVbRAxE9GOS1Kz8HTblkuD
kTCp5FO3qL5dFI7ejQFiac4FQCqzBH5D9g52mCNXH12gqiHnDWUJ+wucZQC3q+7g
QoCpDkTrY3QpkBpR6ePMUg6j8Q45qSYRS7xixXxvi9pCS7vxjRTYsyiESC3kizZd
zHQUZT+D2hu4iYZ1mP5LtqRGi0wxvCeTlS/+EE8tI3Bi5cYJux2NAKHYXLKgWtdE
HQ/DcIevV9NQhJUeM30nbBPuUe0Lw8U8hIMPgWi7xBQ8CyE/1QO8gSfo9wzhRnFq
mj0e3JsemA5/508eHvAXNC0GpIbDjXiuhZrCUM3l/jRac/+0lJ05Ado1xE9Lx+YJ
j1tiRp7kUT3LHgNlpNJRov6y5RvweuIvuBqf1s75DPPSCLOJ6aPfrrmvrkRe1dS7
i4EOOz7FVSTGWS9MSohFjLhEbE9ZVa1JiJit5P/za2Nk2XXx3y2Ua22er6GDVE74
dcqO6FARfpZgWjIrBAMcQeh3lxKu+q/vz95nV0PDsgxlyBs45pnZr3qgvj71pAEy
cCSBJUDkXPswWkXJs8MrlissDwlw2Ci8klac+ajti4q8ZLClTzZ7LN5TIhNwzaGJ
q9BSTkpcKfRSbIS//oYHeFxTqqECkY3LAUDfJv8uxec3+oo0XTtEBXijrtVZpC5O
IlwFytqZ246IFdUa1SQ8LJ2Cv6kTevEE46G2mH9lcNJydEK/OUinsFCK97MJX1WV
KPnjgnaO1nFhsDw+P+Bw7bkaRUWqZO+bvAZdF1DFnIfFkCu01iqS0/tAl4Dp/z9D
tY9N6qnXJy//xrd2rJ9mOLAX9fsu34Hn+7wMZLDplbkluvpvb4uyQlGv6adYh/TL
p6WRwOtYHa2FgOBbwEngRILduP7+4fbhwZnQysypq95CrX2t4nWtE3H3ZLl9NnxD
2Jw9eark1fmXfL+NlsB96nnmIMeX7lR/ZC3eHjDbXdoxFJRP8CD47FZ6DvxOJujT
vwGfR2oY0dgk2wyv3S3qesJ6T7IOlN1LoJgl2u6DqNOWBLo2JhxHB/4DYH5DlseS
oYjZ/4jCLEIWpioIIefQgxlm3xYpFEuMY3agtMnsALNHWtqI5UR98aRRtFYuvmPU
wHMpDUpCCr6z3Db0sRggwXjjAnVxKnJNzvoFOR5juMfWEKZTGmn+NYYS358aqTo8
6I4IPaBHgjETNPCBax9takVkK5T/RbfeQUb/GHNwVLY4y5Iyofz8P6lpjr/35WGL
3HqYe90IMTaQiOjUHeRBgqz0VgWCKIzgdGnFXOYi+dePKXW5T5v3EGjAhP2BsaYq
PbRjRZPsOQIU4Z3mGJanNSyedTYf2xj2rI2G9VUi5TqXmyb9r/VQAUpBhY74iilr
ZjpV/BcrEYF+44hZ5gGnWLYPeOJQsoGAbLF6OxDyQr5cZd8huAcrpIUJLuL43AO+
Nee+EoFyTAPDY91KCYnwD0ehfiyzvljSq0bi1jXtYDKX0A9EJOLCRe6h5jPUpSbE
9n21iD4kP8fwSfORvgzJNAGgUMLltt6e5stWV23/rk/+Xr5KNf9JIaKmswYmln0F
Hbnbz6cNNV4DxENXJERyN7RwNL/0UqYpvO3HmVXKQZJle3Bza274PNpNkiDhTRh3
Ue4enFaMfu3gHIJNAObsUENkflYpKvYsYZl2d0a3jRtjCy5TgXv6naDCOtPhyJr5
T5oWYJaiBSsycATbCZDRwcWpsHQgCJ1oMlOniHwEC7Ev+NCkJZKpnGeaVZvZxpxY
ChC80xHQ8er19Z7cy6BRuR0r8IRW33yckj52ypu8fa27LaYobBMjeQUgw+6VfpYr
oB8PZZDwy3Le2FHfNoSORlSG2k0JCHOsDdYe/fyZw7aNmVndlkz2Jv2IQd6OrMEY
Wm45B49vObGlBfSbuAiPrDJ9fAIu2/+lpDx3n+iCcQLIw6/1GsfUDoKXFb+tAIMf
LVUmC7Zyy3mXh+oI+Qx/fDjTxbob/D+0htQEfcCslzA1xLC3M3cl7WGLuEBIAXHB
+pe1zoDCW9m1TGYT7hMO8T8DKvvPwNFNUEmyMxsPdwdfwntXW1L395r0O9bGtDdP
VlV6W/KfvBc+SxKRite54RlWKQNAobUkS5Wz0chfY1s+m+hlRVeZGFdSIdlXf7KG
mjMwALV3sfh1D017maQiqlYWDwwTq5SsvLW+JmMq7lP29b1m/gQkTIaT/hf9heBV
AqlmsHNgxGA+pdwTmlpob6rzebHpqh2SHE9FcaD2JFyvJ8PvAvWB8o1Xe0lX+Xbi
0c4a1R6/NLMuL04mK7ljtcLjPGvZXXKE+4C+e6SDYAwA2tq0f6h6COjMxAyYx/5L
3VHZvMF54Dk+dH9pBUo36AL07kSSkJE5NjjIJ5RRXfxaxw8Eto73hK+jPDE5zV+y
PKeQS6Ja3F6Qhh/WP4Tn6tkVMafvWhljcptWvEQgkpZD5x9w5Mu2BtSv9L/eh9fi
UkAX0PN3ULeyEY2qTUjZ8zWWPTvDM4heJjCb0x3jq7YcIspluLUJ4DzSGQtWXV5M
KCdgZIyswhibIgzHdqg+/khSel+4frkCRs+CDkqU5jF2/2I9SssHar+7Z0DVA7C7
B6a26Jdcr+On3SPi9u1VYgiNOPicejphvOnRgU/wA+iRBsUAxxFJQWXMQ7Kesojw
DoLqTyCMZBeWNaUm1Ybb8YUdEapEcd48yrID/0gg1gtpWlHWDgf9Qe+PVqKxpYOH
lcncl6DAz0zKVq1RbD05Z2TsAwJ9XaNLqxodoz9GeWFAvOzB9OLdt7/ydsHbNdvP
vb7iglIjd4OFUMLMVdtWwAUk+yb2us7d1XKK0YBObPsgSS6NT2fcs2sY9JJqY2s2
mdHmGZh+aF4rFnb0mxF2y40k0g/giozim97VX7Cw8x5HYyW1siWrNCbKj5GMsOsH
AaA/V6lTPFUat7j9ddfIKzv5V80k7uVeezyHt6DoUiJPzIQe9SfByCPZjUFfZRsW
TZ+hnENGzu2ECBWc8rWH5c228drTAzGYHIThE0ZK1MPz1//dOWqx6Rxr7aiVNcyF
vk1iK5Cv0Pm6Otkqx2YFZbJyKfy1rWmyC1KFBv/kr53T5OWmyiE3BJ4q9uaO/LI3
tRsnRt5J4JAwDiwgWvJ38LdlpVPAhX2+mrwm8nqGlTvx1HpEbItk80qKAB9h4EtY
5Whdp6O2FQHztW1iWEQ8BsmUzOh/XCBeiHsL6uFLH/m4GnyCFt/MZ4WnEKkwTbVr
W0xCvbcSAZuaUrKJl/lghjFV6hGwfYjiX1JwU/y0qSUZy8vyV7K3iG2d0QBozn1U
kKkxKxKDT05r1NIB8cxkogVenKv+bzISH7krqH8M2pc2chJpSx9LukPFsIxy2m5L
6UW2Fxa+9He5Lys2moo9YU6Z4LdjyS9A3QxpIaDy9fyrAeOFogvlAcKXw0+/5+4r
SIv0bNJU0HzHwnspR0cqrRpjd80B7g6Kp8RhvmZO2Gn9O9MuVAQ27/LCMPdg0VcP
7UP7GqVMDCoNHLy6iKOrPqs6mXVVY9VWzWwvGGuu/Y/DenzWH3nAndZ90PQQgmoO
LFXoJ3mND+vdgytQSCf6dS44vC+zRwNI3+TfDnCCSbD+iUmiU0VidPWAfHmSEzRF
OEjBF0jr6yWlkcEV1KkjLXp+uIZmTTJyMOrstW7/QsHGQli0xJylYyPqlO29+jrZ
OEXZHzg8kqxNj3gDCqSozZ0aC+FxSens+drrCSBjBY05vOO8LqmeeCUQucVZbYs3
RW8AUYAXOcWIfe6MdZrGIh7ekXHD7mufS1PCUuhfUzDuNIjWwu98aGuSx00K21kZ
U1mVhIhgchVR4Rql7ixfj6s2Gn9fON/gsRImveslVRVtE+hJIsdmK6EgAsGo9yoc
sOujQylB9BzTerelVjM7dk6iCTw0P+ixHi0gyWYOYFEeTd0p/+Hyxkpfyi4MY9sZ
lxmbp4hMQMLTRKK4fjd3812immn3qTfaj6b37WI2XWAoo6mfKt95IWxnHQ+gs6zf
jw07AB1iX9IwxCHvuJKQtAqw7FC66iOtXOdAIu15+kvGEsJ+Mg3EI/hdNY0cytPh
MEho6N56piXeBFQuRmd+bH1s/nzCRAEolgfcMPC1WzyLAYUzaU39Mj0cGuNseWdx
4Njbw33Af6JSyOrQc/+aXV4QTAVtzbvdn+ZHO7A0Uv5R+qIPhHSReZkIhVkm4hxp
uWkPhaPemmMbWWi2Hnl36+k6ibN5wJ4W1jem+c20STl0ArnFOVNTWYqT90j1hmmL
+C23ZgzUr//E2Vmv3wbHay4NVdpmy4w+xjV40nA0alDbr6AJOIoqbr37UtYIOMC3
yK6f25FGy+DHNKeLwlPZ4tfZgTGX/WeqaEPNmKMtQhDPwRdGxpoaPeAKMbrpfFao
dsBMCx6Ga+vaFp+cGdmYQn53dxhugSd+dSe3u6qXwDJMOMM1LgGbGr91g/lc3FC2
rOi38xnlySrNt5f6iXBrX2HOLASSO1dWgBNPQp6rJrzB2QoGB3zZ4LI7ymeHCYn7
O4Iaeo57ls9NVmgQnt18VP0NpNfqDSe+6g3qoDTOS1UKuVNI5oDbSoSLPPZLf3OY
SwZN8O+qf768SaBAeTKicAJ9etKjNkuKvXh14R19c/cTfhyrW/sx+5arPHNZX9V+
M2eFSQmeEuN2ZBy2LJ2fDZEzNsB3XUjCI9fSBUYy9z0Qp7f6g1PCZI4HA6KP42lE
Dv/gqKJZ86j0ZBu3ZnPD/krNc985KweM3EdEih2GkYPdvmTMW18Iy2f90dP+eKp1
7v9ZUqI2hBaqMHyqNxtiRqgUORR0LgQT8fBTsBhwUGIATRlELfLf+xen1TA978fK
qARrmvXu3/y6xQfak/ocdA2utUkTJ0u+ZZk8ixzy/u6u22F+JX6U+V/ewyQxTtmU
/fP4hlr+NF0ux4saprp/wRpmJ1hnJDGlfMTcKFVRIAXBKpbP6tvqdKwyE6YUeQTP
f3H3PUxPE2cH/BrEVzICM8YyFwBDNbJVr1P0fi99EOfDF/H01MuDCcB1+p6vhgZZ
Hv6WnEB60N/u3BTHz1LfDNBx+M5RsZUdR0n891wJykcyrA/YXCY5giVJ60WjVsyp
QKdEL8EkUZbWi9bKSOdXfNIEA6j8JI0ZlWG3y75s0PkBfGFleyOct7eDPz67Leay
rr1ZZJ/sHlbsnRqlYDjUi8/Y00qacp29WagsDeR/UwpXCARn7B5Z3mT2gpdnQKuE
S77Ue1x42CrnuSh5dsvRqyQ8lwX6FcsKF2/XN79K7skG/faPDJFz2ZfBWgPICz8Q
mtuBuHvTTSktpVtnSK8Ggn4zGeYp396jV5pdcf3stIGeWZY5eOLp6fs0lGKYfMFX
V3rVym2txN0xoRoQg0Vb9WxlUYAx94Bj2ZyTQjghuFOpeNLEAsbKyecwweFKhfja
0oervc0XQBmaLINDo8myCjf95xHj9r8ukS7EbHYXZ/WqHv8ai7S6vmpurNFacZ2x
A+xAMY0jPOpWLnd27q1fRxJzAht/bLK6iKqDh3h0URKjNoAwSlKD09i3SjfRKVon
g5VnQrjYr8rHepU5GIkDp+EUeyaLgQex0pQIyRKXCJEbJrq/bu7OMovJolDHtmuD
AN+icKRqOK9ZAYjCkXKVYsfkkUpzNyARqeITFNggk4p1yelv65FzedtUmkeU4F88
jaF681Z8SKr5sHAXoWgQUuYQjhFP1RVL653nxgA1KrMW30IcoMh5HIpejvW6leMn
GIHLf+FhSK5VSFy2mGH7RKTfMM+N5pSarrtXR0EPo57ZAtlb30ZjMScVB1K/adGT
ZAUi9b54H974ZpTwyXrOtJtgrD1M1xCCAFVv08OLjzeNl00Y86Y5YldQc6qCjqoQ
/RCW57PkcGjZ5TkrhBucQpHxgU6m7hu6Tih2WRCy/EwKgkI5FXhjUBGY/vvBnq51
3W/ZJrH0QjGynVxnDHCqOivFGBHTkrj64E4wo9OMr7eBTff8oL6rTH9It8YHnccB
tHGGfeoKPuZBWFhOWGSTMPbnubPw4767j0ebt3kHhHjjLeDOgZ3KHzwe8o+0OLCE
ESiYbbi8TWuTXoOEquuN3fUuiCmZku7mx406/2PZCwMs8w8WqhJH/JJfDnUEIvSu
YhuLtL3aEw1vsL8veOIHDvFlz1H4Lp2f6ICbKiNWpxFf9+R7H6TjVm2tgDia8ogp
Yqj+XuhdIbOrQ9LdzR8PnD4lQxBuBKL+CZarydhWOJBdn5KAY83gOGUYc+c0f5bM
f+ZJgxSE3z0KOilQ3+OGjZ0wyw/ISpEopIbQNG20IvV+7TMOoSL1eZGZzIXdBR3F
/eOxzgGPATfqb2kVVRKwTv1XsZepTxRCq8T9FqKzZY4HRBN6KMjZx0gYBrSP3Xrt
5zv42Tk9o0wVuRVNpRYgZb9YdPSvXIxPk1RABAoDxqKDL+Xye8VUUXWIBwYOv3hI
uCTu4VFasN7/niOucOXcexsbVV1C4l2VOwGvbCDvhOI5e0S5MaV7aFc31NOiR3+3
DzDYcOlrrq1oijtRf3vMp+NwZP+DKRXmQC9JPmSOgEMmUIsxvh0vmBbDpqVTY/oc
r95KopeQS1wJ9bM3EWKLf3Sw0ADIdH6iotCe/oFgCTn7hkTOh+emcQ9K9bSVbF+f
uncm8tKQHEbaZEOmDwwjEXWhnZV7juitRGBPaAZtC4SvFwyNjsDF3Ns3kSjHNk+N
GOu3ohk/rBHJrvdHEI0fD4gFV3X44mRseW8F7yJjWgWjcVBGfOVsjKw9NMzRtS4G
YOwAi4LAOkoQ/rucd8r9YsLmWhF/UfqfDhqaVxRc3jeYIdEqAXPLVjuX9CI3V1zk
n5AjATRbYR/zhSP/UpQXIvJW/9EA/4x6VTK/XttcXo+oDtLbyaIeosOYo8IbesCo
Ao/Kyi4f9ixOkO6hKKYDv14F0jquol1oTj79YPoQYYNpXAuC5LBAfL/ouP4KV++q
AopBFI5WVkpxKFcT5r6pcUcy1C1ZI88AY4HZKwZcjnY/QRq4pbcYh9wuZgdhCxBy
DhQ460hZvsH4RoVhhVQRq8mXZG3wxl2MhVdo4OzVfNLgo8UhWYA1JZghjB9553/7
STTBR8zsUiFmK5XGWu/+pfOyFwvvBgWS6pp+el8nBDQtbMp6+HPyXBxA7tfnBTQp
LVrE/p3WUDwlnrafNMt7VjdRKzjCo1glo9VRncEkHO7kOYabBHb+t4jYE3ZDpsBE
hBGnD49x9ZIO2KOefKC69kF3cpVlrwZubAl4ihhr+PNM6cQE90rDJV7IWZaQ5UcG
eXIvPTgKjyhNEhIRlTI2yEjxryw2puNcE6Sh6xFk7f8vm2JmjXdlEuGZduhCsRR3
2jgGl0Mi0e2LNkzZItH0QuxweYEpBYUL7yyCDEa4S8xY27uqyasGtgkq6631V/bl
uIDF5r+QSeROB7urmm7pFYRRO1J3q2urJGq2Y2SnkEgt6UyyY5eDZ/Dh6BoODHvR
aF19x839eJsURHQmKSraHTmaAodSIXovoHDR5jTcQ5s/y5MyuU4OovEp1lhtBixu
PLZy0sb3bEo13bPrlMO4aFmdCxGRcAyHy8v8CYJt2nuOh605cgMSSdZx9JDasDUA
PEPfKzmWSXMgcdzUJsdLHeNFkdZ/t3As2rL3zWF6mjfzkrzGQQwpm5IVPDBt7Tp7
Qo+5wnoeDTdHhyTNEOyKrQN7zYwI3AuF43J+xKeK3xVm44sl7cQc9ILC/Uo8rIIJ
9bjRvyIXwcGmzpSuwISBHKuk49ALceynF5aeHIdNZ1jNtijtvKHUO0C7SgM+5+iQ
d40jglsb8na0AdViUFmbxYafYHeogtxJkTLaA4AUL3WCyJJ9F66zAh/YAMwGd9Oo
J1+F+vCFGcpl6ujROVH6MCjXIZoKtrZlhs6i9kDtaO7ffLg0iYW2tWoPNnyySaFH
+KS02JYTiy0SGzLQ7Pd2Z6tXpPKA3YUXRwbupArU+uch/gEVUMHpQC8rg/i/M0K/
bCPbXg3u0A1dXoXzU/6jWIvWQK9cgLDR0OVkCB3pxrknH++rKIDKflQmBnVpG05P
Pf9y51xfEp15j8T5KkwfWWnyFYdqj6tjktJ1P/oK3DZLX0DHZqTnODfF1eCjn/sH
sPuKClnu6R7CdQ+LtuNkOwMhmcg4aIePWGiVbpa8S9ovLLk3C9g7PLU7yztmZKv1
QSc5T3YtkiB1kEHPQu/F8cNBF76o4yUXljRWOn8rkDMWdj8BsQyw4AwkwpY4V4B2
9O2N8gU001ONM+AaPEU9rgFvfxAlNbUW8Gr/Z43Rf5R7+Z5IyDQqb/3htxeIYDPb
2GvtZM1hDh62di8Jq+c8PeCCl993iAIOUcSZLKZHmOpeC4UgpEA8HlyGxatLkuWQ
v1f6b58MOF8Bjnta0X86MET+EsQIYuPEo2iUEyyIpcmN8rRJN4F5s+e9v0cjbbpR
uuHkB//gI26xuf+bLOnfKAcamVHoGd7DzZv7zgdhM8JtLvImuuwu6plvvOjZoGuV
cPbpom7jYOsEuvojmxA1vOBW08njeThsMoB9vs9RSS/oyHJ8bVgGJMrCsDzK/q3+
O4ISkitJ5jlzM+YfvyFgaXFz27Fz5FFfSjywwEcyRLn0FZZjAZTtEWcE4G5An+Xl
UFveKWozcOBwW4e+VqARSoVTp/a7grVhrSpimKE3IuTS+1JSvCLE51Ydc7/MHvBA
OYUKGyXg2vl0qh3mQWFP5r862irozJ8VB2mIxpuL+w+BHOdPqUzSzO/JFvAFd2IB
n8HUCTv67EhRANY/ucbYQmYjny15+CRG7L4IcKlA88HUrW0bk65Rdu/JOsrHpFTE
03WxmU0jDUuclMJyCQ8sJEXX2ptKuUmeUa34wgv2owglA5ZFcyAzjedPMkQM+Sz1
B5PNGOlzdZty6ikGiV/IiVycGdMn47k5+b8Ar8XXoirtav5yZbRSkiENbJLrAf0x
0kULA0QoU2baBi+jmon9XwYIEkE8lrLj7b7xIeWKplbWprT3+RaZQGuwrvzABsBA
BHUC8aOcJX4BP9eaqOTlmp5QjbyiFjc6SU1+w0/hDaGOHKo2Pq20fv4EGLAmFS/L
Q+5yLxapTdJvRsqdBrLnxw9cjlGJuSmBEkmmKUx/iCzNvBdA0gBY4mRAxybqG9tW
gXbx6dMFTkbA110ZDJqNTUWCQQZYyjg693H/fqvNa1q3fAFoNAhWmBWt+70EgCeT
3kN69BVPl14lKY0MEGnmX21BezJ5ZPl++sKuCmLFm0+jJRDq66naBGCpdB4MPNH7
JH1DaLEytvBczh5KVZlgj8tYsPMtkoIiOVPTd0d7yZluNJ2TRULbBmOK71xESJwM
1hHpNqJGtzWrlr4CWVbpy6Ve83DIgGsJW0ga7cRQr0e8UUTQzESlglTeZdMVBBVm
1v+872SzZeW/Hlg90c09/PR6WGaf0jCMBewCWMimAamzrzLM39YN4JhJAlfjtR1d
B0/meq4CXiuhfRqdVeIMK5Hs1Y1nuL6XmSyyZCXcry07bZodO8jmxJB9TispAYkG
wx/rSCH3P6vlAKyPtjUfwvuh+jByFjfAh/L8chft+5k2gROlIMtU1BpawaccujPu
CazG6+GFeitoZzpKBFeElqyjts6EVYJj2ciatuhy16mHwduT9FVFIex3gWgQawDS
bu1+5YCmMeNv2fPUpTFzmSxf/TYllLzLct1/E3tdUGQC6ZiRrxmh8thEQxLM/8Qx
6zrpT/dLl3JNd8NGw+EGUOePTRUvA/D2LtJPSJJwlyoCcmM5jAWr/q8y3PgvogE2
OYW+NwCiHibrhrsC4ODN16jsZO7Tl+Y0EYpmJRL4rS6ePwEFGsYfwyCk34JVIqXI
qkIwztjN/itZ1X9OGz97XdNkLSKAvhBl8+lZWyqIeLYtUjaVwaOPvegqEpz/B1ig
XTilOK8kcflisQp4+qRKMxvWY7kbuDSDJcSiSvgMNVvSkPHE9LmjM+Ar3PHH2FhK
o6UzpvdGSS0ddKoc8LY0fsABldP9b2lmltc8Ud11t9zdIPAvvzzI9u3FLs5fAF7i
b8waOUqnQAsXvAjS8InEOfH7be2ZQ7R1QujgPp9u9LwDEcooWCDkNsXI67MRewUu
IUyMvx7AFnzV4xP8OCAekxTU9ZPK32UNHcnH6wo0ObR/Z3II++r2BHrOCaD9+wTB
3mSJJPlsO6X/dTs7BQQNSqyhOYbKv1NoO03xpoHVwCVKNlw4o1I72K0oPrKp9LRJ
24gG1y5QvNhBcCTblUVES5y9c4a9IWKBsDlCNN5F8gU47cjVuzt/oqEeM7apICqj
GfmqpuhIdDrfX0ErZREaQvHXOORTw92a4rGNVmAhsPkvfxsk6xbmnp0l2nhRp0we
RE11nvlmDcC/V3Lcgoms4damg5AuUAgu9cURv8s/050tPEn0hxYLzrAZ9NpVe7hY
eoThw0nzYKQgQwEj+kks78u6Aei52e6GVXk6lSOpr42taSdoXM5fQq3E98irsKv6
OZcSlOA+/X8RFq4WR7eh/nu+2MUCFq3QMUo76hVkuIU3Vrvy7tpDPj0JgkugL3BX
KY0t2OBL3UnE+pL92yZJKwEmqLF//t+kDajRgLilAW+TK2lCC4P44vn+eMb0UFCi
D3m9+DR/eWK1SVvyz68nHQRIu9DqNO2A1bvF4LeoDrluiSyDcgjKrRGI469vPN5Y
QifD8Tl0npTSmU8yFj0+Rr1ZaMfNKUxswanMEbQN5Gaj58fG5LENTM8gafsUIF4O
JBTAmytI/ixHsqYE6Gsw6bkbZJ2nkF79UsIzG708w96rAX+TBpoCKdjpuyX4EWo8
b1a6T3f+zXcIxbcVtoMyKEj81xxb25n4kVSso3Rhutb7z6sfPi/pPmsKM5XKC8O2
gd6X6bTWW8dVl0iPcXyRXGC3wCDmOIYdQfB4EEpC+0tdRm/f5OHonH7CUkJxaTsV
palC5vlvjSjeK7IYyGu+T2l0dDSG2EPpiglkybFW5gMc40BaeqwsL0cfGuDiXVTE
OGNgNxAJ2Xm04r2ZCypVl9doNU+R0N7WM2+eSEWgbd18yW6MOtKQFcHfd4+ClvsQ
MtHGb1KQa+TATiFLvI1m8FLAl5tFto8CavGawsSXamg7fFAAGeRcsm0a8rfTiSW7
MUaUW/0u6Z+HGFlimVzmVLZ688jhvQRb6TADsxSNRx5jHtpAbGeadLFOTYIEY9Jn
gG0YOxPUDWUfK6TEwAHfw8SetX8gI1o+kBE4GLiOc/W8mPSpKMYR7vhTuHYHZepo
euXje5K6NzYwJRQ7X6T/Oz3cpuqrLf7aYBTa/eyRdwD8TVgRRgdhm3vdr9utMDnN
+c66YoKhzEMcFTP07RTlHOMYThH2gIUrlA/lF3hj9rN7qrA2cUkXfBse2ehftp9+
g9J9RHaL8JUvrUoeiCo2I6xFL92uPnM1jYU1Bcysd7xK5d1cm182pJDvNpyO9Hx4
iS0uYaHIlpqsOAW94rjGXsuR/t/59DGrnjM2a35etSIJlPFAjm0CrV5+ipcjvQP6
5+IKvZ4UxOaq5K1b/E04bSjKzuQW/SA/qUZpM5ZGNykfV6pHfFpzhpR8mAWro4WV
+ypdnI3YHAUrAoReVE2mq/V+uBKoZ7FjL+Wm7ufX784vwtYr4qfyjLhKH7W4XwtS
ff+lAazycPnIrPSbIocQ60ZI7OVTQIiKEs6Eyk2q3raNJOmFDK2bnUr5gMxjWVXT
2XNzBHCExKaY78xZel1onYG01jRB0QrA394z2NKCBRxeTvfun3UVeVMU9MGx/Wvj
YapHPgRD9xHsjFpuvs2n8HszsGPFy4Ce7t7XhOlt0EexEGJlLUJlntk88lPDyDP+
oB1qDPGhA/RmGjeaXvqLc4sRenb0La35A1dZaeRQjbR1uk5wHAsTUUvsttKYlBsP
M38LlHrEBRXV75rKYp7TwCWhe3RgIxisa0sKvq/QJdqVsuK/t6F+ML8qQ4UqCu2X
ezBGnrf5DSj/tq/W0cfT61VC6M8rH4/ndv1WYehdzGZ+WymMPCbl7FYEae0W4jMS
S+ivmPoVDo4wgA+JgH3ke7vkGMb3sCzgG3xuO02Oiiw+/+0N19gzZFobltJRvAR/
zClVJ7S1DM5NL4DWNt/EERgiDynrM5lwTFV43mfrTbxxif07KCdIBeoQc8NM0XGS
chYDDW/5B14ZFHU2LLfyRK3CDDPFaEJUztWS33WOmFx6k5RmycyMKip3ZhTGHgbr
UJKjBfj5tB+/kgw/mPT66H7Jd6atwTYCqTvep8GBctJ/qLOA+l3aJ04yuNKZcnwg
fUHlMmJtPiBsDU4/IhqFZPDGo00GmmURlD2wc5FZsTcwbsBChfESVWug0q9E5SH2
qOueHv7nk48Hnum0McWvRvFGPOphJ6ZJwlEoZerEQO5kjRPhhm1Hez6qOibf2Ta4
wL8QwDG6lvRoZNGmnkNVumg9SglL46J00nVl4yUg0xUOVXKy9FVe/q1XHAKnoEGa
r5Jez83fg98o4vzMqMCGwLI/zp9fSawwE2OF0YIepFc80AKWRAvh1kIYqFBnCMEX
fbKzHA+8tl+12+lnypYEkYD1DJxm75i7Q+ODNZjPuy5ZByLFCw5i5kwaxjhj+V6h
irY9ECEMAZy9G1nW0OMs0qfwiEYhNI/q5dF251wXeW2Y0g9XhUuCBMbEzAY3d8wi
GX5limqUYoQPL86fKg5auKVZd36Szn8R1bZkF1PdwJ9FPdYPkdN/9QlyQL2dYP38
322vtsF7R13t8XVroV7CyCEOn5W0vX11QHZ+Nv+QuzXYmDurIWQ3Sby9/8O669Tt
rCxbIMsi3bUjvwrSf8c/MldSZTb8O9C4ab8ghnrPC4+Rm70EPQQ/T3PkBVVPIBrX
UEXAIp9so7jmfYtAfnAujgowcb8753vxEBOPEDT5KnsqaA0AMY/aWcmC+X4sVrfY
Uc1nCVBwu31UhH6NTaUQ8dyXfsDaYP47GeAv8KynSl6hny1aHOcduhme0C5G4e2D
c2muho8l5SFkYIQUUOmzIvdtrN/nUhlLZK+IozYqVd2hdYxMsbOZuiK0FdoCjFPy
0Mcp/LI93CT6VpsFRrKRiaevMsR/GuuvYN5WZzaVtqD+GarG5N43CqvLql4/+kWp
hm+0y+HI2Uy8nSp8t7hfAKDOpCcSwqisR/jM34iBc/HWdslxJLYZBUihaXAkZ/d5
fJWmYph5XUFVfen/bhS8mQsdJnnMkskAwROk7yeb0RxJsikhA9Vqv8pdMSPtXdbD
NZn7Sw5blYkoIbN1WBIaWyBwQpaVCirWzuNbeEW+6xwYl4015349K6uwPCdxOG5b
tItylbojZ+E07zlx1XnKkUypOIIYvMbjvBiglW/WKLfrm4St8bapTb7bPY+fdST+
uJN6MZJQsfz1xE4rQnc+wsVXR7/tK6JJ2vxGOBeJFHDo21S8WDSoWdyKGrkEvMiU
YwpfrOpv5or7XeA8ShIUHrACT4VZx2b5hH4VwlK3BGyVaWUYku8ChASDfDzu4o6W
JgBsIwytJREVyjEUek1A9wMIYdb5Ft5Bddv1wGX+Fh3oPhd+6fznROZy9M08UdqH
EKkRyrT0XpTTqBHOkF5Y1dlbkpvU5kNlZq2iNBkGhPEyCGyjRV7xs6+rDKruYfeJ
gtHEkNoHbQWfNjljOX8xqRXiAf0XcVxaKmtE4efe57EsEuaNVAIN0kzuZhictRtf
d3S+88UbnShXmWG0hDK6ezlN8M/kLAf8c/i//n1h4dcTTLe4r7aW++g0kS/T7zGw
dUSJyQNu4KOJzfIg3XkHEg==
`protect end_protected
