-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
w0PqAAsNfHXC+BEKe4R21jKzmaOs4BIVf6PC+x8cUdMiSIG8QsdsvWeaRg9hk4g/WzHQtMMDHb46
WhOL7qpcZQOfbkQJGwjhvksgC6IQjlsTKTF2XgwZpjeHll4fgb+UsvR1Mg/ZInimPcO4jWqOaf5J
V5ou8B0q03p3bB1eu40jnZug2RFbsLyqrBMq5EvZ1yTJejAXH+Ygvbbs/FGTgDnJcEppuftLhiR+
nmczIJfZVZNRyTBT25P7Un1OnMYI8ZH8Vf+xbBSiZ3TIfuMcWOO6rbWCh3v/WRl/PA15+tJ9zpAq
SpMn1mmQYo9ZlLXL1FaJxldAKMvw2Kt4hIncRA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 44000)
`protect data_block
XXXqWL3rUDUFfPoNg2nK8YWE/rQ8doOOZVAJG6pZ14sfW74+dJnA7D70C/3F/Wi19i9h9v0R9SQz
awBu8s3ccD3f5+SDxbhHi3wSt32joOidFtSGIru8MhNneZ5iNmlkfJy6+WIX0vjIQarSwy7TiLg0
ox+pLVCGXnV6JUi+UnjF+Lr6GYeSyvqR+YCJKqJ7Rg57kRWG/aO7R/x85w6xT/lW9Z2NIrl4ugOY
DLITyrc7qr4+bstJxdqTr3R03NwMARwAjdUzlH+oMZvwayKOSKTHxa3JUVWGd4Ne4gbff18wRyhB
ueQvwd/eWcy0Q2Jt3rQS/5JJurKk67TJDjduMiiFcPd/CBk7CEqovk9tsxmVCHJVCdVVn2bLNLj1
N3JR8Rzf0IaXYP8qG/9vL3Vf+ulAWIUxC6zcrPshhb9BXcMFEyYwWDCNuX1Gs9p0Kz3bPMS9Q9Zw
ZyL7i8jw+C1q1ATMxsUVJSnVRCOi/4FwDX4N2GTrwz+geDmcVDiDwowYFISYcJd1rsVgvbpJ5KHn
+jx56yBJNn07+YsnS6TfO5myfsKO5bPowVaHS8mx45rRSVEc/5R79RbBWK9dwMvb14x/A/qNVlMT
+QHMbEvyeDd+kg22eWclsgZ7pB45GkeXgzLobv8QKVGEvEi98PzuF30wgYiHYn80iMrnFEasvgMm
rAukWuHcO2+ULH7VofvELV9lsc6M+El7aFc1f68o1yM5A3AswvW5QYp2Z8H/CHWngbyNfnMg746D
dNtYb53V2eiArK6SSoEApYx7a9UMf+45UmrvYVBWS7Q2pY2ya83OFHVGCNoveCi5uRLeQZdqbzco
yMg0lr7kMxw17l+A6+efQDoA8sW5A1HSI/O1CrjDXkWO6GVkRLbq3u8vUXuOJSDPzanHcLrr4TpW
KgSHwIHW5VgPYE/62V91+grFJ6QPcDKPAcGJk58/r8NkaolGfOE5MKgAnYQOApz7an8q087RaYtm
y+APhPMQDdaiRUEymoy9VJ3Sf01qYhRXobkR5nxpMTqd5yTV4pFuSxtmsyu/XObHq2qM/zbLgklI
qf//nXiVPJX/foU284pxS4NiTvas9N9yOo979Eu/cbEbbN5jKsdnPINN+Hvo1teC8zK4YIO8PMEQ
3if9jiUAgCfRuWCHlDx6T9dePqyHJXEbOCW8ymLSB2m6TGJzUySWn/pMd7PqCZs/uek/k7GALPgf
j0mp8ft7+cHopJBDpTp5y9eWCluapzdbIDdabq0raTbS6fvg6HnBtNzT4Su+YMQ07Fbi168jT+b6
tRL98orbQ60HWLxoWno3gXysXXJv/eayb1l8CV0QdKheeEUE5hpCHoZmIY3Elis5wMM2jJoxfQS+
s3TIpfANW0qz/g6Xub9sHCuDfwB5nDfbzFh3cbRLAiGX+lWw9YJoTQwu96Bjm+YkKDPNxe6hFwJL
E1kMKbhPOadN+yecW6+Eo8KtmWn+QNbWSKcO/DWBF6XkTS8pQ8+Hipf/g1GT84ZvCJA/Pn6jr+QF
OphCdeCxaai9rVwb7roQj93IKdvxLKuNcGtV57Xa8bkEYXgjM+K5X81JeLajIvJNllZdgTuNbhAA
053faYRDQVAaWe77FFrDeChFaV30p+3Ud83XUZP156HGjoQsrIQnDCX6HD3YEpEfxRNBOiw2uvHf
r0/ORMRPD9KdqjNBbja5MI/E6TMniv73TMCdacpwAficNfrn9I+GLufzXfznGogSKOHJWQsj+M50
J1yJV9RVre1vqsPyp0N8xknZdXZTdvBUckAh9VeZf6Md3f0sY0qpvJQEgag1QEldtoNO0yoO/17K
he2OhbknHWeK1AELXt54+oB7LX43RcITxGHrFHgGjySBMm+LSqJmLGqeMMfQIot6W8veg3R2znIS
cfkgvUbRuv+5utDuTeNNiSgnZDrW1ShYRGRz+XwHeBY5gwwDnNtZWam6s5xgv1ggMS+2I8GEzbd3
XiwvLOiJLEFktWn7yX+r3UFIVBhA03TU9kfOeMPgEJDhAm8/+F+Sk96Q4+Q3H/e11hZRUNVAi0s4
q9KvTKpghEOv/9VlIe0YtPjtWxWfYJR4pO2gwvK9l4VlsVmrxNj4xRee+ZqZ0IfFqLXA7504G8V9
TAOnn1lMJBrF0AKAjLeArTpUJKRJgsY9+shndyuOyyGx5ykuFvWXjpyVAc01IdKwUPOrzWZdVYEl
aB48Ov9oCN4X4gNvotZdM6NGXyRUlVK2XW40/98ownN6FqJAY/djRPFhTDGqqqKgIaznX5YN46xP
ktIluQpEjdOmoGUB5h9DlzQRWuo0TqQ3ThBmwOUsjf+wmHWE/QRQdNF7GT8kFUdEODwTwW390pZW
8cRZ0CjePSAlxIzqht7dPE8Q0yHiczDegw2At2dlRzuPJnf8pWiMQQIIrs8DzrbiCZZIpETuVBj0
TcO8kLX86zReA87VIMp66vg8qDwMLOkw9or7FGfqxVMfSnTPiOq6vUK2RV1HfrjGxuL94gGjMMbA
yktXjimmE4e4QgEiPahtmxvKp1Jp0sGpW3dNJKgN3YN2wNGV1VCAa5cqwyFM9p6zcrQCe3xOqz4V
CDPt3ypM+9opCOrbvzZePjBwIoNukB/HutsmDRxG0R6ByLQftXNQTgGgu8yuxs+/nhi8n0UfbEC+
F39GciPzDDd2kGuV4Z4ZlMXwZxpcGLrkeomURPBPUv39+dVcjZpaTkwjlLHe2Pmtyvl4jXpL6IJZ
KoW7RcczDel+sErM5+i6QO17CEVNok9Je/44FApH7iQ/tXKhPS516/arUqpwXN+hQlU8fMg/aCHx
PAs/N07Ss+ab41/TylJYlciqg+SrdVUT1HQbDKwLRoT6UvoFHbIpTeL2HJ8CY+/lCRWYAP3eKA4g
jGFcGLuc+4rRJ/zW+lSCYF+uPMIklSD3pPrw1tAJK/IIlF96wNgbj7rCSkkowUAYVlweA3DXR3Yy
Jc3iD1axbGoSapn8Qqcl00tvPVYrxz9zzngLab7SVIfPgYSRFKL5jZtvdQPVnzVSmuUw4lurG1ny
ca63YUAqU9+gCREcFL9voCWnlncBr1ENUSsK+ug7OS42Cxm6y0mM2QttjXE+shrS6XBxkU5rS1n6
LBRnGMdQMjQMsXUB+h6adlA0z75B6kwdGaVW5K0/4wmDDH6eh580kHGE0Az/QUZWtrn/VYSSe/4O
AI5xsuA2Y+6sxD0AAIWo3/d3OBUaAACybfE5sxYmhLvyTfHm+efd30fhTeEq+I6s5n9MWgu5QCF9
eMPf+EtQcW4t3uDaCzWhTD9thEqS9xnoUBjLkgMq8kSFDFSIwsgC4RBfbsJEpokWV/3fjKLA1gR7
9TuYLQt1b/rDxpO5Qb2lo1nvt8RKOFW8fII1o4+ObjFk8jlRFiGsRl2WDLp4sNJfqyArQ9cx8t9U
kksrSc+XCioO3j1zKMHomJA5xwkAZfFNUFk+rexYHkPhznHZJgAwSh6CTEXgU2uI0mgs1XiUAsaq
SdrLdW5GFE41wuHvc6vRYYkyBXAn3tOxr1X0EyN2wQTvzlsUhek1jRwQ+eiqs9wL8qPVOmWICRK/
vdHT8FLBl5mX7tqgDu9oJ1J1kznD1uyEy80l/fM/tfTkBnhguKx+HlGXPHr/iNQHzVE3C2vMGBXa
4XGaTqWLouk3ORXJpW9NorCDbCCi9EgRLsBfG0cs2J4faUo/JFC00ooISBXFr1LmtrfJTSpQQ+RV
frsQRiWFYCdMyh+GEG8ypqecDylZXbSdNNrKIMP70tZ1V8pfjjAtXX+RYohFtXOH5SfggDZQ9V5b
V4CBPmv4ynpum4dQ2wEMWEKZN5U869tL5gwLq5Dx0EXwGoo02GB1ffVgdozcpsc2sVTahV+nk2rb
8Z2gDLLqfSmjujOFzyNZjuydyEQCSLzX5hS5uRhpGgNdoDq8Tk0Fdh0fOnYonm5LMj7GP9rWssHK
vcTXTMbQKsPtmNNlsfeSetTYuXTZ4sMbWYbIVourENBPTG61j3YW4aYb42RJ8AX//a4XDXGAruez
ZEtBkCIjSef/lH5Ag6l/8N+JQipqToTL6QS5feZP2DXpyY36c3JYSsVSdBDxIZoDDLT7VIHpJYpq
7BcxZDa29URG9Lv5sLy1/dzaqyzQuhAz5iJfS58TyD38Ttb0fQ0lZV2YCpBAB/LPpIOxJIB17D8N
K7313xK9URbwi0z5zXf/TGHGGjbL0Pgg7qhidnMFgRz8YiniqFB+YWDoJ9ttoevswRqCBy3n5qdr
y8mgEPAvzDm3O7kTx8pLOw2nbsyQfGBrJGIkPxuQUqccHJwo/MWPCjVVi6N6OEOG7ByhwbxgycM6
JAAtJRxj/3fb9UoUj3YyIKsxvKFC9+yZnSl9bh86AU/Wg3AzBm/bRW+t3viYJfZtt1kUmV9KtTXE
DUK8u4Fs/yALFahC1YwNXkkMplEKa1M4zkTG5wFpFLlpbcVStw8tVxeEt45Jn+Q8gqgK2NCOAOuy
MY1SBY7zE6CrNSDWIYHrhd0pLUTQPzkX1c2DG8hxVTHam4r0/0SXRo640YRBQiSekKIwZUisR/MH
SXu/UxFWQR/KpVYKuIwCZKltmyhRbWnrx/ODjE+0tX7OQCgd3c7VngOIsFSZf8pe+YadH4wwplz0
shskWmURMP29Y19hqlqWGD3TnAgvztZBc9OTF1WnOY6fNLWDYDHrfzh1IKNPZ6zCeQKaq9aLcyu4
8xQqSgtfNHNK/287cQK7vk2gLGOH9/KpKtG7SlIgGn6qmLjPMqG1ZQiHc1Ey5hQ9f/PdSOshqMhn
bbMLc8TmWL+eJHMuUBM0M8nBBBqPyRRarAQ0KTt9muS9G7qgMzgzdlgKkgyzW00fFC0JYNAUBP+E
pLFOpmzl7hzu4zEDHHtDvVRZ80de1/fOG8+qXOadg24AcW3Hi2QZG6CVEFTyxFY7xXSubhQkNf1O
yHjU/aztsqsOB+Oy4Wd38DH5s9bwGC64tl8s4D0T9PiscEUN1DyZ3z2BpBqi6p/Gmp5mSr/Y8LKz
XDGPv9wlffBNsimXVzPbbS4nK5/87f8PhYZBZJC3APo3mgL8R5+L8tGZYdtQHlP4MbxNeSrFxnE2
V/GZZc3WsUmtMVD91XzVTA6G9EulkHHLbUjIWs72mBMUQBJ33nD1x7YQ8fi7NtDuwMA1YoZ/SLuY
ZEbtKcBmh7+zIiJBlwyPPg6T2stUkPnn2tP38w70hY1y1xB0+upMcbzukbFoaGFfMKhOAwpyT1G+
tX2vqdo4th0OoCKR9ozUDVAxJIFOjl3HhQvrjA6rAahBjYWPsWxxOz7qruahxhTKThN88HK2Ksq7
onwIDSwcJ8MLIjn/zvtbf4r2BCY74LdyZ4BvToKB5MEqQbmXwrXmugpbI7naDO1QvjToxkqyjXvX
a6ANjI1xSAs+1mkHDAfzYGVjTzdZsA266xGIiYzo82IYb8bdVQKITXkvUCx1PYlX192GCZqAPClm
2xpjxYTbE2jSqOM9Jbm+Ot1KaUcBKVYHoY5LqDaRL0fLHvSgSusor38oH3tJp/iWHSbi0rpCJuph
BkVxlj/tGjlqN7Mub6t+7S60FQZqvswF9Nn3qO/6/I+YpQSxL2nKWqbDySK+DVWPHb5uGhEHM5qF
63UrB8H4Ahb6tXLVohw+Gyst9lmM8MTeWS9PDX+8gcJyPMUuItJKdx+WLKC3D5zzn+Y7loSTkeSt
05cnmoXezOoy5Xl/xB6kjx29QApD1yn8kS4avsyxePz5sz/nWfI0qe9vwb7z+s5NfK/3XIWsncp5
3U0meZdWqXEZbmCgmQYUYjExogIXmAN88jbqWSWJg361T5lDRujU2tLQkCMH95irjci7DWB5dSxD
LzL8kxd3q/eFIuhx1he9FcYfKwkVJUe6rzaBCP5vr9AaWpBSqg5nZSA2P/nyHqMrdFyBSC4UAH5I
QWddtiJQK8Ad3EbCY2IYCzTzIywa+wj0xDJdZAgSIXTbtgqepSBZ0J8lZF4nkGb94ZNkicX0TGJ2
2s/tI4T2XIIs4X3r4+R6gmGVpw6AXAMB1vi1dGFUj/ZpmIInoTZUOkFan/u8lSiHTb+F1eHlhFTY
VIzmYsX2kFN0dNOU0C3eYhsnBmywxL9jDnenrRcKM0/dvwOwh9G+N5E8Z/5ECyRuJq7wfxFkNCu5
3r/tzA5S2AqiKb8mcl3debzKOdsvLg62gXZeBxu5CH1jFQIfVc81nhXyUnkFzzBsa9DR7CIhwSP5
VN2+p7G7pZLUSojkuHHRZDzoPZSVa/mbi9HEGwSQo5fQjqCrqGj4vBAECc9fXsQVhcOd/F5QhJkQ
HTDxQhUqinexudAmuCgTiJP4IeA+wgjMOi1Yr+5WnRSu5am3XGR0VzeI0u8Kfi9pK41I1wi8T+Lx
fqbhBHj70DQepzqThfkYJYxDjVNEzE/8WQl9FJRRlyGaDMCuHrJthw8pya38IJWjlOyYHX2Hx9UC
6459bUo0l3ebWf0m/VB3QCwkvNEuDCyjtAv6o6461l5dKCuJLjagnuqoVjqArgjnJa1d9aStaPVq
Dck3ThhPPrTkLPzHbCx5UQDx0iUElXEdrBDN4/qB3gfRO30AhuPMUtEuHJBbVzZJFcfu+Cumi0X6
xjFq/0H5gmBuyj4hFILyuhLnb0Rq/H+Mf35y1uV6q9lNudP9lFkWU1xWWHvYb6f2Wv6RNJYVUD7T
t4s37lgJjj97XBPWxdeMm5PUUabk6ujQ2r5uwkz06zlRxxpBHByjNODMochUTvcqv7VYGp2fdMHJ
rN0d5VbD5aEGwzBmQ2SRIREBxP0Mg+/5YutdV6FlULLivGZAq4u15MTs0/9pFMPKW8rMM6c7HEMv
ZqE//lPD1a/gKAxSb/4RlPt45K3ZQXGcG7yTyU+EXlBDFwyu+obNDoqjFbvYV5CLZKSkFOMX+CKH
OXrRKDVXWZQotUn21l186Lm2xIMDhDgq0QYxstrtYYWCxlcCDmzpJTNhEIcRDRCpn+5NGiSa5PXG
vg1p963ywkAzHgCRbaLNMwmoPa7BPfp40cGKA/ghZlKdmAEeCArF8Q+m066O9AjwMSPG/kBQ95DD
9HWEOW+IyLPA6eZewqOMHBGoFgcdDJ4QJhSMuJ92jeezUFu8pjKQvU8FlX/8c7OxCtrXSwOViKvd
27oBrYgpqFK/m0MPfX11TENay7ly8Rwd4U0qXcSVwZf94BcY3X4N+fS2pqQicXuRQU+RIwbj6fnB
SX9QqrpUFixwVIoQIcTkznW34rAjsFs1Mtd3sW4NHpcjde0ycQJIfGa4SmhEfnKTDc7MjIR2Dh8M
eOFWQtRQE2sFxnIPDNuI1Ytnq4h7kxMidPnMthv1nB+TRkhDAlmhVXBlYBBW2cAG5bfF56KgmPY5
1P/kZP1HOMUSZrbDt2JxzD94SyIZmK5XsFe5651NSiZlD6tdZBd7dhFnLtY48moHeQh+GOmW1qRT
Mtlmyihyg1Ab/iDYpoSaQzcfDVvGfAxadSkggpCtgAsug5c5YxFDvf5ScSo5vMDVIJGiITNiaCeQ
HcxPoMmXNHl6HWcwyH/oK6ELGGqCHvkVGtDsEecLopaZsS1FKe0OI+MgNXb/iuhpGcFqUiMwkzMM
f8qd8AJbq6NzOB35FPCWiI9xi2/pYx6CI7P6HnKy6blk0T0/cpUFFwbfY/4FiScE4w5jfLZQ2Beo
NB4kEHh40hJNf/fyXBwuJcB79MRdspLgPcRnmVYdEhaaHFlnz5G0PDBu+dJIBnmDdndJLx8iSnxz
fMttufsgy3Nj2NEC5A0xbdNHeIUfuYyOyiOCgip0Ldx4gmgAPH1q+WX7XyWRyrEBE3HMCaaRUINx
ZwK5n4d2W9Ox92Y4dj5ZROtjzDle/1OAlW8g7Bnl4zCSk9nFJwsQNfdi/6GUHjWcJ+ImrWLKp5hV
xlKPdBePNWZesufvRUiJ+7jgXrGjdeP3XOEE0GYZ46nLioQYahjWgzckbyoV1aR7L8pgnEFYHg9V
eAwUqgvT9Gxtvon0YjaSHb5l+RGRU2PIq4Fn6CqBNk+cnO+pCKuT0x8F1BNezH0BqUqQ2wTTQgSj
ivKC/EWvIpSnluJTaTRgjPzTIoQu91CrLY3vD0jHgN1CpgW/WobXrR2IyW+9fYvucCIyNN3u/GPc
yb2JRBLQscTLfO6izw1pUeIR+0Vgs1D2jcrkgEEtBxDncTTrLk47LDg3J2rF43Ux3mynxG7VlO/B
jI1zmPP+Vr9DQcyTOv4tXfOE7t7FHipgXLCV/aQAn8hsm5xNWWko4Tc0IJjEQSNJ85291nx0OB+H
/X3zmeDe+5oBtY60N24YP2fxVTc7/ebeP9xGKM2s83fnFikqdakClXaaC8sbB6lTklaD9J5NVpk2
GEX15aF5STeK0tXTlf9DOF3KLIm2Nir65pUYQvKqE6KGp4GKKsevkHy5Y2DlEL4FBSM+9+78qUPv
Id5UxfqMo6Je7yKv+o8O2pSmsBcJXqH2cEwNbf7oXDF/x5HwHnB8OQvDbtxzpBLbMdgJzmtobxxh
y5rYnFc2hHJYw1Wf72V59Q1+12zIPMPTr2YsCW6hVji440TLmhT2YUjC9jyovywmI06LgHvHbL3K
epNe7hDz//iKPbBUuEcRPPGwTn2YGt+l9g0FXl1CCf5S0KIeijPYMe9PcTUX64WWrY0d6W0fortl
g+dob/INhr5Cl/JgzAvfkuuD4pnup3GqXbwFlje3FgskgeHFosQ9PTT+Rb1o7b/IeLdSD1N33GyJ
9KomQkkYC3fwPlLbHMAT7DDqHBynvJd5tUPiQu4foPdXbIoZHsrXgDzClX18+XzgGV89da2KPR0S
f5BpCYpR8SAeSi2hb3F+aDVCOpwHNFqU34K/INKTYRqr/kgv7SGNl6qsrTDup6/RkYr6akBBcDij
cJ5kQOYLh7gq+8Whd23C6grY1yD2yFbkJM5eenp1/HEZds251FKZlPsqOqybbJnuq+BQsG/T1oRI
+c3OaLAv+9L5gOJbKX/iLAvZnarD2UWs32L/0pWiZxpjqG4j9MB+zK8/BOrkp0kfUNero65O7cj+
9564WKJ7pGBKGRdCh/Q9Sdi0xo0yFAD3pJMoRaW6GumKYnEXXqMsV7t+1rRtzoCh2CmFK+2WdLVY
dUoYCX+qSGfw+5QK2Lg7Jv37/GfLPrJUAr1LzFP6sfH4P5ZC9UaY2mKYxIrjAroPHWVHeX1by6qV
K25JpsptVqskZmttL1jcLgRNcSUKwzOAVPtCdgDIZ5co62HfR1eaTcIJJBTXyzDF7KNnLfoRRZQ6
fDk1n7uvf9uDdeNADSM6osOuNt8N3T1U7tF5jdfjrFO51opNeHUlstIdg/HfqBL9ApoulawJneTx
En906BpbBAdMP4WTbDWIuRKE1cSUex8WL7pbSsPhhVo4l60AJbNSaKtPnmKf4ylQfdLjs6JpDi1t
NOjgrfPptgi0VL4hQMRGq71LU0LPk3lB0VMxOhf0zxbfUJ8TVOFHfoVTamYIqUBKbO7pKyCNoygi
F7G12SXuZvNTSO4kkF3sz3EUHcuVcKbMmyah1p/HZp35sG5/3aDqJOn3SVOdbr89IR7r6k6lw8wW
RYJJ1V2gCZcS1TG8BmuYyMwjEXbvdeFF3/YXcqV0gwOZ6+1AmBlSnTATtUx97szT8i03/WkwD7K5
UGjVyv6yBmpedTjKOqp8IzYiF5RtMXWsn4et5yZiFXCdAby5pXvpNojvCtSicQZ7/GkDw1UGPQ9V
atTi+wx3OsX/7czO2SVzGroNmXnF2UERV0JiDB4YZMbigiDfNBQDb6HU42S/l3ry1fgzZT8eysXr
XyRwuLKhJ7fApy0X3qV5pfEScmPHkvTE21SHTp3lru6tGdfIRAdlFJqviOmPx5M6FhUEG80d+LUS
aBVThFevscbOLeni91fMztMBZn5ogFDAYEEwPmrvE331b0T9x4crIy8murmm+NJEh1rsnAprdocK
y19gELcnwBHxbTHzBGUGckZ0nL2Nfi0RpZh2cIram3T0IIGnK8wUvziS4euCU9Q5stmOqUxcJXk4
ponjuSyOi7Zxu+/SI4ZeY4sPO9ZAdjea2vo4QaFeTDSXTrawqW5bS0zp0dzN2a5j67sYfNQdfUR1
FMs5TVO2jDCe2xtolg+9qvWZM8wdSDYC5dbmno4H5S5n/UslagnjjLUQHGrM+LA+4CTj5wtFUful
vIpvz+mjsxUH8J9yPIX8hhKpDoipmNcZqDqGrc7E1Am5F/Qhmo7/8m8Dq2npQ71Siy+qIZ1VznMI
KEeFaWNEbJR9nz3cSIyUUpqipF/WJFskAHQmwATJnS5ezZrdNlWY5hh61qgAUjNuZTh6yKP5cEf+
LbI5v09Ac73qQ1lSHp3IKvEzR7i/5OVJW0fMCBhBAPkhDmrw4h5BkoG5/1WalKcOJWWtTFxWY+HR
xzntD/uSMq4IPcF3oVEgZ1jib12/Ys7r5d/sisx9VxtJN4eEXBEmgjSQXx59Q4thQSThBo5ug7sX
5jiy4v/I7qZVDdEFdrretY+fKsoK9XqAgR1w+Y1aOjJsj4u6kqlc+2R+lVrCH76BtHVqbPKB8ZMG
QclfTuSekZzHQEfZDaVzmPltqV0V1c0Ix7cTXeK+mTw9wybUiyulBmEa+48w0rYivItNm47z+ABS
ElV/5+FI2AmtThsqpW1CdQdU5JQN96sfQkvPmdUkbFwhmw1pteuw/T5e9qYvUkUmjf3ul+4GIf4Q
EmAmMgptaTjiV75ImfMrp+TzFRLfQt5zeOuMT+wnth2gFQ4tELD4XjCUC50fWnKSs9+uuEaFjHAV
2rc4z48EnOFDWwvPWBYvqXRdLy7j33reRc5w057CgK3uGy2OhtQgqrL7DUKp3gMwhdrjiqFAT+tE
+Lr6ctvsAyvHjrlNackdYX/PkIG9tdaQfTkSX5t1whHQdlFsgjiv3TspmyYyRMqeIMkp2lcJBSJP
CY19P3PqYXkXFNsp+XNKoAA2mssxnmrwTegbpzT+ZmLBfbGsIJk3dvyHLq7Quon1NoIqQECwbvaO
4yZzaFJCF7qo9l8Q+7yYjNnlOBnTxiIuLxynz50j/jH3Y2mKKPv5RxfmQyfgm/mSuFu9L3BoTZl8
owBe9zPM2OFctekpVVmTNCl0ly8DAi7wB6f7x3f7R9v81zo0qoe6vnZ6VYpB6j+Jd7MVgsdsSMpc
pYLBBfqcPrYCxUYhZD5dBRJy58APpLn/bzRdUW5nZ51YCt7pnRZ7Vs2r8fHGZbbjVNGCNul7Y02w
BQOa/yo5ttlKDec4X/wUbKvJGQTuaBlOrVcS6U30qRDknNn5ji2JDL2m8AMZABjCFJ5V1HcTbKWB
DBwKLDlBl43wkI7jeuf84fnPK2winF69lj5ncmbBQ1Pkin8K0djh0Embbl9aXH+ihDdUWZCW+uqY
JPqslAkRaLZeAU/juVuLpdWl01clPEOyB1kyxBzXPeijRv4hTTiEOtvwdYU2Ra8Oo6hNZoZSnaz8
RwANfsg5swLaNyEFs6eqddbOkqXLlva4MBOTj/zPNjVN6NMDQKiClPYHTN4Qj6WkteXAUqEi/WI+
GjQin60pp7tm1P0o5hlNuKxnWkeTwAIScdRWv6v2FYrSjnzu6qTsHiN37t1koXpD8jO5Bc7H/Orp
wQFB1rpdeieIBO2wGw6eDeF/ggYNK8VjiFYFlNKcATcioSH9qqRpASYoD14T4UrsfFNzziSqVlHn
Mtex3qmIicWGVgvFx9K8s2jUufT1xZC8SmNt20bG0Cu4ZkqsFgTQCA6z1ZTOePrkwAQ9uZGZ5uOj
ASUapTexIiWRbHCB18drprHjyTX8/U3uiN54w/zhKG+1dyJ8NACJBsuuHxHtJN3myBwG3zFHvVTx
iNw0t2taQEz9lWRkoy5ZPe4vSZjgJw81bVACl9S39BobE7bdqXWVbexPAcMjTgnT8ROlARqN/iIH
K1GA2OEPpWrUx4n0DZepueHpMgZa6SWY9RpdJ6/KB+QvegaVKNWvJJErO2RmrPI/T/58X9VcxiCb
1OvuxdwemBVa3GEk0m4z2N/AWosPByYbgxxo0+UiRpB8s3YS8tEYYHN13Cj5KQ9zY+bJ+zeCa92F
vWJ2xz1gik4WY0GnPekPNch9Q8BrbqXENVuwb31kbAnt/qO8U9rFdUphxP5IbXEgo4Rd2MG4Kpzn
t3MENeUVCxHDV3qMybJj2eCMiQXzUmAeGD1caIXPGvf4wQx3Uv5+8m4aKEjiruA0bqxNon2HE3RS
Ctk1ym52r+g+IRcpw9M6WAJCpeTJSVFbg6IADoCBGOxNfbLs6+Fu8+bozeQ2NevzsW0HF5BAKZ+8
81Rfwd1ppBqQ0dWFmXTqacW6DL8uZZUsSvSarBxcjmtI6c4V1nHkvS2XLDTERBbm5XOMyd6eXskL
SqNrceXXUyuGvCly3h+g5BRY17AbfSMbzs1YaJuFf5gm/l8MK+8cRDjtew+Cw3P6oY1ZNRjAvF2O
kssEyVdkTDf2vj+sYe4B6nc14dV9FSYWJpCp1Oq5ZGMEsSSIuSAuDpir89D7mlDvrNM53RWTq4l3
dEcb8TxbhC81fE80aKdP5xsUL5icLbS1o5jktZJ8t1/OMYzRj2A8LbIN9XKHDNMKyq5/aqJG3+Ua
t7aQPso+q2rZhd5u+6RyzcOCvpZNLiDuGsEX3iKRd5m0UmgbDoLTjEZ+G0jilFTcXJBhCzPPei7Z
hCW9aQq7fjwwFrRKvAhRYlgBcjWDSiS27nJ8oQ2s3lrdUoiu9PUL1QhW92LFRzxZWZVo+7XjUKMn
uOoR9foNA0jvf9AVRwrJJ2Sba/XVjninyFY0OKv0QDCb2wtm+gMqCwuX5uZT5hUXRwhM+ZPnaB13
LDjRqhwgNt8Cqenr0wLL1SM6t0geDsI0rPXbEqHdCRO02CWyl6HtF/s3je+Lhl+xNQBM9XN6XNs9
zPxu+2hmc/X1xSlP8VVf167BiNEej9tDpd2UG7odwfOiZxHY3kci4KDmqPxa65b+kSFKmIdM/Nqj
UyvelY01OcoXEaqGM06rdFFY+xeybMIX4PtQ5M/lpt7Bj72gmVjYXdcGXcG5GvdMNkZNCvJI4K4L
zmD8VcvOAsprxZLcc/wSpkOiEllJQAXWjUXQsZhbMGHLawvgFCJKdHUzsp+15wspvCVPTLF/IB+S
z3ZUTkdIsR6SGk4gK38H+VbSvShWNr06F9qo7fz/+INuoWgCIseBlQAXOzn/c2X8fEw5IzySRkE+
maBjvmyff+oEvXZan/r1F+5YgAkjumSb7UI5XQONbVsJKgXkfOOFmNCMADQHxHl+wLMpQFU7WCJO
YQlQF433IA9eGH8eNva9pUpTp8zOlzhpYLm2cBdT21EmRjfJ272xmSZc+gq7IYPhWx0irF43ZD44
/4bGwsHA3RqZMQ8SzZBIWu9EAHcQlIEBjau2CqKIy5QWj+2lyrDst29Km5/ZdimQfiHdxKSTC7Y9
NngQMpul2IUw3imkJqP7feE/HYNd5QpJawXp+4xZP353y1cvvKYJRLS223rytRbQgzZ8IE5wC32H
az85YOcYWgFhCAjKPm8p4oyKNnoupo4om4yfQU+yn3DxGSHx3B83DvU6rxhdYoguDKpMCpv6O3Z+
3zEvadxbItNa/Xqjt8k1eFtcUDGZrahu+rAiJCNTeHBfgkVZoBxKxaLGTwSA4AkBy3qDaUK9gWwH
vMw7fqA4I43+igT9bE6cx7sQsq4/rfYH4Cz2i0k7juvjUZSjFgMSRNcwgxewcAT8S4Zy9lNR2Lyl
W849Afg3Rydgf9ac651vFtl9HxHumQahvgZy78ocvqNC5K184LUaup0MktPbjAK77qhgpTfkq6GV
nWqaIIrE58cTcugVcxlkeLvPmqpaPpN6S1CaNfVPsMUDpkQGNrJnppPuOcHi1q0ysukWLPQKdmHe
u7eyz+gCmcWJrKq7a9MQQH0HpWO1qTsqqhRkvyJdIiMKMNYnKqEE/t048obcfaVCTOmVGsuUOgKL
15axjNzBvHBbTcbOG13SdaIRPEoFX8M6RKPDhHoKCaIT6KSakU1sXkgtkzyPmxBhEvq4FpuEmKcU
skWvi7a7b+MNYLM0Y6nQFOFafDPAfA0s8AhC8yZ59HmbaV4lWFwhPEY5b/O1sSi1dz5IjF9uJC4n
fSMXXHWXtqUlEqzQsIZx0CNu1UgmA1q3Owj0chnfRuG/nqKzomTJ3IrJwQczCeDtA9Xm0RVisZA+
in90Hndqfo4kTjkQvduKKe+IRUZhT13y7PLBn8RwXUsMd6eaKCb35y9bAaWSC+RRXYbcnuWWtGit
qzFBiujrvfRX+8DL+MVypABksVsLCh/GN8jcpTzfrj+1V3QnjH2rxmefxl7OOi2i47B1zf2FarYI
DHL54ijK1hfxT0BP0wl7NOg7hPQkWMykofpkZEO6xT1pschC9V0lavrTS2WmhiVi7d0OTaUVWmPo
Fi1FXqW/cu63wlQaHm6tCMOX2CHup40zSageoP95p0EdYzw2r+/xwrmqcaZLNEMxjJSM3flCoJzs
34cjgXiyF3YZID1zVea1HQc1tdvpt4tFhLoLt/Gj344KqIOQQo5A30gXsKjhAUgo1pUXA3ytc92o
jW1ogUfrmNFRQc46d+0ZISJdoM9OLgyIGJqzMWEHVjC/sRL0wdjIOpP76znUw2NnzCL+iNXoVV5P
IpaURUXm/tkO3s1EI4wFPMi+iEDZy8xvW93PWEhF2NiGJRVp0I9BW/x07aL+9C/ti5SY+HEucB/j
igIsXHUChlpH4/Gk4nVoOLNb0WNhA9sj7G/QG1W62TycM0wTgBB2ji6x4WJtWdaKMwcKGaCZmgvl
EZ9ymUd8zO3ZxV4dfe8h0H/CaFOxazQBIPAGzYvIXA7sCWXfoB0Z7X7i5NdECCGXkE/CC8OTbO6o
agauAJn2ckEfOCpt1QBQt4bCeIDv9yTNy1yypHxuJvAv+WyHKqlo357iYA4IOtg7ZcsNWVuDSN6n
CkGQAAN6gxUByG2PeDtNzu0NwdGS4wL1/r/QhFYJwgj476zLxGM9krC4c1jGlGrOduG8hgB0yAk8
z4q7ZJ26kl4FHJ7LejEL2ohwQVNfHrfwdYYOZtqhABhkiED0gjG+j8+a4u6rPcihG3hQ0GgctqH/
URsZa99RZtk480lFPYMIWtzw3CB/OvrMvEw5wK4HzggJHwQT58hbZyre1+nVxkPUvrEUvpC0VoEc
CptBJQFjewhXhnqT2c2KCbivSkXrn1pfXZS5TQs1XF6cxO+ZXmGT/fBniqSCzP5tHyQV5/ThoGxr
MzqV6M5ql0uLuOlaNqC8WkI/3SakllJZr3Q9thHbFq2ycJKaEpPggwrod1GveYUSOz8sWzUOCp5Y
vt5eMNGQsUTYcF44yB2FJcRNd1Go7CB5Cidj5JYAHr0za1afBNSWRVcYWzneYOKEt0lmIplmAnhq
WCZaJ+vT8qC9yC/FjbhvNG3gNl0n2olmCiFvUDuQDOf9L1tW1nAmiMKCqBuSO3qMznb/GGnmo1C9
VX7GIBBWreJfCZHXb4g5S8RYYkuSL29arldPy/lKLoCuszcPKVQUzygSbfuKTFEj/kvoyX+o2v0Y
D3wTP/0oV8Hd6Cee3/JkphFCt2D2/FR0cZY3k68N5A3kO0GgJ6nrdO90eRx8yxHP+L+jbMgicPJN
nzkrvUruXOppAwB3ctlYy3GX8FxDq7nISOPhgDV3CXmM2FExf5Zs/lQHSc++abZRpDveGFPESJok
sIXzPEf8X2dEQsPyqY1uF6rxTn2DlGQrbSuYyONVBIGhAhc7cDdOVhx82ff4OyGdkiDY/dinIxWg
W5DB61Fp3GbwGwiLMVGJm0LVadULvJWVJkG026Xaq/GkIEBPNM3MERkSxadfDotL0EVR2XtFGFG+
t4hUPM4UTTVjCZ2rgS70wLlVkC3c0SXNYFQqcjyuRSf5kQORlioPjJL9gd9pEsdPTctxm+7pq7F6
6cG1ZX9dfWjWdeK6TjOG2oHjI/ucNxT/eGyop0KhhWjLLBDW8aixiCzrsdfAHWruQ8gyQ6V92yYg
z+2G0uiZ9ZULZfI0zzeY6QExJ+uM7cqfZbZnmUjVYzbCRyIowXsw2YoqhhhfXDIaO2SsftLUrq+K
1vqsQvmKPEn4c06Ha1Snd6zsL+76QBPxQzb2Uo21M0r/A05Nq1eqxrFPlmgCnGXcL7zAOA5JqWDL
NpXy19kPR2ynQXAFJherIJR+T+UTMWvgqYnZNzZZmzwPW2TuXcRGFB1dUatW4/D9/4cJNSRPV84S
Hq/ZlL4eBKOucwHMbWTrdHboPaq4AOtsjznVMiRgeYQ1DtjG9uI/VyFXTesq/0hEyuiNHsmle1Fn
vppgSNi8t2GATpGiNwrwDNMQM+/5eG3Fh9NMDW6rcs9y5DusrDIeZOheCBSf+Ac7pS66YjXFIdRc
JaXhpYj1Fafu7z3t/1uixA2H9aN6P/omqHzW67mE6Vl1wOsFiAAuxpDZ9SAQhCLHQvERSQ2b5CjC
SQN/hULCRwmlIl58jziHhFf8kPqeHzNHJAdDeECS79xGCB0uhVO+S4bu1GgNC5IaJ6Rewj5YDYcD
fKnYgPTAxW00x0TdnC0ICYUWIXI0hoB3ruFSbjr8TYYSyz77387YMTJsxfj9M29bLap9MgAzI2jX
W/1DoWY/j7H30M7od1WyIIBdZ6xfMWdyTsMxmVCBSydEdz5MILrtEPksojdDGYdA4dcOpENUwCF7
xaFC7tevc5adqA2hVDK1kNMuENyqcwaZECYMy4lN0WyHO/XzEMR5Hq+b+jPW2ZZU1vQqcmzplm0C
6UWvWB2cVLou8bg2GctkvqB8p2SN4Nb28U9oLYxeQtO+EXfm4dQcmGgOfc3gNquf0nZTmG/sISyl
Rx9YrWx1OETLjKRJHPHdUlZ4rWNnpVl/0Lj7eQlFwTsPdJZxrGq6NhjJDIql56wpH30cEnVT0t7v
HLHnjak8nS6N96OUyrEssGXW4PrM0li0vFf0l9vRs/zRutNpcNmeFljXjVxYtuvflU7+6dCVXXIo
OuSitl9EvyWoTKzEzplqgWHKeEy3/8s9olFyZEYVq0kvtrYe+C0tuj1YnteGmLejuHWqbDU4+nig
ntzioD0H8bfl+ez+Ku/J3r0We8oIjbwUUEMbcYMWnaRJDx0ivUv5k/9CQ6TUCn5hLkZw+/rUEa05
Uc+jCwdAuLqCEsMNEhD19dv5XnFj8NpVHLbsh0AL66JvbogWjLqFItMFExOSKTwxDSJQgVUJiQi9
nju8u5jSnyQ6S4wWt9qdUCc8zlPcq59fi+xwcq+Kxc+eX00PSKz2YvODUSEh/Pk0/qKutyNusFVY
2LGgj9Wzsgl2tEODYqJsMOV/GLqRS50p1CTGRPiN7LuG9Tazhm3qYFiRmrMWw4RstZIWv4CXku4U
eqSWE+C7AhBVcoT1ZPlVTsawWKaHXofk0x9SkjrlNZVA8XQV7nDE/DHJ/3uNb4Vy/K79bOA+jVLP
xiJwKZh4q8d+9MlQU9VwEGajyomLgEJGfgI/aJbE3TGuvuivthPpC6Bcbj4ugkrgSgSPhS6YL1NS
k6MnZ34fp7Jmo2evV2Qk51XQOkxzHpxKBBHzm5ABZ8fFXUVxiovjhPfe3MEGLy1bbBDzwowkPOUM
DL6C7gLKk6izTZZSfc7pbMNyW6wV+LoTg2+kphSGI6XW3OuICP5Xxrc9+BSzP50yti4iTAMq6bUV
RtjqsljRvBL40a7qfAIXjzTjCy2ZynwEGcWywY8AdwR/BlqdbEzfxSfhrh6iu4kQl7YLEPquhHGP
VujHRhUfyNTIcjbEVOoqSOE6y6HphPC5EUf8ZnNFN4tiat7Rm/cIVZewBeX066/1ZchHuGRGVXHd
+zUSfBB5pvEFRjjIU/W5HFXcsiXh4MUoETLTsh+F+T5JbRwLIm+ocXw5bqcqWQHTQrXMHuZiTKrq
wd94/eklSjkt8v7uXq6GWXqHO6cwcrQpwDR49zaeEbdYkcGAVdaZmtjrLq2XK9Q8Tko/QRCIU4LD
9NJZbbY97bbSnbXmNXxzpSzTStUYPOEKMVxE/yih43R2XHTEY4TSPWu7UtxHn0j/s8JN4jF+X1BK
6JZXfeVPK/+WNG6E8aY3ToF/CVjFo9eZGDaxvKOPy8FbKrv7ZfDcZ/mwqV0IfxLd6iHm5gjdTgxa
5sHkIXn0Pye/fMhFzvEohh/5sQfVpezOW1pYwd2SGVcMaMzqecTnZyag+pznw+GQC3X86pBiYFx1
dEKL34v8+C8wL3vo1BJxWzcxVBYulkpJHL4H3rx2QMNR4PsdOx8z6D4JcT0nCWsnP36/e6MmhEaw
ENxZwP0TCPLT9j7XYfMK37whA/5wOz3WdK1lo8ZCcCYOlQ9/qxmiGFaQlIYvOe6zVQUJGKmOnos+
gpsgtlkWRLIgpdslqZeoP/eDdVwEJJgHdIwqHprIIBK5bkwx7kOdQh75n8isgQ5hGVK4vwRlhlx8
82Dn6AwWNlvF6TJ3iScX+RkmyeWo/YKOXRQPcdfomVmfu7O5gIeZPYiS5JNZ7JXW5DmLBSi0LCbK
SOVlIXBM75T7S6HizQFb2RhFNO7aLI7NgQe0F83GoQMTbaqV4bbMYazlBo+TYdPZYLxnEfK4MAGQ
rJWDR4SN1NS5gqO/NLURHqdeMK7+3BumyPodsM4odtQVY7sRUin2VoWhqYJ6eWG7wGIOwHlNLWvZ
jkgPtgg79kEwmaKy850hQPwK8NTUvs9GlHcy3G7easX8xSQh+0Ks+fo2Oi9B72tsrY8OYeBqQPf2
GKa47YT2/f90MzXc44CDFVr84u0rGkXpl7qg5oE/NfU/ZY7IktihdoXff7U4x5mbm0d0y8R3Nh+f
KliOjoyXStftlCRWQ/SqaXgjurVdtPKJJE+/FiAJkO5MjlK2nQ+ssEyBQlnykkIE7LhWS4ov4vjm
1mfftd61Z1pxKBwAfI+ZQYunkM3ZGF48ypgNJhuuW1N+q0Tq/pMFPtd//IAcdZMIqRtaUb6+jhSq
Cp1P3xAwUg/ZP+kePebbeZwIC1xqZ8g8tyhAMTDpt75vDRB5yHYgHYaErZt1uSnE1eGV6M95e4vE
KlbswhzU9TGVLe54LSLQIC8uIaOWlxtDWHF/+JnH0ozYEcxk+l6jQi2F9abO/zo5EWl7C3mjUn3U
ExCI76PbtyM9NlLW5tga53i2bvBHaE9QctbDoyyS0Lh/INQksWjS/w99dwBq5v7lRsccKKBg+QtN
9RyQJ6GJKmtpY2UvBtL51U3ydGERA54kp/xlZ7CvALzJWtaaXKvklXTe8R/lShtUjgn1kY1ni8iY
MzU0sET7UorXCIklU0BKIeBfqKpr4jaL28fyQhIb7QP/82rr/NUAm7j7MtcWDBvBIE7fPM2cRRZm
cV0AtwU5oGXJ7iXyROggdmQQvgwOmyhzqoyB4rwuVQQYTOh9Pmu/QAE6wcWAzLW1BRi0Dz8s9JJd
fDZwsCUbnCM0IgTcoodOssLCXHU96INlJCrtdnE4093i58FSgN7XLntoZtwRCZfDeOQzfRWpVVaL
noTYu1CbCgteS90qlp0YtqV7TFK8p6HUjsiEtEx0uDCYxqdg7oIe1BZ71abWXsmPn/DdamqZsVzv
YAJWd038fkP0odgAaUV1PQED3P1i+k+oTh1edJO5MZTngk4uXTxY9Txe9j20bPxjDfx8Od9lK+Bs
xkSv2DhabVIi8iSTfz/N15tiLp6sWD/ephYJt8oQXSKRUez6OmpsIrgAxxG6gFY9a1Q53VBLZaDj
NDt/oqP12FY4GGzzrB1MgXYiOns14OGyKdwKKMjDCfWOde4PTLIZbYrIvyLIoS8ywPjuxBR9cjGZ
3uGSpDlOlx/73CGbDbY6i9mjWCIadsaIu3nqf/I6AEorRXCYD5R5b24DeH8o2wlVWKRjqfAXvJGn
zP7dLx3MQrLZ57WhlN/TR+ni/7Ja1abBak8PPC6snQmmA1AKiImZ9Lzpk6dkMwwph0zsGOTlOXNB
NUczJgBYLfLs47L/f0mjbLVxBeDnzfHsziSIFkss3st1Y58l8oCvsaBeLrGKHX/FUbQJfRvUeWXj
kriTQDdLCvT7bqwZwjRvIQw3MEbcKA8qw0CIBGnwgMnmDQVuXxFEe/t4o2CJ2EeODDTY3LoJA2lv
39EKL+NzaLnkUgSEexBuKi/68BqQEXjneCr1sOLClGuxSLUPDtUx0YLz3z4qEnRdSIqS7BWE9u8t
v8skzcyWXmEPWw8bMgBVIrgSTxlXoLVT594HGQgaMa9KWkW6ShdTgEo6eyhPE0LMbz3HcvvZh4yi
r0OGS7qa4dFf0jWV5KOshCaQNfihRCqUx5z5rlPlVKkAvfvaqi9e2bjr71GkxcJJSp98jgZStowE
l4dRuoqHvQYNnm1qgDYvd2RkKJKqOW7aWwN2iSZsTx/N3qKBB7jJhYLQupqdr5Z2CnhhEE8C9AFW
BIxhj11PryFARxlU7Vq66zcbq0CTlfUhVQ8Mx5LL1FK9lzsKDMgPTZM+SPp45Aaf9H4YZDsqPQZf
jeVFJe/uJE85ocSGx1DPQcJocmaaLohjj018+IkEnW4AgSAEXa9Zc150OutX27VjSCwJ1JqumG8y
x10108QuZZg0dUIEgLNAFpiVqiksDRRzLGiimI7C+BwmnsxrHs9XH5YRBxYsBRioxcXRDjGhR8do
s2aR8VG/EnSn9SXR/18tvOb59I9d6rQEFmwHGcugsbaRGZSpYM+/azTwt7FK8MoDgzzkgGLtwPhn
Q7/dA5GdsUwWxzg0rX7JkuvG17D32Mz+ZElMmeVPz2VHLcLs6NZzOFLb7jpAbakFxhaGjY4mLFFS
FEDrNt/L6Q5lGs6NraoNPnkxRXit2O+zG84rWiSZTlRwSXKUAdmEqCHrSU+519iOJ01iNiraV90r
JqMGVoalvFdrVh2n2j5AqY0K4/DPQo+cWiqmB2FOQXjdUryzAAJWNzGXlAocU6tuoaluPQgKcoO+
gs9DQ2k8DdSWzjUfd3TwnxvzJHOT8sie0TUpnUCaJ8a+WYYrEOgreJfgPbiZjUioxR+CtVm1XwMI
9bnAd5SxsXIFUyxggPatw6fwWZGlWYSUncpRtl6lt9YcHcBG1I++DA5W54WPHxHGx8C1O8xBUVgu
vuqW3JfJSKh5IkmgGFzsHzHmZ3siWyyLoWRAAbmMf2Y4eM8VumhJ8k7Tv1WIf++LgDJBnIfwddEi
fbALl4Zy+jf9n5ijJNkUyfEwq774hWjkZzAxZ1lVLIqTXGTSu3cWZ7g7iZ4YbJdXqTIgJI1jpi5o
vitk5FpD1j76ik6gj7FOEoT6mVsf8es8SECY9IgX972rQE8uxjXuQIGIrL8Rol6apqJ+TFfaX5nw
CZcv0V50IaKe4AOsXzA8mpTWNqirQXiq+P73IldWMbMls4T0LGfuHWgmCB3EDMw8LWP5X5pVON1V
lZruNGQWO7jK0YS+WaPwuzr85MYMGbJhLRcLLzzjBMd+vdRuKRL9Is+gnr6iyYVrCXM7NenlT/oZ
giIqfmtim623CbSt+s8vo8/UCVFjwE2OyKvbCDb+z/+Iv9ZtmLRrn4rtnjCzNtTZ8AbbkV9Auv1j
3vWLIL2cJHlV280Em1ul9tW/I4pkf2H5JFLZ799Oo/SHn63PKyNLp3NCTxw4S5d0NbxR8w1yO9Dw
WVrngufSe9swYUayPipULfNq1qevo7u2V/PQO+InkHXb/EfjgyMknj8t/TLkXLc4PSbGhdltRrVS
eJvzVBtWrYr51NfIaA6iUKCQ0XXGaqbWnml1MddMyx32BSXtKB6lmklXjyl4+ipQ5cP2n55GU3ym
Ukrwe0anJZGicg1HqgysnOQOdmpkp0g7SYSVdUxVLnVwhbmLooJFwrSCZsDXT57AhxT5NJ/iPyBy
L2JgnrYImk1J8su17tnL7Pob60L6EAQEeK2rwpjptCK2IrH34fIqCB3rI6UJI3uwNorbhQk3+YGA
QlvuzRSXfLsrN7250o0zvKPCKwi12EgSni2vtr22XNLta73P5PQ9oV4rYVA0dMbE6Nh4z7DwcQB+
sPiimcaJj724Z+V0hfhhFSQIsDP6jZp1xok7AIXsLc4ePJzEVEwYF6a/kq6ykQjCEvnRsnk8Ox26
XP+NjtozbJPgG768JSR903McpgrFtoRnvZsObK8ZCyzEbP1/r4fKzGWlLd1c3M3jKHyQVLiKBnNO
+RvrsemVdoMCS6t4uQlgTpQxgKYHpri2VRB7eM2Ud19mrwXKm4G1ShGaZGytYk3NAJ45KBsOT9sC
VmtgVxRS4e5HQUbKwRUXPU1gCnOQRWv6VW7wRhmnKyC8hZ8/StGtv5qYbpKZHw6p8AC8waWlalnT
kjR9uPyx9cO7g2tyXa6ry/QmQQ1zl1iX5VZdoCCqRYHX71h7s/6TgDX7BQFeyS1Q62sTzizWNiTc
fgo3ehJLGv72R4aMPpmCxabCObSWR5UWOXjYa3HXhF1dLXCUK3IvOuzu34pKd9vw0KwB59giOdVU
IkF8ieyGi0xWU1s9DuOez0e9wbEM/qirFK0BjlxG7Up5HR+BKvhZg/xVORPstzvSSThNANkLqMzN
63xoHBvKd8T6IpvIeazVCnH47i9ZQQUX37TwIG9y/DLyMcdzldiO3G55Nnfho3BOSg1GPcjPyRcm
cPEIB6i42AFdsEvpQIiU9fFszpyCGpCm03lQfl+kZjyrj07vvp+8DMP2dayIiyf+VYzZYA7arurh
AD9Kw05VwGFFIR+NQazos41jev6R2P0Jn1dYrsXJAA2V390rgyWhAPBy5IpxuazIkB5WXFTlTTW2
fWQ9mMOmYLffp6Y5bnMeH3FJpswuu94x/D74k9gQj/26IJt4g4p/QPLejypgXTYVZi3pa8DiRSNr
Ueil8pRCThH6J347oddraLJ9NHhACC4jdYfwxAMGLaeYNAFKqoJCUwui+WHIKA4Bj42R5G+Z0ju+
S+bx32aEHM6cSWjULn9TIvNrH45fohV1eWYL4LI5jwYCgiRFAcKxJnfHJ7jiWOquUDS7Blad5Ur3
taAEQ/xddopjYA9oTztRb4QFPejLdaSAKsXWJKjxcMYvFwFOzAwm8w6HwaBtZ0f/IKqtb/3MRoOu
32cumnS0+Uai0lCwKkyd6WpFrFTR053WBaUvqNogCWtshlNZ/KGRQ/k5C2V5qaLG0vDCygazQppg
BDXpztSVHtLEMtzB5ekAmco1jI23LA4FK2iNrePbKi/5ouAflmFfFhobpp4Q0XZXXnV/R4HU8e4V
dNf2cQb8dQSB2SJ8Bz518kX+0vRSkeGH3u3ZKVar0PRPX+iwf9lLVYl7JFPF+g5jH5nG4uwlF1bn
xHAOj1avfYVqXb4ZXdk++qYEm8Lk9rcZozGA8WyAcir8TZIbxmREFpKsicbqadVEcmtMak9981Lb
Yv0SSWNvVFyasPJ0Wuug2ozhwcTSYNg92oRaiUlrLqRDpMHBFDc/CZoQMVEsaqxHmoLjwoljFOS5
HOyE5xkhKvp4hepWa1vGNc6pldF5Dah+fzcHqyZncFUEkEWXBkb74aGkVPg3paJ06/Jz0I4zFzb2
DHIzSZuhQMm+2cviZtPvssEu9QeAJZv3rwCN4GE+NA/pYTFk6kCvOYvmW1AQyKJ16PoqxZl63O0p
PL6Q70VQywc++c041tX1it692wQjccP+uKsszfegvsKQAa/BRapfAslX8QSsykcrfObZoMh9WBU+
3d3H3aXbtvQrcsQw1oU7CwGcSI9Ds+TfUGVH5Umsls+apZb2o7HT8YfmUanvg/3XDLEmbCTvF0h5
5wlz643IEESYGvxbMQTVhdFqt56IBR5DtZGmuaobJ2f0yab0ZPlrdruThP/lodSAR5P3mPNNu/RH
LEw6HntU6PCyMUUkOFuRxE7l4sYtnrkWMa7a8aGZjc3pVYzmlun/qgFtBW3oosfnRc4VwqNAULyT
YfnZQA2opzdRsQ2GQIHV02bxTqEEs83P6dkHEvAjW4qe1MTQx2c1p1U9bbry5b1KDDDW6Iehzjd+
08NwcrhT8ysJU0tFB9IV3PrpkfiLhS+RuTRqvPFmqsp88Ai5QspcSm8aMo6IBV59iN/5mQXyxhfZ
c/7z9Aq3vPD+qlJ0gV2MpkBkgtbajiM3LmxVAc18yaoMoF+AUgIArg4QneOEmGkUf5JVxM0pILt3
q21Kv8Y1rZJrIcLy9dO1ZdFQpz42R4ZZc4dDiDCJlmIbxBb6+VPNiFzEPlUUrhbpR8c75cS3FpAV
wc+hvFiNvbYogqSzWjzb+9dFQ4YRO46DmrcCqeOLUuwG8rRIK7iv8Unws8Bp78z+6Znssq2kJgPh
+W4xz0vKxEccttjU5PrTVmYZCFgIZinYDOsCbucMS2DQ5x43b0L1QpFzliUTPjXGrUKEFWuuxhdq
QPs6KvjPU5bjq62Gcwyhg4xjKs1i0/9qh26ZaRdESbWSntO3+ag+XgVRQPnQQWQUqHeelfgf+mS4
I052u7UDRJiskEsbjRfmSNV2e77lXt0TvRulAne69iaXBjNfrYOrsVauG119JYvMoo5dIhKdjX/r
M7D78GskhURS5EVkibffCKTr2qaBubraWJFmWXSjl9WoSP57O9Wm/3aZRlEklTqdrr/48JLYaV2A
sfK/1dKicqBcNyBAvNgV+ypyNBFjRGFTZMr2iwNPV/kp/v9RHXHeA+0yU1G7aquIDTEj18r3lBHR
fvUXZk+xSfK/GuMSPHjcHVa5Mw5EWYdTFCMYlJhV4/SrfF0jOjpgd5zp6shqTphzYGaeN0VwEHvv
mwOf/iBhLEA5dxuZG5dOSUZiMbrEj/rg1GHWUzJqmCiZcce7Uzaa2YuSNbT2I1nLOSMLZgV85ER+
A1Ep3hg3FI8O3lqCdOMVUVIbySNXZz5KOrnOPiQ0yzCJXwNS94Hls3KE8BPR2pwx67CTbySLteOO
7vTGL/slnV8M4/PEaBd93HWPtUv5yVsYfZT9upe4oq3d9xOqb/vEFFJSzAgfgF4ltDEffPEkVs+v
MZ37WHfQNkQe6b5wgm+E+rNW1sXXrlVt0V4MyBksEB8yAmukhJNRjdy3dLHvZu4u16ipqooI0ty8
BW94j4XTmFh/yfIwBXKqE9qnWqXm0wUsvNY13Dl4woHixK0bVArUVZNJ/A+TsNexSagz0TNsfGDN
wwVRx9Nc7iulY4h1WC/ZOpDzDUL8JLtnkZaf/qeaPOBWkgW+/Vj6/0pbEH3q2KdQgttYR8EiL56R
+LfSnLcXkIPtt37ip6HLaTCpKyLqh1Ix2pCJmiwINH1hTILcjzh3XuVBmcqwIGVa5g0fu2OG7nqg
o8x6qjgxn+YZGGgtIx/Fl2lypF3PF0rPlBBafi7A9DHQwVJgCM/HjNgnXhcY4fFCZSnfoUGNoBj2
rATIMsVCgNzoVGk0eVM9QbkslhIH6OLg9Yro+K/Awmf8tj0J7o5mDOA2xS0toOqUl0ewltys60xa
45ra7EGEozl3HnXUPcn5Pqfcc/7K4AaaZmKdh3EUpWbpTv6m5fk87x+uY01D+5wSRLzSep5hTXCC
zLGfJKwAKDOxTiW5eotixk+CKfGCzW9Lm2nNPf4WyA8ObbCdNo3Enc410f7aEfKWF4219QTrGEFJ
G664gOWqn1dLkw2tPWQxxGvNkQute6orKBGNDEwk3p41LYq2ZpEabir6GGFo0HAv8PNGRnpRuru5
9N61XcPn++ZfhBX2h9uOlFXEzVvZSV4tlNQsWB+a+vkOiDVGeQkkO/vZCA9LDqnPCXaumpewmbnk
QXTjk+5s7gkRaAbSx4a1KpvDEwvI1iaippgECG3dwwn31NsZBv2cI6SmYWDivxS3RxqX55cew431
qxVA7ix0m3OUXlv34svjrvy0rowxrMxSbK704vWBd+PpOx/3hcIpHCB8znttnCEjV3KkXtm9hpC1
klXYR4MqZEZCVwwYo6HVcpuXNFe0qlxJ7KryvNaZK2Bywh6+YBD4ZYyymrdbth934btbkkqLWi6K
oxo/0szBMcehlfV4N+UmnVhcucXnSZ1U6Ee3nBahNGhKJdQOp+WvCbNF2LnLfftLby9M8cfOGyuD
IiknJRaYq32UzKE2EjIlPK4TPxfq7EELIhEI9Fqv9R3/avMYvpvCtNqPhVyH8+Rj/SdCXD/7wML7
FfepEa1H7rh8wD0HXEvDkam1ZaXeMHS7VdctjLpEBs4858j08x9EEmt0MmyU6slnzgaCp9PruI5K
8KFrEfsvgcTdqlZdqmylHS0Tzl7r7EFXSlcxdhvGjnuWjEgPo3gQqBRxC93zsQeWx3n+oGiayheg
vWUuSRAbixPWQXizCpSqZKOGmyj46fm3JQo3D0I6Ms4vDKl6jhhq9ytWbmb8Cy7An/pg1ysQ9O6L
ftPsCGOi7fO33EYFjJXvN6iieYrHULXAnAa6mbKh+42g3lIqIsLVZLO2ghgnJQVW9HNWHWK8a4vx
d2Pk1nIZH5QSod5Qd31ch1/gNEueHI6Mpw3GshOis1W2UEvT0yqJLxS9sRmkgtCXQGaVTwOhi7+Q
gE7E3rCAcnAEiHLry50Oim0Zn+9R7nhE6RAaa0FwQcDdTLimlgDGYdpZu+e56pyWsLL2WoY4hbV2
vs0M8gFa9+TdB+xABoVHjWvh40ftNzrN2cGqRiiJ7mBtG4zDCVf8kDRgSg0Qhya7BxVRZUlequJT
eVhvyzIwVv4UBM+qtBqG6AiqEdzfuLoupDyRnmp+KXBKzQRr9oIadyXd4T4JbP+qEVXzLc0hC2i5
UKm+aZjp6Aha+GbV8xSQZmDdhPdPzJ4Y6w1iso+Vm0Tv5wAllOjcwb/f8WCPZ817Ti5iiiMpHAky
8fefyXtcJWcMjEAU6Ylu53Fc9pJEBEW0I2w4b6svsp3K9P+KqM0RZStoh+Z2218r+9STCHXgsJED
f6PREOVmU1pJwwsQB60IRCoWjnSt40j1iYyU6fJN5LTCy/JDFpfXZg4Ayssw0QCRiVshFqi8xTdT
tph2utO8mXAMNM76umRVENbGO+hSFxVI1OgQlsAK7mXjWC+bAr1XwvAMxpziVFK9B+5QfmTwYoVs
km3Kfb+IBl51ZUx7H6aL1Jt0KhK6Wif7hFtQG4RQt3Y0HCs8wlzgMFrlEVlZTR4oyS+DcI2lXv7b
9g5W/1bC95PNNPLNoRk2ceC2rqMGX4hp20DegeQ4xl4dzPRmNYE4qdM6cGgy8n8+jz5ltZ5tTDUz
T2v9QYsK7J5aobX3+iNwq9SGjwr3Pl7XyqCjOWQIlXd2rUHPUa9v69EQvvEcIwgWO/9GZiNr1sUp
RvMRY8q9LQTGJBoWxpfoehY20v1VMrCBzUiyIgyYN+g0trwCeyqH38lbThj4eWLHzHRiA4uCGjCw
U9GUFWj0jG55sUSrXtqxXUiOSMWrAQWmtFzy1w0updc62AaftAJB554n5GBrfrFd7TS/GTmbbbCU
b32+nWJj+zi4HcA4o11Ag3JR1tuFjDXiIOrqQ7aiJq6nTup+ULuouhBmR8V4J8fp8xyy+o+vHX7X
fr6OCg0WV7nSJohG8DGBb/5n/N4gRZcJkBlItSHqUNc4XCN3R/xwJpMhtPG++4bhfSsCnFk35/W9
mXjodVZyPAcN0oq3OQDsV+BOcjxiHAul8DOwXVSY/JZzg3QHRrDQqPc17pQ65kupT36oZnQwoSw8
WRSGHjXMVeqjh6J0X0A9Yt0qvG7kYNfe7EBp3gwcaBtVZtrZel8FVpv/HXzJxifb+NPIu+HiZ6lz
Wt0mpF90JbnEovRJON+HonQLNXt/z3KvJrFnuOoufCGTuC2/RNiO/Ada0Mki8Hoso4OhY/zQjebA
rbwoqvig20MVKpshvNZ/+BPRon+xVyCXXbphqjrbPvLcD+CI6kulz/qgzf65dVV828wkEYnHo2ci
v4E3XZ+1ma+D2AhiaFyGIorWCOsg5fRx2ojV899umtVQiM2kw+5yE7OyZ5LCgeaL+qLqB9cQzkEp
4ktRuCXJ0Loq8qLt6mg3gChox8LbaiGW6VSVOTz5sQxguf9tozoCN7+mjK7mqGwJaUROgw+ufI16
c1KWlH+ESaZNj9o3Ijz0WAiBu+T63kQQ1qu3pNCBSaDgbIau4L5aROb298M8EapqAxxZLwMZ6xuK
qlrB6Jvm8DS6W+jL8jZ36kFHdJ0UWEFnmDBQl+CarDulNMwooiFplDbOsynbFOlISJm5W0l9pwux
jqpPjNrOZ+JF3/nCdT7VnpXAVQYQfPrwgXbZT3tmDn0XiG/qSKQV5G5rQSlSSYpK1zk1SNQv2i2z
jbkvgM0gVLiTrNUmuhXwzo6z+GeFeIDPnbHh1WKbRby7/6BAVCaIdi8YBIbGHuuC45owdeT0GVbT
ZAxLvWp4ui4nhWDN/lTIfq72DBdfwUjpdGVU2Aze2SrZb/mv7RdXzp5m4jciP8FLtU+wQkdjyNbj
WyxtKy9C+VIqsf4I8qODF9tljLNIxvK1aTQGO5qZLrT8YH3vMrzIOcY5XeePs7qkTlCkOS1WMCFn
FaFDpfH9vSbsWDVIxND9i9MYm3hPGw+C9DeVqU6v24Ns0gBcDwsGzPY9qVQGpBoAYoCH4hIh2Wvb
CQmiPEFGoHAcfs+Rh8SQpaZuq3vDRCTjyDVbrjnTUdC3pC2x3vU1/7rhkLcWms0mSbPCy1wuZEHz
dbloh+EYRuvfPp08/vji55aM/CE5NtEsUaO5CQ2M16S89ReBXBhdszESJSKHHrc3eMeba22kWVw0
pcIQIi6LE8fCvwP+Gbusz46Os7zEfj7nGm2KlOqO70ZSSy8mKIdnhZWjaFsHBoyUwvNyFM5vKBSS
qx26abj4hyq15mFKuGzW/hlthxZnU3bclQq/F0nV1t7THPsLz4iSynlsy/eK+iSt2xr/Thcz9nKv
rbT0r6LfwTUimLWJcvAhiRKu2camxAnWLEmwiUFax5vg8LAYmxEe+b7uVUiQMMnEwcc4msiJTxnS
9TJC6ygCLE0ukLeq5UfsWLOHT3SDg6vep+kMFDojrsrLO/xODE/vIOKGPFxDOGu2K1RKmELjaAr7
rbJA1SQDtyZ+qksqCxp+WrmdbZQgCOP58Dh3wgOnJj9rp3UWXVnU0R28pitwYkdNv+AtRMujV8Nd
fQvUqADHwu2dRa0OQIjFdBlgbr0+EDgDuEUVor2qavdTIuAF4LE27NsjZ2stNQ1uXnAuwri8BhPl
SRdHuXsTx2+oBek2PE2YFANFkSRWWeDVvKS2dc66be7s+RmL/O3DYhxOIZ9d82zCiUxkmcwuOnPN
F28DWln1kqPr/xvgoolPAhaplDGNM25//3JxGr/2PptRjMKvsRHP30ZkLfDDPedDh9W7A2oxO5Ky
+Zx8dHkttStQX9Ou9N9RsqKTJipJu79ZsjkE1aaEn1U6ayb/HHprW/6LBScbY3o0um7gVzkpbP46
vFkyXnPa3EyhE8qqzbqEL3n5bUtw27O6Qcni09/q+iXGxeDDJPk8ck07ZmO2PcPe+cGSaWoyQS2+
dB2drZVZ+rlkxqs142eHDgE/zSL5IgmD8IbC2r7ENKWWEhsyUSRXCIN9AF5YcmHNWRPOW2iPpYBt
G/bGsen8Z9Lz28EGcqrv9Upr23S1vubkR7GgcF969RUyX8KU5g3Z6CNdg+25Z2/+XBjwdw57kV05
DvlLFUGAbAU4QIuL0yclLI+Etm7Dwb8M+cLHNuoY1ih5AyMhXRRK4fLFVsZd42PK8hBBjmGVW6Xl
obZ+FdyasxS/7ed1oYjzNPuI1uHcmzRIDeXPAuoyCVXITkfkaN+mWCHEYDioB6N0vk1mCucJCVk7
CfROkUNIlhkHa5N9aqDCoDFgz8LbCusm+CoFpaeoA8eXrbdwuXsp0GC8KNzA98iab2VITUpXXj3W
s5nZRIyr65yNBLypT67X3flckD7k/L3LmMsRahpjzCQv5IbbbGMGcH03SUpIYkX0DT3LBQDcP8cB
djJwl/pnaUpyqEqT2FlkfBConUK4XB5hDLNDVFw8t5K5SV2Ei/wQWqaU4ClGw0Y3vJAQlfWA3tXT
oGgMYOTBM02stLD5GxiPTAiUs7Fku5tDcHSz3/7BfA1wJgjfaryzOECw3Mc+tei6oDLfk50IojID
BsworG6m/+BleHNwIbEuE3RerqRJmDrd0jFsub7WyBNceZu80MBAOmGNfHv8ebcDc0uH78K6728r
Ezc+mWhmHlC1IknPqNVghJ6ON7b1yLe4vmv4cT4K1h+e1WDSlknYMy6tISy+84Uf9GqF1OQ7djZq
cz9iDSzFwmkero6rp76q22+pcULbaDnivDDxKojzQ3OoJZ8s5s1FjBS0iYUt0IQ3G7GM3b0Tx8Bg
+86F0kyksubSDq5RoRx2T1vPXrAouwwQSBFhmafwtcV6idvIiD4MffHuHuBF4O4xqNxnix7+NmLo
9nWiffL5Reg7IJXnN5k25uU8aFIgqG8/q0AGGWarSyeRj5XbUt6MsMj4WtwuHcrjdZY63LUolvwb
VlJxqL7/SiRIxCUq1zxuq9AYRkGFIjEuK9JQ+HIcBJHfGZRdOAUktOzq1yTtOfKvYTcHTjwpLoLH
9455Hmps0m7Vhqm2FxlzMgf17t974g324xjCDc0Y3Hd9KqHmJg8Mb0hD9rpREC47DT5CFeazTKEN
Pus8J4sRgqoNd/PkI6Z0wZUsldLIH/nG6O45Wqqd6c1uEGqWo96149hzrO6likJFFJ7zGiAl9s71
RBBppBU1TJ1mWxotTOj1tQXoP1JlKzOGFFv1SZJE4PG3XawHn6As6HvWGI4SuM/6MeybNRQjx4gh
D+NQajZP8jGDzly4cbxHmIjP0bDVrBcKk2P4euDc2sqEnjLP6TNGJF4EKO2GfP9BDXNI4qXzsWmq
Khc3JFtTfS9Pl7ctrloUm3fIj70vxgimZL8cvTFZtbihFZikFR3IWR26L4xGOvEd879iYS2lR2Du
xqB7jarvvzXsbOrEAAAgsBBi2TRUdUt4SS8xLVPz4OQGuxwANP1O/09bE+FLe/xEKDf0r0Gj6WkF
DM0CZv2/MKzag8IPPU7fUIE4dI+lqbUkcODEY8ZXGnU7DDXuvIFO4uvgJA0GC2eiHBkWZU+9tJuL
L/WwvCpvk+R5zexxNejgZVczv820VovAIImIgFWkYUXGZxrsy25/i1jdMAixGiD83si1kOYXNRGf
sA3LMjFkk30njtE2FzxT9w7mnpHdzrLO/NNTImI1Xe27+J4hIVJoCEqvTkXDoqPDiGQNS3QaDkTr
x/GLXgleHq8LiUZzli2liGrTsBUEv1IFc3SXkJYoksehtAbB4haMQIInkgW66EIobu5aLjI47SHo
YFVibG3oa6bQmFg1qKhj77E2kJpTMiPBrZftv2B8yUxmlcWBv9WqEbXpz03fK0+mKIkDXKHtmGh3
zVtFpiYNC1TteaW2dq2NQI/xBSOfgR6YkqtAAAIHbr+6OQVuHF9dm6orULqcB9LtRNEY+qkh/JqB
fX6fFaV3DgcuqyYV0zP2l+QiGrzUt3MCYMpfXD9bRn2e1Rmq7THHoHRSjWrkWByHSuKLFfFisOul
13bVNdUE+P18m9PB0VyF0sF0+a2OM933Hu3H5LxsxD5+zUq8aRwihVP2R7+9q0kufaRwf1JHj0IF
6yfc6tcGD8umNVlldiOxW8FLTU7e/Vm9xzmRa6LaM5RUDP3tlLXL3ewiEUwgwV2iZu+TPWA17WRe
ek0u5OUoeWfxWh/AF0U8UI1gYrJKxn+pve5XV8NhUKKvxvSdHzY+D3/MpW0A0yBoyaKAHQD7Va0G
G4iYivXmUYfLii27KeLwccgiOoX8uEPtYxUNhFP+lPNxP1JHp61N3ZYc+Oal6z7W7LzgZmHKcMu6
SLcWpNWO53PvFMa5iS62cCqPtCOe3fivaPIu7Iz1lzc2c73JhlWLQ9uh4PXhUzfTWUahXHA/qgCn
ErtZO190ghOiO4xjDXocl738U5tsmRO9Lg4sbf9hY18MfV9A0ty8mST7+nHrAR7O05JJOS5N/dxn
LWRsKXT5P21oAit7qXUsOtc7peGbcEr8uSDgWrm0w5jK+8Zt5+757gC5srMYryFaLGCbwy5ew14z
+lObJTCVk7X9hqkXbp5HAYyQ97tGFsahPgs2VQZ+BgZbYaiEvsI0ttnGw3DW02NwqSQxKce4WULJ
0yJK6AKxz9boKV7UuaKbpB7HfxWik1jg84Q/xpbJ1ocvXT5G9/uu4hWkqGc+80uf5QwWSiGvzlKh
Abld1+vWzgpVvuEGs+KjE5NWdG8r/hvdtYClOuuZnf+MS97TMwHNaHYTi3ozu9vLJ90QStYwOyJx
J8ujaHlPffpAHey7X6GT5/5tCO6iYYwhHUyDLW+dnxF4lGUlyk30XJg/wlMJcG2MjO7nTUV4eIaV
yUnXidRhgJZ784n92jv7OYJjoPc89jOy2UTRX4nuKK4/Gc+oefAUdGohbu1qujxPT3YBz2v1QKvd
b3dEUxKIaaEM7aEJUoz4JnsvecIDEl4jqn46lN2XzFB2agC4y7wgGyM960IhvJH/6CkwXt/TaXuL
9V2kkdHcLRojR3a0pCygrNkxI+bKJjbF48q31XaualgGtfncDO3Hxjb8R3aHVLllopLXge+dLUh3
r7wjEXEgUKZEDVIPiKaDphazeKwZxSiRF1FegsLdth+HT9cPXBDvO+rjtMI+9f9A8/DKrEwIt3f/
qTVRuetCrtpAdgaw2186do7x+v7UyoEuQ6TZ4oDFttJA3i6iOS3Ecgml8IE5uisybTkPsGp6gJxg
jHBUrfmo1Xs2LIv6dZkec9lb/fZJbhVC+AU4rI1QzpxFu6kT17iIxG7oRtNuHaL48RdJsbu2Py3g
mIrBaErh3Sh1rk8IY+JfqCiQdeiFZwigaCyIaMSuGfX0OKIPvBznrjDyTehuBtl+FnrOJcqELzsr
vumeP3Y1DJ0YwahSs/1NdLp5jHHikYK8BkcGT6mchhLwlbdryr3t0pj82QVsVJAssG+V5yHblpCv
DZ8ekckikAsOJiboxCpO2O3HINmjOVG7iHEsSxUe3DNGNYbgEXatSod1oa1Z9RoKwrpWkGFXPFxe
3jqcPeUKpnObWhF+T76zso0BQy/JlPZoPWzzvPb3kmSyQx05XI5nz94RTS8vItguo/Ais0fo/I1X
WbapsXXCA+Vh2ppgMEemOeawKGyToEe2pMFYnJ+pQyPImW00koyEKXD9Li7PX/egd4fKfuY/c8Sq
ed4ZN3wwIiLw5IAC7jvZZU52ZVwm4gop5N/sC6NKD3DwFM+3wA98K33mUdSnGOcG+bTehifqKeEP
kXwvkxtYn5Se/L4/wn8LLTtAZPB2sRI2H8U8Hutx8KKLz/czofJt6l2i8v+0k8w6QAaxv8qg7nvl
tK0ixJk0WCcjp/rNZmW+Oac6N07m8R80IttjBdCsmefjOFmTxwWWszfb6ILUgvdZvERyP8d/CH34
oy6vI4hFDj7QUJOHBxFRQVtx2PaQQMkS4pCuNEmvL4J38fEjd2khbxu40K9/t6gcGicclG/tV5wX
dxhVW+6MIdLB5wEW1p9MvbdndvaxLCJ1VvgSFMErPQvvrCDThvwdkuUmAnj+Fwk6MEYJrQh2E2JE
3mPIYn6+i2UIkMd2RzWfEy980SmHWb6zLgcres82GD6alTYDKbpg8F8GrXneHNd3W1k2cZhHfURm
+jHDZiI3lMGUO/VdGR+eY5ZDCqnWoZF3fhJVopUViX1IAIjF9AyTKpACopDhGfd7V2wnI+VQ2gBh
Grz3B7rW8tPEKK1GLqji19RFe4GUKnAhzcsuEFsSgVNQwJFjU+idUJOPtscESxHmExjEYavZ/NIk
VAiF0ZAENVQajnu3NnFMwpEYzdV/dd7+6dZjdzVuXic71z2DFLMtgxSKCwhfpy9wewcIMwowXVQr
fDHZPRK5/ff+Ha8PV6emrHcbiM0XqCrpB/Qg4jDB3jJIY2lvNopX6Ts1pVh5zhkm9UBhgokN25HQ
kHP+NZSWqGOtO2V7zfF9mzzz66Yp+o+3HtS+qcex5z+BifD32GxcZ3C/6pTLVpgWPwdpmoQhVYl6
WhvE6ydOw60UHjgT3lEcIi6aNPHwd3xYVKX1vtKP2sX4Nu9ndvIJGsONP0/IJXskyvcvq0QhV5v1
rT9cVGjMqsTmR6YkMx6qfpz+BTmXfiljRf5xOCTNpFMlcMiFYBqS7pjzYF9k00NAwMTjcF2dBEN9
fFyOVdeykBw2Lm46debZK7sVvJpE2cRK+mb3DdY29Rzmvi0cEnedgEN7PNEuF+r+4suOkGNiMuWv
R1TfWPL/0vqD4ttm1jTroFXT+8bixlQGxtHaVRfv6WWhonki5LOJdIwFcS5zi8fUDy6PZiSOm0mP
uckO1jEqF8EBSNdjgbLrfTTe5KmWTBNVsiQb75fWWrOzDmGcs+WBdm6lRFTI6kcQ6gMMX2BSRd2G
7MHBoOld7VNQwdMiekv6WZwPjpQ7Q0qOI8b4MuT1T9b9ZwB4576CKP1vVTfxfAXrxppjHT2ck+eX
L7IHT6XwjsXZTPtBNPmI57mhCg6vtm4ihq/XQQCKF2XxZJlbV20yvFRne3bQh42zqfpPaUOsdP/m
eziorsz28tMcGVDxT/7T/ElfxMrlYlCc0bxmRLwVk3oy3j7eyTAy422CwDDBB9QBWacj1GVceLO+
ugaihrPb/hSaQ4ksm8vn/8eMXlHa1rSx7PydqhzuC0Sr5FKhVEKqtf6WoMvmVI9dD/oLjswuSpMZ
YF+8f4NEKefzxqWmiv0ktYfgu/zh5MnEWkJo7fJoRITm12mn4P+wy0RihkezRSutc0oqB4HlGjE2
2nKBu2MDCBUPaXW93pinWvjr0VEKQVPqWI/o2HEtAljjxMN/sSimluJBaZCuYSBU1J06lTLw4ahd
OI+PYDtUNEdAR3hOEM8NE5tGFQcF4IiwsRwQnrqMWvjd2g4y7ODCJjLlQCrSdKIkwAv+K+oihnve
rYj+jR9cp1IT4lZM43KqzNW79iPIayvcJKUpyf17R+Q3JG5dICUdeO7KQa/BeB9LoHKaDyrwezds
B6ObSb99AF72+C4UaTxt+2QG/Cpd8yRjUHoliGriOAGtSkb46C2SlXVP4Jt+HrgCyhEy4a8FPOd4
cWIZXXwoBCEm5Laj5fZveSVytlgqEcqci/OcxHfi+kME7ofzW2qLFpG9lxIK1nR7DF8k5wEXYEvP
941OLSMjA2c4iDU8cLouPBCulkYiyl3/Lro/LygtlfXD+2CoLXhEHIM65ZPs7Yjpj6zMmA/WDqcv
EhRcMjZ6Hu97vSj5JU3xP6mSqedz090bJXZXDkabeTDbzv4AUXupoeQ/gdwT+xFZbXqlxebiTKKe
LbW+Q6bjV6gkKzuvm+cKAkQCsnmgivC3DRWpe+oXXdYW2hoWcIATwOGtnnqH7eREfx/iq9qV8WTI
055hTkGiLvCeeMv2y33uo1sLoSDGtXN+5qNng8fL4Jpz2FUzHI6cFOZdDOtPtbwVmQZ1DVNPqFlx
SOi8OZ6jdD/PngoAddCvfc+nk/8OB3TTKd7vm4dtHCYRi0nQe13nlLjLxQkG9KY5T2feNaw2Xd69
DQPJIo0t4Aj/oK/VYU69Lx1RjVhVWZBo+4hWKO8cF/6QL81WBFPIRLwKEIRUoYW7NqJCk6NYEc0w
1aDspqUcb3aBS1dr/8S/5BxgNOKZwE2ran8izzcjcw85a9ZbmIixIgsCbsF5LjHLOKCFwmrDlGjV
9xIcNqyyhlftrx4RQFp5302JQRd8DEnesJ3okvOW7MKbzraUzLyOKKxhwHQsN+sI/lwv+iYIkdjg
R9bxreQL0rHD0VMa6W+eyPFSv7N2nYaajM+Bk93+jv+9AfpmGzRiXZb0zaiL1FrfRZmyugFbIhDm
vKOw0dfVPdI6PFnxybLXgIyjSpWf8rcKQ/d0zv3U45BLlO8sSWoFU0UJobXMiMqsjqqIcUdAbzzq
cvdgfUCFOhMXNgUb/vPMXT3w9JWLwXdFZ+6+OlUp5K7qAi7V5C2tIxET8eYuTR1n408WB4w+xlxO
EXoZ67CgL/mr2mlSpOdTmgPy5Wi6+DOURjXNd0HmjQwI9ZVNlalzyBWRcUNnHiQiRB0sjv0CLF+W
Jk634F5K1k3arb0pmag/qrVfhAya1OFtqBp7dxSKLkbmbDixVs5QbO9Q9q7bWCfLbmkLPWf0VJum
+ArZDL8S7p9RXZOxD/KlSDr28FDe6wyGo456YSM73y6n7rasBkb6tZXdLbRkV1ktsO2hXuWM15mx
gEC8FFj65X7Ua9Fqg6U4neyjqq25H5QVJHE859lGecVX7IZx0TFVzESlx/2wbKywBemnSjeyMfiC
xRJBrXqgyLPWYH+z6mcF7c+9/MsuUmAEBEYXlxalEwdTSw3e0IQU8hdd5NNsnYJWi1R++QyXR0JW
j/hmSjpewAuOM2KHLUBNZxR451pbPRosBM/XredmeF22fV/g0Uz7gR0+/rxV3d3UGyLkTJdz8jZE
F5SP4j03h7YpF+1Z8jzs3iCwb1eafovHbzNs/KVSjamuUmIOBvxZN/q9F3mz4yqWo3ouFdo4gGmW
a9+r6mohesF8arNDzyXQyKTCLsTfOpKDUeRkOLUumfbG60pKPXkw5YbLh7OECTJ6SivMzZBr0Vjj
lJ6dzQwsXR/vrPmwXS9DoV1+kMftkXTsuhVwmLSrXYwKpkaWhaELKrHTo9jbSbpmon4O1aKvufa2
2O91d0YqZpPbuM6OmlYR6rarZVupdMdWpnrIFgByHPNWgSqUk7Ri9QVfgD6X3AedT5uofl7EYwL+
zRdUWda8NTSoEkdmRM21NekxgobycK1Mw60u5xJx8AQA/e1ko2g/HNXaBuCalkB0/W6IwPliurYj
QoFR9I2oY8/SYJdMc7gyyJ85jJ9d0kSPKa4VpqgVlAz0jqhBjuH8A7ghiMwNPGGzTMpo3r+/eKmU
igLUb5B1RK4/hGX0AZvi2RbOS5z+Mt9HFoSVrJwMX7m8tOv77/Fh3jXEjRPDpVgVqE+2v041/FjL
qsZJs96NzA3OXGz+31m7VtJTLpYHMnbSQYTJpuruF+FawSrliXOH+3YaOwIwFqtWPr9URFzDqcV/
1uIi7oZxJZ7b+M4MFOA1DE+tLGoYWr+fV4AZaKGFSzSBIIWEvzSkzz1ho7Ra2L5MmIoaXnoiGyB6
M8GKHi6g64pg0JNT3DBB297iMSKoR0q9xvJMVmZqmYvro6zCgxgu0QuE17RZvKjvr6hHmsReaxBy
KrLef0jQgyYktBlmAGNykpgEIZbea2vjhlkz7uN66/7/ByItGAnk1jTrbYkc5pgLDXI6YvV0kv6v
ZNoTUE2By47Lh6rx581cDN7Apun4XRdTTdqZNumCc8fHiqI3wOqPtPZ7XTPeszMCfjkwuVAEVNoa
8TKjWlsIOuZKTJtpholoxzTKInD6nMiydPDkU2fzq1J+JfSNCdHQgHpizM9N36viZFpyTov0JZWc
hJTz6P3eGjefTB8aXgO45Xtv5zlsvgw4IkJHpRzmOqMEQS4v6QmXkd2/Mz+OEZGuDvgHLU0DuRV2
h0RbaabQn6LWlIinL7CcCcAcEuH/2++xsNpq5onOmwHjIO8aWcbaRRU9cIZ5Tuya9aIZQQwBn+cr
DqZiTTuOKoPsfgfsYtFcuoTCXkGLfXuREBhba7ZOSFx9/JxcXmgY+pqGSEMuWuPnRYoXoOlG7M5K
CbjKz9cML4EBqbBV6YHjmOpMhdBwIwa707turTY90Rjg8HpgCAuygsU7X54FLQzSjUJZmqQU+VMR
OXBRoe4KkU+ATPQRHBli7FYuonGmR7Ib6LywyV73VJ1LoZLnDUm4viGAoY9xfn6IvXIl3ESb2zEz
uKlkd4KAvezy2pEqMga3mJVKD5oPXF4J2IsHUmXc4YAEg+NhdWegpiqdjcnHxSmVqLJ1V+vDrVRG
/uZdKzVuIClbEG9yfOB3w2JLvW09S7Dkq+PnLuXK4sOOUtijhy3c8zgwfSwK9vc3kNs+w43tqjqe
0H1K86Gee/W6QiZDFFOgRbst4qfsjqNule2E4yis+No0Ey+72HtcoXyoT276+Wm9alEzLB+gU/HC
4C/a+AkP6FqhchQXJROMK8LC2EMRXwc56vMOARGzpY8s+8kVfDmIZkSrbWef+hEDmhr+ClcDbxH9
myrxvYA6fdQmzGDQJFjoo3K+KhLRTUhGQneHsB7yhYmFJCb7MoPKSUpEAIzASpKdP2l+HwGza8J1
flylVwD9ivHWtIQPjuq8uGrod9RxHpoZOjpYU/jVJhNMMy/0fJqpiUEfd+LE/p52/Tf+EGvNqgTb
3G2bDMk0pDS7BipoyIweG74bd+NKbrlXFVZMRQxh7Emi+DD+pkyPIFi/UiaO5DNRiMRRUvmOCBLq
vvHDLLZNILoYXQJn9p9PqzfujxJWeXytzg3F1+WSxiMq69EkA50dgsAEcLD/L3jABjonSuFlwHZ1
E12vX0Wj1f6axZkOsAazKPdZjiWazbcSaoQ2dIHzkyTespTg+0iHnv2DN8WKL7bMWIexuzwHkRJ/
kR9Mp+2PUH64eLjEr3emR4vJg81whodXBRo3PPzkZdwhTxYR0E9lHWwDHYw5A3TZTaETSPKFejSz
sJ2sTRoYiDvUl5XTfW+CLOLCGiRqcCUswz0EG43xwaIqKcesrXRynzW2w24n3QDyL4LRScBUluKn
Jm7NTzYOzkRsMh96GzZudGIRPsVXlBueHb4mgGiiHg51O30bWljmIEKwFgHXCrbU81D+bn1Czb8b
gJMj8yyXEF00QtZkH1bSDe6XUNTdAsVjon1AMsdE2U0TR89WKmNYxqJKEDcgZqu6HmK6o8jAWkKu
3ATAml9GwJnqv5k3lroP01O1I6rvyYjoPLiQDpzkSZQ2Yu6CYWfGPK21dK070WMKW3a61ketLFwF
kkdK5oClUTjHooz82l2usTmkqsswPrLQS8Uy6zadIBXMLU4778cJcTjxMJLZ2Dnjo30Yl1LyFk5W
PttBH88nIpTpTTFJfD3IWxyTfW+kogFAkDRy0129HOkdXtFTEUhjqAs1zi8r8NNtY0bCOodLIN8/
4LqEWPBy7GIBYTBA++zzLmVDxFLKSTaGlsAKfDfsvI0/G8Kumd2k6/OkXLREbh9ir4q+CL0CLrGk
xdYq+GXaPy5T+6idq5sIlgeUcWu2Ihkt1oGHYuHhllr5MC/QVS5K6u9HiSEYXTKO46Kp2HYKYa64
o02R4nFzNKPHBdqxA2zM5+JnxYHjliVyR2Cz1rwZIO5NWghLx1MIShA8pyD8AR0ZMjCuBhX2x+OT
U6mJMEcJUXNOr+6TANd0N2vV+7IsowXISA43BCjRnE/bccH7ZVw2+1JDA26WUZWYqzNApgu+GTvC
24t5Davic5ddy29Mxi1D1kr0qIXzYKOkV+X52D5OwJHtxIH6p9CCjRuUpMuFQH2dxQYMHdOdIyjH
2D06fQMIuQiFr3FIehHMrfn4uLN739h/io8Va8k9r9jPCdYNKb/x9H2/W5+9SqgYWuHsCpkFkeU1
2LHDHAdeQ8RzwBm6cMBFrv0yPk3F2XLsGNQiV20F2G/G2atIbPzdRVEYN7PIaWZvUKUdJTus1Pi+
Fzse5+y7FdUlCWRAlYvCp/VyofSCrCol9L3nEePK4PhYpLAjBLIG6Rka0RTXcOrWQf2tSmpks105
Kbj5yn9arjvbB6N2t5zV8i+3fkdvv6EsZIMaFZtssA1rDaIXp4E1ga5ZIiVTiV/Jy9AuRGTryPLF
6XTkB23USfnay3Pe/miJGFzV+n9gBmY69A0web+b6TrReqwSzYO4+D6A4osGOlzKkrMN7z3XW59O
flDG+LbIXaGBr58EzWccHaOO/4ggk9uBZ3uWc3+NpgmRDhKyik3nk5iCp3EXOJQC24IMywLuDYGL
P3wC2pxQizddXtW0UbL+NUEWxoOfxrbVbkAIFJHpxy8uuX4i4LGgLGZT5/2SyT20vud98gLn/nVu
BbyZ1VBnBtXRQnts8mBeqztoamSN0F4Z9E1/z4hWMSmqCG6gVf8KtQT3RlDZAhN0ft0hxD8bauVO
/YT2dBAIcz/9nAhX0mOQWsjyJzmLq3Dss8B5EazXNzGuiplemEnlZ95vo6YJjtIHG4im3lay/qG2
isU1Js9psMvoexte4hbqA6NGfQ2u7qZAK758UkMztL1O0+RjhZz9lK38DWInYT++Z9grER1b+3t6
D3jqoyE5OChb4q4oIgPw+wFwxJFS6QzWrUr6OfqAYknQZSwqOV4yKRk6F2QhPhS8Znjvot6NgTwG
PzHtfn8P4R9cOTg+PbfAA1zgMw5Uxevr0u5/iBPCN8h056PKGOnPXFoQbJVLUeKTprFjS4tT2Zw4
wTlEB/sKox/nXrA3LuMkiQrGDuKuhlclgwu7IcV7FdDut60KcXSduhmzQbhMeyADMGQSPSbUZosp
T0BF8cxYTPnTm9vVQaBRZIMbBhZyddi7R19SfoFengXRCZ+kSSP8ec5F1cyLA9hPLzqa7zy/43gc
+n7Au1CFzd908Vp/EtrBOugw4oL+tSIIcoXskMUeikdWgjigY8d6khxSMsHte50FmUeGunG7cBhN
hvjIXBZ7/zr1CHjSyvteq82Hqyi3/cU0SQ0JkRnxU+aI4HvmkuBNo9rdYs5T0kVR3j/UeO3qgJHO
dUiE1Zz9ZXDE7QG/8IPuwz1dvEMc2C1We2ckNHHQJOvEk2pztMJrT3TkReKA2wKZJfZl7ZDpf8aK
j1MFSn7GoJJjeWWWj2FpZqZ+wjAI1wg/EucnF6Iu5jAbnWDsNN2i0kBXGAuSraUdxx+jogF0nkgk
oh4wQB6JLqwUdPydtz/q+WAj56+ZFtIXZZ3ubLWpSc7mWvD+9dFZ5q+YQ6JQdmAbb5Gft16EBowX
uumsi+znn8cTdnxDGuobTrq1IGDlUKdjkQJgDxc3Jyz3d/sxYvGV2Gdn7VOzggfma5Lmoa710pX3
bWrb/zvpr6diT+qSYmkDBoy5cvesA9JQEgdFOPbzzhq4cZwfKJvDXUeYSMniMU1PwKC5lMT4cArP
zjqchb9h/05hjzxXaw0s0xdoxxwgwnHGgRmHsfWpPnPP2SGxN9Ghyc/CUyDHOShkQTpMBO9qyj88
RVL7ZFBE79qb5jbgAbwW7LtLZ75GuLP8IDWGR29Uwtzt2RCpQB7XIlE4KT0kLPzB0GE7apIstnIw
/qLEaGxg31zjJ3Oqvn+1iboSmG4HKfsW3GdlYHe+hf8ubSHwGmKy/Dz3Bpcsogsb52CHEn4oRTlj
SbawF6mZbenr1YvaV6W19U31SU26GhPehnbc/8/L7nIcSdLV6LNVqUnFTMIgZha1sZ9+lMo6tSyw
uWGMtGjzi7rxKLtfD8FKKRlXgyJ61qa6q/r87/kY0sAj3+qY0DI1C3EsYdm5Cuv96ML7rw0ZSL4o
HhvlIvnyF7s3m9+QFX0AkNMzoUIxrfYYfJw+rJ3MuQHQWzVt7Ns4JPrhmiW6alqOjlqGZXOLK937
Qa+m6PXkkwTED5Q/0FEpIohvyQ2YmoMK++HvUagTsgUVrV6ArWC7S4UK7kNmUNvLM4PbhfFnsBxq
EfmPSHxjtUZ7bQ4g6HU4oQDEiQTMT0QQqtx3rG2IV5d+4VoUXCggsgAAZnZRgsMmjs2CdA9gy9Ft
vtUprMChnuaCJ1EaW8ECvOF25aXi2mRHFqpO+UtGcic2PwqWPbG2fSmJMfpRbfDLrvP8jzrtQk6w
9Hy0mLeGQPTqMmjU7+bjJWtcyD4qQfLvulibBvjlRSmEPmY8sxF+L/8ioZAMQQZ9qGK5LwxACT20
W4/4xLhbSpJKo6u/1C8+gbpUWjYfjre1VSlnENMgHGdAfA0uO9BLtYIaBNa72mNe5TwqYMjr7g3G
IXQYLCZO3/NBSpB/SdW74QQ/ERJopsQMh5W5ERivGtXR4aF3Gl0C7xjXCMjzBTPKeSm0+76Coe7y
P5k9MgvsRmWelo1IA2MllKveUE9L5dA0DZW4nyOdbhJDvvbaAak4j7+RwdqDBB/Te39lmRFm14sE
+7UEhDBq4MxksA9PLtYSJkrzmN4Xy4ba/2yhY+MnRYKSvLzeGmRSI++/cAZGvifr6R/gIst88LHP
r66eC25l1COubn/4auj2Qtv7E4ds3i4oW0Cj9jCEhlWZJ3lLZlz1ziOHozLrS3OriQ6+w4kOMPr2
Nd6Gnb8yS7lG7hOnYEdRMspLQ6PdoB9/i4fjJi96oPd+yhg34p2JjxOyu4jHbyV/4k4rJF3BOVLm
ilV7fm3SpkHaJ9Mj6JQJXHXY1KAe79dTj2BWkmF45pgRJFPxSSENuA3t3BSNFgh9KVrPemzd7gFi
Jh5Hi3PyfGGMN6Rbu1vm7u1gTLDV6DdDs4o3UYxruI0XjGhW820EVG9H2uCpTFYrAIpa6IgI+9IV
aGYx4bR1BRDMXF+6gvXnRdMlPspRUz/HhcgMGR1Uk847Yky6OWB9AOTjqL9ZoXJAOjc52fbCO2+Q
UK4r8HMhIGg5T8+EEsimpfozsODoUb5pyVQQpCxIZ8C44ve7qXV+3izJ4+5cpZUMoy2wFJWCS0Ub
DAyWhLIioifUYBMcz+og0I/rL1541/Gzpib25+3rfLHXF/qG5x9fc1fpbJESJn0FbzDXnCes1dqn
Z6NG7MNVgW6G9tkBqu7MheHLm7PtZI2opQHIuDLMBwkxjqdPxvdH5AcRtHxW7x74l7FacDAbUA0C
nogbzgk0NFaWa01Eapi9xF7jCYC8lHv+mPJ5FF4UYwdtEghcIUHltRrJ8eVMTZkz4DQKdyWPdFNM
DJ4oMDY0GAsYxKOmO0nvcXrUi7SJuHWXY82Ljlfi1U+ULNzlvf08jmrTggAyRKDD0T3HXJ3FCYhr
KJmNWbbdYBtcEdTULN/15c2UCNpF4STxPTdJbtywbL9NTb7mhOWcCffevV1Yu5wMoO6hpxQugVAh
UaRvOwMCgLxYeVpN/etE35+v69xV4jJL/uxs5Ym15siS3wH7GEbNr6S+a85d3tkXvwsCeN7ZhlPF
EKGufDhuzZZRQvUN5us9IeamCJ3VHkXIt6/wXH4c1lIchh72gvk79I8Lj/fpZz2zncRk71IBI9Mu
2I2iRminhIFpJWUHduog88yWYfaylqal7PF4FBiD9g8Jfkj5a6axl5qYT57owmoOqgzpi9Dosuy/
Zaa0oqGB9gY+ynFH/sMOm7eRODexKfuTuhh9gXz5IlX0dWpA4N+ninUNTw3cANnpQqvsIMtkIhRz
Lz+BQnAK3M3vfv2NZ/tRbbHb4nfzTtQ46wiIqyQK4qDc1wFXXdpo6uWjIVjCENhqGMuM2WwrGITK
XUj/JoHVaxuo/xeq8X2pffxM5Uh7njQemENj1iYocTQb7eYL3KmZYHPcJi0ox3VTffTqgQfdAGke
tf7/WhDG34rlSWPV5DSRjm0vhYyMBlFsPdX2FBuHx9JgiGwlGd+L7agWK0F1b3b9dMujt4L+xKwz
ONtvGhpklpop1UEqICXjlmQeV8Ee8eQGJbqBeaLW0dZyBfGrFWqSNzsaO8h9lnno/DHGWIiEQ3Oc
JsX4W+bAVACbjggbJXKzjvlpxPkFMUDYnnyreuqx2a2q0NWUo2G++8vISrm5c8DUZYZFbwXlVHej
SaGT0P5o6JSmvNu/2vMa6BUSdzRrqvsE1p5zuHqO5XOSy2dC0fKBchGxBEjMMAAn7uMp/K6dmpKC
WLwPVc77s9dKZpk9WaMWBCLzOuaMGCvE/Wnhq/8D5UKkRRaVLENA8skLekABDs6l7ZVl3aLNqeXi
I1/1OWhoZ9b6gJAuUwD7/K/z2bu49vMtP99jcKfP1sQy3feNer2EuPfaUCQfal21JCOlUDwMEKkO
htjjf2hq32JdiKRLiuCsWfgeb4zVXTWmUjLCIUOnk5SVUrse1EwuOj+ZZkSyn58tb8Ce17Qm3r/X
TwVVD3a63mAganyCrUPmFJAQNgRf6XZby0hx9KxGanidh9tsHlyb8KGki/9lKRJcGWR6w71SAiT2
8LdjzteBf2RhnUiAsHR+UDGKiBzvMwGL+W6/oL5YIsJW4H8H2E/CeGSRp7I4AO1Bn2/7NKUeS3Qq
WaJCryCqNkv3hmbe+VVmqjqmsElrHdaQ757sdnlRyl7rL+ZKIJnu3Ekn1kYDQEw4lmhSxN9u7HpG
gf4Tkw9CLisomRu/iDOk1+s0NwOVIjME/Brhkpg+1biIbR2h0NLEeXp4EhaiSnDdyeuEH2Mf+fzY
Y9vgcVrLNQF7FN+8Xu4HnYDnBn6XfMH7t/zXz6IP2MwdbfzJP8AZ0Fq6Et/XUuFz11WWfhqfUdcU
Iy9vTyeKP275B7skLJygKdKIFmIRV+rhCtJ6LGhMIBbKNtw5dOjLsFRbxeZzWKV6S/JQKem89Vfk
tRpVcEjRuuVT7mfK/GI75rRyNWBiYIbVk00eVtiigUPhjO7FSKuduwA63DW/ZOhiGOLDYXpRxtZW
Wcd6G4nzj+iAg7YnPvmi+x6BGx9HSHiVMU0q94AXIJ3hlMY1TyQ1Gd1uBNAfIRwmh322DFReAtdp
ST2CwjBRhZnk/iGcQvkVERtuZh+LQE9SgGcGCAB2lp3raxHZ+aX+41fqtx0K+DgpvEcpA2lhTOLw
ogW0VO/Z3xQq/dig5joB/MDJjZFOF8i20FMw5chLLexBuiZiAy+hprU92jymeSRukjAMzPcApYx8
jcTvnW9/0jXnkO4oLdldNuqBZfbpttl5d7b1RgAquJbV6uje63j0cPc2LtiYG9HilqcFaVkMogfu
uBy2lMXsAMLL+VvIR8uyp6z6DdJYVQAtjxZlpoDGbDjY4YiWkkQD/AbGlMTX9fKLyXsI9GQJUCat
95gcSqqM4LUzwDGC9DjG3GaAreSW+654dbwo8PO6nG8xOXNK98yukqGD7pCK+KJT5HXz6BkpcTRB
xN8Nz66LGU8Ss+h/xR21mEJwuzRXcN4Z44umXTuohe/5YdPdPLsebcl1W72osab/MjFx0yg7zO/Q
tvM+zy3FTzg9FWMhnlPTzhblwk15ADesVOiW5eCxxJvVXG0bRcMjDOgWUNgvlVLV05D4n/Iid4Vq
nJ4A8dCGGrp2H9RDo2DRifXkIV6BnjOnzpVrtG4tOrhBILu79vm2ZlRjmTttslI8G7Udn4rZtnZF
s/eGwagmLmOfuQS+g9o3GCGUmbXmnhZteHyGlbLSrsytmqCJBsEtYKtMDMbDU66d6eo1q6HCdubJ
oo3j83FwusJw0ZF3Lv5I/9GGb/DeQIMBMrTX1t1cpp52udL/II2hxu0FC6maEbXtcWkrl/1RHnrJ
1JHj+mH5h8tINtqsxW/pDtg5AfPv6J/6HHPi1ti0Nt2uU7t/R19iLYWQ6r490uJZrFLosO/b201G
J6KaTgEyUHfHoY7R7ljoXg+kP+N721DMjRW9egvVY1NdEFixJ8PRO8lW+9FPAvmB0SpcQ1/S6xRX
8UdwQKPrBOZ1qb1z7CnMBoJKtwZ9YcN9opjGG1dCIxL2A/wwmKicL1oAjH9hJaV1O13+LZOprUlQ
7i4f9iK5g6QvdLmhyA9iGZkRCeLJHLU8w8WpvfuOBK2phl1pcdEohVknWFpyMfIpJIY44VszLaFp
EH9oEd3vnZpjhiksM1uJMhKz6QHO9MtFd9gTOoYp6ZS1bxbHNp7uoCbV8Mud6NKwuKOWiVT7VCv8
mCeOUIxTP6raZ7DV28kY2dVQJzAfsWbqBOdAthXCitlLQvhqkmRJQrWNEyLagOAhCuQM+jqde2/o
6lSltHVdIqNzOcd2liABeqA3hjHj9wTNx+/13UpBz5JBtIG6ppYW4LGlCDEg7oAlDTaLUH0NJara
qjoUp6tFJwY5nOshnfSPyEEmFpYRw9dDaqK6WqEpWUJUyfBM1djDlR1K6YJLio/BQsaM5FgxF1C/
MGZE/7t85g29pMvdgg/gDPmNKs7qbF2A7E73X+o43CGwJESDm9jKXpL+gt7X39NLt/NVmaB+h6mk
uJCwG9FhOj4r3Z8OjyZqUF6W5RZfvNdFxndCMoSLNKhc1dFp7djRe89UorchgKpi8rCYAf/vuDMD
+bLaHBRISuLau1aIhl3dB2hEK8TuIqEyx9J/YEZ4top7P9kJDHgYZL3MEduiTG5r+DWSM+bpgiwg
0srtqHJvKSqrv0+xrDmnbBiTUSFUfOojZh4Hb0I7H+VnRkT7h92kw96KH1GptRSsLrTzK+lV6gkg
uqF6Cr1oERcCOmqm7UVqQ49Mb3FQD4vDhza/xkpq7uBiSLEBWwlmwlpjIlwA3T7nDNYAY+R62fCp
8OBswKx3FkB3jAAX/kuohM/fZTGOkfzzAOyHWK5u41MlHFV0Y6pGPaYtgq/iGF/7c2E69IWSQFEC
o5czrjdNfQJIKiBc8tpJbcIZvsZTndU/E6dvfyUxpScArybw1sXvKu3DX/rLK1FwdS5mI6aD4efC
AglGpPYQ71dAjJ9nHfT4YWADRjCfRXihJjd+uaGv4d4aluq05HSnDUtOCEyuot7spIL04TonEnEC
HOJuXp9kD5oGAmHEMldt8xWkTWkHKzuvBCcoi/Gpzpi62+kBoohBGGJpj2u6s/gaiQCVlVjJYOsT
D7Xt2IrIMVwez+j7PwucOQeXvHayKYAfEfpjZyuQH23NNtlZi4hIzjBLyMTnonpQbab89I9TFkd6
txblYg6TbhtogjZLUXYMbeOxTBYotdKTRKdggNM1S+k4lly1fDV89ZLxfI6UZ6LwVli3clHmItlY
g/8goEDUimrC+G0Jd7Esf3TUjmX/7fWET90KTiS2fWdN6hJGYHoxhGhYQG+5GutzuVe6C53KUEap
GLhNKiJKxeY2F+2qGZxqZVqqw204l34FIsCFySjLNOGwg6WX3McIzyeWW2aCy4QKNXLB7cCKa1My
PqQqkSloLY/2rajRcvwlYdYa14q3yYRUAIdY+LAAUo4gr39O+pmlqYfbIqntaJf9HnByZvw2lszW
ICouXJ/x8NWvsXCBJN33P4/E4xaAC3mwbFE7QbZ7CozA3BV50DPcegpDy+am6oPSm0vQ9yx/dNFr
mcYheT1GXnLLL6cn25BLlpnjMhgzChd0/OUx6K4KA+8N+H5AwtdwbWa2r+zwoN6E95W5OKeHtYcT
zGKkqeh5J7LPgiHyhdfDmCuULkMXeOphRQqjBdB+YsQKOf/xUKWCawL65melD761YErfOS2nDR+P
CzgDkbxsm18fxAZLXzTgvCS4tQtnYa1AJPTkeiNVYZsf9+zXE7cWWZIrIK0AK2St4bGojcuFjSb/
YGHUZfxtY/ZOcvyUYhKKkhWiFEsXRxzaI9zx7eGHwqyO+QqLIYxqxhhbRk5ex30IYAK31xwBwKqn
JKpt+APEKe64P1iW1/y6gthAQYXirTH0QTU87hRRM9F3h2FclTkZRO8X0+m65uC8K/XrHQPtPOmt
H8FWTCF0hgVEvbAnh7nKBk5hNht1rkiKwEAfbIofxdi1uGXACv7EEatffqYmzrggBtHa3qnpo5Ux
kO1RgP2H6COdRXBruNB8hWlNlHfdl+c+ap+kyK9twJL6SYUxZpnk7r0q6ETRDTbPMtkIt71t1oce
eQNsvkgS3BV7WG4LKb2L1bKrdzAUDMbPRqOnKpOtce4OQDhPKobwQP2yYT8Ey0QupDcDnbtS92Hj
7/kKYa7zjQmrgJOvkaVCDVAahELEcplEKELZOXrg3qqATuZ17pRIUAlXb0fFii4mSfWlu+nmAU0f
eL94U/ZeaSKt7E3oxHSA0FOtTxK9zBbXe4H/E7nAgR2QPhijKxbiJF8LSLo9WkvoWbbY9LOsl47L
cn4UOo+iVdfFm9KKv2j07rsNNCK/zWBNkpew017+KIFevl8IH/7Qz4v62iPCcif5o4mzbsgkrHa+
iKPmuSAie/cD7u7XjY9Snq2OtFJ5QlgEdIRpBeoZx6noWQ5BsgCXC8TE1F2GJGazKrI5gMwqdUPP
jq8RyDkF3MDFUp1vl96PlQy/lyZ9jcxR3hsC6nFmFG0C98aOOuV8abWql4BDUJ/PnDWRy1cF3iyu
6GD6MHic04dVigZBz+Tli46K0YWL5ArDjr6EY7a5+oHQJlxzidGA47ILs8ld00OFNFAAcp28R7/x
fYAJNdS/eJOqFq3ugu0eNekrxz/fLap6Z4xrvD7Z++mPWk5hWYK6LM9f6VOgzi3VDr4yYGLNkGbI
N+GdhZROgyOOtux4E3dEujAJKlnvcKRWyxsyjuZuBUiWoip+9IbJMlx7dqDP6EU7reQSiFHAVzBs
GHoWmhvrdp4b6uv299ANyb8wrz1+FWtjXb5l0TAue9rYGaHZ50rM7bGIP34uWXDUV/2LP1sgMGUh
24VAMkC33W/sSVYEAaanfi2NMpBvVfgnKziljjukqdNUDIedgzuOq2mluNKE02dErzFtCc52/LR3
jMRu3eZ4opzSd+rvrsYrwNoZM0thThkE8i7+1GdMALiQ1el28DIn8yEFSjWB+cFwnD+5vpwj64ba
TNkbdffNMU5zyRVTee439ZFKqJdxD/hmE+9Knu0yhyoFI/ux0RYUm/vNzcppzSr+AGssWQ1qyD4E
8b1mBy8HvjF00uvg4HE238Rh2QcwSrqt/X9ZfkCs50ozYs/HbzqHrtw6RtqHB7CbGP1XuOGYwRo5
1Rqloj5VEwin0I1wDlZYt6DrTPbxY+a0WcBdLkWaIwq5+DvTG5YplCbKBUoZ0VPzywhX6kIGAEXt
kT4weXFGSI9VKzylBwyEPuniEM2KulCMy2zbQF6YaVHeLMAvV2/nPxrsIXi9vPGxN5UDa826lol1
QzUxnve5LXdeoTEZQoT5tqG0CU7GGF+Ba29QZfMfaJ4cZYxUqttBzQLhk2SKUgahudR20Ol1qvMM
6TXpJcqeRI4KWMneKf8YbpsPYl7eotTwuydlsXnR1oL1xYYbFm0A26fkN/BW0lBLkl92nIWblgbt
9B6f9Zn4GVLdoGMfP+k85sVKqelMWIU8PvrEPuSjQ8YLD3sVnFQp/2NGmZvUqmTArnwDc+VTlf80
OEQS7YqlZYpCzXA6j4WvAKlxsOj09IKu28Zfn4YCbMQFiczrB247prgeKoWtgfHp3S9YGBKkHQo7
X5MjClrfZvzt+dUhwkLAt6chvtmCphEkAk/WoLMFrqpaxrcJyxvlCidrE8Ijl42avAE996S81Lqo
JPuq4TkMp5QgEhJKTZr0QaAwJISvueV+T5a34ST9y1Dwr/sfrs3bx3oI5fnnDr8hSr58Yq538WE2
JXN5e+HeGq6lDKTYlzmPLNhMMCKLV+fdlLBysyGgKQ24O6/1JniSzn3HeX4pckgFDhy5FXBG1sH3
6gX5z+Di+Td1IVjb1sRg3y9p08kx29L9laA1X8FFI3COLwicjqtqU54zdt3nSJQhCxcn9XbcShSu
PGQ0ij4eNI8onsXkLgBOkFYJWMHp8OGRhV3vUzDrwlHDIGZOxggecp/c2wvtUg8YyEVzUEg20mmi
Yjn9ko0fx03wauNsn1y+V2+dljwTrv16+ILuOM4oPtgZI/x/vnyZ+CUaeaPBXlZ8HEQ/cmFMceu1
A6ebFVOirLNnvHZ5kp8A5V00TwxnYsgLfA4P+FuDMslmGbTtvskWtn+BvVleaw6f9hLa6BRtqXMP
DohYK3Te9DJ8IeXdnX5wIrTwb2P8CYIdB81dPIaMkgIoIrMEp1YIdEBWo/Z2HF26Ql3/4gBjgyxQ
8qkl1qw5Gr///zW9253WiIldPU3lGy/cTE2fb2jn+ZYda+F6PuuJwn2Pue2jqgBigeR/5zVJmJkf
sHmn1I9c8V/Rq8VShwubSiefO1UPerKMeUxDLp4iaUAopP8ZJs9rLz6O4KEVpLffIIZQW0nfT26h
GP/eR7zY4nwiy56X7njxGdsvLqOJChqLdcRSQL7WTcXnilO9YzAVN04bGkRgCYcUAbBnrPaqc0w+
MuQZKd0Ix8VWFmDuioOPmzNi38HaiJToTvsQAspS5BJiWGHGkD8iDQlYEwPj7DgMNw3S+F1wYzKh
bUadN50HaMpT2Ogpn9oPf7w+ejlVA5gSBvNM88gbhmdFEMYNtQtffntd62949OcCnpq+aJTsmyvU
3B5tsz2+V6QDO4T9nePoOgIUpZU3tgzfWdV5iXu5pBLBUpr22WV0Yw/GNRjvk8bffjiWOCJYuVqz
E6hOXYFfHF5eDo6sa5rPNHQ9zdDrPWwA9SJ23KbaA7YaId2H7wkuHbWQnVjhU0Mpn47HSi7ns4qK
fyUJ5B+Xd8nR4lT37xsvhStVpZD2aM/orSLMCpa65TC06eO62hqIAHOcZZjmiIOnTpasQoIUSmIu
tbpZmj2hqCrHQVOyKrZKrzm7FQCu/pGZUhyFLpKegu5G9XpWGJRRF7E2ezJj7lLT0h/64imQT/pQ
Y4HdHSDRrWry1ifj7iiMy4FEGDH6eDl9ujO2ujFZC7EFboNT3EjDO2tQKaKdI0P0HwO+v9OocIxY
AZU54UYJzDQyhONH7AToOdEbEIAuhONHZcBLDS8KmybCyroPo3L0Hamop03qgUEt5FVdBxbovxdQ
ZFgJ7x2PdVOoagQnAAN2qYrTmGDRRBlfCWQKVoAGv9XVs+nnInA/g5FGoQUFXfyJjh2ea3lUBfcx
XHCN3fc985dOq3yBjJyIm72lxTU0V6z/VzMGCKRt8uiV+eGctM55xfUe8Qc5+kbouIcUDGuu9+cA
hv2oJCdw6ae2Ya9ds2kn5bBpfASfuIfpUuHHS9arbEvecZBlOc1HrpnWVsSWsA66ju/1AXnGlmLt
bIn4fVla1AVGrtfsHuouXCzPJHgkwEYpJOlVFKfZSpkX+jD2fm/g+4NK07qtDrndqYdfZVJIDC77
R9vjYupNWhofuSpDp0Lu68/CL4zBSK6KQ09Oy9QxBfVEfwSHkXdKd0phnb9RTwPK5TaDZUjhetDb
jXow6LMlGgnh2Xm/EDtLDvpBcOxUm61iHCkU4EgkL31I/8Jdukg0OM2jWT+RuI6klMYTGKME7gI/
TFxZhaenQalJX6iyMlc06zzWwEcPZYC6Lub4elFBChkUdUDmnhXlS2JUWfJG5IF/SXnzlGuYXYjj
vP0oiaMFt5wD1qO+Qo4TVjN3BfUNaT1+yXu0VCsbHq+2BCkBIBGYdM56hQ1wAHh1an3uXoxCCV+I
5K0m80tpbmarq/sZ/ZQSAnSd2up4LlT4mg/giS+RzW9S1z2NTKfb+gC9w+bca99QDBk+C6qNZbY7
z3xbdtkPN9Jvv3LAY0vworDXXU0A2srTrFyZRu7ZUIU+4DEsOST+uOyvsqx+4iP/+FqwVpknkzJD
6rK4z2s+kJdS0UoAEdWQjSS8UMKt4HCuHcCqLl225py1i+QCYSRNOtWpZwt05HTWsBjZOvxTb2KR
n15bpE2LCyE0wRC6ad2XNtmoZINLM39edXQFgMUP6Vq554KS8zqlEcVV3aIZ39GOTj6yll9INyzn
lrpCPXd9p/dRZuP0flTJO8zMZW0NJ1okncMk9EH8JU7WJJ0m7wUuxjKGkKKNMwqvCS+zoT0jOR5p
jfwFUc/NYKtjNGXPzK5RJwFz4jlAZ/R8BNJOVvKEhTdCalef14+318Gwwrm6nVYa17VWUpiCyzxG
e30IojuaoFUKNgFZOdt7WAVYfT9cGSZ0DoPDbyVzFbgFA19VO+wGV2BiXLVaiQxWkI1uEPosl4GI
EIb4CIfetrDZq1kwkB2ex9IxbuYm1nTIBSPRChxBon0AnsSlyz1ukhvhYEN7RfHZtHyhB+N7Xhrx
O/exbtfENFZetbehls/JPZT+6LQFDHIJxS7IK1yK0mQoUIMvCfKfwERwQENrnH+YlcuiaMHKxO2v
zs7sijuvXQq1HPQi7cy3iSNqqOIrGg17mfNMM9x2iclAzyvuzocswEsGGY6kJWlwj4+TICMwTe/E
E3D386TG/nHXEznrfWvGZMPUhy8rHFk9IvlktYYIqOkjMcXkQyPZ0ojHFKp8oZET9/OF/mQnkhhT
ZSWwnsb10z5Z279CayPjh73GGRuFoDSm0Nln5Mg/F0OuqXcEQDr6iZYarzC8v4ZlHm5jqd3ZTTfn
h0Qs5IqD1hQTQ3G3OaPszJJYy8lYb4+mfmllN2vV3ci+N+rIBTTA8RZsmjjSbsSwtxJWMwPQl+vW
XcsF6CFVUxUldVx9H25f009e1DWRDbpVM9nYqUfJDQLmOtAn7IEOaeEm/rePJ4d7+p89xyYseiHS
AE8TTFgOcF//ma2veR3r2tQMR5LwwlQUgUbYtU+yvdz3X0iT+51eHfS8+EFoYQwFnd6R6S831+Z0
ylBwf1kj9OqtghtraP2MEQXK6MaAmt1XIhZSFqnlGCaroMeocWwK1/dRhx+6tBDX0pSuvvdPJGtC
hHtKAPku3B4vm8Sr+8nNl71h9g1Fz53DEmYLXmSnRunYtZSKrm3q7V5O0R0jgiEfrWdai4fG6p0u
bVFEjmGIhWvXOsHb1T9nyP4XMA3pxz6+J4pVQok87Fp5MWsaWwWmUy70PSmfpLUuAkcZMhe4hZMR
25jV8OWNEKFhYUdgRl+mU+unq+Ip6UZ8P2X0erX298JQy2qFr+AR9IVVoFNGHzByHAbv1Pz8PeOd
LDJuvcSfN0tZIl3NBajlT2ykginBWK7b9Z+ZplRrkuBKDFq1E7m5NWwqLxqAw2PrHAChfBKBJeV3
2g8fbHocot3sf9fiPFl3vocYXp28aHutPAgFzrhyQqdBImcdmJwDB7x/mL8rwqD1zgZxsNzCI0iD
8IM8kX/4MkqsVDGeGf3VOmng2OI8NoDmji4nE1YjCsJsjFcuinQmuVAAQGgiKhQLMJpp3cTvt44n
dnPsQzsW27LvSzzq7Vg0DMcw7RSFBf/tZkFdC2NaKsQcgcv6OBDlZId4JWGf7xsDQXy+gfv8d255
gKkOzFqXv9joCjOrLpqODN+4kCYH5zYxToFTTKj0JpTKz5uLFl4JkTKWxD2EppME+cg4TmJm5XxO
CshiuBmC1KjC4U5YuPpWhnn6aCbFYUdaWw1cBVePGbsa0Zfmpy90BLNf/6sznkaZSiP5oxBuez1e
0JBLeIVH8cqv9yZH7GAwN5s44wRVhZlGFVBpPn/Wj10sYz3XyczkWH4wJmwc/6nP2D+GGhRfIlzo
Lm/9Lzalgd9EVq8p6WSRZqb/MI7hLAgEzeYRuP4J8+ivT6Ggw7tR5BWcFjNbxLVr+VaMwwJtg6HV
snGbmUWdEycRmSHs1E0bLJABSKxcKWqgjhgFoiQpwKM0eEKA12Q5OcUYenEUQOC0Ggvjwti0AK92
NPp/QcfqF+tKVxYjA/ffca9O4UlON2BqmdxHA4kKPQ1A854mlh+E01vB8TodmeM47RZVC/s7cwf/
bSbzmw0QeRXJ1092fve5Tta/hdlte1MQdSUte6elSUD1GDzAtZ5UkP8wfW7OhfVrYXA/p4OhvEDt
PU0RwTidI5+e58ueE76zl2Utgd8d9Ga4gVxca2JkBjHQxbPVHWWsMW1aA3vGSC/+I+KZU8Goc0fv
d0WU5Y3BuE4rD+qwLXP4BPWC5wxConQcIY44vWWaPSLOzdnvXuEesdVw6EpU7jQ87ehjMCiBSjPF
dT0LqnmGo+57pEgPyqNFAAhw/R3aeVJ5ByldogyMcxeZkFQzlgFG285rCbq8z3hrhgHyrtaKPX83
tRAmbIOtLZ3Tm1q/05j/IqgWmA3NzpY+WoUIIgDv96/OyInANs/i5btMqNMrG6pqpm46xx/ekocy
NwEa7R/TsanZlaQPQvqOvob+y5HbqIULizxJWMmG2swbm3ZGz85RsGqOzhf/HXiAsX3hUFgmoIK4
sQPxdTTm6s7QAoRpmGggo0bfl0xs2sCeqAYByBpAz8v+CnjpJi98SlR2oIPiqXRXC2ZVgIQym+Pe
RP534PQgOWRz7XWADYvc3e0EadV+vKAS2eFRys6sM1k8kNM2k1GJISulZhEzed+OUPPq/s9r9GvN
IzHVETe+hSD0fE2vzsyjtQxkr6fQmU4r7DVt+l2qygDIHv6rAmNYVD30+CDrZf93cTEaSBy77Ntf
c92jGKlW2/jE8jYEm1/1y3vtJh7tYxGn0ri8CkN8CyrUNR5caQWQbf7qam7ua62AgiLqM30TB6Mq
aDTiYhseTKxN+GAmQ4gUSzUKD1jqbpCS0w877oh8rLupiGHeaOtsLIAX0GOdiWzLX4DSz70iZ2XZ
OsL8JCghiSt8pOVk/BFLURo2Qhr7NGgus6q8vMrCx+PE+WOFAHnQb3Q6am3MtKFfYcZjBzFROTnQ
KJBbjDgQfGeGLUcUlX2deFesDJT/ZOuY4in4J4zHaj5fKR0rLCuPETpsdZldgeNtILOouxvm619R
iZXPt1+x094VicAnTG66TqmucWnbdoADeQMGt4Jo75eJhBb6zHoPvTflqwK0OAAsBfMe5AkuxOAz
JHiMNCAlm7Ebr7Xcgh8yl18UIwebJVJtTKXbdTOsocI9szHmtBKWdmChBY/oK8XeTx5bNOmYqPFq
rT/Go6jM8/Qv45HZLxN0IZp/lUOJvpb5LxcUfcsyzUaVU80R6UmDXG7m7EkTHqS7TxC3VCceYhaN
cJVocuXbn8XOJrlq2B3BhBBvU9glDWv5c6YRVyI3NWDkh3jIH38f5g1TB0pkwyhGFpDjF3iuHo59
pLzSzU8x7RR8swuAxCrwlMOKT4hyql1I3up715cQCLMSqH+OWd7suUYlmToYrgH/whVs5sMPSPrF
NzDwEb7GIivtJbq47BSLOz4m410pG4rZRaXv2GzfATm8Z9Vd78kDCiZzvJhiJZcREBSZ3XTlJAh0
aPDxhUBpc4BtSrXPqb+z6MajKetMPiuUP24ne4/ir/UQg2WRRC7EM3assMB7qjG6NstoSHv92Inp
Xt506Wqg9Yrs6bzNs38xo1/MNuRbZhgDmNYZqG7hILj3tMA+oLpFF+mBIBKcs2pRv9ad/GuRQZt4
qIh925pRSjVbJMmoCkxODb81PUNklZyJtM7Tk17unb+GkE57XxRHkpwYfklKs3lxpTbHLCGCDKlc
DeZqWEyCzfr+pfv8l/Y+UL2IJ0WFgJxYXW4wG4I4kc+OK4SH2EO8xyW7mkCQAA1r7cGPYFQd8slW
42QZGesKgFWjTQjBBLePqMr5ayw3JMi6T0xes4sW7olO/3yOvtRRicDznUxUHk400mn0GRgGKITX
GlKM0krAum16kNMiK4jrczRjqVSmE6foBdH4rqn9ORyz07O6PAQu1syz78ZMfH8TnRzHpJF+zQzt
AfMeRGkqA5LH/0w9UcLIPwi3A1R3x14XTr05wZRkNlgT1jt9/03948JnGhpnSAK4sgXmmTHZOINg
x02z9gV8WIUa1IzRMTC20oUuqwv3JZPVYyysMwWcJVGce1OgN9zqAFM5pwRKMVJcvCvbJgsLeTIB
jVxJyrcnw1FX9wtxM3H/cG/uOAy0QdOttfc/Q2YcrmypGJHY3T++5khJjB4ikmU2dKtpSD1xBxPm
J6FRtQxrKMapjjjcPOo1E3aRqptX9UXjSCi3e0HGclpe7JzA7/cxC2QyRXAtD3MBZYyQPq8rDPl1
uDtUwmPAB+QXoeyj6wr71ZDPd9uUGyKskG9YKCyKVgDL0udEXwN0Fy2S8Y0LESgL/Xn6otS/FXUU
im5F9V40hTAoA41pGUnjkzuJBMvEEufDzM84DO9pPKhmXSs4ikohL3cqOqsZwna9WD7gYe8N282J
63MhGmW8GjDAcregvihp9EI95Gz+pim+2kkenDh6w5Pc6Zr/O7RiBYGBCgytnNiVL/VY2GXQwtpJ
M7XVQNnlM5orZLaUJ6TkcK7KNRFvkWv3YaD33yVqWP3tcjR+J7sa9i/lgj85Nb++3EgO6HpcA/Xc
ABFyt0p1Tv1wUXXAuQ5iGUGkTbMAYUuQNwPto/1pKhjK9zlALXo8ufMyatVTNnYbs2gSylEglUw3
UYJyvugTFPTsHwZRv0H4Q8vv3aEY08XbDM0C1YZYun0XLBoNNu5Ua12bVvSXTI/7wcOHX+codlm/
xk2fqTYaDVmamA6VDzP4KUBblKu+k4MSyINSsWPZmfzZ6ehhxgNkZcsadG9UySnlfj0MGoMpn7MP
rQ3I+GtzHEY/+LgZ/DvfPcMpQrVZHXHfOTyyiiQqdKKkutAMHqgsT8obfnyTNcElamYKxwU78tEF
cKaw7S0kxqE+ct2lVn51aChLnr9qIs6DPgGalKYDAKquvb3riW3dh4hPyw1MvhJ46qu7Ph0WAt1Z
ToAnsmu6UqHCDEQtEUmylHI9/TyBQw5OVeDYSINEWIMLQ3bQDYJABUKD5yalD3O4CibBL5RxwFWj
d+URA96qYQMWS9jypIDX/Hbg+5gqoc5bhMFRIsFcpvqq4SqIuexApFaPxFJvD3sLQRTZV/Kll+3h
xiGlZQKX9sTsrhcZFT7yYKADZeOYea6FJ8XDtoxbthsBG9E4SJ18GWigxKq1vgzXnYATjf6kvqkT
+pvX6bWYHF1yvmn74R9iWzOAA1gXKwJPpZaK7L/iV9+HBcsMCmVec7huNc1tgtk5nA2osps8bIqt
TrosLnRO0CzaPeslj3Yur3k9Fh1eDFYxJzy/0Segm49fEZ55sqXcMP3gleyemE0LrLikGcrJdpUp
IOJ0INd/iNr9Bo+sX6pPZ/DvfL5pQ4oTHLmGiZkPuqSgz2J6TQvzJZRr83ZJNhAyFm1tTJZEUK+V
LZQuqr7+JHkDNyhi5BPIJeDScmZ8a8isIfhJyj5aKyrgMo+VXDS1M26rH9PVVOa8BvnqdGOwAFbU
E5XKXZgmbbWZLQ8uJStChkw8gS+KPHOtbd/+JP5JX4r459JvP29fjI2Vk427jfERi+uGthvbwIfc
6wQCdFy1gUO8P8h7dZ3H3qKbhDtAi764bv9ZBvpf7YUk/Y/elPg9jxswBa4dc/h4Yeb4YWX5YajW
Qn5sgtk/MmV08Oo9DgFwFHXOWtx6egxMSjwayKXag2JvaV6ljDRH3ox0ZUv2B6P/TUzK9ptAZJGw
7Nsi2Kwp7gTegR2iO7DF6MMKphrsLF6eRr4fia47Pw7Tsn85y44//vkxFM0i9ImejWeGUgIYhPOs
1wT2aVRZrBDuZd63k15IqyDnrA+5r3g8Zu9KXKmYwSpuTQ3/YM/++CLkoZQPXI9geTREeXzb06tB
HwdNko83X8aruM3MkEZYeIl/9lw4hRGlgUuQDzvkwxr+2Rwj5sf1KeFCXrJBBIOmHW5DdnBTFB8w
FCH5dJadxsFh08CVZiKbqGE9vcH4jXbrkEHwdZk1vcnxHpvE4dDpPj+Y4fJ7gur7WLQcvLec0ql0
wF30Z5rKeAEZV1Mlta5OClzvFy3DcsumdaD/xk6gmdonvKCkhBKwUgR1ACw1QMSH4uCsqbN3akSB
/zefy03cMGIg6MZJs6r4M70juwZJtYu8JYdXxDEOvN0VlWvNHXEKBbdsHx1jIw16AaEOaRcKwiJ+
08AoCaVTcFvlYqLCMsD2Whvh7YHfSTAhzcTAmC6F8D0j69mB6smBR/5qgwV/xEc7ESCf+7KgOaDx
HVlYCQ5mUPy8mTzDmRetHrR3AQa8Aip1sePEPwvTsUkqv92G3fljZuSo97KySfLd1tf4YvB+5my8
ft9zuq6W/H8HA5pcAz48LLwdvqmMC03hIljsuZGHvLW57QpSpi/YaY5VZMcGe6BJSi0rdv4qJ6DE
df6EtygoJIPfQLeLHhxfuNFunjpBRfehXNP7Uu8ey7NPjtPgx/INSbzyVFmPlzDuHMkPUIVhglZ9
znjn7V4YVG8vi9iPT2NKBeJY2hyewzW9dmazn3DipM6AntQU0liPCAQz+pKBgk/5c+TO7T5apodM
OJUhg78QX+u1QxEYPDsTqI2cJgvPq9oLDFbnCRUwFoDJpWiC8zZS3HvwOTkpof42nowfl7cNJ+Dv
8DONExOA6I+fHcJnm5b56QMIJsT6O0/1E+253YgEKmL88k20EzAdfQPa+tvs/4zFvVa/UPXkZejw
WEJ2Q1uSBW3HlKp++aJ9hQGm4fymCj0MB7Tpq2EgB5cDKXp+TD7p7B71Bp6Jmutp/s/ZodBDSyVs
cP/RzgamJ1uBMcAH7bVtnlXh6vEBq/ajJJycZFEuSFHaZnAK42HGZpV9qcI2fVEViV2g/p6se9+B
dS1ej7/91bcTQ/4Hg4v+Fgog73tLMnNDrGbj/TdMrdkffVcTt8Oj/x6KlPw0CSMiXtN3+eCyVwJl
HtWYhWiicxVmRn8/3mAITvo2gmO0akyUZEPQY4gnuu+WZf+SRoYvAdTyusvdPFozx8PwLXNiBa0R
zeY8G6orQ5qTFokZ9BNcn7QLqyBjbQk09TmO/f62GecfxR70AkqHemmReuBmU2tONm9bkeBuvecl
dxirCUmwuBfZA9Fd23dFoRQrGnaQZST4syu4B7Of9wAJ8U68bkKkSF3SGUze7Ney7L4AG0CeO/s/
2xFd6RqxmTuewQsTlB/jigBQKq51P83Stu81R/WjOhwmG9UxZiAA2ExdvRU+A70TmKKMT5YgpxT+
yjRZDqGDHMcNkZ0S1XqxRyfL5dAmpyK8IFjRa7s+Dedot0AKSreLgNc4Vc157cWyIXRaHnjNDR0q
T0DKh9SYOngAQe9Igdu1GyHYEWjGAg/OKkUlbtYu92bAO/MIEqHTCTutKiBl/0AMcEFhxw4=
`protect end_protected
