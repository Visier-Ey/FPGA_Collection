-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
bf76v1OPUXy6AMEaXf6fjOf/hUHapaRJ/mX70q2TgbVqIkaocFJ0n/uC8rBZWKXD
ngxts6zvfV5wzTK/h4BLyc6i4oDr/zVz4W3Zj+RHSznhQH3aB5MhptdGQDfG8WQd
mTbUtcHTwlYKMqkl7uGfTBWT2oEBBZChlmjwZ5YuIbY=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 34688)

`protect DATA_BLOCK
4+6u+QQf2gD3JPW+wDY2hn0IVuFiK4fdNP9vRxwdUas0NP15mJGKewRUZSy5VvHe
Mxk0/OpRGFT3yDOIa/yzAo0lqsHMUSKEZvagrCMFZdGSVPrJvAikzYc+VQ5sE8pC
/g9/3diZX5eZjhyEuFx48Q9/vWu9vTHx4yzXlNTJwUJoaA4qBHDfjBmzJmB/AT9W
/YDehL0j759yg6LBhAdfqo60Hs9A43TonrFNSjA7Q1OVmLjwui+91Ydo34vwfejz
cGfB46K03tIYvXp0xLu0QGM24p/JpyO24JFUKr8/pWTsfJMPcwUsKZcMCi/GaCf7
BESX31v1jNvzvKvEQV59es2Srrr46dYqCNzitdaUI3v5farc0obGZpWsi5CTOC/D
5BmPnyFIqJkr+TzFlnDSRgVH2Bf8BUJG+ektGuggrgNXZzKVAcniKpPHR22vSckG
S1Np/KE1Q/FyQklGX0gGV+ueakU03HO3xJVuS2r1MxqGmxHM4HP9VqaEUNkzso5P
oFhYkqFogEKMEnCxh/tdAPD9djqbTVV7DiMrC9lxhXapjbSH+xn2UEtx47JW6GBm
tMjHLoad6NF1lC7PCC+U//HH3VRa2wUW4B8SG7k6gyXewYVKjy8hwFwnid1QOUFo
pGywMGKUvF0DZbl4qyJ3tumAIF5Pxq7aNYJa1TDbUb1qf68aLzyoCMjuZncosTUD
/YOusYJpzWbjzxbmAvD+oxfYofX5AeJnebp54l6gKtW/cDlJx0PxEZIUQGODuZtK
dhakwXlfiPE6JrzWaTKQpB7ekbOi905V/Co4pWDpS/gkE+PD5GYST/yVadLZ/GCY
dRKoU2O81QlG7wos8XG2SVhkoPhSy2IcfGd7BV+hcrgeJaoj7RBOw1pyzU74WkXe
BNLv7NV9cubtNykokfx0N64BNm5pohsWM5hn+lOJbGTAZZlpMsevMkW3UjaGf/eY
tmQWZbM5abbC21wv6f3626p2xbyFV5RNx2dqQEYDwGh+7+OE381UhmVioCTS05OI
HhM4Pr5A15z2/oVL+PgKjx/70bgkI1nUOFiU2pXmvMRUlFLpmZGElpwtcsGTVbde
v+ovifs4oCoa6mV+BniiqWcronUc4/3ESqIopkW6hJNtudSSvW9k8uz225WVkhdY
eoYYs7KfyHALiWNz2zc2lrxETWNFN6UZDgkr6o6Bn3+G6keslSHcn9Av72fGAJKP
MoF7CMRNFmN0+qTlfbB/zXLGWf6uQJZ49waiO9ciA7HbGTDC7HoQvwUVP7qZDbX5
UO15tu0ohCUJdtUeMQqloLqFmNBV7P32OrNLu0p7zZnikNxLt6H/NpK/Rk3s83UH
ffc6N706fTPrA4afYgNYmrV1sKYMmzY1s6howr2EZEWfP46uURmt3T0vsx+nFKC2
4fWVXUruREDdsY96yzzzQL1yL8O/ZE3YcC2xGV20oN8SUCGs1b3zcq5DA7C41kz3
JEI+6B/HGOP5wd9Cmc+cYY2LclXgCBOmkD945/fOR9c1O38+xBHx2e6Ye07ogwcG
DeLqQrEbzAZXGOGUEjqNvk12qbIfPXe+nRPhLuyZsczgWjUpFasD4VpLi1ETlFXW
xwAMeduikgUBqWI/m2QqWVXaUqfVjc7mUSLLe0po5Rzo7OdwpZvF0hxrvM+wmCdi
FC+dfOZ+3vVqjSrAJpSyRg4SCfJuhMyfIU8siclqBvmF2VsUzqYDwZnw3ReHGKrg
P3OPVBqqGsPxZCVKwoQ8ULVKvanFGp3pqTyvSV8VxwE7AIvOc1w4PoKgTrmDPqyR
FCM9OV1WE+5G8FXDJCHMw9ksjeZmY7WJe3Ms8Fo/BTWSCgZh6b+d+YWODCbHjIrE
8rIA8n9NQ5Ih9a4si7opcsFx3F2GtupwinNsKiCYmhgODZhy4tys10r5zvdUvdli
Nrq+rn7U4IpiTrdDZv4ujWfD/A6uqUHico3lVyPvpmcQl/x9wlxhCxdmnRY7wxHV
ShJAJFE8h+pfIL0GIAKFBfIwUpQ7pgd8HuWWfSzo/QYcxjz6bwkhRFveE6XxAcuB
fjT1FgFqqTXjfRByXRJjYRx2gcjQp6+l/U7UCCZiZtSXD3Rf5lRXP6sZdIyTp85z
+YtIQTPBpOJcKejCtRGA8nx40Z4cs1OkgJZG+WbGwDTsz+BhJjbTkkrGN493YlpM
cuHbV6n8JZ+/Ftb3Tpa4mwOTw0dNYoRUWOES2oN+sLkBcb8E87LHklr/xz54AAlU
PwUOO/95yBTuFLsEx8M3MsKjyYmJhb0c8WFAvDpcv8J0o7Q61744RaVHufMycw1S
KY7+OAM0uHFWc16nlywh/8JfRSkI5AikTUm0l3rJeM+mbNy17GmcxcNoE8uXoJmw
hs32BbsBepIsEFW5o6+BMqiOFaMqd86flvD0OLKBBd6MyfdP5zXlJa3EJwGoC9Yu
cak8V5qcm0mszJp+9j0qAVK0+NzsYWb419Z/3umFdN/uTNtbVI69VMxeR4eIZGJ1
qJlG5fySsg0sAf6p7fUuzIT1xdGMkxMHiw0kmiSnuPgbKm3lDYHSy2bUVHgXP0Jp
TGeRZ4+Z7Uaj7LRWw8kd79Cn9AUNioBEWNMgSAtgIJSQNovVfO60xq+Vr6mw8oZr
s6xLSRGgg+6rhpHri+OqlLW/v6kJCF/ZcYlyn55/OAVx24qtzFxFArayITJQ30B6
OUr2KtfZIpZF6Jg/ElJSc4CilofLu/gPxrE1jgtMWRbTLShn91mvTFJ1THBka2it
VMQ1tC7506CBJ9Mr9dkMTaG8xWP5805aoHplCQaEKtceaWoE6fo6ZG4+4Dbu2xHU
gkHux3JqlfwrmIxpayZ9Gpkj2x5bx12+2GebuBFflZIo7FFML/hg9jCgfr2AbcHh
6R8EytlqeUft/ccmcxmc5h+O6FeirTcYanoG6uCO0ZfqyQMF5cPl/pSDlK1rEtiw
ojG5eabb40FRw1ilc8niWSzlrvSB7VgGjNQTwouSPCAC0cM07tNo6UNmFrkZLeCe
dO+ROXJogE25gbKMzJbzwfoI9owmts42uCrrGHwq4mIuoyXdNSlegUxKieIno1UL
MeZKrmxYE2sUKkcwLNYaBvg8boIVMFtVPTyD25d/hKxcLzrA/xuF/htsNyE3PnD5
cq/8EW4oA7twY9KoODXNcZ5i9WMNrFnnI0BnADLs/OQta4/a7wCgn2JTRuI0zVDK
MKdtlhZa/Taz+qN1qLapikD0/JSFxYmWJUzOmG0urO85r6vkVVLgqb/IOE7vLrig
gXpTRAhfynHEixwwlsUVdojTbHcNQYiggwFkYExTzYYTe3HzSTVmmhcTTk0E7RnH
jzaMfEjo7WkJQ7eyq375Pk7ZBGG6b8XiJlJHCiiNuPk529R4FQP7Nm19CEtI83qA
PqChzGOCc35TsyKnRvvDVmCQ7kHRCdKY1hrHHqn3uJXuqaqAX8//z2w4o36YsISq
++6pjWN4IFFP9mRh4K42nG/ZoetMYeVgvYBII4Mwwf6n7J44IYVA92Zt1yu1i6ju
4fEiPKqCzzbzIoo9XXm9cu4X4n+2YCOrqa18knL36ZEOwOEwjfdTqKKhBvFyWYgh
j5wc2QhZ9ZRwFjEXGeA2xWsBnld9eIxFRBCDdavhT7dtvGoCK6wGpU5vhv2qsliF
uF271bWqtETu+aIytW6+wIJgrQjai9BGL4kDUgjzKmWeBJvkAvDwT2MRHk0WP2WA
udCG1pILGt4Bkf9WIOoru/g4/IJfWipMae7F7d5xVyjqquJp6M0YJW0uceov8unT
Y11Bd2wUMAVlA3MOlIAsxuS74+HL3Mny/QMHezpQU4DIOkLIKkOgHKzSYFHUeXYO
j/jyMD0Azat3gpD+T3b2FX0I2Xy7k4n+aQTVUQhaRdxt1T8zF59v6BUMXQiB45fK
9pngY/QDKG2e/zJVD7nR9D0tCp0gGI2q+xzlu640gFUOtnrvyUsfZ7COOYfb4Zzi
u+ElE2Y69LJZsV3LHtO2J/+vwS6X5awfNIUb20Du7LhGZnjMpH74gLqa6zcbHrxk
Ymy95KdnQPMK9uD/zCYF5w7q8o8CebdPudM2SHKAuXa1UsmloFHtnfD/Y/ka5F8e
lC/R3tGoj7ELDVkI4JGUkYYjkBm+ZM+6LL9ovXFZbIMM/AiNcD9Lz/FWbfDgnjUZ
PV8MBJfEcJlrB/kEEO/Sr/KuRZsi1Sw4kTwNP+b5f5LlY2grpyCKHRnqESieEO7L
/1KVKVKDxrL4SQVOIXEr6beuX4J9k7s0zCTsd+e5FIOp1veoj9FOU6ygRCgeH5RQ
jwn6sJ7OPDokS1KHFkXK25w2iClJfv8RAdjruuVoriCBclQZeTZlkGyMZkMz6HMf
HIhlK82cdqYCqbP3x8xKlTmyx0hNdVY32M6zQImrrM+/HhzkXyLCpA0nQJU6YAGv
7MgDeeNXRXfEuW4OkF0us0HJv+TlkAAg45YBJ4MIv9Cb0soD9w0Q+Oa8VV47ww72
fSsHz7qZoGyye/bsf1LXnQNtONIFDdapG7Qqj/WG8OWApH2VG2AtxpY2wkr/4j6L
Zy6l1IrEwCH3s++/DnzSH8QZ/ML/Pa37XB5Q0TpkptuCYf70/j9vEkFjWXfZxb0q
WhbqXN7KWVUfMVKJCaBoM9Qa/bHlrs8NwRH3KfMwa5ICKUKbD2+i/1RC/hYiqVfS
olSrTEO34px8TgCQMt1TxQiRVuN/TGcfJHDRJqKM0GBeqL8FbFMpTVTZJVJZjvV5
gNF0F9ksTre+5jWP1H0pKJqUNEXakdv7PoY+ALd9N/RWrPH1G6zDWbYGtYZLq7Vi
UWkw2MACRAS69rox3vB3WVbAS+zH4c4yH9gdiUFix+IK5VAbsYN2VobfwoYh2Awe
rF0OLUaexK6IsMFDmvB0jTDx42Byx1E5KUE8azjLhRCRt0QvvgJcMv+JWREEiagg
hPI4y9Mj7Dhx4KF/oNKemjI1wVE0PYoLcVW9FG/m0J0dDz+zhYt8MO1vjqvQ6m8X
o3jlZhPxNAMVEfHKPbTLpP3Cv0zYqRs0VKTxz9M5+nth8uN9Zlr6gPLxCoDm7KiB
sxshlj4gRV8r4ANp16pu5xMDYY2TGpdJ5ogMvTsDEwcSH6ZjSJ45p/qwlf2nDSzT
F89NfmJobU/LBJmemJDG2eIc9eHq6ejEI50kRWoeQUNofTMNrUL+0S/03V3+B2gw
hVq7SQyl5GeE/Bykg2tOp8YQmRUpJhlpbq0OqNM786Tmv5C/aUeC3njRiSRV28z7
+QDJaqVJ3Zq8I4XCwiH1TWYzM7NlxhJsIn93SglBrbUu5PboqozaBZKHksZaK8lP
zNVyp4THZ20hqpEodeDnXBAhPBFJn7RFr+BKP4agrBl/zXPO98B2ma8DOyR7aMBu
Qfqfset2iKb0sos42pjwmSygJ+ttKtVF+XgG/8C2cz+a/qNaJlBvkcMTKpNiG4cf
iGXQv15eQA2vjy2188mk74fKkPmjMWJrQykE6OQA9tge7EF9677pNZQ1i+pRPcCO
SFQ5b+wSmzS0BJhPJlO8MnbJkYcrKy2qA32hKGszABDDdT5swYbY6m6iTLqkcriP
efslbPMmJ8iBxC+mq30IFMUv7EaDF/ll8F5YeM3++PLh9DqStlT+A+T4ESNsrvzX
CmwZ8nit6eWAp4S23G25eXbx51cWjK+KYc9e7sgp7OSJXilKTd1yisTHSP8vguPw
+UcMIJbfMLxI9dVEh2A2z04PA0Duha/OnVtLkZWUIJfXFeLaN06JsXg6TjhCPvKC
zhzau9ptx4p+pxO3YV2RfSdD3rWWsTRsixSc4C2VK2DSFjB6Te6o7kZ/FpQEfLQj
V37InNjkxAhE+8Fs4c3awnubIXbwHjDJXDMLXqGRDJhIE0tfAHrvdVX529jwxp7u
G5eUXzmStWdPNaIHURAn8DDetIf8CXPTat1llYoQWOvHmbBD+KK5iHIdIuKwPeIB
Q1AGDEN9h1HTB2CLGFw7XhqhLhRIA/JzdimfCCUXeJwWilmthsG278jHHc82O+wx
D49qwYrxv3wVcpdn/Z3AMPoCqRegI/jpdPmzCa1W0mNVOecFP3L2L4l0s7QTxIcz
DuqUinPoClE2gOyQ36p4ysqErQcUEEJd22bO442Y01POtrBI9mrcJnPdM+VoIIvT
+KCrEO6T7YjdBvjhmTIi0dP2WE186mKBAM9vgEn012R6Go9rOoGhhmx9B+DYTWnA
x4sk9wz+uwI2BuUHzQNn0UG/3e/ZrkyyVXNi+++x3M1As0piHuGJgLKWiIklm//V
igPpFrj5x6Cq0srcfC9dBiqeQLHphgGu31x7dpd2q6USLF+MOiPzYPRa4bU8s8g8
jLstxxsUT5KgEJyZqRdyO0cLtCDSkdy/XH3l027JQG5k1UiEtqQLtwi+KaklglWb
9qIdq7UIsQreHx9032acB9QiXKGjFCqcSbDEf7YFpZFsnWcOhEkN90rRQJKlrvxZ
nMrlAUT+GATbISpBiDFq2LjxBwkRXenj96ixTOIdqZXI6cek3SRAG17+9MLlWqIq
1CwcSOU5pASXSpoxmhCjfQS/HNe6Ye1zHpR7IEYTmcsX6D5dyQXa6J6ZaZ63kBYz
xvDW1kyPNAxU1uArTXOX9E6DLYj3K+51eZgBkB26DNshZZsHeuzE9Hd2i3SVwog+
nEhYgQ8zqObmtGRhAD60O6APxPUkeZjN2+drM6IxRQYMVSJuBL33DGPZCA4ujtUB
ZqbIU2JZqoGV9TlTzY5DsTi9jlhUWFZ22NDPrSQFrGv4D+zUTDKRzRaxUHcPM8Un
vqAksJT97Xj3E7UUpkWUX4Mg91sl+OP7ZZj6fpkgaDCzISU0rULLZP08PJ/MF2LN
A6L3JOszJbG3hgDNKjToJ2dYfQbHCiu871QIxM3s78Ob65C2arT6sy1zU4nO3IIq
7XRCk3MM+3wFrJvTBecGqwIrvUp8Z6sGx9+KG2ROENlaScCdyqHEIurZawFiP4ix
TSamZhnht1XKJ8Xs8W9y4b6PjzgxzDGMNSzJFdYRPKXjs9mxud1Rj7Ar6iMJk/1M
3hgaY41GHKF6OvK8qeZteDYPpHPGXq/gvFDktOcaszrc9Lkkp402mYDmIjpCoN54
lmrVXMI/W/nHFhO3TInVoWZw3e2UU3o+pqCbZleDkbyHzIW2v35r7xCtiD5b7691
uoXRmbZeIBD9AAKm7Qm6aEJZroCehzKKYUaM5JhSiu/0wFFGJHv0FjUuVRwb3LTb
RXphsAxC0qU11fSIUczPkGyLOOYZlux6Sg/mwcMURbkrXjgMFhPh0/ytykrOY5W6
ISyqoNNKhdbi9avjVjU4H/6U8q3sLJA0XWoJ6g01x6VG6zlq531UBgp5njsH/sTs
JvlyatLSoqg7Ot0R45VboukYKtaz4RF0lEpH0Fy+vyCgiYMt31aYDsXc8upEAQpR
eMgetyf9p3IhCH/uF+UWJXnLTwwcyZX6OnrbONjKZ1Gs8+t3YgLRvzZnt7SU/avp
ggMSAnRwbDCPVJzeOoTAC8r80bkzIVAks0ynGwRtgTTRPl2Xak/txqKTLzsWGia0
RM3GhtNDpbiDMl1uDJpCSBLpJZiNKB/L8/kVXo6BoSbuEBm3CL4CFcAYmOtyl7le
O41PAM+ZQCOlNWmqHl/DWDApOSAc/GlmBdcOeScn6fhVbRb4sle0/KrbmbzqEA4k
ZwTpRIcOdaahKHACTcZa7TxOhRZIZXfTG4mUKZOKdRVF4ID4DZWQQ2v12OO6P9+8
RlEemGeveHI3K5EP3yzOOgYayxy81kG9rdRKpHXkv8/ds2UaQs3FQMIzy/6XRy4L
lLdhHd+BniIlcedeOba7mDUs9uwzlT/kJZxS6nF6WeTC/M/Cs7xytj319YgJqiVj
gDQym3ZH/IlmvqB8WYvxOdqiXnqZRZsMMiCuxCJqUJFc45xDhFG/+V6A9Q+9CCSm
sh65b19RfUEAdP8LOmGbRDQCUbpPNTBU0MXaz4lKj6TT6LRvr5yMwbpQMHaMUqpG
lyYWPrLJYyp2l1tHzL6NaeZCAhgJX8ip1E2oqqUZHjdjkwG2m/zFBVWKL73PzymH
SNeB//Vb+7lXkYSuNiU4eaAmkNOES73ukhB77ZslYomXpPb5fMbt0qpYhg1YJQ29
6BZ7s1zVPv1QvLnyiBKGE50co6nFu6Nt6iGhBa9rX/zYBlxphz3iUa0ykxdsA7aI
do8wUH5+dvb52br3IFE/3EB7l2IJltMsdKKuWL19yjmwn4XbppO6mWGPvLl42Qj0
4+mcTckbnPz3YVwh0wVnkQpxuMAl3EvHayuX7DHA6X6LdMG12il/5ORi4JV+6/vI
HJToQrLlBXR3Id6Vhs3d2fHwq5189KkxbdyOhdAZu0eEqPHysfWAhUN5FHgFPoak
7CMc28I8v7U3pPD/QIGdmUsZMG+gmGvgNHNJVaTtY5bwrjR21qr5QI9a95LRMcbM
V/qAx5MkYwUOPu2WTdU5hZGYV1aRlT3MeLxh68H+h4yQccAVs9SMNSchS4qeN5v5
izYOhaJqFNXj5abC3V0tYNWvqgalcS77wCvBPAVw8QhUD764lQsesSrcTTPD6nlS
kZL5U2msEBJ4qcs8TGiEzRKXJhmcx4Uv6sKi00CgUWBTcATyymK4JP/EYK4pJbjY
D8WZLG72DZtgbU+MXmGIbUPuyyUIuAudl4fIEiOBfmU6/ENS048zluSKTfMqFcLX
TT9p0bEhl2ew1LC4HVsKuF/Rv/WO0kog6bu+pt8H+zjU84aAwV5pv+cIHQkmbYfq
Vzs/gbXcB50kWPdXdjukvdm50K+yUTnNFCP2sj0jMGG4Ed0kGSVQVxlG5c//kiQz
LU1UqEP8BxUiUki+fSpKNL7lJv0dJ5LicW5z074ZoKYk5dHl2IfT1uKlw+56S/QX
kyi6xhb/GjM649hOptAodjAul/NVBjN4DxbSe4z2dnvvcGngvn+f87+X+W/1FDT7
r03hVhUrPUG6g8l3tzjLYLHJNQNk+icJn4eQvwH+oH0pAzpGhqHYxtkFb1XHJrWI
5DnP18LT+PvVct4nWxz5DFCbEfc7c3o1uBMjpVqiH2u/FI2QoDAMV7msg8UvTX2t
7qobzmKq1WzfOnj2VFHhv2Jp3g9pVAq97Kx34WYejEzF7ON2Ipgft5PoL/6bCcWy
XlOYcsY7mybyUihrEaGT7lAKtdbgvD+J8fgjxKF2gQebrpWToYN3tOjAYJG4Y+77
FmcmmT2rJjX+jCqUhRZU40HrX3X7fSN1ofpyJR+fDnH70i61mZ4DrMNA33SQPk67
s952ZWisXEqHNgcm3yFJUQigIpOTJfCtP/lnnvUdRK5gdCNCpU48FQv3rGYS85uk
JISaxf4FlDAvNIzsrWe8eZqFPmYv+sN3xzNBtallvqX3yGA38qjjtWXBdwnDo/HJ
uZQeaN8KfoW80f8SLa/vnxfIQiV48pQr+887tzhCcwngAAbVb9QQGVEZvp3FQhPj
PvVFNoQBJTsvCGWm/CX2tIWvX7uTed+Jc4CQRzxDP8l3Yoe2xKQAY3eRRlv6/nE2
fIVtP8j0rkQ5fl1NbupvwnauE8sSVCJXDO8O/ABwb0yfPniWTIEpdyofY1Qqm2Mx
h06ifSGldMO18Xbi3mmNcAKzeHA4A69srcwfGzgW7fnYQYf2PYtHuKK3JYi4xcat
BVr+giSD8BC02ddUebq0JQ0QVUQ6wxDhI+Wc9H9AWi9ISIqf3Se++lFZl81Hwgbl
mzRn7VhcAuMnZ3yDosGQ06AyRRRmLUEzuPd8rpTDIjjB0WTgoUMepGTr5PunymNC
arNmtJjhvhIa5dGI2IqqvWutKIVFMJKbSMPvhk1/KO4bj9xUTs6Mtx3j4K3pF1mK
xmtR0opq7HiTdOHNOOMZpI/tECIR1zYdw2lsZmPHqsslVW7zNCiuIP0So8RHBF6i
KjXnkZInOwrM7l3KkypuGpt8yTH662rDct1Yg4Tz/NWqjC58DHPzI0CKoNCg6+U+
Mo0DK2pnwEjiep2GHuwDmahAG57ByPSk1gFkfuAlg7WPgT6rFpWHl7SNG7KEX1Dh
/EtG3YJnLATrLHzI1sWVWwDaV2hCUSMrh0jSG9dS05Pp5jnFuOED/K9RDwLRS18+
Ss8pXVA5Pc5nOKKAeUiUkfT7zW8ULPcGda69qswPhqycnn54Zz7McKxBqi2fDbfF
R2JMjl1puB0PAzrDEOW1XAt5/ngIWYLhsVHtWMoq3/7pCWuVRO6qXTzpzK+5Ucf2
QRGgGdMVwvPpnSPo0iCvPYe94HD4kqUG+22sVmM9qLKsVNjeHjTr8Hu1rpaMUiKx
JDtvk5RHoIPFOALxG3wNSFnM1MoyDTg2t/jUURjwT8dR8XRRnoTWTDVBq0daDvcr
G1kEz5NqICaTKqj9WSKQJ98Vwb81FwLEWbjIlfCPAhDgzLWjnBmv8LQejKgxl4EF
lYdi4tdBUr0l+0LZ+ELgt+gw3hEgRdcPiIs707Alu9O4tJuhZmKDQYqJfxfe7wug
/iKV+o+0CeElGQpKP6ETWVj4jrSeI6MWAILcVhW0qm5Ol4NsI1XPPTp2CNO5Uo8W
zGXn0ALqT4uY59LNIKa1DKJwS4898jOAVyqZ/8sqJC7AevcqoIXtXe6rG2Q1OL/D
8mY8XmOhXgEUBxWbB4Q1cHmgsH7mAX178DDwktrjdDrnWgy/pPXkfTphXaJYpxwt
jbwxCotMdupNRLAXznc9A7BudnOntixAWSit1xj95Yv3RH3t/tNKB34aqPmAgcJJ
A0Oe4CTba5XbREmlc7ZbaS3JZLiqQbjDnBVQ1YB9CUMBVuKR5YabeGsuvTiejvGx
UvqeucltDcfJVMbP8zEsZILH5vwsiOSFIiBI9uVuiI+No7raNQ2r96D2iaWVszsf
LoHegxWv/zxweHYP0TOmBdnqhYB+mtAqcdJ/WdZ4wfmZnVzi/nVAmlqj7KZ0yfvU
A7zMXKbw7IUkLSBaB1O6a4e4MkveldwvHIR7vApFwOEdZEKAuaxMPTPPN/dUm0vE
L5JRFmxR0D6yGajEYDo+7y8KB/ga4iy2dYFFifWNuaOkvw8q2VU6FigxtIfn1WTE
Uc7L51p8Bmya0II5sz+EIcOU2W73dtlQD3VNrkz8yegArsvv3SpRkvpgLkSKulGm
gI11mVDddtME6W3HGpeTQS1BIElZIPv7E6thTGegv5b6ZLihoq+XiH05zoHJJ2B+
B0qAQb9x1K8yI35ZoCzYNF8w5sd9HfAyi5Iy/msqEDsPsh3lm2Jw8bhvXQ8f0e99
dySE4oOnLkulJSrRLqgqiJm571SrObkZjBIWzQ4naIXzidQPP/hoOsjS/UU5f5C0
m3t3nPkSJu7dpnvbUuUqxdjKopmfngCgvzWeI5fXmTO/RU52RmGcmhYeNgVkTIjc
3RAPvsYTtQLa56ZFeYyQUfzN6shBLHXiFjfgHJLUFlWjyETCttUrSR2I2NjdfRHl
cX5y87VTsCIepVVBlovR4leyAmpejJjvmP48i6ZoXasThs4+HIXxxf656/ymHChJ
mbdnxhHYvBeS6c38kCGGhd2IYPPHZYdXd/Szk467uClK9i2+EF+TJtGbb0Tw+eq0
lCUbp681/NigS6QudF+hjSP7ZPgxVAugOFpFtDYwZjqwpFKUOsO69uxcGKbWpotO
tsmHn3lu+RnO0/Ar5pJkJh38q9TSa07G47qTdaMaoJNmyf8Uydu9K3OausD1BH3d
WZwkvmU8t7TGXEMzAKKrQiB0fiVY34IUrlK6uhVF7RCh8jGcM0Dh004JA/6Y5Pgu
DN+92foVlL1aHCjxEvi5LbK8lkCDFmBIR1s3rVZkPeB1TXiF2BjAJIF84QVm+536
AJ72M5gfm3Yj4JNI9WFMjDUy/wW6cI6J67rCKlrpMZdR/QUIzRgRuLp4NXMvYF8g
8nj2LfOP5/HffyYrHvtQk73OY/znfl6RX7IPyEq6ApfT56b4qKY2Z7FpQwK3ttyh
Z88Q6GUZ5REkIMbtA5JcvSANTWQmd7hgVAPVLE/WxdiOyuvAQbwI/P/9wduuX7cV
E7Ef7b5Q0eMrxgfucdveH62myvKUIZqpKNKuEVlC/yX7J/gCsulOvYlkSRDVifN3
BNScGgaDiEuVifHNjctkC0D4q3qOJot3h5LTlFwG3v1Bwg/WgL/GuGeYuGxNzizN
OztRRIlsPfSujh2GMgvNiLNuy08gB8H4RY4zqwuuDyRhPTrdGSlVPbeV7gEXxHzU
9oTNTSr+aQJOAuiWmTE3PDm9QSoE0LFZGk9CoJtfONhaV35QTc4RLNqXHfmTuNl7
EEIE6njmLNsZjj/4h20RarerALqLmyaytgwVd6sfaPA+do/UbdE0WG4Qn7GAn4SQ
Exum3X2E3W/Zr//FWgB9L01UffJ/7YfSE4NET3/MKJOASxRRJnQN6cvwaSJiEXQS
wdw1ly4EsevWV7v4Mf0vcGAYsv+wQq9qQpAd2x5nzqMAb/tBVe5V2KFeqfpV98sM
NAHvCDnW6/Z6MQ08wNctiw1LXbCTvqXD8eylIaeNxT5hEXtamZU8TPTca5491mJe
P+Ujyj1N7kHhFM6ofpPb2/OgQFx4bXioeuiXh4WMR6rfL254M25hYDlKsl4x5aFI
FCO+/gDHMcaULRqZw7qNt/evyqIIC9+Ge9PXOjqIepneTC21Gd0nEghmh7ft/77i
6S0UH11YkIXst/qGIb+4iXB1QBP3yto8hlYHqJvZ7tqJ3EIcgJAmUUwcaS1EMFks
MD5IOPyr+drl1h/wXDypphv6Tv7wCJfYM3i7f0/Y3ABoT06PEn8t7X4MJHS50KOC
ghHecV/wEGfLSApqobdauDCdL9uDYbOoIJpjX7WPQqVWJQ4s5akgo34OtcsYu7P/
FXjoN6c3yzsZ9k2KnLyRjgLkv6CevkIJP2HSbkYqFdKuzKBJhtwSMyTkaUF2lu+o
8FVoXRyD76cNGKYdYDL1QKVgWu0+5WofLYe9xwpSag3D1M4tGAGp0HNqH++eC4Mz
9fcI5N5hixRdzeFbq6XIvv5sjpW8sCg65sPPUWsi6lLuZkynuvlw21AxiPhnXwZa
Pe2ne+Ja5NWOnegS9aBwDLuHzzIkrjrkypTAz0jLqABqGdffFgniuIY1ZdpJLdVD
XOQCGDq7jkDGWTZIvymxeoCR2XhEQ7Q9Llu1u4YVKeu/Km9SNsbbxYpA4ToxiZiL
7eZf94kj9Jmhk/Od2ALf01T/2CbLx20uFdeEd9Ed72Ta3ptXhid+LKMZB54eTyU/
6FxMIE2FMppgC+sD/zCU2jn3xp4aQqrtzeX44C1AovV3YjjBYB+0viVKED/4U+8p
92uIHjVB7Ucil5S8usirChx7D0zz0C8ZFIzQ63CA2qunQxlCYcurSZsVfmdV76wD
3zYimP2pBOO61a2FHIgYtV8owI6dJZ8mfmD0LedP0Ykbbql/7p+A0G34SHMnlJRk
UPQJwxnarLVFIRCwmkQe5ODv2haOAYfdqa3UGUWFoJdoJ/UBQiXA7B2h+QR+XLZJ
mt/9YKFxEtuuYgUn34q0wzsFdxLk0VXcKp+LeKzHt5pc9mzUnO85CqOhWmhqLCkc
Um4Hy1zsKxVqyAdZ5rlQ8QLr+vvyTdX+UBDcG3hipeCscspk7eFw6+4TT036AFGu
mTOkETN3Y6CeMIt8DJR/rX8stdG1yNgreyGHLOGz1pIlR+wyL/xkb4Jb21z6CEhs
iqYVV7eae0l0bxzZYAK+HagmFpYHHet5VWCiJ0J1Qwmd5U2WW3YOC/1FZs7yEZ86
cHdQ4thgzpHt93ksMCy4AxXJCysjpxUVwhQILP68Dqx01G41PllnRIYUZHWO+OW8
AVcBKaNL7InDxSUJuJb0C/RmFjR6Hql5K392x8CXTCwFjcEbEFTPUcslYLPNjLzW
UyXss25A/1lK7MFaNpiQgoXBygQAc4CzHQYxuUbOhWJFnbtwyqEU2EezgIfI5bRU
a+KUFIW9mrpPc1++qcSwXksYe+yEt3vc8/SAaRufEa9Fq4mrqz4HMIkPzMgEl0Yi
V3/Pe/pqeOEckUlWL5FzPumB2/C4c5yUse1kNowdnRvrlrds4ez6sHuNqG+Mi+CP
YnsVPSCSo1GdQ1u0t9RuCfzrNDNc2Va80zx9tc7sisz6AeCMmgBO9SK4Orr8SVN5
0+ciBEpNevIUk1gpbtnTnw7OxHDBAPHZKgLC7KzEqQoIHxqdnrteVIcUjpdCNSJS
3eTGRwPETS1WewUJ66jMPBFRrAdF304zlkBhFJ2inyqFLfWwP0Glz9Tr4ssvbYzZ
2IMBrUAB9fhEUjCaxF3Khsa3UWi/rmiqfoYiO0GlTDtX2+bzr2aEqQMGUCi9C03N
XPbVFL04kMNjEUmLmWOxXVAQzaZ/16Bi+OhJ6U2XcmxmaBG7PtEpIa++ElPz6TXR
dSkI3QGLesq1UoU+wMlgHCCctaHuJ9XdJ+Va6NdeJs23SaLpeNF7hBzT0NK2C1Q6
xZpRUt/IqCTEjI9So7g8kCs4VmWsehi5hhwISDV1nTLbdjaZ/0S5FqcjO7DXTl2E
XjyNAVREE8yh7TsgUqLMisE617HFfkhtZd1KxBaPbhkNxxg7UuW7y0Z+Uqs/f3Tc
LHSVNzP4vbcmVTkBHa8w8lQ698QIxwH/DTPHprMwVnPJSE2xqLTntILaPZ4arFs4
AqeuPrxYD6JTu1o04z6Ll0+lf4kPxfJ7gyE0cK5/UlElVW/c3wBp/KJWqEj2R78h
2g+9Lur6gp/4pE02gQd1/TDj3Y/Jv8jeCCpdapRpz8myVN2/uylCGErUnkBQSRn8
gYBqNfFv7/tJYT+DFwEPl+lPrqWH8Z0JeDcGAPDv/9CmM7YPe++MmwaZo6mV6qvL
ZBYRk7FaDZwdy5modJeQWAaIBThAcVZgOGL8AVsBA3afoburr3tyjPKD3YQ5FE/q
25e7U8I2ej+4m1NWVVL4Px8d0pd1vebvcYDlkz5KNRcAzsu7zhssclsnMyACzSra
oDoCrfuy9aCf5oI0Mlj40nLKGh4R1VGTEfLRXZY1kuHhqePs5VNHx5rJFsIwnCOw
LrMC40ekleXT3Ixev9t+sLnm8eZWoGe/lyRVPrCw57Q1edbMy7r+UB/P73fajDxr
e0u5QsZoE4/yq4M16YP5kJuq2o4IT+iVXOAwpEPbB2BmhX1hSDZuECF3MTaZhwjw
Xfx4A232OzYPBXagKSQOit4XAV0OHcIQ7shWLpVOr9a5FyeYi9Uo9rqVr6/7bjep
bAnwWxW972j1eLorOJPBdj3iF1gOKgZGwkv47IqJsI96Yfe3iDsH5ghyJNEt/hJ8
lOnQXquBzNyrybzdAgH7svFZTPdmr4rlGaj0nekexkuQtnIwiqnpnYaPDOIsBdzD
c6tGsFx8bJ8f+pxmPPYYgU7cTqxg/0AaNaM1T7beAcEbQt5BnwByFGiSlj5L++hp
PvSSq/tnlMt/6eTWuZTTiXnpaDPt4Q5IEZz6yGvsy/uMdoNx17GONIC1/rEZE6bX
RsElmSRVOw3llO/EwzpaCUsS7c0Vi885wREVR+GNR8lji6GQqMmlNq0M+kQ8iYJT
p/DXl7f0r6IJTx0exUtg/aJBtLLQE7O4xdIOGn3ppt3c3ZGlfQ75ngt5TjJf28la
/KapCchzDSsHhzKtU05a4JthDo+DIUexJAaH0r9Xe1epVf1pRbmSssrCIdmpfBRI
u6/tDAqdGfZrJf3FWQ+w4GGL1C9eeThSamxBP4mP9Mo6GvsvtoMozJdNVNz5BvYz
uu4LQwcOVaPZZQu2jec9iOyScVNpeTRqTzkAJBn1TzBpKE35lujNDsjPTMI9CkBM
F4wgUrBPNsz1yOXhXzNtdD7AFzfSMNzDsrBJ9gPYKQC7RYTkQ2xDCTFsZ7XW3Qux
FMYLtlCauh+5yFwE5TmkwlpypJmEYk4PMAiSi7Pe5XxOEJnWoEt9CIMh06XEtssT
0sbZg5gTb+GPqlXssQqGcE7aPHvlx3PsQ4Z6VTm+soqXKxGDsT8zjFTdC7xXPHGB
Zcgcz36bn6Wzp7Sk6d2HAM7eV4n29M6+T2riSfDAm0+rmkfHAMGWchoEwOQRnOUT
SpDrmUfJPXZnqHUKVX3vsq0fEG/eSOulx5xPHGqlaMlCwgRxZjRJYtGQPYTOvkPE
imxkPi2s80I+eS2GXN900FZH1iFG5jqj6lygdkRqOmH1ZWa3sRZ2p8rSf8Uck4l6
JawKvhA58aYRRs/p479o9Q5fQTyFqQjdECEDyunvrGwuIe/QbQxOp2K6+u9Q9k9i
xUhett+7NrBAnYZVGoZOG76ntzAcMCmZksi/gGtfFps37yu02S5NbR7frJ67Dlee
eIGJKDPRwdw82k7QQODKLzAR+DWF5bWRyp1zCQaHB0fIjrbg2nIi78Oyw9u9h/TA
K2ACu63dxQ2k6+PO/Lv4Beje+vaUfe3G2pmzu4kewvOtK4HJRpiuQu9zCt0TBcaY
N2Z4BnCVzdGiedZwfh6kfGcziFZgO2hp+s73artKNvNtDTRFlJOxpMDdQOjd4bm6
QzD35xFtLMbAPB9fh2ZhPwf3hPmzWoSSKC5Wu1rONwLkxKiizHYxpVJLmbYXTaVS
5yeNqUJnhh4XHRNH43d4LbG5/h+e8sbF78F+gEl04E4klknq9onAN0pjNpJIdH4N
51Y+SexnBDzC0T3I9LVMqUX3/pLLsNPp0xDsRb0TUq6kCRnVFDFJCSrGU6L66Cnz
YB3S9/ID9ObgUDLmAbq/w/dYLU4dejg9mcEkB1VW5GItOaQ7xRB/ZLsYw0jM90s7
LLsPrOcEO+PpijAzQH3X8qPgWOk0HtnwJ4gCi+khwdroUDhkN6u2ozaXB1Y2yKNg
EqkVdMQkSKokzGmdCKCIA757c5loFziJnsS7z+1Fxqj5NGvrR/47r1Ecbuk6IEL8
X+WBLRu1VBQyBQ5Ctb68I06XoNZcAii/Ob2jBkFBLTVI3d9iRNHURR7k810r4MoU
NqTf7lof4sSlmxVn/14EybN930+YumcyQuP0VmNJgNKeylBu3ZMVAkRPDac6vzYZ
JKQ+G5dddECD2F+yezwH/bTAS6ef9LW5Uz1s+Qebq+xplpsCVZ+KJ7jpNWLI0ly8
WLiuDJuqef78Mws1B7lu66yWXZ9mRQv03geZ+KQu6NfSrclzEPMhsGnhAZUgorRb
xkD9PnW6puRz3/UhsI+r9QYkGWURClOOssZGYbQS4mWgJ5FJCJARvDeZa8qNnBa2
jJTHOxj+UNKZ8gvrXQpG3YChdXv2pNceUISZqfmB9sbnqihwrN40XSt5Qi/i5BrM
/AW3GBqrNDtEgZYvD3VNCdkNcRulSHq1pH3gSyl0KniF0UbvmTKwYWriZq60phaY
xaQ0Mb1MyRupIz3RGuEo1LdIH/NP9MTiNSQHWWDZ5qkhpBotBuhh4H2oILQJO16S
5pXu8WhtiAR0MvC/xazPNidBFv8LYFEIIgkzlfaj3UdpGhZWdcYptaQqmNV7USMK
WqLxwZXJ02fn/BnvwektZXIprmIGjUx/Yv+lHj3vzuJpwxKaTihcpW8cb/d2VeDn
6xNXiOI9o0D8P45pd5+F3I6I9+dBZtyNixjaD6T4xEhNkwFCx9xJU4LyTV0M7jHQ
+hqw0WmTlIV7hzWaS4DJkSKHAmbSka/dNSeQBpWYnx9k/2XjHaoEPerGOJux3L+f
a7PaDdqaa+W1KjSjoxQHjbde4MQJOkFDPgBw/QN9fNk39YtuyexnKmeArdgFLiQb
l26kfF4k5s0Q1elcTRsacZFiotsLmfpDIJt43dZKiE3up5UF7otpZkqnzgPrBF1+
pFCd3eaTtxEwVZNbp+paphUveYZsg21YVF99sFRGZI8l9/ShuuhmOr1D+cHoPRfT
iaBjn9MJO4B6dIlfK/CS8iyXssOqTH4htdfAIz1H2RmVTIuE95h8axR5YAU/iwgN
nCnm1TNYpHet1/na3Tm4n4kJPazuJkDB0qtYT9JHcv9EI78QazrA4ZNXOm5nVIjY
LBnkGYqTF15u7STEoiIDdrTI1v4WYBeb0qO3wEdpJ9JSWI0zKJm5a5mj6zmPKD0p
wCuqv1PAzI8CzS7KV7G8C2qiYuFvt4sdkrT+hyrSURNgCK93DGYPoag8iAKQzOcL
hBhTI+utd6bNaD/qvVQBUWGrciGp48Snu8TR7gJ9EQemXtnFYCr2o6QM8w19PoOD
hcSpFJUM5h/mqNvRvw0OZj97NHFFls70vG6m0BxAVdYmLNHCgdQuEnViqnbQUkrE
Si4NAzIyfVlkyiV5XUAJ1fWU/3bLD2uIJH+wZSN8ZgxuSsGd3TPM35gwF7PZghWb
aFBb4XB5dBrHPcydjQPrJHS+l/X8siq4toassH3ydFpqjKBbSFa38KAJxR6ad1uK
uQHC8jcB2zEoU4c1iqJjYn8JrsPd6bBxTvRNkBZvL2sl+xvSQEOnUlEtpbvjk4Hj
mpPIrZqeQwujtUG7dqrZi91p+tpIl90wyMqSB0wsSoC1sTZPTzIfszSG4bVKLQ89
vzdHipAmxBVDv2qFO27gZV5C5h70+uX/Y8WTj5jBMB9VmlLJCshZXcguoSjwJcCx
TIMHVqCV3mu9u9rMxFVx7EvyzA5MmT0hq0IMmrZny39Gjdt0zyBYwhrLJSIpWA+2
9a8WhL5VHRm8iXK2bV22VVCfqpR/xJZYbBy+lgkGQbXKaDNFwbRYS8rqjNE10+qM
pIMi/i1gEDnbHy9rX3HDqy3lxt0qEFj5Tg6o7xCGLQKm8hntaJPjsAcb/If6YmUL
oxS+Gs/t0Vm9b6lpTGNLs6vq33ox9wh7Emlo56+9Tong0bZONZGJB+nlEObzb6f4
gLv9p0G1raoW9DZ60D81yhG5SJSqkDjXXl0oApzVaVU2d3uzDAsTVnPdpUYJpYqN
Td1wu8LnGB2N3UJU7PLy7x8myuh9pchOWfcZlaNOYteVgk4lVz63Q3c6cKLxCFOW
4zht0STululS0N8wi8bMEYeE228WR+RrMAZCjGAWKJzWKoUFJKsl1DJbHFFhzpIG
kZBCuBsfPq2Sbx2C03DWbDx3KXwYgYJtlBa3c1rXdn30krPkCkh3+WE7T0WdkauJ
yS7LdhULWAW+A8DxPYR9rmfqGVLflSdXzQiw0wWyZyDP3JOikgsjI06/ARre9qjM
vD3AdCrCLrM/qzfmYtR0QF4HjlL1gwB6ivq5uM9ZnbamIaiCekjwsR/4jQzperYn
WF7aBd1KlY7Xe+7DISBY+J7FT9Je/Jo3Q2a5Wc5G5LNMt/L5b6oM98fhzOHNV7bl
ixNOnjA0lSFmFkhyrxkYN1OisH1WK81Df1Gr+1RjMd3KidAf3UOxsBT7T/QAM9k7
Uvip/xg98eT04bfzjMbJEjJ+Dfu6vHfWstWw811MaqROEpL5BV94zjWx4np61WMR
qVVGsUZE+WECjPteou8Wse7ckLrOwiOxvSag15kBFHTTPmO26n6HFEwRYT8/mD3H
V38dG8oBnga5snJBmRg4BdDgkzD4tHCYN4djcMHA1D/NmYVBk6RH9rhojMF3OKA8
QEvRJnzxOhkeRwfDNhLWuHGYexw7Hm/N/+JI2s21zpBVcepGBgc8YkDzvM5gFC1d
dEIcmhGmVQrhgOIpmi5SGZN3CE8dnO478tF8Nh9mDX6MH95eVBQRfQsWL17iumEc
mFQt25P71QqYHVQ6rtw6vLbBGfQHs5w0CpdYZqUtsPRkSyX987tWSJNRIqdy1F/J
SPpNKzt6/lcpV/s8n8l+bm2k4ZiH8ad8eNapgKZ8ZaID+UcNix5KRNm5ypK1d9Ds
biNG4cgLq4uoggm1hQYPCcJrgt4xnlKVjHPuaPyevijUEz7z5Jyl7hisvB9KNXam
FvIG+e8Cdlg9SH1HCFh1TUtXw6mYbDxgyOQNTSb4K8XSVBBz4Apy1g/0q7YbG1Th
urVUptxmL7VTfxI39nNuORYp9ZaYrRco9oDRP02biWgf+IOiXXacF9G8NM8nKjY6
eWMZBINuyqVChnpKREecDyrwfhai9/Rkt5uOH4aBWTrM1tyAsgxyiCw3KTXmf60h
B6vgW7Ql5lXoDeSYuwWMZqL93MbuhOgmVN/Ui1tRYLgheVDr46r0mJ28LD1PZLWy
uzGykgt3kM4FlwdC7Atas9uCDJsC+cgHeayoof4PCuKdelE9Jo+pJGz3LOCmWkUH
mI3sR7Nl8m5+optrMtOH7gzwftXy6av5ti6vsA655q7WUPODnfStLCluxQRQYnLq
Ckf2aaZ32BkPSfi4eUCouFLwTTyqtr8QGcYGErq3hbwqecoeUOyExY2X93QXAQg1
Y52d+ryMEU/8F0CLVwc8VHRu3XeRDZ6CLC6yEiRiRT5vvPJqHhdnWpsrtFjyiI4B
gH4ZKHXzr3nz3Xc+eFm0ZXI3tm9NCAL8r/SnbsDcDsgp1u0i73FD8tHE98AcIxOi
TXJvZsCU0EarLFj/9yh5r1qBjDf4vCPTk3SN2ifPGKMNVFePmqj3YI4xXrcrNS7s
P/PekNALoHH3Hkv33eQ7CzjS/fuhP1qlSqSK/wqZ3hNhTgG6ZsJuNUhcHthe0b/J
xJnDnS1D1xT/6AddsIzDwPRzEqBQyXxnOtySzSEe8cNP8x+3HsjKwtylZKFDfwif
K2EIDl7/4IV080qQSG6YtI71VX07NnfCh6Qj2tHj3R368/hz1GcYM72VrjgdQR1U
Sw7y9mmhKnDy42WllGcK4eQxF5i/aLZCQisZcDq2Ymzgx19h4jJeQHctyzU2/eju
87ycUmZYkCUmFc9JkdMcJujdGZVRoheAjy6EdJYCnVvAa58BAmT1VexA9lnUZDsS
Fnp7DoK94X/oXg/Ud4doZA1d4cKRfYtCRamNEfv8uCOSu0JKlAiIf4EO4RdI98NK
/IewWMfNZcmw/jfdQxtXNFlBQAcvBsP0H1a/uhP+MxyInpC35R6qLZ4cnEnyioES
qDT4UNbE4/VUx+1mzh5a11DAnkxMS9p4xd4dt4S8h0KAEkwadoY2Dwya3pucXep8
ajldUKznracWBzCdSZjbjSsBw2jkcH5WMiXOVFLeoJEybaGqNHa5loz+BkE3B+4J
tXCf8CuPr5pEwor2TMhomHQGzdovV6QaJtqKjf6Sho8cYvTxvlaiO27CmC95nMaF
W4fe0Oq90btdjfYbrZ+WHnJ/n9h3tf4pO4OvRpupTkt1E6IDdgcnn3FZ5p6z1aMZ
G/8Arif5xx5ldRiW40SWGCFs5dZufAJ8f8btwo9SwkqqHqgA/zk2KsZuKsWzXH3e
rSuJVtlsKoYVddBU6xSackG3M19KD2EquC41vHt9n85oc0ObLYbg9BVCoeG7pfK9
j5GUmZvEHzPHOptILt7bFUC8dUQqcZlk1Pzh14DDLehBTEJNro5SW69s7vNLMm2t
hT0QkFwO47T6BzjAlLrS01EvjpH1gXzHCOtkKNhKqdxaIr2wo9uF9RcPzQRro4rq
lb8xYxCvjJXDI8IDK+5/zkT14XhHFQ7P4XJDKS42PNOuTj1QOD4O6y+76HNKRmFv
oGoBHDtFzaGzYiMKzpicAWeY51A/4nDW6123KaAbDUI9XM7wC6b+POYmXEAvpRxA
5qp5k/hmnfPVM2C7qiGuBPBfj7KrCED83DTE2Wbch7IupdDgsUtkjtp+6W8YJ/kj
3rA7YehCl4N30clOFyXMzzqFzgKZVTe3ljZh5o+53tI4+QiVzl9JYAop69pJ8Pj8
OQGZGT6m181zMNY6P+PPo9TINLR6p4NZwbua0opjsOWx0JCCoj0U+9Gpbz0ix2H4
7EjfSpB6N8t2wQi/St5SEPYrX2phQhbvwnFReh2IW5zxmgTq8dEx2gjorgxr3RLK
C8cQw34u3/b3V/ZlAKLPRGTf1fYfewV+fPcC4BFv1kROHi/VaVzABl+kG/C+meC7
JvGLOc2eV6H5YzYP9x3cXbUrFVjLz5aLnC9CMRKGw/3oRFTRsDRgSQXE+mfppMqD
EZ9uIFwqsVpgxIij//S8HuUvAJnTzh5+yI7+Rmd5hYAL4Tj4DKxs/PA8e8Yr3BKS
aFL50EHWPt2T62Hv7lgPvHmRqaM+bI7B+/hx74mbm+Stzo3pzgr8OaWKk6TZ8PJH
zmPaFqsxK+kKkVyrJxoOeTAEionJ7oHIv/SeV1qaJANeJaDu5vVpQMT5XeQ61blI
WM30wl4z5E2o9PFlPODVvzcAvk7N5hU1rEtDoAdhcBS2xCrQilSUwrkrE+AsKbvp
F8SC1X7QXXPjNjgVFCUunRqjJGR88ol3RQtnD3ffQ9nn+3c6csl785awaBDdE/xG
+8+mrG8SFYgXOCOKy9Gz5H8FZo67tqFxWFasD6OWwvsWB+8jDGvfZIyzvohlBMdU
iuOjGL6kuFgbInc04jx9+8FQnRubFOXELU90zZ0p2BKK+HzJi3gLz7owFuUt2UC/
xwxQr4LdDqYGkPvKdG6uOyYDFi9tpBMI4W/lo4EVvP/mgqLC7DLnmevu5Gl5DqKB
fXMamVplba88+UiaeRMJR+EcJJqA/vDdhAkAYVZvWdvIw7cGmnScFDLdVlHdp7cc
hsFI87BCxhic+OrvqePj22W2g7ATSgOwKhLDEtjXFgwhJcc2KJ4aepZDndubuxgZ
BBud69jH9o9TrjeFrVEsZ2O7lzbBMAyNV8IDKlj+N19kwr2Dcjoe1iE1jDWvRTsz
6X2lcHEJtMd0B5wDtknTKMhPzEtlK80IIPsX9j8Ipe1zRMuSNRfAsmHogLXmtBL3
CkptBabi8xA4pGNWqiCwHCRcbWQNs+MdKNoWhSDp+1IkBbsgduL2/j3CIUATW9iF
HFvvFwHNLpdcBYwY0IggrWArSHxC9xX88chhrbiltLobI1hZFYk/tlrZWlWuSlHt
iobQDYscrmA3ZQ0xrDFdp/IHmSyS1ggIKQ38eA+LWD2xIql+3HsIhXoXV6zQPqTr
upyolIKrKvhGRouY8DMqAc2dDsdMJzTeBiuvS3hMy0EWjDPmZ9gOpIBXhPypw2Sq
Ld9BdezQ7vlB1euYHwmkUeJCtUaGDeop6yrfm9qkEyN0LdGRUWszk/Rtk8fFPEQm
yCRn3JeCpXGFZEyslPaM6ThDOwo20WWyVa+LfJasFQi/KFdLOcFdK8gdvJghq05A
0kKQOB9r0Ol0vLWOQ0oY2b1H+RVjkON7M7kQ1q6AyuSY+jBFLTiHn7RJz3p+7CTh
equn2mS/smOOkmVy8T09as3vU9GPOBopbrduwvyVftql9VYZ2zSTWKCHmCvKSWzO
u9O5hp2y8Q2LC3KWjw19x1HUjrCzIz9t3mfdVV4ewfQHDqb41GiIWhqh0azaDTO9
Dws0ixLVFEpwTdmEH5PW9/ZFKdSEESxgq6JULO/xUtSd/cUF7zCgLtnt6RugAv8V
soy99u8EDoNp8gWmpyte3gVxbNvgdfn/NOzCIMGCkcegpi2niYvAjHns03DRkCfz
7SFRU8yE/WyZ93FGFSuOBpIFweyvgUIAMqxaCWut8MXibTapUkx19mN8vk8tDCAm
nNdZqmM0TfGcrixUXAmPE5V4znlYA3O5Rtf4PiMI+VgENtdcHzUu1j0BBBWUFdRR
ilflPhFROmR2m64XJsXAd9L8WdWAqFbHEDI0xzLWVXVwK9x0NZvjDA4LnZI3SsHz
myjKV+oc3Xy5F35ITmVsFUKuH7WpqQn6OJ1wGqHcpJA2KHwCCET4ud/vAjRUzzxo
yj4rNauOMTaaqH0ECt7VllMsRee3qX9V/j/pUYn/+AfGEUOElKpuxRGPavVOEpoJ
t1QEzBe0VzSFW4+TcOGJZSGCVLJZFzrpGKzoiU1JtmmkCi95swpM840va2VtZGmY
0vsn/btbHG0vT8HQqdo0B4KgOg9SHSgR7hkznvazgf9GrmSJEOqtJYlwLnM7W92d
3cBGC+3q2qlpBtMU2gHLcmRmiSy4MwOOj6HWQCjUlVTcorXEdkDIqFR9HsQ7lDdt
3KumKwiVv3mPI3SRfBNF52yBS7nzc7bXW/E1tNQobpFmAoPqwnDuhbKCob4qx/9Z
qrDb2CUDMTdIP1uO4ioX7N/+kpGPiOhlsZPY8KId6pELSJPfHIVh+XBJBcwbxqRI
bnafy37DiH+tOXZsK9gNrMRmlXR/Jo4z6eYKhaMybcEpXoqJwXUTi5X6hNIzR8FC
sLyCUnD9we85C25ai/wIzT+vpM/xMklT1ME87vxQ6sJ+uRd404d4gSdXwBaa/HjQ
Btu77zkDhCJwMzMdpGtOZA2Nl1uqK0FYXLl0H2jWUddqJsSk02+uOyHYqIzgyIJ9
Elt8/UMLgdhRKgPLeotIBFmMmshyFaPNzOA5OIaC1Nm1V42dgjVaDRYo0swGiPuU
9FkGB6pO4hMh/RTk/QuNIMB+/i0Xdj27tdCz5hy0OwnWMvXKFd6RJkdqVNON5aP/
2Sr8+MB2LDDBh/6lGmgD2MRZzNLSy0zPBeeev/wZDxODMUwIyjDaAx7tt9NJLDBz
Vc1xU85RfA7GoRsYI9Zg9QaW4SUh6iKF2somtvGjJhnFIOFA223fYTxSsyzFfoab
cs5RU5tj05z4E4oUR8t46i4xs6fihRVMZbGT9o6k933pn1n4zVKdVIFhc5Rotawi
tTpCbWDYetqLvp1vakid3Dsp3YXUwTuNe0Ie05f+nOSs/NTspOGZguP+qyt2XpyB
RECbgozVuL6rSm/N++xnRAUruC7sUZr68Yx5ALsj3abbW0TEx8NYLjS6g7dS+lml
NKRP6PEkTWbNGH8smEunucxKUJSP37U0M20GGoewNxpCA1YNEcron17sjX6EfHSG
cYFgJRNAabMnB5xK1dYXZD/TgUZR7GudyzIuKq8XK1BJC1VzKX4UWg5g1ohzcBqN
7FDtYRPoBhvIUw/zP5rjWuERmS/ioZP3TVTdMJnGD6IHSLKVR3mkHn0nKjJwjlbe
V/vXr2nLKCfkqYVocakt1BqaPNSBd9WmCn6BFrt4/EKj2A10j1N+19s1W7DxDKsT
ZMXlNRNq5HfK0vyrIPQ9diKMe2SbUUQGsTck+aTL+vshPV6QZHMKgeDNNq1Qkqs4
NF2jKS6Tz/J1QlaVjSZHCJaBAXImxgP8fPN02ch/bBIPwHEbArdQ6DuPNCZVgk+a
kR9B452X1iI2WTZf63V8PPQM9U55MflU2hEyCVi4rbHPrjeQZbz7WFtQsWaDwTnB
9FqLuhHu1N/Bk2PQVFmYxKAY4YjP9dPToEwW1s9ktPHDoWrjqMgSc9VtRXafq49D
OsEnodr/ervvTgqNu7GF7NFrriLgqaahKAa8EaoHjEdx2cPQDRD3mwPCum2sjLN2
ja72LZovdc68CFzN4dFgk4mT1OVlzfG4mzlDXrb9HG0HectR4uVGhCVGX4VwM/1H
pVDfxfYVjUWXxfdlAqsodQk8PBB+W8/sy+FqOTutzcpiTSkvasWKyhvBKJQMqg36
plPOQVqWwI+2l3qk2H9/dwaXgoJBmOdb189wMKrnRo0gV5sYuH/ypf1mxOD9nkO3
MAikf3D6QWjaC2FwXS4KkU8p8x8kmc4X1QuAbOL4kES/oA996ZvvAjZul3FC58Z5
4Sq7FhfA1Okfx+eSlcN1/Bcgom8K0G4hGhgq0xOmxCmCoaByvqVKon4YJ6S6Zekv
lR7XSFj4c09Y0twAsMe0kiCr19IhbnTMHbNaHqu+MZN0GVCiu41XBR/UFu4Bdh41
IeHecGYTY5zpKkyDPE4HQq2Smo0v6ldWKE1jv3QoXHd4aljiQhdNdkwXQbBmqlpb
iVfNDxBv1p0mLIKbgopiT2TrOQbhKIisiesyJrv3Gfu7MPlyp++rIamPOSN1odUv
SyCOhVfqtBdeyCdLE6Qtydz6HIPTpFCoTyHuO1Q6o8lutGqFQLZPl87eKy3VXiGq
rFPjuvRAltgXNz/0gKucXXk51nOb5SPXPjgkYAVABeR6fBVkbhROvGT5BAHVB4Yv
YRaSEQVjOcUZGP8wG5k2hxxN5TC/2mJJlGf0BPOPZ3iklgYcBTd0lDVy8kf69cTk
QDmoVjdP0O6Rvj+Sw1lwUZCGWTu1wsVGrpcAN9zjdtCICRSil1ws2rdna390/G55
npS/NzqYaoyzbRtrrY7gOP8L4v4QpvuqQbS5vAUKGIxWPDvG2iEZ5Zsu9uESNhtf
C02HGTvBEpOeI4GRdho/7dIQufg9+ujwHHUlWaX8bBUD1yzWq3EocMH8ceMdS4ho
kl9+xqSvV6QnFf80ll6I3N1dTKi12cQyAtwyWKsSBa75Cgwr1jVh3PqrlV30vIMy
BJzrpCn39EwhpBaMDpNNoDkQghJFigP/lZE1WCQrtY8R+ILLuFyZAjBuSldpMdYr
3W8ya8YlLx5wQuQLDRAteki0lzdfI56psmvmXMUrlQ0zWJ5tVScKlJnUgQ4T3/y2
Mb5oVh+j4pznQBEsB8hMWXvnueTNBb3La8eJaA1EQ3FdHwx1vpkfdAxQ+ik66scV
oBBMV6VwQUbEd1RJhXL+HxhK0i9rhUa76tg08TNrrTbn26mxuX2tttgUp6aldtft
E1pDYjVOZfJJ+z5ffK4vFfMYphbF3W+MXPyUwajrTnDrShTSpWiv/s5bxGIhDXLd
c3w8doTEJQPJoqraCwsIUO4smhLVMuquIksnLctr0MnlU36PwJDO+TjWXJsdH6Fe
AVJ0M0YREpIi+k++8Ovk57c+J1MQvi7z55DIDmI6feK2GktWgFCctaK/PpCKehyl
LCioTQXfiLdKRciA1rwej8+kRrOfcLCvKKcHR/sDEs+SxNbojrxNT3gH2smqQBFU
6hThuIRW8odAL1ndP7713qAJdRYnxW7dxMgYAfIQi+/+kegvkI3DvDhZ2tHHitIb
LkMFu6VZEyo3Z1gWu+DYmzfc6XMe2kI2uY9gjPgBPvm6ar4siK7krgwsbRiSGJiJ
OkAU8yK1ZcAasVBg9a1jkWyp+n6DFzxWvoFe0aDqvQ5jy2qPxRReybYRoBlImZ1i
4DgGMKAejNp0o6T8ooWV2vGY0JvfAQcPW/4shS65w8x5EFpVF3EVuyjkX3u8nok1
rdRr+gMEahDkEcgO1sa0R8gtXOiLg8JK6ughcfx0htsyfme0IVYHW4blmWXD4nGE
eke3J8WKI/qQplH9ftbx7Vv7zv9VXL3mDAmfMl5Q7lHaGfOif0J/12u5QhZXlX0P
zIHLncFLoyhmiWQ/FGgbMfk3a4gOTs73IZ6OIVKJ/bCB0Uok8eP1t9dDXNu1KzF0
KsE9g5dKeMCLZVwR9Q9dpx0wSkMAlGbth0Ne9KQn6AdJQnnNEGFxwaH1AO5fm9di
qSvTeQjoyEd3reHhlfYPJU+csuBE9Cs3aAAB1mLfILNY2DsH4z1e7vTIlLBeirGd
zaOHWdCyAkqNuA/poIZE7x8OCbRZEei/qHn7HVx/0Iu+4OFZN/PIbgrXk4QfLoiP
/JBKLUE38gAnl3uIvsUVJSloNtLfIPfi1m4QXh3bovp0NkkICab1KxZMZJMu7pnQ
/edEDVJzSLMQRDeqcvcMrzJJrpyk456D/gRC0r7Zz5e2JUJkh62MQG0MKgb2Pm+D
M0qjumDGDNZLWbXH/ybib6y5+RRJlIdKDL7EtgAM52wlL4ZNJEPmnaD0FA8+IiUq
Qn8Y8DYKyfhRuOx/jPPOjwuFaM5K4Dfin6m6dBFB9EvFeB/ERwdoqyvOYuuzSv6D
iAIt7Qty94dbBM510CRb+avQGN+BAFdz6L3rs35iOZMsSYrzhTVqahE/Th94vnWo
GrbIchhlSrTD9m967SumEmBKmw88434P92GZ0mF4agBluRVZimhJmp/6albUasuv
Y1B0IUVNHSopv7dYyw1c9HSQ364/uenheKNyXdADS5/+6Pwrnu76zjS8g1EZNYja
C9wqR+4mU+Xl/M+Gq+5FaeqtT/gxUDv8QQymGNQyXYI3PgZrnVGrItiyQ/iCUrUj
4w4LdE4dkA6jOn3EyMJfkKX4Lg6YYtdOIG1opCZC078k2VlOJuo1ZZp5nNVdbsBM
PALr2I+9dDzT6+NuyLdIDPOm3a1a7gMYMNIlZCJ2DASMOvOZMJuibvPBgviRv5qu
hOQi7w9m04P/Cs/8fW9mRt3DvuWQLrtPo5ElAjoCPH91wv8b5ndvT5qw4PnhDIra
x/7yFvn+XhAhLzli53hPFfAJ9lpPYcesU1TBbV7m82bvJ54RePEGDEbo3iioibxx
6OE6qdRfGAYuJGnJOMIPFZ11U4uIiVQJ4OZsKyHP43HKViEHJxqYvVF2X4cGp4Tv
Tzrm49PXIQ/QmMZKwwD+c2gIgNr+2zSj75N/7jsrf3rcn1/nDZM5Wq/tFLBGYJFg
tPrG4pYYIqmDcOLrEnh2t4m8P4Y83WYp3yZwT6dSHXnfboiyjCQUVJuasCjGaJkO
QQ1p7yL9O5K11sq7N8oaU5uBxKmQrSOEiMAx+FodmpVJ1ox49/QAGlwrroRiZPWY
wpydLCQ6zxi92KNCiIyugbnNXqoaGd2pAZqLWhku2LydH0JQ63RUI2CeWNgNJB+w
SivCSbg00eLzhbemenZqq0Dz9oHeiIKJ6xuRBet9wvPK/9dAQ8F1yP/i+aP1wfdL
LVO1iWMnDGcqbhwYoJ+yN2dxBUdJGynADPCeJhMvyyrBqbBF0EMJVGm3+tOR5duN
84ATRTGXgzxUrkIwBZvnwvQk3li7raibN2fUuotcoUouXLUMvthffULlILNoCNLf
faiWvTzbQc4vZc1rxO+63VAUBx/oCMXvxZHT2M7KnclKpxJQIM246DR/Lh9gipwi
oy6rP4PMJ2hmtREFESc+Slo/aOYJVi0Emm6EMswUZXTDws8ACv+aq95q2NOXnb56
HV69tjQ1ehscJp/7StpWURwcoMQAZYPH2qhCKdZ2t11PK52vqoSiIvrwdsOgrVb8
+Okj813PLqJuvEgAJYrx3kPWinZpw1VwWkG+C2SLDse3r8Uw2KzsSHrR8Twu9YC/
UlY+DHY6oeclf/eIBokWaqPSks+A2RUXs1W0Eg1E396u2J3xLUlNWb4gm6xgwsgQ
0jtmvu0Fb14s+5arY3uVBrhFyPrFrCa7qkzJXdBAjaUovrxbKQkweRYRI/Z9c4NK
L9dlQvIy9rLY5RNU0PqDLcGCKOh54S09Z4FOiDqJ2+HDi8YFasXb4Vg6jpED7+Vi
aJfrI5PfSig+C1m6JW8AcwIb5agOvjGNAzCMVoGJQh+VcM8K/Mdlhxbu17euFe4Y
G0XtGhAfl1ox3uFRkjUD9Qwi6exgUjnbQWbZQG97Fa+E7y6oWxvta6ppmt2SgYYp
gK3nwyTm78Ino1jusbZOqfMZw12q6JBuElhki7iAezbpp6FhLCSenH9qWMYRi7mw
VzD9bfTW9Xo1Yd+9bJuPCtgsIG4Fg45llr2W0YNcmVwCswg26vCTqOm1zzHHiRbr
2ToIAIpsJHRz2uxMBvRBC2nDw/JKNr7vEfex3i4nzd1yE0uIoLJRjuhhlkYqXppQ
Th0iE9uguwVG8WRUX/EZmvMi7x3WZiKpw9Ka3F0dpBJ4oM29IgRCUVtPLpLyioL+
y3ZCKIvo3XxaCWTteKsIUfJ2lYNYbYyzEbDQYfYsZjnB+FCL0+AZCWNRZbKedVHx
9UjAxQFqzv/6mKuQVKniiDR12fT34szGtqLQW0NE2Ngi8aR/TLit+eZhJYb8/zAm
j9KBMfzafq9zsf+fAnkmYOofCxP81hpOzoqsnxljm2brMvPhZXogKOKww0u5MIks
p9mzSP1NZn9RbBcrHQaAyxbpAA6D+bNo+kpa8At6kwklos0OfarY+uakTkKD3wyZ
05LmGUH6wbrU2FmugkXYeGNaMO3TPB30ROk9+iuS5LmPDwH1FwQmK9cLRuJPdovy
/2clJvu/Jg+HlTJ3H7R5IZSUOCk0VusVQcbaCwkIzQ4Y4SOjzZRXBaKi0qOUTd4q
38x2Epjw6a25JCwPcSG9qpt7gybPKJ2Kx+aOCzTNKwdyc5xahKsDJjpdAhC8+ZPa
kBM5KNDdR5iaJ80XSqGjbnNqkpFrJRJkbpSZCjPv7eS4MeoJkfSYn1PSXgW17V6Z
F/4jSbE/il1LbTJGIXoIRqz1pmHazi/hmahu2uP5T8zcjQTT5OlWu5buIretBExm
jnFv84twPmzMVkr9WzvUlarwn3FTbswMOWw0PFK/q3fkCts1AGjpKzHwUD4IU33R
soD/39Mfwe50vPLQwBGTRkFQTAJHRm9t993VzU6+RPXYMlsbBXLzWf3T0rEmGJjW
BpT/8KaNFPzh9hm9O71KYOIn1g6lQjUHgNv/eylXZYH8+opbIWgaPmOoRapgExL4
reZXmi96I4UgdWEdaJRQp0wduw/oqrBMDpfhYVhR4ZAwNAG+TGdEH6mPSgyrWbN5
es94u1xofh+jVcDyDXbpaqpxaOqfIgE4iBVTxUWPgncOpwUeMxt7Q8m3DMetaFIn
6Npt/tmVrIS8gWPNknNGwx/pCITE/xBfPRSFwGjKs2wErzRxF00EbzIfrkslyWDJ
Kv42AXBDKi4wW1fnnL6TIlcZXJiSv04fxjeZ3FHrCoLWyYBZSyfGsBJpQBk2bgj1
OEeclIz/arLCt2t+7NXWbSh8CrGPYfZHuclw3QibYAMiICsClJq9KbNY7+7TA+4R
56u8IRJomZppZpvOcU9LePlkNmws3sfKUqFigU/FwE+Zj5nhKkmek6IjjwYJJ0+v
pxapXqjLseT/7ler1dC7psnmQSXfOatmSdI67OOn3IXuTPgFXGqZwq46GPgXUfsU
wRTStXZgYuhqkueR6TbYzrHORw8naEIf+rXjy4IVWSz+mjYlIwbNRIAhWO/aIj10
WzxoWHbeFKgZ2589wXvrGABTSDmrxTwmbd8tFJe5xXpWF0JKqirXQAbAEUZqY7vU
M3sXabJbdIO5jca3pBeX18AZuJGt7iHHZIsiOXZAWvP3uN3Mq2crxqY7b+zSTUcI
QxxMloaiDCZPyJH22rtvsgy+PSz3Fx2fXJG076n+WVkO3JwVv1F2iRO8W7ISHYeP
alMMJDZlPuaiA60zGqUUIlCI+W2P5EAxsRswYbe0r/6BefKYeJSaxA3O33fNdPcg
O+PzFbVMuO6L9iKMWm29UzXYJRURDrbAdHzdKohoCPrtNMx1pBsLBVzWCxbsNkIp
cPqueDgUVHBE1df540cOZFB0LMns9nsdj70HF9ujDAxhtJHKWiMCl88rrWqy1PJK
2kPX46ofKlAmwi6fXHb0xTQ9mTpH/SvYFtgP23Bmxa3edI7cv9d8MN9kKSH1uYHt
Sr7uyiIs1RygLGBISQ/NxTl7mrhlLZ+DDOzCdLnJcN4dTMK0yny76hGCu1kJq3dP
WQB3Fmj0L0H5+6SnzfYo8a309UeXyHBev+/kNnWCs60LJZqdmJSpsz2RWk9JnDnn
8Gn2lX/X72LYCc4omAxqx/Cy5vEpfl3JcBFqaDXJY7hGoNSfiPUJzrpWqgnFNQ+O
Wzc4EZG5LrYqsz4Vxdp7J8qe4ugSUPFyzVKgcZVFwmtoRKZC9ltQrQQ28JgfV9ZB
6+m9GXfi1N2TLhjgC/AjdQi3w8spRNN2BniBBY+6kjfNaaC2uk6/X7jHMpnTiUZj
wtVvN7HTHrXKiuCjLE1VGXm4f+X9MSTKwGl+yN6sAQw8s8boqyZDFJIDVIqf6CAK
T4HcGA9F/DxkOOBij45tG78tiFlqlaGOnuGoMvYsIMUW2B3gF7dkpIf+L2t4QRka
OgkN0gBRs7JZe7kRdL5iXzJp/jTv4szitp2CxktFZ65nGk3R3RUqOj/0m8HPHWAm
9YnjAvS805QfRA9brZIWhERu2OoAlt6h6BG6FWzTHjf9Vq+oCmfdYUgKx9NDJSNU
WwzNgmRfAFw7zIOZh0CcE2RjVMOqqf268Dr0yi6PbhcY/0mLtF9FcbXUTsXyMHLe
ron+d13cktNvVfic50rx5jq6Nrz0Uc0nFVxSHgIdlBQUTvUe65CwNuu0atF+HE+Q
ItGKGkFKnV2IMwvdRg94fdjcUy33lg8amR9q63+MlJQQZ30lkaFY/3fkVaf8ORUS
3cOPTlFtGG45zOWlR6xyahHK0U+l1cQBrjMMzEwcNjooxC3wt1S3McUJIjc/hnIY
FWAWLJKzGLIuhctU3laCwXUjyMijeK1we/AdBA0E8fYRDvy+6JlUFJASFBZL7y4j
0uXgFz6JPjExVLi5PVBlXjrk18bSmkvi76p2CPsPLTAh5mM1caQfYmfyBM7xrJqB
kF31cQ7jMs6I5gaJGD0ns7jt8HmonxKRZu0aUglzfCOu/5bnWEX9ZNK/g3n57R9L
aIppgZCgO7rrGMfAPrnL8kIRKscXmUcb2ZoIG8Ht0FJ5jVNtO0XmQUw8McFN9KIX
nkmhI8u+nstTEYjXbY6kFtZt+1KnUPo0vlIh7Vgeb1YW5bE/gfrjr+8QYd85hixk
kQUd6amYG+hjYSrIMMh079etJiX1XHW6Vxi+XD4vr+kdHrrCaCg5fRl/hS2yHn0y
Qws+St7w2V1fXVpAp0ohhkwqBqQhPfwFlIxyKmVItHfTkEYGV/En5Hbd5dVAv27w
3yOk8R85SK3/8Mb/DM+9hU/rJHVI/MeLBjmxR/EbChdFhax+e1PlO1kr+70xpoaa
ApiElUQZyGtnTlmJyJWXwMznhcvQHesrS4qJcRxtI/Ow1j3twClOPUY8WwQKke2w
xIZf5mw7BMOAzSAAcagP6xd35EkFwVP1s9C0uUpzKXTdoHgycQd2+KiF95mbleam
iz0O6g4KL5OXJFeKsluojKAKfO/nUNUwnmZvMf7t50SjJUZ5PJ9xMCEbPWkNdrEp
w1P4ppJ3w1fuAXhwXb4BGmhy3PKBSTWITk4Cnp6okXykLjcPOJKmKRUb/h9b+ppC
HdOV4cEJafrZS+U+0xuCPMssMojBaIXA5Qs9aaOXyUHrMwWD2bN1VkyejrV9OFe4
ntW5MHsWStGpKJ7B1TRH4H9/L6ZtcOOcppGwh3AnN7lg0juoh7pcTooonCfYcRzR
8NwHRpUzQNCdiWHqDs9XXZ3Fs9wPCqvRmxdspRqOsaGl14UkMEDZlmkGhGkW35dA
xi6C5SZU/2+QRKfCn1Uvmt1oSoLm/pmpar21/psyrF26tjAZiov/1a/E1u/iSi2i
ExGp8tAgPgTgKPY1TZtnFs8rjigUW2903nSf+aYHCC0Fha824WLxVE935h5QAVQE
SzpqD7JmiZ/zyJr3YgzB7faIF8l6gX1wjcvCtQ562+XO8WtODrcViHkdDJUXok5l
6tpwfhFzd1gs4j7uNICuHSMGZBI0pjWLoQLyhPWb8inuvVdlS6kJG47QwnOKF3iT
M5//ATJ0WmccdqCzqheuXbzXemmCOwhmq10M8cypCDM3Ydj9vP7dVTGY4Yn+oxBw
nDGoU8FTIzhWWcUofN7ypSa1o+HBFNV4b207stZeEaXZt2dr1tewu0ISn9nl4zqO
fHHP3cFqbzeTaEfF+hQGbmNTdvSqDc0RMBclyGsft7FvDAgIQryo0g0JmdYOGHV7
zH6k6o0BY8Db0hAmW3HnRwiqs1kbmupWi4e8K7AdszURJs8qGiIhs/h2gYq0a/ZF
uM3lqcxIAYd1uitD5pwaRdv/m4XOvDnsaIfSk+KR5xh5VsnRLhLLV3CmmILaZeiP
GRBnefjz384rZ8FdRmLeRoFuEULhrYhFzlfS3xMQyZXlJCrWzPJ1tZ1TnB7IiB+Q
1ms/a1W9ihdLVmxZViwpgcBOKabg/2UZEx3ULFcoQYkQeRro33Bk00RVTH8hMZ2f
RKFwPgzNhJJldZyT/VIEY3iSCe+KBfSIUsmDddSiTu4D50fGgQPOLoyYu+/xiVK8
T0R5YzLM3qdJagpEJEGKQaX2LhIGZNDhTuZxvsmllzT9YjXOsg8/J3uyrFAvNGEz
Nbhhf3YaFx4A14DNyx/Kq/uRn6f/KzCF9D5CisuutgqlA26gzy1Z8GiwKBCmas4M
PYdLPV5bOC89vQTKc9ZfJqkihLCchBtol5LIjd+ZXfoRfOjKlGxUGIk9PbGu+Q0A
l0prW3DwqcBaQM+2VL5POwB43Oho7qZCNQZ667ky1KDe1sR5HuTKXlTfKrbVImrR
Hsdt5b4CgTzV8KYPCSFgmtp1jkB/iovf7msQXbChLwFQYuY6xFJ4EWiyQQJX6kbk
1yEQn5DCcJ/OsMV1Cg7izEtDDIDLPkiAMIjoh7faeim4tM1LFkDU1yroFSmiNstP
bpQdMu6rPWjeAbYoKHSBA8NqSr/fWto2KajRZX3TOCGkPEttP2OcEqYldqwuDPMp
/g0A0w8MtI9SCffMkP8bQ+94+Jmjw2d5loSxmtzDT2PekIUhtnw/YOIfELH3WrDp
8Y4956AqbnbFBC+3dSs7JfSlDdMh3LlMTVWAaG2V9IIOBpQSW9jWy+E+LDUQAQTq
1ZL0Nv5ZHSGPgYAQ5EydpADeuw2ICBoP1ojfpJ102IMcsv1DgP7DRtY3IFWWvQwE
R0ESgpVxuAqGPoO9FWM8hs/KPq8D8uzY9xuiqd5sRBZ73uL7ITzI9p4EMl40TZ/a
mLZL6j5OjIRpQmY/3D41M+WDSBrUEYgZJAwejv8foaIaWC2JzuhBkuTnUSxkmFCg
rM+NGe/UYAxr+m8PrxwfJbbKbyZ1xHbEtKvb+OgB39i5QmE9eSHVCWzrEMdgFGW9
9XK3O68J0LIvI/r3rhOEutj29DDhKx203Y1xVf6UdXoELU5zusnoll8ouSsv4qBi
axuF2K/NKwgvz8qfo9PZQtUi/dKnvDnBJEYV4swxWQ+Gl7iDwFP4VRVl0ZcV9zwR
Y5vfqvDyhnla0kkrnnHDOL/9NJNLMenuFLKYSMpA/O+w5uw4sHnc2+nUAvyzUhHi
Q5D7qkZsZdEQ4ajrkRICA4kQAKi04TziZiRRJ0zSa8aJ8yfY/7qfQnn0J4OlMLp4
WJNCuJhe3SnfbvHi40iLjIWVRjTsZXcXaYrww/qMDfxNtIySzk4PH9FfnLn/TSq0
Vo29gZOTfTCSaJWewciHCC5WL4mO51UHdDiPon255ohj1CT9he9LTl7bOcaiUIBq
XIMfys15VF7nzbpas/rfW6a1LpJDy/EMOT0adRv5GQ6QFYAnGboy51NuZV+NE+jS
rQFsalCP8fsFNQ9oeRCs8OhOlGczxkMgfQOmffmWBG5nmPNzmbb1WNksBWnqBWni
9UKEXlXbXNON35PIyZevFCC9zCcVNXqF6ZAwWdzF8VnpUFTXj0mblEsFPh2kWs1O
ynPPgvsH062zsMv9YPifT+aHPMR11Jy7eL4NLjX9/AM4Q33nlzziVSXJDS6zENLr
SqSZcdpkpYIB1IJq8C4xuPItlGzRY6Avwk6cT/b3YQK2xSNW4Fm6CfbfM0SzJJxd
BqZzlG1PVr8S0TEj64uU1bxtW8hPWq7YnLAaGUY8wUpGwZrvmNgjpojnbOon52xn
Zp261hCneL27gFk1vGg6j9unu1BhUV7tfEVJ17dqTKouNSiNBAc33EBeVaDo8O9s
ZClYYgA3Rceu6/v3mKdFNXX/KhqhlR/d7rYLDZKNFwr8JXCfjlQsjd6nyBSyziI2
TyFGH/aGYt1pJeqI33SKp59m/9iQNPfLtQ+66g7fuVRuhqAnJ8/mwd28jx5LOq+F
vs0gMFvl6szf3qINQDv3NPmlA2CKCV2KGPABAIMfXp5PX+B/eKIb5aQa7hik8reF
YDGrJMbMEji5sbBrMVzBoTOppVGMjeIa94ZE2s5jsQVLzOV95vswyYcPlZ21ZWG9
ZiNYQJ4IB7q78/xln3OSNYbScfFi+pP4TnJuCk3Yvhr+b0pVkPwPAr7AERFi6PcB
T9XGk0/1nbzB7LuFo+hWDaY61pM6JVpCUdK+tExhHnxZCh0uxrK76NgJxvoctkpH
7L8mA/A7ubQ4aZQzDs5+WIxQPI56E8ma9cssL3E6QMuGTPSL9zDHHbQOFJutP3gB
zZybemL1ype5W9X4iZeQtaesr9ID+rpoYmv9gLGHvDQSp6HMvDbdtsG5u/x7xbwC
2GZ0JK0egqDIahImIdF1ShyB+Y/tUnEUvIMS6ASorJJA9zHcyrxviHIQVL9WSIgK
6gZ0Jatob7tWQ1EEBMefHBAnFGrgVuEwpFenH4dqoMMW9nqHuw415Ug6wfFi7E1V
Al1fLQUGghtO8rv6ucqwOCTx6pEvMO4xnOefYnSyDRkfrVMWxIkpFl21hu7XzsQR
ZBReNnQ9saeeFUWaBRRHs0fTYLtPRFFest2gM1jtF2NLGg4c0djWtBXUOCON6qLH
m/f7BWJuImFyea2zkS0EDgsX1Q9R9/NTMggMmzQUbWMfKxpuJPTXlSwMU65PkiFS
FQ2A8faj8jEobEoAfbEnn2VWKMS5wZhafGVzUm4NbdshGqW1c3I81n2NmMxyh8+r
EPvKsdSxwzN9e7afq/Eg9sxaBozAXIjww8FZORIkOB+bzxY32La++VnXdPmY5wsa
WmO9NdkRniAzpLCtVhEqi9y6OyqWUcVJjMEfs1I5+81L5tZg2uxa6q/pg+o6uUBw
sRvo0EPAnvyy7bOkAYT1RukkTSAs1s3rUnqTW2xEAAMU0MHwCNvkvDi2pHGOLsRU
/OK7gNGOhbw/+7kygqwZ8SkW3jlMV33J3Of7WkAdBm/+XuJvSjP4yPDQoTSOmrka
AbUsFMPbGPFPks/6XfH4k8IEU7fCfUe0IMVW3ICe1sUqTkUqJBNR87bCoCys1us1
VgHCaLRO2Vbw7GaXFEjxACP2bHOY/8Ly6oj+/qVkNtHA+n+EJE3YATX/+D3MWsBH
yGRKySh23G2ei+q/uq8KM7XInEHcX32EyuXocIeNv4wFyA4t+kGDWghyuBlCLnlz
RFx+HUEkk7G3pB473+3R80Ndg+icNdvJuyUzfytrxj/m9hDq72SwnIr1b62TvU6Y
WMoUHH13tZH1SvWh1Kh+zREe2ruUC3ekOojLoF1GtbZ9LAwNWVCx4UmOi15y6klz
AChUx9zkbKwAcNk4orbaF1rz9cNOTtJxdBLDXhB/m4suwJaqHvO5vHqdc80TfzvY
NBGxJBZt79izZp5KKBLPfbBfAv6oRjFIc0O7QqsSW5PLcVqXX3wx4rd6LSeD34LE
JUtCH/d8o2pS7p9jCw6KNoF7fdnkUz6Hqyd7KS6exdbQnwYtc9M4VJEjbw8Dv+x0
6zH8DtBrZijcrtx/mEWCG1x54Sxn5oXRya1BhVOaVfDdXHdrXCS0etYq8S9Wtm0J
s0vBz8AG/xEOFN5j8CQcHdUN1VxL+hJquX1vb7SGrQHiDUPoOEedrYTNLLbZI/9Z
N2mOJ1xR5XZ6vQeZ8/1ShYuHPcnNyvMvl202eFDKDifGGBU11gUPLFtz2AZiv+Uv
TeAvJ1fD301WY5mrCpXAZkICo3mNC3Molvdb9/NBf4/7mHCACshVph0gvpYEkLEu
bLu41/P/YkKuRkQB86q/QtIFoFTcCXojQeWxk9uyNb5BISJt9BE2JemVRtNceq1X
CTQ8xK9LexRa2Ov5sS/yEOSsJ6OBhrdOleKEeHnkxDSWtOgBKJLONrUu9QMoZS0n
BrgP75BpDG6jd5TAZcxrs1hnSSu/FPOs6nkWvyL9/ldxdF4PdKB0G1URE78ts4er
Tn0xH+AwU1m2dH02+1okJlXysEIWMSDnkZRsOailPD46vxy2oyOOXb5tOXybQ9kb
sUleVELC8TGoNT4q5/MM+qomuaVn6YJQDJfPq0EJcO0n4TKb5Ui45pjUFXGCUo5Z
yUoqsIASxSg/VwFOaE/apvZ3YAFZEMKrcAKW67PomWVnlKFc+hIZkGpWBw7ujJlb
V8gqVeggosbDwXDH6sf9fOceh+p/kjhVsilZiE0Xx4dylH1LVSD8sdISpjhf/T9z
bwvkye2eX8dALeCeTSvcGs79uEFHIMjgl1HhnD7OFr68uwUBCvBgZIcWAm/tCX45
2XvNrP8iqxi33C46/TAiTqTazJRriWOsgM/sZCgb7nr80xf+bivP/4HAqa231tKx
GU7ujl2+Qh3ZecKf/zPHWcNTCmA6RQISnexYOfC7rCUf1y1neaOrAXnAn4L4r3QX
Bo7LR6CsoYRsymt3r7RDHgGF2uof4Q4nYtFLVGKoNP/xeQEzypbwd+Fd0kQ+qVGl
Z4NePdhgoBHXH4cNh6C3b+tp6Kiq+/lyZlep1J1BWiX5bSNZkT0BRBf4YdbfJaIm
RZuBYxqSDxoK2ToeOhIJjvqRucTaG6Xnpwd1D+1Qse/iU/NU++XT3D4sGYFfUyhx
FpcoAC8Td3E+seC+pq0gKfaKG829i/Df4JpQu9+QYV4aOcVaKxbpBsLQXc86E10p
MMATUnSFg4xw9AqOaz4op84T59BzbbovHtKFSN6uum5bPE2cyRQRwK/j3R8y11he
Sp25v3+3Rh1osRctidSXvO6ST0PVbKtUgjSqisq06BSPncS/BTqZn3N2I2HKSWnm
tE18f52GQzwnWt0INaGDPerGht8tOeMhNeGHxRJ+YeQlbHb0mKVaI+Q/i1ks04GE
jUoDIwGML9Vue77F4Wac3BXsdtMUK1zNmx7r2T8q5xeDZ22B3xeTwYyrI/FPMmBE
EsKozqYq45vPy7UR8A7ApAhrhqJ5NjAenvu4qWZ6r8ErPBH6uVVa8cRZbledwt8P
UNUIgLpXWOBpjafrLiin6kpf1P4n83CjM+5L5DmAYxYRaJPT8Lqx2Gd7YpUA3CO/
bCsJ4fE5Ux4vFhccQHG3eHucHtfaPJ+8sYQeUlx+MMdNWKNiauxu0eVKRlEz+VGB
SGkzLT04WcY2hMSOZPxwXoLevGoRQEwxy5lXa+F/IUpl5OnXUyyRsQ4OGzTABSM7
HgXWp0oMbL+ae46c9DjzOyGZhnfyD/+wRV/7OJ402eUD7NNCm/VzMoE1+Ozt869N
E6kvh5dZQkC7+k6nGKYVVz18nyRDe0hZ2nXBhPqDhhmIHz0+XGBaAhtN8H7xbAuk
75SrkFNEWC2ps0TTBEqbNYipWAAxTyn1ZrixSR4X5Jo6AMXIZcfOEQI08Pex4IN7
jNuWMm2aj+BxY5RJGp0dYNF7uP5efpSCyGpTGJPYI0+9tBZAO1oguyaGptU+tZvm
ptoTYoFJVnO7jI/hIY34lAwvlMBLbck6T+d8cfRMtirj1a5bT7lX8VGxy2oQj9Sq
9b2OKt+7v5CgP/9iE8yHop7dms0QSYcZ+NT3twqOIglNwlaeFJ0mne1/RgvkC7M+
196lvCv6a7BtAAPD6cqLAQ0SnTnlwMaDmFQ6GEzoHv6zgXKrV8I35OXiNcgOIiYW
kuAy075D5EiCnJGVC4iCa91s2T+FDZTIzLFXSgAUaPUwrIzz2F3jzb2GeFBd/Vgs
6bf5uaNapzzafviRYZjPsErmuJHmTCiuWDgOOKWL5Ddgl8Ka/J4weZEDUgnO5W+v
8UPGmNE97LEB5FQlc/UDzNpX4YtvnBoJ7+fASbc5J8Yh+O0BeLvd/bubcQ2D3BPn
5rN84WwZ7H+6A0KzCmtywpaSEKUGhfhdpsxpbCv9w6UxfuhOOsNnz0LsWEV8P0o0
BXuCfQVjQ7JE+84uLzEH/7792pSHS17uypV7gkO6JK1WbnUKJRLWVbcS8q1Gu2kG
rZ/Bf8kQJNtbG/Zh3jGGDTSGZEEiyuzAcIjrF16jUJ+cT1EDbt8Zte3Hu9A9MVl4
tXoYURNq7x043mkHTMWFCr4fVSuqEVe/gmqeI2eLTYqmJ+VpF7i4zZ8DMMSWYMyu
4J4KXaiSGq3JVbSjic6xnxEoU0UrzaFi46TS0P/mKPPBVtn37UfGVT1KNfZ3Y7hp
LgeDiTtP4IF6e/BzoejcEBDMDF0eB3QK9Z1FHDbR2KA+RFXCZ2fnEGpNPTP/Pa7Y
HcNFcd7AhOfvCAbMQ6EIKc02vNFW4qk2sG3WvtdJERy/jf9PATUi3nAyhh2fkofv
EDLP+8EGV7hvSvsbREr6NKk7cuUxjxlj0CmoLxawOj7uGp+tqBWnwhac8EcMXY6X
Lagt5o0hJdIdrVOCOHgJZpRNOiuYjYlZsn9uszUsRjPUfzqJBn2guItP/N04taOB
g/Hrwnfdo7aZfBUrraLnSobPkhd28EqpuXS0+gs4Ubc0jH3BwAlH9VMjwyz4zVnp
U1FUdVrLXo9v1bfYtyEEjy+HP9ixZiYwOgdarzwiMdumGmfmlWp2j364RjBsWTO+
y8g4tfg9UUSkP4uj5ZFUd+z0UmkR4rPdkXcL+UVRxto/O5udA14m7m8ZpdwnAAZk
waDSvFctDCnQZPfGzEsdvZsdAFszgxn6mnpFVfWC+IFf0Ju8R2q+ILz0cPtr6YYj
f/nz6uI2baGuhWDjPkhVUCEbjI/B6YXjP3h9rxz1QVypJf4dyNr/Vf0mvBZFsmeK
TUnKU5Ru2aw8ChVb/QDJB8Tv7DRYzCdf7I3ySgZHahWTkSh6MUYZ5L0entFiQETz
rpATppOapRt7mzz+rfR1/EubZhfpHs+gvQ7KrxHzfa6BTSl1cVcJuKdVboIQvYgo
6WkJuOQZJ+FWDhtLtoCH8oz4ujkS4ckNKnHLwsTn52R2qzIb90GSkibZ/J3HJCkR
BQkbsqPaRfIkJELo0hhvxzCTsRt5Fqy0AS1XuSBJIx3a7M/H/Oc0vBnDtvTXbhrl
i/4X5ZImflGNX2rnD+mtWMDE5S7y2CJ+Eg0lWDhSKz6JskFt+4GRY8j5FcFiiEdi
Z+sQI83afEgo+icMelLivTqdMNNLbFLGjFa8XKMCOfRjMxuL5t0ltjY7A48hzts6
H4z7IjAfmtzF5clNKr7vHETRsVXc47HhA6lh+LXC3IPtCwWF0m7mx7+zDCZlj+VF
y2+fQXC8ITKdtcKb9LoDbsGHDXvMPDsE6O2riLUoqxA+FKH+yN8/Kvd7LneUfD8x
sXaduK5NBQ+VOgIL7X8eOMLKUZD9SRqlXVCt+23KbpaA/gaH7zXbvFDgkgMT/Be/
NpIW7UnOa6UqOcJ7gaAZZMnEUVrHOn01jPiSNipShAwEKT5T2CkcgRoqrqSzNWWy
RXcMtbmWRNbeoF2W4I/mE+JsCJvnbpkDFYVzRZ/W6hTac9eAMPljM/Z23v1N+wDi
dRsq5Q+stcsBaoThIRzaB4epu8+mKN8/ssheULX5aY9LaghjhU4tQzELBjmLILof
YD8jzFdGN3XORY8123xR2eegAUKes79zzyxLh64ARx4ht/3FbN0cXB9sp9cEtMgQ
vRQktzPR0vkPst5Vsx8wYhHnoqoNynruoyGHlmwtzSiejLs9MxWAxLOfYfLCgI5g
ZLOwFF3agQ6BymFyCEZADNlGcxSEEquNm1K8qBLYDXQFf2nETIhMCrce8lzjiyNq
fl//mHhkXqWTyu0+WxBVeOpSvfmhKqU/BPTC21UDyNT5ee2zV9asOByXdJ6KYLU3
4JZxqPiV1iNYQ+fdSlnirj+MV4HV/23e1etO0Sxl8OOlj71jFDBU/f5k3lsqWKtS
lOCYC8szny7X1hoKYqDXNdMxF9YQANb5RYZPTuIr+8/EyhYmhCDvzVZ5pvSFcQ88
OjaRcY2EfmOTSMnhO/MhX3tDQtCh+5PPqp6uc2wNTFVyqEUD4f5AJYEubWBQC4qR
C65PV8iHe/qRrraMHEimVOy1MX1Qr4F+CfXO8u5NBVt5txCMc5+CJ6gCdxi2uUt9
CSl8QZZ60yigcLHE6nTE/OvR/sP7nUbxQgV3HcBYv3pWiYV6Qpcj1Zg4vl4G58gG
Nd61YZzk+yc7/rZF/m3LU6EDwWz+55w+roSkPn5IFtF4CW6nARd88qUKifc2IE9h
WKbaj98OT4/l0yrLHo7w2t/Zob1wdTOB1OT7OHqNcbUj9/klxLYyHtQtK0y93lWM
XA7xTUIWuTD7hXx5hE60Gx0/9V6ZzZj1VonCULnBOdiE+aKy0yTERFbx2L9aBKi4
P7WSQJINJ9YIuBRUBcRRdtmqMKxSvnnwsKDNyTp8QvVt2xsT80rNZmTiDLmWEkfp
j9cZf28oOqDlyDu7d+nL4ASmOzfY9DIyTTZJ9wu+uj/3/cpCjTYj3Mef3h0ROBWd
IG31atHb5JkntmAjyLfpmV5ZXH9KITj5ddwszIQ3kSTkdLETGmOqWgRodkiBEer4
XHqroKrR9+lNVVxSZi7CF90dajJMbsVNyks2kEopQq4s16psBb1OaZWL7Y3l24Pa
IbNC3P+aM3v8KWhuic5csM7GF5tNHSSiRKgQrPnhKkVmD/H8udLqhERJSV+jfKty
NbOGn41iadbfgUn2JqNlolrlpsEalKWrrMShDO80AVzeBl0PllUvL9roj80con69
h7gqj4z89A4PmDUVoblVifcdgDmCyOtFCMwPC0p5WRGQ9tNjIgzZck1gBCc+1bLR
flh9zc88Tat7c6JnqKK0gnhxjhSa1dyvyyUJW7NInO1/4asCbR7mOsxnKe9+wLto
Abi7cwLw+CGgeb8MYJPvJPDPclOIal07Hze3LPrjzmgeNHXFo0yBzsapI2+USj5G
oSxhKd4m7oRV5Dzulqt8F4lilgkdjePl/yb0H37zA5oIlzHh82EgQX3RE2cUJez1
wwkCZHOgdgGNcYXluK62QLAJZSn44djCSHfrIOVE+VegZzWvGkxoFEuIpnLS62kN
5jv629BTKBHvCZr5cb0z8amVcor+KBWhuQSZdjUFwg07fzTCN6bfrFngdywD5JeQ
eNkdziZ/s74CN5ILKIkUdb4ilK8hmzrlKicTPLafWN9kXW3IW86FeKEch38aZ0ax
pl0gSU3GOBCF4PcyfRkV7454h81r0LzPG424qBtv3lD4ZlBjS4f8Ypa1XWvXzjKw
zbx3ZjS2OnRaK1/0Vqd3uXvnC7rc4LrdlK5cai2VbnQ8j6JeauMjRWt5DHMJohbX
NiXKs0e8ZBsN6PXoLNpg792vI8Jwah+HXEQ5JyUrbgtUH1sPjnzCv114ihgDCzXA
SvvWgRswwqkleAwk3yVXBTMaKOAHUqFNDLBwJKv62ybA5nAo6FvCixkMRtoNFpjf
sXD8pl/f+jBB2gTI/eTTgf4phdMhQ+i4p9cve1PHt2UkcZXnQK0EOV/zn8lObWCn
1YxJpW0B4qyPa4qnswNtPHLZIJfC4tJ7ze8ApaNFKJEePOfcFoKS+NRj7ChxKvQq
TlbHd2yr1rWM3uozcqsvavu+yglVqVH30VQY2wixZEGWp9DZZaNCAFADoWIGbYVv
PTEFmqRQlf4gH1mI7s1Mr93HrlVgKvI2flDc7Uz/iKk70SHVzIwiCQbB6cz/L91m
p2gSe+vpdYCxfC1irChA0gIGiFemG/Ai+fyywVg0UBPAmzH0Vrppl8n8g+AkxGZN
YOjQwInbFU4nfHH1cA66n88cKw8by6bNVkfqR0J1vsLu1fmDAbsZ+u28WQp+X8VC
4uueyrv934vm+FiCOPjS+3zB7AUjrmOstINdlhNELoHqhmaVp9s/AkhjJgNNBsIV
KPPeFfKlaIGlpqKHpdR3BDQQ0y/Lk0S2g+94qCiK04opLJFc0G4KiRv/nLPBWncT
QtY3z7NihHoHyicsZQa2OF6BBeOucJ3+ICYP3fwhOlqQtblYSxqW9sEKJ10tzZx8
qbiITTbD1+Nbeah5gq1QpwY659m4r5Hrv7ow0l8KVPkOSxtJFw8rPkP5PBp3apgB
Cf0BPE/bKzp0Sj51KlyWPeiLV5xPToJoobmr3KWoco5gdqxhj1+ttR3Yv37/+RFA
LXh0Gh4VHRZdvlvt54/h3deSzhXQ1esVIzIE9kErmHHVRGbMLhcAotSw3fd181U8
UCYBmaj6HtVILojMGTgxFIo0fGc9XvoNRiwRT4dbzVd94+ufAPHmWTYU0jmrbVqn
lD0Wk4vTNP48pSl08JbOQSk0D37Efn6sm+uBhEju6Cb3AVQLFLPGuwgWA7cAx2qH
qceoXtmVfLZ5I+1fJ0Q6wEXFRTF8qVKPIxoDe2EhsnieY9c3auRG0hnPSsCSWpR+
wCcWGKKbU43nDVKZl3bUFuyeQ1IaV0wHvVZOKDTiZaAYgW0BVSKwy9xxMpPXuwXP
vzJOWjR3fCTrhKZpsb0QdnzRVpW2ZCgjbWAy0UAS+4kVLJrgW/uPN0P33SwOxhTE
F9DR+QVKxl4EyT7/7AWZAhuu7AnUxtke2/OLrpxRnrU6Xz7Jw1qRTKyqaKygg5hC
nDZAEnsbmzzWKbiwoCZfoRriFsiXuNBl70lN9435kCG0jdhKPw5PJdiFXIgcAkqw
Um412Zx1J3oU9bWWOqCymo3nn0eG8ep8lcYnpacXynMC3RPPgkzQNtn1EHpfuD1/
rimhKygdKT2mERfTvY35WHhTcFjAesq4u9qmFomZBPXy7b5q/uT76TeLIL1lFZ5O
S96/U6kfKSUaOZ+h7m9P37+auwHDB/3XLoMcJ18fWerHdY2mGQhzQzPdCQJe6j0R
i7p+ku3UjCKET43r28CyV2ZVa7Kfv/kJhaaNqdJ1wyIcyMkoYxQkcPk7qz3Zd7pp
uG/wWmUyzjkf835r6Tzkg+24LNRRBrbfrsLp2PNkETXkQuJgMxAo0dcFasMQQH0Q
3dwKs18uuuWd3hL6K6ZfP1MvpvdaMLbxFPdOuYgRidllF/eCy7L+ERQQHJLTACgo
HM4nW0fiMMhVNPvkVRzD5/fNpCobq9wfh4s1IB+cTfAaB1pDa4IyoMMfqoKZ4bk3
IkIsaiX+1tWcpIEP9pBNNrrM3wMSrXNTIX3YWE3hkaKKNezyx39m9avziKHKi5mO
M/zOGqdbfbgqK50GCKRuBUeTow8llNFyngQIuJmQEKnoVM8m2Uj+iutZl1Ig8jgg
v8G160O+MBJPDsFDHl46vflUNNLId3bTQ5zSR4IiGBgc+Ds0vIUWNfeX7FzujAeh
VqzOamOyhi8gcbSCkYcAq9sPHPokRx8oK6Vp+MhQzSvsVIoLwPAigRAhMB2tauG3
mk+WBDaYWzx1NLbnQL3m4/WoPRTN0qEkpHfkQhiIq/rcnJ99W9OB05lF/ee5Dci5
OCufP0nSj1dBNzxynez0BQJ+pRooFE+/JmSypOzb2BH/D63smIxA1hQ0Sekf0von
IYwOoQuJSg4vWwvLQvOvUGbPMU8PSwIYgIh1Y5JsgdPlMVVEnu4EJt7Ay7F8FI8z
HxFc2YsHdcgNjZO44pA4q/+0WayfTyAapu0cbl33dKV8+u1xoXF3q0Ke/8Z8qYYu
zPHlZ45WzX0jaROLo6uJjQqHul8SVPJbwyqc6DBjKnuxGw+tOg9LlmbZ7DgJOcSa
yFoeOhElCcRHg9D1I0Zs4mCHEIwpHEqOiCQCRSt3zUGTOQ8RtHb0w5eK3eXFmC84
v9M/vz+gmh4Pp/AsdP1GlJ8Gw+chMCTEDg91JiuvMddjO/yr0xeUzf0S2xty0fEK
gVaU996F92PLQZ79cyGEI4ysbqW2bnsGYZmTwILguy4pHRsPSNxJYp4kAImJWMMJ
Xlc4JICzz4ZeQMfUtIp2h4NdBaao/vM/otpf8huRNaIxSNi4M1SekmTMlPeztohP
Qw0T7QbmUzvA5gBwEczOjGal/UU/gczUbaYNet2p/L42oP/DkcknADLXZimMFxek
Pm6yiG7+1hC+tORXt8l2TpDie7YuvrdcyqAy1jOT9P3BDtfsZIqupgqGHd47SYXY
lZGrtgauoNIPFaoqzLl1op6l2l7MdP4trYD8Yq7PRQB7MY2XiPozQSZX/l/XxjGj
AyaaKrWuQOGBaJGnd0vHUsLP6Rp5X4L4SnX79s3wGbzW0zGp5w9ZQ/bjwrJ0M+Hb
d3qX43h97h49feyD0KGOQcvLH6atLSPLjtZUy0AJS6ISYiNUP/B7nVL/RPQ88Oil
cSHOROFpekIWGVXz83ceo8o1g77+GCj+eYvJsO0a/Jp9imHppvQDhgrc7G+M6q2J
0kBsghLEoUtXkEbI9re+poBu/rtKnff2aKzYgYmr7COugtHGjzCJ6PKNtmutAePj
F8HeQVcHi0FFKh1wjDrCiMEWNSnKjGIGsm1WMSLSyLc/UQPGCGa8jgSXQ+CSZEU5
DJSTzaAMLb+o4zaBVFuYru8Tdd17HWcC/8/+q4EBYLKFilj4KLJ75MTvKw4pqswT
YWbNTck1ipHG9hWD8JLybR0FSrc+frFUP1quhTyYFJjFjssfbw4El70VGLJdvbkP
M4VcFT5K4Xn/gXfq6gQZ3BLfJ2ujbN/VLzPq5kVzp9TDCvDiUCIa7dpN2BpbJxSg
C4oVleu0f+cYwYniBrvMSCjRFkkUT7sfjl0OHMUe+/k+os6vL6p6Hi5vvyfTbQw7
QWrlIJNglK6eZlZnc4PnQnNgWo9nchgikpPscCJG6CnbpDfqqxIQ5zQAqGOLavXN
WjclB4iBOl4UwWF3FsuNtw==
`protect END_PROTECTED