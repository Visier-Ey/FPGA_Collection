-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "N-2017.12-SP2-4 -- Oct 23, 2018"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
kLk+MlsI16EmAsiffK0MUMXciGjNXrq3hm5xp/yVwypK7Vk0mVZlsSGIBsuy9i5E
9mBMnw0KVayPdqNaT2rc6xoDV6juCuCiEYN16xhsRC5JGfX1O3GHxZPn3Ub5Y0mr
ByH7wiah8m4FIlrVjr2QjfrSCIwuMdfQ4KoJL87EXq8=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 7984)
`protect data_block
5Ct/5QCUIhpF52/1AEgzF+2k6sw0uD0TnjGKnjUiVbEgG2V5rvRQD3tNL7s5wvpA
YC5TaN1R9a5VgFgt/i6PvrJ2Amz7KZr9H1Ha5Q715aJqL68+6gCnGYd4F7d71eYY
HTA5ITqUwFfOEd7jQ0eGDPWDIr7ZdV27brAeV8jPve16bp2t3u3UY72N2lFl/zE+
bKUnrU1oRVCoD9Ystn8xJLbgWAGfzK1zYfztbV1XosNEy/Gp9q71d6FPGKzKBC+9
69HsAgBn3V2iU1N4atYV25FY4tT0IDLS6PDafyp+o+coVbY//lbGwKCjCwySttN8
OxG7LFrslNYT5XY+A3tYi/+1Gu3v9Wl+VWt7GkyKu7ZDdU8zL0hm0C8W873ke2b6
b6qqeHXSBzI2Arkb6j6xjXXM1zf1xvToiS3P/6Za1+wHLr8X8mbS0BDTbVb/1RCf
27ZA0BeOFynP349d27ecebwhu/WFGUgCaQqp0E3X6fhBGyaHbQzzTjB2eV+EAPq3
aJbQjpFWOIhNueJYE74C7bazjXEeftHesjOX2r1oZ5iMnRNJx1kWjorYIZZjt/Tg
sahHC6jVXAYUOaovgExK3qkiH44/yU50Cs4H8YDkO8Mc+CCejyxu+rGTiG0HF1KC
yhOdwansm7WkDCMrh2sQdi2HsQkekWTAyNxUgsyBOaTOdC3bI29AqikVfxW4PAHo
yI6x0rs+cVD+BHm3AohIUtDmepBi5zhSCvdYBiF4j0GRHPf8maNpk4oiJ7WulILw
vhbdU5ZjFMuGruX1iyGMREFW7ELl3IBQoZOx0StNgpy99G00+3z6ZyRjvKsgV6qe
wRDRRzm9QlWCrAPlSBuQO+Wu/EKgsgIjTODVyKK+gQDj0+d1dRca4myk1NJOzpGT
nlEqJL2R27nAufd4lX/S39LiA/G2f3eEz/L0gCXjiuXq5cfbtKl449HLaAFeW2JQ
QPFI8LCkUXnOTjNYiLI7YIoZzsfbk8UfAY4B+aauRuNQfG5qEQMXuy65Pcwi9AV+
D/cUoeTNff6Jv8CmBIvTU9iJMxsc3g8XNF4vH39JjiUz0K84E0Ia/QcQFSe0u02a
1fxEiPa3gPZGS35EA+Igsa1UCTSR+TWQQwH8ddbSXlqT9pbFA39bj5hd9xzms8Ah
8wVGcRyCWoaNZKzqcsUhqnOvx6bRZxO2CVR8jrd7bTseS/1yym5RHRqMuvK0zK9v
5QTRpTHE18KOfFK3EdiggK/irnEJCO2sTaUG4WubxglodfjnLMDz0wuv7XCkN11k
1lWyZwnoVYPBmUVu7GKmngerjWgzVc4kJnrAh6jEvrqfZ3wb7U5whg7IL6spaeR0
Zy/PqJUAvQRpePoFe0b+vMH5BV/Npv8EJbDlppoLS0dj4g0QLx81wWGU2X31pMNY
4A/T3HA/Vt+hnNjbGNdxzxUtopcz62VXDQbKmQN5pzDI/dhjfd0CI1ALZR/u8sps
46Dd9gWpYm0YKN5ARzrHMY4oQuPTcrS9enzCNQw2I7KE1Xb7lrMm0udyk/c/8haA
HUkJRQqvSAFw1mz1LG/xjy1QZypHRBAwCnHVXDzmFS0iz6cYXUXl0siX0C1cniKy
Hi0pDr6lv6LzGi2zFJ8xO6o/YI/jJY/UaTFpjcq+fDT4Y6emqjxk+D+Bu6y9TTFA
DU+YKPO2LKbZvHnGfHEfdnTT7Cp183MICHpwAEgTB2+zb5sYUqEeRCX/vxKfoTbF
QH9XiAdJb/raxP7edncwCY39dFDabFakWj8HzGFYhoCDOCxIst5kUXJ1AcD7M5Ky
ZT1lci03TIV4EyM9z9kMVlCAh39tT2wOyTZoUhxehkm2294SvPHzOoYeigMwSfa5
WG+v37cI7aZ3QhYLLr2/DdgcWEIsvO/VbCEEh4puVbZKAHxqlxbmP3VSlyaZ+TbC
hs1LkoMTgfpSygs60q1JE+eBVhw3wtZzbE99H/38QXDjWIpfR0EqXFzLpzGvhaKg
CBqSUpE9VppsFI6xR73m6W/0OSrLDDvM35L29WIryO+wXiRQo8/JWnVhCRIXT7v8
wf5NIZgwwFUIN8gy6qmEikNLZQPCEQqol+d4Hj686a+Gf9GWDOVBFDC1J5grhDyM
EFRms4ePNoMRwlUUJlg57JAU22IaPYkJKWZdQJ1dcfPlR3nHq70EQSVy8wUI6Lj7
t7el+3N37omcxf2fhcsSwRxtDO/AhD+zVszuhhvpJm5eWz+5xWDyHjMqYJbfUw7m
DSddM23bWMwzSL7mI6Y3geQe4uk3SYmAN+Cxm9WS/F8+fO9McraU6do/2ItYt3TA
UYpWsilF1DPTsIjG6wBNFKtZ42gBgnR0Jd/6FmbT9+D6kabPDrWXqsGZ3oFhV69i
2I4wphp5EOH7bdPkCWcsg2MflDE/14ZryGXDf/Qw39VqiD0NsFNwNKIHjXGKIkNV
fjufXo6DObL96QqEZdVPlx8hQ31dA88PNVyJx7YRZr1WcRUQzgT+OW1IRfZSbTVx
Kkg5FC6jAdrGwdZf4uEsmGzztuOCwIM9Eg5MJShCV3tly3IRYz7jxqzirjZThoWa
bybgNAJ7AKgM1WglrorSLG6o7Aky4sGgLQHZ0AcjmWpZMQeawbUXUlS4HZKxd0rL
gUs06KuD4/+BUeG7SvfSCpr7+OKrNDuBaaMuahtWcbGaLdt4gvzfcYIHbEmlwBnV
IDBEyUm+1jxf8Wcy5Lyj2V+VDBIsUohyAesXYFh8LyXJumTAvI/WfuTPf6c0cTjr
4scHN/sEz1mV4jMxoU3ybc7eEcyqfWWAp+cMuJM+44DuK8uUtC5yYNVSy3oqdUlQ
ajGvit1BRq/32YUJ5S8KALW6zLZJDKWrgMI408WAfy8oI/lKdXBWIRfZAiN48mQF
ezS22wXxiWobp+FwAc1or71QpveWF4rUTPAB0HoUvVggnbJZMSHzS1JobjuiD8/i
G721zLxZhXuB0BW03sWitxS6YeF3eS2ruYZnaDWSwGP05mGkvXn4XZ0PRMrTfkFS
snQ6lRqtFEKFer6/lb+rYjbq6kfETDU0ZUrlx5DRl/SFNNpGwewo1RPHzahpCPZ+
JvnpREcXBEcI9AVLD1EqKST7R3tgVP5bQzmByoMiRvmuM1tUFPbd2veTGFV4jO/x
igTW4NxnkkMAyHs+3/o1g+G5DhZrtngevsRDT8Z9POYy0KPK99gT9uUYqtnHtDsl
/kkkfaNJg9LB4H6Y7nmaWPr0REqxCkeVmaLDXzVZXusqUJ53ii3u5IFEd5ZwS8cs
otEmgCXyquWI3HCL24mQ1a2MgGJdj+EUkzUmaCj2Ia47mNTnEExRpfutajux6Wxq
2EnsS6vBpWfEAfFThsF0ZT8i9NnrbxpMEfjUzBUxnqQUcmUf8yMMqeEGS/tYeP+p
gj5ei95ooRobfSKPD3Wxu8XIjdQIgdMLp/B+JGcIlvpdMVvkOYfvvvGhsJn4H2p+
pPhZnuwRAtFisHHmlS3yVgNxn+hfAulgiKMWgRVR/QrjYijjT5DNnQZ/e6xebry2
UDshK9xuYFUYXgVe0Q40czPtouAHuuWRQTj+0DqjzsYQpcw8aBcrDUhg5W7o0f0F
IvkwvkBNwUFKt7gStb4HPmWxHOmaVdmygwcAdfoC9UsEh39NfxScDSmf8InHJ840
mNwcU2XCBDWhagiX/JFSTUBkIQcQrUkDsXEGMIjvd+KbLB/5vKDzEYaDq4r9Ebtb
HlxHQcaTef3ORXpqlqhsjCezd8AwRXlOaV+0J5RCcuQyJelDmrycaj6n8nPNf3PW
5FE4rVnEzwOeXIMV/gx8pRjMMPCEz/k8vePrRswDnfXoCFJ/95YbrnUdguQdvfqv
RUmgsskRr+cXfvDhh8ohPTZB8xWPp7fdSUHca55Oidw+2cGAUs2F2U9fPVTGbRCm
5whKVJvZ03a4oCFoKO7H/VNdNv+INaDbxvPt2SBKdgB8VU2gprTreY9Pz4iNm6+L
ClLHRMtkjTS0Iajn49asZN1k8XVUL7RLD6IyfldgYmt+9K2VDjidZ717khB+Dlc/
JFyQ1twjrm0pgscQu1zb7FxmWZGhdDrKqgeJ6FHnQN/QrRKka2uVbH2UD0YaC3Ju
Fi/q7oHWdkjgPT2Im7VreABPixHNZDdQ8AwNwkalozwlRHXryx2KgN8NNz5yr5PN
uMYGCL03CBAhIpmfUkj1+GySnmMdkI2q0Z38QMSkyWbGFGPgqtwsN5F+JqmJaVHo
zQE78+XxTP0m4+f+AvmaOtyywePk3Wt6CrW4NPZsETkt+LSZkenBexJ4hZLsF4pJ
rHXW/DJYqg6u3vf3zoR4oiuu1zX335nUYIGJU54i+ulH8Mn/E8hI/OVoonspWJez
tzOw1PTVgq2oyKMzWEFY5Bn3CEPoBB4j5wbfRp0k2braOXKwKGfNxCja3569mchL
3kMqCdaDrsAECgGXg/JMfOAvgfZ0Tt8TPPJ6A/9JcVXpcYXfPUOYYCz1RQfF2SFo
lsWwS93nsx7Q1mfjuPZ7mLilcxjYhp3kXam9v4xwVU1cU8Cb3lNLHt7Iwb4cDaDu
62J4qD4yCEBXyY+B+mIpLGkE0jWBTIsxvXQ+46SbcWpc2JgSg8MtVDhpGw0I814d
ZUEl+e3kNy7Qy3II4wdfa8p0xRXgB6XEWdTz/va0GYs4d1ojbQ2K2xeZJUnR864R
Wewr/Sp53aurRpbiWarcXrdf2wE3BLlEPQAg7GqGxm1kLc7v4IGb5kffFTFGAIy2
wcNaZiFxXO5eLHdsMMwaTa76S+H6FuJHSHx9eAXjXI3aWyRnRex5uCDuE/roHOtP
3JQdK297v74JjkrIDjbafehqMFYXAntHIKnWacofgO6x4l3pyY2YPKGhnmK8xE1K
O4zrCLIuLZ+EUeIuDjH0dtSRsAGQha7RQkzrzT/ayUuSwHyEUjMxRkCP2znyIubi
Op2jA+G2Lo6aTeBOchBI6n26Fx7DuvKKNA5h7/vyZb+jv2HUH+pcT5tQLEVOdn5l
yYbBv+gBFJP0u2U4M9eDDQkaY3nT452Ki28dIWOzZJhpnY3O19uBM2293c5nus6b
c2/h076Ku1NiNZsmr6GhBREBbMLTTe8oTvIe52sviOnEkvD535fiW9U2Z3uBwWx0
CnQHDQtbFrM8lE3IR6u/P6rlIlao8nVWddsAlvOdtSTaXJypODhC202NgR9FLJ+J
lhBBo/R6jVPNP+zTCxOXGRtb04TTPzB+6xwGUNyqFC2kIKt76y3AcSgzkE+4Nnah
cH1on4DqRe8iTY1IwXP9yCnezcgJrQpywnNivcmdxrDkb6bDgBRLG2j/jN+xzlvn
W85v6wbGV1o4GqonGWMUnfPWLFNwh75t26QfWp61x/tUtrfEADQeOzX3c3KGI/fU
wHR4GJOayXMsr3IMJeWC3ZRSzbd3rXXC08Ds9ZkCujx1Q2YgJaPxSUQSp8uhFo2j
v3sy9aT7Gf1bzAdj90WOZ/zgzp7UymLxHTKHJzeyZl+UmX+eBvaVW/a5lzJokK9R
uyyJ4bhpwmiU1xHYW4AwqN6oLsMq3wj41HDzt45rZfGHaBIg/rgeCdK9Cmh/7TmV
cB+culwA8L50WNI9JGBYqzDQ6NX21jQDPG2MoIoX4cqHyxYsvcLNZ/0w3T1bD9m3
gevaiaa42Xw2Nx24/Xdz613NFUciA5dBJsftbeo3Z33F+weHeZ7edEIMwExtr75E
hvVbCaBm385mu3MwSkJCMw5mzeX9D7ji63SyZvI7dJpJ61Qdb4Yt3vHa8khihbs0
wZ62Ul7fwOUwsA0eS0Zhdpf79SuS0lCXsbJl43yB7IRy0goQ/AECjXI/eOYWkkLn
xo0KeKHOs3fpdCWFrnTs/noqT5aEsWSLmUAuybfaSpUAEQJxjlHJ6pKj9StumS5x
HwRXAmXzDwPgBdCbIWBCqOUDBXKMW8Qf1ZDu7M6IfwO3pAgasaqaalS0XZ8BOyjf
1IaYsuNONFBxnKv/0IlWftZSC+yNx4C+LaBy9k/wIS0LXmRmncKa10fnhX+fJ4A7
FTAbxM5uoRzSQjcfha1yTxvDOabqbWCNekYnttCeb/TfSpI07NTFpS12uV1tUJrx
qT6/1oyTOFbEdzDgkDFMG4cuajwkM22HxoP6V/M5WMVByx7+lvE3vdjBhBMxyOR6
aHghN8G+jF9F++zWhUwmp9BhB9kiVZ74fjosYIUmpe8yrAi9HFC6a3GQTKHx4+f1
WAAKV8CDVYXJmAvjhy9uWChVn/qgcZEiGrRzT7CxtePPny2cSV8KhEHZcYBHtkKP
VZ49DX1y7lu/Fpa/uUouUkfeCwQWQ23K3qZFT8qe689ReFAKnon7L7y2N45zKFMs
OfV/A59Bzx7n88/mLZBDJhh9//SuaQoBjsexzDa5jGXMphFPfGMwLBB+tJoBg2/9
RcTL94h9mLhcxRGyBg+7ukk4BXClJpzZ/7E7fN/uPzB0AGeOU+4BAL8E6woFI7FX
+zzrvyDXzfiP0buCDqho1NFEXNLIDlYXKOjiSJkIFrtAi/dTG1OpInNQ3Qj6O11l
MRJJ59m6Cuna5155vDYCuVx15533wycl43vHD5vVc9Z2qqWl8IrjnjFIeMP7nL1B
KGSa/eZo12cspsRN+ml564oe/LwGPUMTj80hW+xN4NC9r/1a3z+35jPLJWikq67x
XgwuxjGiRXTrumpdgyHjc1t5euUMqTougLwgUkIEg4ynGFUUCkYr+1P3LrK8TRJd
UGFRI83/QfYN0nfvHXXr0uzjAcqgqNGlyaCsm1NPau6Ineo0xFkwHQCQhEcnCjr7
caYhUrU0k4LsAduQEuaS+dBUSSAnd/t/Bo4v7BwU2iSFkd1Uv817VDpssVs4G3ET
kGsH8ewprh9o9xXwn4R4FH5Y9h7vxPFlC7mc8+qu8qXZE77z5HOT2EzhdFE5DCP9
isRF8gz6kjpYTyt87bHt2Vs7pA+uihtUkq0/DJ61xDMt4lIAO31xTNMuiWLpsMEp
Cq0mayKpnq4afQA052RaD1lVlncWr1TO0spXLc/exji3ksSUaluR8gzFQPxsS+ba
qyzfYddpGgkp0UFrR0T+LD5yN52Ghz1jkJxzCOlu6ecBVjQ04BqVdPgOibXkHgGo
i+1j9T3WlbIAPq+9URtifm2U4TlHP0Lz5EETAEqt8RK8Mf0irBKnd2EG9BMODhDI
pvrBq1jQoyNFx0Ue/Qm2SaJmjOP2Nez4pFM4UrYkeQADdvR9CtAqsNXJM7RgQ8qB
n46NGnrloaQb5zwPBWyA0zFpq1pVsrxZqP9W3mVzbME+ZNSW21kuhPapt0Nf67ly
OS/AnxVdQ47ArlJuGCYS1d9dHrMg0gu6Vzq1UY02Qu0AJWaD0/TSLfGoLGStPO+h
JSc5z1fdwlo90HsP6fowbhhsjpIYsgjfae8w+YoPhgEZSTEJ8qz5EmUwN9w+AARW
niBbO7kLAP981mFDn8NNbC2HyChxWtkTmFJcf/NnwQKfew/aNowKqspeCuKyha6w
Qhe+PdTFbF5+Tyck1DFWw0ARQcA38IqlxTwFqkdjAZ9X7X465WUcKPhznmYQ16K/
psgrHcn0MOUJFfSX6z0DfljFNos3BjtvhzUasYk9Dzbn+3XYZaJ0c5EUmNsibEde
pt6YPk3McT4b3quSm6xBsCWGzTpI4Vf2kjdezV24CHffMsPVXpilsTEa5PcDhL/S
b645ueKuaWmOuW2X5PWRlOz6ibJja9jWmlC6/SgWeBuAZG62jsZMUICJVwDoD9Me
SjKvZwkkXqhX/6unrxqMRCu6n/qCG0MTcuDwPzyLM63Sb4d7YBb6jV+GSeOlofYK
O+bs3uzXJK5xCSgr+VLXq7LtcKgE6Ts07fFy+681itHzwN2+PJXcOiF5tSumSMbR
V0newoJbHDAgjuv/5IvEu9YAJoGMPGW0b3/0snDw7605ZdltCZM5TNcggglyjp2H
u4MQu+QTzWK0kvx3LatVnsPATbtEDWfovW8M21ZJQZVvoy2X97574yI4kyfBexyv
d48gK6Vw6+AjK81IQLRCnyrxb2Ttmo5njieQ88MBm2828C47dkwqAO/rrwI6FMCv
KC6FwUhZ//AHW9CSV3QSAhViG+GTCyz1biE4AWGv19H0oEoGIBkHPg1rwzqUP1tN
UBmNjbNQ7kQNbTXoDtMO23YNczIMKZAgiqBRhTT8g2lStfxZo6McXaOkJW8iJlAH
PKGbD53bZBFGQwESW61FaCs3xJJGbtXAfqDTdr3oMHTPbuW+mGi3nYtmvEI08hih
3O31YnJ2hM1UGWdwpTlDudFK7+osFsnAw/MiLKhh50/g2hUuAshUUxgKy9IhuArV
UN/z8ZwzJCzJFqbA2h8M9u5/Nj+lyOQfw8bmVPQm65ULzltpy2epm4f0LL9f8CmM
p+ztxtGCpUYgnhJJFzduIzgRNlwo5sLQfldiiyWRbzBuRPFbVjvrlvWbEfVLJh8p
/cpkPxb/Xv//1kxHYu8zQvx+WSD1T41rJrdbdBphWWUL7nAJT4c7ij/z8UM6TJH7
vAA1POLu5fNkz/e5NtqEAjP91oBPnW3y8Sd3q/TNUG/Q8/YCzMLkql4o8z4CTUPW
9zcn8c0pk6JntJ2PrMPpQxi78+gi7Hi3CNoXiEAj2Inf02cI0sOLy8o6V+FFpNLf
+WfLg8ne2a43Y1lyR/sj4VK/nLnxfyBCRulKbjB1LjnoHZjiA8GG8UUwpzC783vS
3IKH9Q+1GnB/p09A4TBDt8rDmTe3seLlc6XSliUQHdxJYXk6oi6Cg4q4f0DrHP8X
RznXk77bMtpFT6cZjl22bXDE9Rz2Ncn+xvexJUeHKpWR161cr/PbkU3AVhboRcG4
+xZsqXn8zI4yJ4aIRIM7h8CCZFzVG9Hy6ivIt24F4mqUiWknjyKcuoKFrB5T+KU4
zJdLQiGoeZwxbx9T1i1ZDdNHWyygBh51lBLFRZ2isnGsqNXrT7mKf/6nM3FY1hjk
aaRN5bXwL0630v+l8wIq13LHsGPJpvqFMG1bNpOCqEjHM6gCFoXpxt1FZPdeNzW0
0AriRy+kQ/HUrYYYl1JfcHCYDqP0Z4Ho54mBZD9Gj5ILZnF4VRrRzgv5bsY6wEME
5KMnATO3vhujWWzAkeTyKQ82HdNUarE61W2adI2xBR8hTIcvRzn1mwILv7S3vef+
IWqAB/DA+aI0mIGWZfEEFImHPYb41UTyYVtLklgMPb43zo5590AHiloS8iSKX+cS
VmMsVs0+wOag2IBMIa2hmSj3GBvZ+wZ7kd5OOik5tciqVk/lPAhZ0U+aaWDTKN17
ls2Gi3x/3ZuBzF6lOMUG3LH4hcH5Q0I1n4GGJRpWADH0naHmoLymMaypzl5x32ZZ
sbCrHxKNt3JdDZv0J2tL7FpqdKSxDODUOsqsJ2Uc4Chrei6UaZltivB6HNf2ugOh
nLdooQvz8DTVnraenpppuGms8CRalyBfDcnCibEujdYI/pXqrEgH2OeUK9INYjlf
BMRbPjTV84FW130zyijYrHM/EppNcE50E9eHzyo7qK6r7BEh4Aq7K7N2gxRfn1lN
d6jupiUsHE4mYvAtiF9/CBrebQ2ZpBgajcYi7544WdI2iAFJSSBe1+4t2spjcsOe
FN2STkjo8nhx9OVk4vHUKszaLw/WlUJqOT67lb9xXl91VchhTCCKRZbE8stCI/13
qha8/0Mt57FZi7VwOy7Gk6yimCuYFpfzFEdgXoqppbgqiYB3/5s7YYeqz4BFZJUY
otAqSHqIM9H6VoQfENO+Ccy8cpMHbxxTiOYLVjIofoL1fj722hclId8kkdOTCVSM
MCrwl8OKPeRSVh2hlmD6AGXDhgJ0BADbcSXHFuM/E4AIDgT2XmLqdTpnZ14q/YSU
9+MBz6XgbLh55Sj9TF3gtkjVwR4J20ss/OTTrMdUp8279oZaZjmG53fPlvFDzrpx
SODlSGv0D+Hr29tA5wkSXwTvnYDxpYVdes8Sskd3XEhaZb+LHNY+Q1V0vv6GyOjk
dY9e5wr6nSjIbStZhtSOu52UnEa3bBJjfccwWyjsRbpuJgP+LW81oDwEM7yFkowg
mx/59a25ybxPeEeM68y+IKKTvBgMSZ+bun4qra9FTReulM3Egre2E6LsbLGERJOq
CkS2B/pK1+vqk6Ct8f4+zuax7gYrVp2de1wXBSo8MIySjnyAE7pCu0Ke7FikdWnS
IdaBtjdvT+VtvvaAKnXd7pAckmK8mRKFt/J6teO05gKKH5+KJ5MW0+cxdl5iHFHg
pJ1L0cqTQ6CA2ip+00XouWNvMUxKZJEOI4Cjb27Q0dhETxeOtlkV+ZiyeX2WdhEl
H2U7E/xiL1UeZXYoqPbopGuo04400bOvlatWHIVScqYtJ5h0UBo+92T4m9t0Dpiz
QHCLk2S+rPD9L6GC+pLoF91vSebijuw3i3rGtEOEGtsu8aPCfjdoUyUbfN2VAKHV
Xn227l1QiqX0QkUWow2uxfuwbfJ1ilf612z8PVu0B5nZIysgOR0XGdhs8UHoffb8
K1y3L+2NYn7EoYgximsuMW3oLPIOenM2Xn2c297zHn61KNt2p32YJCouM9XGf1Le
IHlOrjyE0vbkLNwR81VKlZIAhd8Vq0ebyocin0f1kYMcGkiiP7tJKfsR7KfNvMti
7kmc326vVNrSNb1OCFcKWA==
`protect end_protected
