-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "N-2017.12-SP2-4 -- Oct 23, 2018"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
qOXTS38VTZISYT1NXuVZnJ6s0NuEQTC13tdoo1B/VGFYS36Z5nRWzFk1ys7pW7mc
qIXhaHWH+CxAUqVgG6t7Gyw11Cf+T51FdH/3KImOLvXWAkhyazANyUacVYVqdqpK
hDmR7veTfDro2KczfNdXYWNwvg6pO1PlMYkvr7vdghg=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 1040)
`protect data_block
MWh2Jhfrjz2Wb7QfavRgLmSY2vsj7S5TKcqlNMCvSxCepNRQORA30PieXz6kYqW1
DvinVfYybn3gXslm3ctGgPVwXZnZORipnMJJycx15lD1EWSja98mWySTf09N7tYf
/peYD0H7hUsG8RFqVIONpfx+vXlL2JbaguYqKRjiniV1pdvywGVoZZHrUs3a4yya
of7Ic7G/C8oqH2BtHJY4C3+D7dONrvOQ2ESGZZGaURBgtKHrwJKyP0dj6y3mGZ+F
hfju5NAIoJIiSbkQpYeTp64aXBBAEW9rF7V8cgIIkJAXEldUJBGTKVYflY+Cxb8I
fLoT6FAzRRedXaLxW1kcejWv/XQyqT7ML7bkuNfyM2yn597Qfhtwox4lchA4ahBU
Zoec0+GAfGUthDH9Gawpe+gFpuNRnBn14+a3E0FeojPdygCF3u2qXA4czTMaV8wS
XNTmoWZJjBRYKc/HAxqz7RxyBlnDgIhdJb5CHvCrki9pDwazguG+8EQX9Z49PDaj
i/A5ssqchoWAAf9Z3eDO4YXNsyfpvQoysab2JJX9wxKeUmPLGhWAqiwzDhsNBqjj
z7TqhgKtbmVcm8xw16f+dKbJsls7ttZRIia539uqlJ5QmwNdCzo+neawNOqcHOUQ
E+8As5K7yR0NrApqLIFGKpY0WnO8OuCjJwTprQ/eQXRPblsq/6Kl0lwf9DAvw5Sq
U3dwNvpnr3sIrsRFnqkONKVVI+HJ1eKKo7yh+ATm6HjVf42E2OOB0wqxmLglskA3
k/Iw8GHao/OzsR7prfnS2JW+KF6RGQFtJRqlsM2J1pISnMZzzQMkDAOPv3arem3k
QVIj5CaBohpjzhn5izWlmLczaSyDYzd1rKHiea5sKfpN2yO6IZPBHzMaBDS99c3Z
5geX3XxlopF2dwNaJoNIjN28ohqMiR6YXNFReaktD+dRhVdgoZC6VGAcsp07ifQ4
91Ec7GShQE6Q/vu0ljJtiRA+9Sy/LqOr/HVR7/SueYkN0PDHaHDIJ27Cnqc9GuM1
kFzdKSfljo++s06pluP3mNX6hQkcR2BgSxZFkIuVzYSnDFmuefq3qRnfzoPziQ7e
QHPXvpqf/Gv7UklNRnh+UWq7npQtL1kwa4IudFrndKlsdItC1Qi7fhKOc+waL8Zv
zl0Sk2czqpjXb5urFzF6CD4yTFiSNRgldXut7wKuzhNUqS/h1lWgrFLK89gYhHhS
GNAJ/hZMcP+c1T5RyFpv2mwLwznJlXXTg8pFggSfLiG6vxsbuB00U2Dt/BsmVSui
W6c/zmch81jzOSIYlkCm91uhthAIC6Qxfdc1oDoSVWEs+aU4tmbDJBJQ22VNANQ9
NLjtWJ7e/i1nwDyMHGUsBOUTYIicC1Ecs70WtigIcAE=
`protect end_protected
