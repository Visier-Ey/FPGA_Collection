-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
--pragma protect begin_protected
--pragma protect encrypt_agent="NCPROTECT"
--pragma protect encrypt_agent_info="Encrypted using API"
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
--pragma protect key_method=RSA
--pragma protect key_block
bd5hghpPVnJmmEYYexQjd2GpCQojYqpbcJMC7paSYl4U9dzm+cUKxVlW7ZRA7SgN
bBziW2WKyGzpuYMnLZeWX7NQVBkgPw7kKWHa9o6GYnPckwnNHfogLOPGnQHVlU95
XKLYbfmwaoLqlS9tb03P4evHctjnYSxFIjPBgYjnNz5VwKcl8fwV4VToqfMit79t
o4wML453AFWdIm+kLPDweSnvQZGeHEI+WnvLapICNGDIoZE98ND5TFqr4xslNWfF
Qv2Ji3WY5c+PQ1bhRV16RS5mTuUQNtkA26w56JPSIdA5CELI231lgorYsc8dN4iD
sg0cTBK7a4aAV0KCbu8c3A==
--pragma protect end_key_block
--pragma protect digest_block
ecZYrNM1O/yl+8AstMEUhx/5HL4=
--pragma protect end_digest_block
--pragma protect data_block
xtYstqFNRh1kPEIwQuA9tL3fa9mVjXjbkyUvf5DfLczGdstGhz8ceKoDoDJupjtz
oJNMkf/86Hna6M9vzzS5DCiUGwYQ+in5aVT5eTTHNUi22rf8gFAnokI5kn/LVQLU
g2W0+7EWPCicdR0kQnTUl3b9b42oP8biARaknE/U7d41BDOY9lo2n0fl8wOL2KbU
/MSLdi8KSlk9brAkuWB1q5ZuLNc29p125+KyG4AfFzHGd9fJhTIKcl2ftz9bkIuh
37s8N5+WmMKEVOFQvhqA+a/jYtIWf39ukQ2RvAza+qV4FMMIC+aSthQBv3g9sgHI
16dLNZAm7eYwTAbFcvgoLFk4oQ/YSvyJaSJtD0/uJymHKS7XmSVqmtqA4HiUhzMf
q2Mjwwhj72ziSLVopHVHtmMzHL0SsnJM2/2UoecDsMwJT4Dii3MxB8+RMl19OV6M
n5rvoz2WjU1XX5oAPbtNtEs+aKksx6YzEJ7ZDuW7tDpJKqfpk4IVYtOpKs5mw9mW
RR6W1l1J/dd4kGL4JyFPf4FUHxL/+yse2bwL0reQd04lYe6xr1VktuKwuiKb/89j
9InjN0fB8Kl1mS9GNdk0DY/4vdeW0DpgavdwgSqKDrdY5jWro2XbUuhSzeaSfL0q
YjlyDe2gnnOswQhPiuBzTKF4ARTuuoy5Nmpwb8jmbkMr/HIUtvduZq9pLJvFWiG4
B6rqFUhQQ3nlhDNvaug/Vi1daTOi4tIVqkDQsuwhLapMOYHaGlDfQOnj/02Wn1Jk
9iZiyFW7mZ+4JOWSgwEnfr88btrBFluV5iQxruSBC6BhcjCHuk40qkWANG9s690E
BXOCDnxHGGWx+xKCu3KBfQ1+Udjjr9ZrePAawb6IP5saH/uSmmHNrLTbg1JPtu/A
gK+dpaLb4Rs+6Q0Ryll7i3jDWUI8qrwpZV9+4De5rfZ0iQog2O+TdCejj3g1Pb4E
TW19iL7XsKr6FxTNu5lxDDbpiP0RqThjeB5/fYumBKnxCbvzEdTbeYBzp9taoMdW
s1hPvKD5ZGftoxsoY3FjkO00QXmCyDmkZetB2cqPKi7VcR2DVP2nWMBy8cwzEJd8
V7tiQObTIiPoMEDgROM2w4G01VQoO58HyYmXwatM9R0pQ6B5Q9zp7dfH28pUcFM3
qNmEkGKQRnu0jOzxceJIorR+AY9THEy9anPkU8nNQr3HxXmdJW0eOIEDv4rH1qW7
pnn2PKfojDPYA4R0lXciG+12M0xSoTWMOwwHOLehSp95aAm/GR6g38Z6sg5z8N+0
VfJXBusLv5FfCzayxD7k7hg3pPhxGu+tg82WhCRGNRHY/aIDuccFc8L5cb+4UuFm
dFpSQtneu5C4Uz4LgpdHiqnlfplxPavPZiiBK5QSZdvCU1siLKDaGOJZ7fv1K+zi
0NWsmfDT8rfximMDup1kQOqTAhIjtJU8U3RnqtGL7t/ZqFaFKyxPuXIGuoqh0bno
vTmGqZmdLuOZqbSnTIe+jkgH/oZAXU8ni48hIDPNJ0v6MG75DQ5kNcZl2mkMxhSy
F73mNR++Ya/LTM+W8/1RHy97cfL3xKazLfRXistCK845cS1WNGOiQxjco76/9VKk
kxItCacLZ+i4d/U6eHoFyb0cixCdVxdD3kA5y7MCYK7JV9B2qLNoE47nfoA5AJ8K
+33XdtH1qLefpokiOVxGU9jN0jUmuyQMRzZyN8XJB6uZNiX3OZtSWA8NONePZzWD
nd90p7k5mPyKiiyo2sMHTQy8KYq8FSBuBvjh3dkVtMFAuOGX8ha5yGlagla7Y2qF
iv+fKloMxmi6Bb2SN8dhzD54j1p2YXYHWNfi+sEK7ClZHW1lkwy6HFNemspBI+P4
qNp2D9bLBlw4IJNjf/wECPktY9fEXCYXwtdCLqrIyLOU4qUBpn3DZl62QZISbcBr
8gE8HluRal2aAGHAZIFVT1OHNXG3r4YcXSG6NGXYE4cRkBJrFB2AKeLrtDGXj3tT
E5SGj393be225bpxMsM3MU/MMDlFANJUra7xbSue7PZjlylnnhCngd86ZlXW3ieR
hwnXxfGsnRU9ve0ILm2inkbnCygKg+ujpq8DY28loNl7r/9l+lECIEH8H7IzTwJs
Gb+Ss7F/aSS/8ao6U6BzCruOofLQrkSQDQJN+vKWZkwpqnEYymw7OBaS/MPgnhWv
+1CMbmkMzBowoG7gJNtS23KhF52nVr/7LgJVnWhq7xbzPoun7+rTQZZ8LZDSbP/8
cgin0RnNNXQWvYSoM6rEpt1AMKvYDchTNdzQFj6nVFDPuADOnJCRKJA21jZKJTgD
hHM1TtLBqnGOw1whJ+Kw9GzZkcNA/nY3y5EVb5cOSMe/V7KDf9iMFmwE9Yk1bNjW
qRa2v+W8kCFgPV0BkDvLZxStiyAhd8bvQ0Qe+hWSLSlGKvtNoSTb6xwQAVQpPYHE
0/FkkG+zt1nfQ82iCPT03atBr8/gMA8OThIth1r6X/Jw6ZcFS0LvmTqnBwJumIsx
KGmgQZ5hYiqOeSV2a+mVl7wJGgXmwug4ALTAMEJD95RK7+GUFDpFqcvFxkpKJgKg
LlVAUz43BPcf1s7sXODoG2uEYDkY/NEZ00iCXdXJZF+wNiaUtgrQ0JjJM1WhbLSy
JaVnYYBIMKr3XNu0s1uMpYiAbf9pSnM9ifFxE3CxGN0Qmp31lhTKHPOLtwG7aXdt
vU3yoEPfNNe7PyC+59XxTiFRMty22P1+xRN1BcaYN5YkBGUrU6tXQsis4NPPi1j8
AIxpTYlZo3R7UnkY+9bN6OfqomzllbJHaXm695+iF5s/FdnisRRXemnS0vCt0pdb
jKQM0IPnPxurTs2BCam+GDSZ84TCUhu02sRAbl1y7ZSu36zdPUvzgFzzl95Rhd2j
EOH3DVRZ8kalejB4MwGKI++826bj1WzB3NN8Avf0gJXsrZEYMvd6E48yoGT61ypg
343o6d1W4UEF8yFrZVZpD0aahYbbcOiZPaeVZgRks4cAWHRGYNalgnqAIuQr4hRZ
78fRQEqV9JtPnpq1rKz4s5xU7eSFvCqCA2ze7u2V3S2ttidSFyTRRq7WrSqe9d5+
6WwMnN9H6OVFhRcs6ujbncObze4LpR+ipvYgGNWVayLITny+JS5J3EXwJy0Oxg41
l5YUSouSeSK51494oc3PkpAhnTYnKWPCPimBDy0km8MMP4taQjmJN3SSe4CNsJUK
LYGN6/spHKaBTLPYOe9fnhoeBHC+J7j8oaJptYxm/T33+TITHAZNEVHPTLbjcv0M
fh9n45xgcwYFEPLRr0+F87h5xw2gEbMGhhA8Qu1JYuSn9o4ZnoW+fHOU17D/gb2U
NAAN/aw1VoPRgogFyUMkcq+cB34mPUuDVjRKasMKiUkUkhdPalnLNW2hd4gKTXPm
am8dU/iCNR39481rk+awjFIRX982wURpOIn+K5fn63vYPP0vpOXZ9EzKZ+rKG5zT
IotMsGd8s1k9RJ3yxmevnm8lVj/T4C/DfCivkrlRY11oQs0Hqkh/uriox7MrvVIm
tm8aO4ZwuhknCUp6vRqMeKN/H1B/hmofFTss5QABUUQ70nocHVJDicW5jIyYnJmX
z9fhdzk6HoHjnXgRBjUMAqw9GedFoC9e84WyJlGsiwnWFbUB+GTkR0UrLgw3qJo2
/b6JaPnMa1gltChm9FLm189KWeO685RQh7QMWNsBktgSVIYGMwF578QvYH8bVXTh
pS0YWYu215UOZFgIOa3+kPYraQonzvivGwonpNwEja5rLhTdD9I2cAUPejdDr/uR
YBuz4nfp4MIxGxXryM9tWpCVx73VmMLwK/iw1PK5rTINpJC5HjBJAkzEiaUHYpDm
uX7t21WNksHoeehxMcrEUjYZpgClaFLgTTJ1OcICczS2rmtMKPKgcujFUhMDTQUQ
BOudcW83PXsAArL2dgztDswSExXHdqG54KBJNvzGxoJ60WaifiPgDtCqsKe8I+Bc
jEndQshIlv4oCcZ+lwrnXbi3f4/wc/1/Yp2y983h6t11O1xy7GwNNHXtgBYlD5mf
jvBearYL3/ojjTcLg8wNnq7J0l+DZjMulKYcT12L9h+sLaNmQTUpuo+VcS9AsY4W
pkWj0gipQiILA/Y76ooiNrZMjO16K4Q6qj/iSfKVsWSG8Qa0OAkeczcX2Qnb2B7u
FZSYnBWEiLknz8rNkvBNps6xIuQvS9Ff5AGeM8uJerxHo0ir7ekTVcZk1N+iOuOZ
AqXyO2hjE06VkDH1Ou45UuD5z0UNjWjV/Q+j7+oFDT4KgRb3pxj9JV9KxJUdIkZx
/EQLbIQmGS/SY97NPsML3NBbOwwxTJHB1XzTUOBPB5hIOO+qiHu6ddE6QXkHHyX4
uuSDfmWDP8QtuIeIePWUxgy9zKSQNP8Zm0JR8DMR03hJQUiAwpoti+h5WTvMkPMK
Z4AbEHkUpKtG29CCZvuBHUMfx8tYdPwjr2hjM6TaO+jRTCrzOEI0zLGFnJEdrcke
gUYOIAz2UZHWlqBDnN72tRmfEs0KN4xaLGcLoHKAthsbg95yP6aWnhM+2NTdSXu9
o4HCba5p7zwSoW6clAXkxKuo2CWII3C/jEqpTLRpIZku0PzXjRhtp3wArNtm571k
aVc7f+h4uWZ3mZi4qRWDJiwt/sRfU+zGDER1ZbLxMv3njPqPbxM+qSoKj8OnykBV
mGpyMU3iFEEwYASZEyaQjeDi+ACRxdJB3qk3XayVJlrwgEbII7EspNfvfB8GwmJw
dfBqVDWoOHa7QgIUOm2swTtUz6TU+nRx0nC1HL1UTlkPTRiyAvN+zwX02tVoIk+h
VHQzypRmvngItEmLcuzvB10ksaOMsh4U1RL8sapIF/FVuqGPyjWRI14MIobei3Hs
Fi/LUaSyZnywofMZ6KrsJFmSIINv40acNNqUPDeY87na4NICVPQKWZlY6EamF6Wk
O4Tjd9GsC8hc/ELV2Sm8olPJaubfaQ6FmCOtGc/nYyxLG7YAQglVqhFp73BpTbcZ
Q5xXD+65V2x+IvVKCL+WwkVEbJFp48/X8VmFmsz2JQ62+0dU7g3LrhQxpc6loQMA
jE7DGsBCUrbi2PPwXKS3puE7OZS4ukZr9b+YZwyKYie6I9/YIwxpvO2dealOb1U2
XUGa7CPXJpRSnTze0QE1zgeTG+HK11TrS2dP7IBNZQzELGS3uPsQy0aLuuY/yspm
e18lQplwwQsIz8bpnCd61osgOY0MGvkDH7J0ss7X+eWdkwUy5nye9JcU95NE+Lf7
eTaF+r6kBZoDIb8METnocSmPwWc0/J+qsVDwdH8p52wUqMNYkztmmQYXTPxyHX5P
SwGgbqrFq5JtmAw5wYbJ5tBaQXPpK294v7XsjE3tPnr7SYxSToByvZjKLUIcHrPW
RcgoCuxZr/lWuV9yEHIw7Y64NdYz7jLwrh7sPplbaQpeqlmaLEdZSnJc8TPNzwmq
IcCXJxrU+lOYHAadc3udX/I1ptHmAhvg4Q6WNXht5LuEDS9+qPNIqgGGfls6m3Qx
mhDn6RAKHkNlxuKWCsrhDpU+PvecuBJyzAKNMgAzwJCW7a+egB5dpgjoJA9/6JK7
KdhLgjN+x438GAY/q+E3/9FJ3wBq04FzyKZrbVWNJUWLIX/QgQZ5g3XBwYYjRdNc
KkVBRqaI35avhQN29fU1ssWgTdqb7b/ZtD2Ti+TpOWp7ysXlW4YR8+gYYSmuefQA
vVD6OA1Xk53PyEkzGzjZfxEoRpAi5ANFy2j0ihVvS8lHSu5tsARpd4xAVKnZCV4P
oCQ9u8NxqzedGhIKwh2Pqh+h2+J1n4Kb8PlLL9JXn1a/hmchJlSoRSD+Q8XNqno4
Q6oIAbqSzdyQ2+r7gZlBIBc+WojUvMhRqivtRVrKh4UUWLLr7abIUavJZ7OcyB0U
zJrh9F+Xf8ItLm9tqhNYaat/W5/PbxMhsaEWhUJGc0xodPWgVTAYVs7QDnQ7KESX
n3Gkf6PSAFp1/hCQXo3mP8rWrhoicSFlB1v2LKrZQJ39ytQn9UnIqOmtxrAc1+j5
Fe7nk3QFkCYFpdUgjaOi259vUpnmt6dzw1aTOiuOrse9j6KXNKMqfj6Hcc+MrMRf
7VlVJJpwwYoRYo2MnD5kbcBvHJVIzpS2cWGKs1QFq8EOk3EJ7VB9wGBFIzE1jUvy
Gy3mcpFG3w5dGlTMJCgwi2O04eYPiJ//zGyNDqc2iS35BrfuSylfGy5JHdHX3Bov
TGngAvPciRw599QThhgFjX/NTHN9YyH2pVmAA8dHuuaNgVEwPsKfG8gMZJsGUzjH
cPW5MUWfeI83O9ncfRDV6iqPgYmEoC4HLGZJByrpI7l+I85mgPPCOBuvV2Wh9agU
vIkr3FpdRzx39NoYJTxh08ebjfEXJxcCFr6n7nFZj1yp6QDVSlfO1Ec27yQVTQyZ
paerjGTOZZFMHYREMMG69yjQn9rC9EHCO8yQPU8YEH4r4fITg5pDTPX5aru+8WxF
uT4EG0O0OCsVNKiDH7/Z6sWX4UCUvemN1QVtEMwKnMPztFtbzlH9aMmmE8jv0om7
gR5IT7mkbvw9YfjD3FJ5x9+KXphUGk+Hl5kpYHSX5Fq8qizfFpuX3LA7y8dtbdU4
YD43Lj/cJUnBoHnnQAGVpxfhPi261vsv+W/bv2MCuAn+fJvZw5FRwxNPG1lww1nt
wnoFgqiOTyih8spJiVYrCF3pvxuqAV5aDGzt+r9zhTBcDLVQRkaZ9MKDoVDzQU4y
Wy1pOMt3/bX7I/UTGRGoXe0xxY+MuTgWETbJr29cmcus3MoQNgNIG8xH2BRI7OxU
TafFm2dzdHsrBQZXhd0F8TRcl6cLW7tkR75Av37RAZbjHfbXuG7CsFmgE3Zj48PA
7A9JQ9Qpdul98xohg+on6yq6XfFDCpCouJQwIiCdL+UguTeom3jgtQdcsY9TD/vI
hUfRyxof4hnCnI0Qk6p1CB/PyNQHcLjF2DoX6S5eCHsDGX+D8N8zoCVPY8KcJyAW
zvNnCpGEN2hw1OEzK9YPzQkpzRimBz3xlMY0clryHoyGHJeaIDvmCV2bG8zAod/+
SOwoPTv3LvVQXlfTN3XoPm1VSxktFnWgbKb06BJ/OMvWjmOXGwDFNYXiKPyMK/yB
LHs8YCtSwTE96svOAujcQBab+4/hNg+Mstw5tLVq2JI628Gy1ZnB7vmg7lFtR+Jo
uZcnTQ5qmnrh4tbCS2YgMjhdQX0wDQLSZwJeGLzeFVBT4/xxXdQz5/8m3R21+XR4
rNIhtkEQMU8A05+Aa4xuV4z3/9EKTmQ/0plTX5CIuWL5nSa3Ig6E5VJ4tHEDPDBv
HypYMp5JaNW8yvEFANC1r81jxOlGwo9cfQAmtdjYB34qBWfNOkJeSq+3yrTmnMyA
tnMP1hzf8LxUmW0VSOhUpLOurLwRPvr2UzXebkJdx9H6f41zO1Ox/0dmQrEBQ0jr
1zTQvjiq7x4T/tFH7wTCJJGaqXYYSFkCYAIZQjm/GYRqkxTZdrfIwPrJ6iV/VcER
Tc8f20Hvnw5cA4GkJUKNuRuHDm/V8hGPjHrzM2BIr7uHB0Om7pGJosj5kLrkZWki
FsmDbMxhth/5sw5l74Zmnx2L6f49f0MPHDPTRhyrzBYucCtjO/m7d3HIOMoltEdA
brpEqK49Amu06lmmAJi15pdyHzdbQ5EoSq71sPB2B2LfRyCvXCIYJPxYYkjTLXIa
Mewy5gWSi5gEFoPERg2jIt3nat/2WqfSA7cMiyIAXSUtT0JkujPRuaa3Nw6rXMay
FUyeQ6BMMOPMGsRPmr+23+KFn5foNLGh281SkE3UJstTW61B3mtgq12Oobhzbl/v
KNrNWpmA+ByVZxuolZ/k7TQ4EMoDQzjNRMU27VnFiIwQgfbqm9ACPvod3WL3E1HR
Vwzf8PNuIgViRglCzX5v3QUcFbOLixBIkmIKnXAIe1EhSlFMVa59ZNKz1WQQaLd2
Is4srlQwKsrcnbW9lKHl2Vj/Kc1KbXRLCKCrWMwUxOr+VWslK44h3eYMTLVYt1u/
83MIUYVE87ukSKeyx5Fms7LwbrL7xfocWhJ2IRX13xfkFtBF3Xq8hqhXb57Ev2ci
HPTYqKF9hmDyVMy76QwaL7AJgzf5xyFOUvyWIU/BLDyjtXYN3d0vsEdrQuUdtHXF
sOV3wULp8A6+9V9tv77MWuLW412m7CxZ7tAoFGlJ36G8i/EFUVrLna6cOre/MgUE
i/OQ3+hOuZ/0pDeyMVlIakQm9o+0WYOoA1R1QqURifjubyyir+9bNZVABVDSl41W
ozjgMpiK+nO0hxXW0d1OcI8WX7x1jAK/WJLydQZPzBLKp6QJMZTwMJKuiMpD78Tg
Vn1pTRBVGXNkHi0dCpPHb9bjUUhWT4Wm+JG0llDImondzuC+2HYpKKn4rEUqASpV
1NXPLPZB73RtXpAiEY+9r35NltBYgCfd7nND+4bpBZbGoKLsAXsaXpIucEUqJ7GW
R2SbHku4J+ov7Eq0jXSuPWQEHnf7vfWPLcD2mgxBCfnPheI+Njn4afDceSqT9s9L
itiC0jLZkhnoyPtKBjJ4m7IUDow7VZY6SEllmHaaHZNLuoEllGCpy3sflopfelXS
wjGvJgmZlp1X1UtptSdp9Vxsizqh/dE8VNGL7AA3ZY54BfT5cJxq6+sL846P/QNA
jys8nCE+Mq6RAkerk7IPI+0rklKDQ44Zz8TBg00KbzQkfvGcAwUWlqn1jvVqlpxV
d4pOZ/gAdLZMopRtgJ++PbLStpfo7luykg5dCmfrFB0/6NU7YbnPHJQxWdLBtNUD
RgbKuymsmARzjORFWX+Wys7sBr9GTtcYxna/T2ot6+Klv7678JxEaHsnX6ij1G1/
plGKjOaWFb5UFTpLrlx8w8vx7eT7mOQMPTVgtJt4qOOhWcuhkmeoVSvmY9ueDVZB
0SHC/Biypr0Hthu4rkojbtI3/Nneos/LhypuRzdrXCvWF8SBXwHkoV+MszrJF6e9
ecefK+l1K2f2a3/g734s8Of9KyMOH4UVoegI0M6nIsfvicoAdVG+q4k0zTYHmBop
xFGkxvy3nvPCp8/nyk1+NeNX2NOhAxB9OeMFNGfaZA6BhNUKs8rgTMVGg+9k4BVB
vdZ/SKJDhJ8ysYeqmnRIUFnD4ded1pdB8VcqGfgYw9IivC8XKOWPqFnZ+ntP6gi5
TZmAzk90xXP2sjXUR6OXtUILWwJiml0IHrE/cVvJsSm8XAv7sm4yIiB8kAj8FdHP
s9sjHX0pjMr/j0v2l5IqTlpnIYSh+XGF/apr4b73FGXfJeXQ60LK6RdQfX0bZLKE
0LNVXEp2MGACs3vTOtEKKtWs1PIoHG1JalUX9AYcBSliIMkIb/z5NCC8OAW1AZ/3
N77sJuGXCpNGepqmvHua4AqbhvJS8CHm+In63H137LyggH+fGZwMThGN75V5x3hG
HPXC16zOGjLU2AmwKUPseGjWeil8z1gmZKvJ5NaOCxTog/gRczNIpmClJk7ECqq2
xRbqLsjuc1gHb88DQzdR2POUP0fzmB8GX7VmiyHE0bKdj7UDoSIyrmQCE7A9R2hz
KpYTdBIrTEeej3W4JPu+36hpqElQRB3vHLij94+nhAL2KTdlW+QIu7Q8G7r1urMg
AHQsZYBOvniikSCICNsNoBltpmxLdD+z0mGwc90wGzMBE+zepGW4K4Fr8/fqBnvM
+2nhnQuIGjJoc5/8di2qr5bizs8pzPRCcY297h695T6Fmoid48OREV+PcArvxHHU
qnK/f6VOnUcblJzz4vw5LKS5hhW3u3cYNyjHRHK6ZIm6V6Dfl4yQnJZh9qL+fWz8
bKmK5nWGo4oi7BsfNK6Mk/x+FD+IfDB6qGad2iLhFFVslB3oj0vZ6AkHra3oVSyh
ZxY9GgRP1+LfoT73hwj5BgsgwJFCbtMd6LHqyP9gmodLZUM15S1jKt1z3xEH2LNu
0lNo80G+BaF20heEg3wTzviCFtZQ72B9JdMShlh5IngIX+Tet+V6h7cQ/mWW0bxn
zhrGM5/HI4SkUSzK7zaapQyagHM7zHaK97qxqo2i8nhfpvYRFnbSEUzm/YbO3bLE
5uhfLwWdSZnebYRvLg2lJFa4OEwNtvmz0gXNkL6UyHYYBGQyuEprk8DXx7D+oKKH
RIYVheqaJiqJ+A8YHsPeSkF1P757oBnaZzn1zOd60Ud/ZuXPzeJbQQ0Q6+Nr9P7l
70YE5fuyKYg8xmr0la84xBYzI0yq71kLYGZQzc0U3dOVFXpupRrblzGTo+ToLFtm
91sSnGq6bHwwJarNWMUYI9jVQy0IZy6cPYJnAqNN4ic91JDmXFWqqkgKMnJYg57i
d5yEtk96zfe8gFEvc7L7sbbSglmbJaMqS4vpfbav/LBqOrTIVOqrL3Qw3vQsdBUP
7OhLlXdWujhvIHeC3+/NCtxddpFuO0MH4uaZEVtyshiaA2aeUzBuwE9O/ZUV0QgN
jLU+RV+Z7xauQO4OwXSPyII760OUeX99bf0VLFxp/TWR9ISYxS8n9w55GR96wBNq
XNQbYpyzWmUWwuzuXyZbr8o+jmbBg11kN/Oh+5yvvmosZFUnwSAiKjeUpqXNzK/M
aP76ApLLy4epSDlvhYlotAMTmULm+iYEdDr6TznwHOkXHVKuAEtZfSII43D6uK0r
CqZtxhX6gEYT7MSgo6vW6hy3yQKLd7b4s+Q8GOSRpEHX4Rz8skoFlWoyXKg+1T/x
2+DqIjsV0L5Gu3aLcHPY3Nx1GNuNVbSEZvlaMyDMsbpoxENSZBwf9F7W8eb6eb3p
9U8/6SoN9aj50IQ0+Iy5vJIFunUj0keXLejuY1N6VUY8f4JzEo5yZqzFW6IPoRdw
7A7bjD+T26N8al2uEiTPaqHQMnQ/jNf0984jAnq/6QJlgwJN3Ci8WAapj3gq8C+b
WiBq8JgexkgKilvax4tqYCPvp8+Nf8Nsexgcna0Pbg7ZGsx63NFXacKDNqfOi7D4
je3MX7Xuo7p4QIT79NYFH38g34qTPp7AGijxj4MazmQiqplqAg021AbiRBSLnncU
04bQeGJZEsf+nnTORO9XwDF+m7eCtWUPjLDks2UNhYuRlvy28VFWc9szJ6j6Lz+t
zwmSi2CHqZhlKEm74KmEgjf5BRQDp0XOZHbKwaS1Op1BuuVtcVHajIiT7lGJnBKT
nMTmdtuAutQI9Aw6N7AwAJmosO9iHIN+SG24Vy49BMLqDbD1eRmueq25O/nS8ZmX
V7DJgjFtdOVJmvzhBq0vUJlbae+LYoMZqW/9+ehoyE1/J6C6K0Pdgf7a/LiEOSkn
5uG1CtkXYWLpUrNUXQ3swL4eRi9fsBeDf8TcwvZYjZYDcsq4upXsK7L9eTQLAhWr
PCjNy3hwqU3amdDRlLwA0G12sD25vukX81zN+aXa2/Yx+sXOvHD1NpRoWh2Am8Co
B7bTOqs4ffMpH6+lz8sAErlQ3p6BZwrHSKdZ0BlBoKf8mrPe9nuA8S88lCCIQF2k
ZTb/iJuPiaFFepvv4pSZgavugmDavTZxKb0yTR68hnqA/pJNHcgP8czzYWWqsLkG
YvoFT+3LVH3YrQyckCSrPKpL1RsNx7qYUjuAS7JINuvWIbkDhoRE2Ps4V56OfNud
stvfow9xNUurLAe3K1lnjRXJo4ZFjq7rlsCyNYrOh0WyKmhwLsbPKBwEYmSGJ+bh
WOix8L+I4wz7ZInSjMK86z4Wi8LM6gHzLgyf4uDvt2YoRAZId4JsF6+sNPhX5Af8
K8JF2JzgOJazp52rXnPi77h544lh7+mQuV1ONcd6KkyEbemWNf7vf7w1a2VQUZ8D
TDKUKYPM262rl6iScUWdQUgBjuP7/95qWt3ZilRDcNTDhq+VtseDrXxeAR0nXa7t
drbpF9hAlDcYpscXpyvi4ZrLmmvZoYUTgq9RPr3Phkvk80fa8jjhRrSTBVRJ6P7z
W+s46KGb9MttZjmFnbOV0JfeOOoCc6kg/CJ67oKklcBJvkEEMsifB23VI6I2jt3H
+UFhxY2jdErH8aYm6IfQdJzIHhB3ldDcbp6GBjCOx3ElB7dwAB9hOSjeNZSLxIde
ki8Lg5x0rl1GlsZesm98yGchdlBc3YYBWwhO1eDdPjlvo/LLuoEUYHk9OwUBhT55
IUZ0y7DfmftmQM75+Y898AAI1+bJJZcj6mn3gwyFvq5z2my4rXJT1BBVOuhNSL/I
fHmAsLqObeiYTjMj2z7Y0IfpMz2RJITy1b+fmkzOfRbz8AvjqNrF0QiW1W7P3L6M
QIJVndgUrntq473XDspjV4PBfXJOBwXvYvVAFbXeF37eauopx5O65K7VU6BfScz8
rgg+IS51i15U0yRC42ZVX2hFLkx0mzxZ+5DnHKM3XOmeIyBCJDYpM8luOknI2NC1
tTZVacfJTu8YjJkeqy+AmFGFLLIR/o6EC/t+doXPlrSQTRZqiv+uLW8CF4xLFw60
gQczQh1LSs3ZoBy/JpX/f+GrNOMijABI6ir2l/5xRlWtJndeEq+5iYHCo96FOVmh
mIHiieS0A4wdzk5g4WUSkhLKRQ/y6T+vinzxUSyQ5bQMUM8EUn2ljYUc2iufxVyL
2/ibeiunA/j4b6xnMplo+Sgd83oE80iftyuLbkMm2D1/HsGWdtbzrGH6/pRUlJQr
8roZrqEJN5ZpcpsoK9fnNjSD9FJVnFA4L4jzKmFs1XWFHxvQCh6p9gIhqTHk5d7u
OvryPPS4xn//lC/Ev+JzjeswzOYGtiQ3y3PdB4iwXSdsZ2QCMga8XxMZMTok3OXO
bcpZq89CTCL/wGUlv8GC8mRsjEf5C6hDW2vt+9rVGacjve8WV0t3tyjCvetJvqWB
wMj4Bbez9G+tc7ZmnOUmMqo2BwJPSyyKh74ncwJ7B1qG5zrIDhNd67AzYnTG4tud
7WEqGpVcyxHC6Af61SgP5vVBE4n+ZAVVJtTepFj4QUx24pPxvHhU79PMa8jFv56p
pjgK9iGlP/OUKnKgGrgutqUwdDtXhNa4gW7SkyWFFHtEZHhM5m38xETThqPHehVS
Y84Hn1DC+3qrD1OrVYRtSYf3c0FGL396uwslHe3cYIk1L3Xxn9/SP3v6BfAU3WHT
sPFb6qgpHBIKDw4/A9LIn8BgRBydr3Uuhd5fXBjnlHC4Bpb6cpb5flvhf5nBzDXd
+bh6enCHZt7HTV2+p21H96bXKDXVqzFV0RZDX+a+07ymJ+yGG1cw32oQY9oMaKGH
uoIq24e7ACUpif8fwPakX6+IU+JNIX+RS970+50WA0Cp/JPuL0FvKn56mppzUo4g
a7gxqwjoX7by3dlFJCnfz8rOQjlNjvK4/myhthC/sPMAI1pzkmtyemAAXb3iDcT5
G0ocGYCSEijmGSHYHEZHRuDdJ5v+AcLuCz1FlVvv7N8o9e4/k66ha7OD/E0bC8vy
ljI/jtFe/pxLhnsHh0ns8vcUG+8H4HDef9hft6lpbzV1+dXrr9/ztzxOCKqvGaQv
Zxo0K+Fhaq1lg6L3BEpbj9qeu+ehJ/0MSDJiKfSAjz20oi5stJorc2ZjgVBu7K9Q
8uezBj3mO1Ba/OF1LXg3QZ1c7L6VVV6Izew6VE0KoHEV+aemDKNq3/JI6+9YkPXR
yizeiwjoDVyvABIljBvphpDNS5M8+gW4AKJAnX7QINPaKCVRuiTVvjpAEjmaumEd
81VAcQTAD4wAAz6tU1ed7hX3l4a1krEHr4ADFxQtCKeOg6iAprxOPD3NPM4jI1UT
8J9o6nxqYam/eHBagvB8huT19CSx0SklsRFjOpw+ikb4WNGFJbWkrP6d4NDJocAS
QrV45P44psXEE9En0lFZV6V3sZB+6mQ79myUPA9pFStdFDMPxHz3XY3z4PdFQO+X
VJA6M2KQIfX2IxADQB7U8aGaizjEE4TUU0e8SRQRbTz04L/rImS/fFgFwk7D4hzt
SbBGEyyKcmr4MLl+9AoUOUhrhhKY4nLoU+bwFGRu5ahTd0FCsyqfg227FW1P0A9X
f5h2MTGzxkazWDEMf9zITPV5wrW+HpSIhrcH43qiZD8fGkX4YmlKbrPd3SanXRLf
zb4xSG/QIP15lKxhynf2o7G7H3kwYjsQ1IXsQxVxihCKHZ1GRo85x+NjeFQEh2jq
JhfdCqZCF54xMhWtx8Ze+GRe+kAtK/jqK2kRoqEfN/NHYCcAwbrunSX9w6j06ZXC
Oj5FeC3NEAqBeueo3DplmpkIA9gGmfpOaaj0FFwh0NctdC9uMlED/nLa6mF8OkSs
ZnVC1ZNUbDkLIZKwx0eFq5WkbCNoZBxlxjFxzyLsSt2i646KcMwDsi+8Ej4DkWa9
pJ/z+JaQhkjITld0R8OBpeyacsc5gJRjEu/P1v93iXP2LiALhIeY+IG79t5uaLCh
EVG2BkYDI9VgzqqkPuuyL88YLz/PMX8CgVP1aLcghAFT7y6ou6Ew8pMovdPR8gFJ
BJk+bZcwwpDNu9usV/t5XdaQngFtwPpxzRPHbkBqKceaaCxGfF71pdJJs/Aqkmih
Af6B031ZWTqNdHWxKkb83nMekRDmwvGx3EU+HQAqrKrqgV+OwkbiL4MCesk54Bb8
A2PwIvkBqcx90xnT72BYCZNVZI6/sIrFDjRNIjsuJ+NlKtYq8LkCu1mHZCMBk766
ZbxlS6qt4BCkvUwudibdscRtDef5v/r4NrSwWBApNrAeDTy4ojYaBhTvXcGPXoIU
1PNG0dJe/Rg+bXBmtUHRcnCASXdWQt7Ig1ATzt/MxqB1iicUv0RBDeVI7Iffufw2
w19bjYh5nUTkQ4ynA2/3Q9whMK2ZYPIZ30YT7FB6ZXUQNqNGthRN7pgnJ15QYNms
l7ICn5wBiiih+3tuPdMh65m5q0iVdfkCePbXoniqT3T3PP1Jn0HEmUI331quKK7f
/ua6SYHDtXahnx45YUnH/Q016M1PCdwkiYf3rUiHXojgRCihRrC1z6DnkzqzA2P6
FHtAoxr4mV9R53wBfbNFDiHyQMcJeKr7NggTz+2GVe+y2s4SrUFlUmjNht9fKDFY
F6VzATGjJwxSnj2/9FkRfY0IDJ/Geqg71E5uH7Q7bWBGJEXKV+1QSo4S/0EKOffv
w0aQqR5m83kpNRAt1mHl4Dals5AtpYdvjIeKEq+gueaY4Je4M90/JWPRULzBZ/ZA
OsV9ewxHubpppE1cNQPGnNwXrimZ+UJgZXiG4KKJRN6Y/xFansy2Da2RrAa2DEmE
De+Hcst8V/YX928ShFgDVLSheJR6vesJ7ThRK/NHi1Bf2y3uvXY4FthGcQzBwyhZ
lldaudCkngc+OhK7Vt2dDvhXys6IGUBfb4XQAKdW3KHyI4nNBXspXQ/3sSPJQONb
znXUZCTMMya8ZaYVRTqzaZJuzN5P0yyCPhRCXwUr+ryAatxjltoqjfDd2fDONljU
xxeY0N5mW5nrhH2KJc2aMAs+CfsANrMDzxC5XD7x9hr+fcPxw34bYx+7g97SsXN7
knenE8jYzO9e6jHwXQQzvnvHuRaNzjZn4HPRZbydFL+/D/vTkDjHDPZBqjIW9+fB
Wm5YVzBZblHRWCIgHy3ZYmdxYVuYrZxno91PmBStBJtxlgA3nYzXZzczVx1GOsN1
Zg1S1v48z7CzMGLNeh+p4Y8jXIytS27sied4p6l2kGxkH9u5pxFklQlD9Fh/i03m
i3CBItxEJt3ndmuVhwEbMOmRzXYf0DSCatfy47hpAGeo81pH5W/f24lUQgnewzue
WSLUcF1VVfcPhwSE2eOfTq8n9KkxHB3c470EoEsDOnrBLl79nCHWqSWZAcP+kbKv
ODHrCWxq6xlBImD5EQ+Dw3WiDqWEOj8HbvAzjO/tgjnXMjLdQ+pn3z8b6Jeb2Ama
+RfX6sDrRQImgb8VPllue/BDOPs7/dzP82gdcqBpsoXkj4vwa5c6eCAJ9wajurpj
gzPR+N6GJnzI5J08YzSES1xiuYcaJpSBx7ypTfsfRN5UqseoOEFaRJdZa4OEZ3XL
POeZqr8GicK49gWNAbRpsmQQ0DZhkCNdlQTNXeGsV1A0hBvHn680HjGveFcjqJhN
djz3ffEdsVG7Zpghm4wmu2fmXin725MymtbTzUFWTtaGdMPBlGr4RLECglahBkIU
J7CXGLQ3bUTnuj7TvW+b//3s1f/Jh7G0j6LWZLrHk2F2QjbJr/Kfa28Nek7pX0jr
uJV9+zgVnPNMVjXc7UQR6HAIIKWOaB67DLZtYirBFwFsrMdpayDmIMaoBysktn47
5VkzGouRoLN8KRyuypwSkJvm8RtBIEGjWKoU5MfsC15ouWkxMgHsZdrO9bFCenAx
6CydT3T7o5Hb/gsbXyumHir58+sa204Ypbg1CvUQ7BA6nce7xovThRstiBpVfprv
Ia2Pgyl1lS11cZ5FBH7ehRwj/mmnnUv8UryVSVokxs2grIiBGKSkPGgfRAwZ+DZE
AmnJZqRUsqUYvn8/RWfZmL128eopwZieIRosvAtvGPnCkKzaacCOSsqUhM4CQWJI
8LnUanN1WHTMnZys4H2i1gWL+F4vlOBitIjp20tgMRgucQn4msHxAWcKp1v+0C4G
oOiPOW+FGKVWlo+7KRwu0cIut0ReTaJ5IG1wg8ZgBczEuseqjIzjoR4/dpE56nYx
9H5LUsi+FLLNiENNSa7GxGuO9lvw8/7nZZ9AIZxCo7AAye3nCu+j38tejbrZ43q0
/cARf4aLrl/cGvgzj2KLtRLhiYpxlf0TyGBcxsi5Q8Hs/AfLPXtGCWZziQmRf2ol
8QtyJLVOyFGhg2q7e0UyEsbpg62ZEJ93jpE/gUXp400T8I2eGfRAiF65fIhrxf3j
kFX5lEZ42XshZ8L9Q2WiO/5sMwvKXhLe49zlXrUvXQ3nAJ9yp1GZtidq3WKRv7Te
8JOgbXh8t1P6lxe13mF+B3B+Jtm+Acm2/TueCexX69mOf+PImsy7S33SC75Kj9Ie
/x2EjA9TRZbyLQhbC9xqIIgop9OfeO+o4SszODCZfaK+WP03NsWX4yDpzcEvS4JV
RATJZYHNn/1M7gybV2xm2ve43YiUL9RH987H5rblzvWul/ggGQQnaMowuSCRW+Or
54f5+Ws731nbKRhZmimgLwQN3Uk9r4c2kWiGPizDwVFkga9Sd5y5yqqGiWERRa7k
OydN40VUZDYq1Ni6kf/yC2yuHQcJXSjWHAcH9YnmLWgWsxsMfx5WdBt9OIVJHqUR
3pvWBffRw9Ddj9DaWCKO5+PledwAH1FNOE4/OCKBK3IVvzjfO+caOY94U/yKTi9M
UjmeDj9VdSM70h/00NnqlEPVTjhzCRNbX02jStc4Jzo1le/5nSRQcsPhwRNTTs7G
TUOVtOKPBHOzHkhxAmcR9NDPrkClLbxlyj73zr+EGs7n43pGGEaUEc4OkR0wTGKx
Ey9O3Y27j2Mv8mpbt35yHn8mn+9ts03Xr6dxqTXwSfTXo5wDt696UsihxZhpj69M
8HdIpO/ePKzdYbDTS5jO8YzkajYnFgmcGzfTNFTGhuTnzG7xc+MnbKOPp8ovDwwh
qFovCx2otueNMHiXGZw0YSraJ9Spg14XbEKWw2FzqW006+HwQ0EN7PqhMpxudmax
DgFnyRxs+hFYtZrPjTEXYHnLP5dq+Rx0Usv1goTRqtZBvo1aBxQLyxWm2/GxPv26
SUMi8h9G9Wz2pCnbte31K/LfXmQClaKV9WyFn9GIEmxi8WffNwJdhkJlPD4B+6pD
rKK2z3y45/Q2Ap3RL4RlURpo3lnhmYp1kveFW3N0WT/A5WjG3EHscuktUsF/H9T/
XEpnHNo4tWPzniyuuEnZERCJb26JQUO4qoqSwo0ZNM+hz3VfWY+ys7yBJ8rDGxn0
AlzY/038HT6Ivb9ep3pt5ddIssLl6NnHYOq8p0FTwbR5v63gZTkouJLnQcrtjPqd
69jrKIoIgYWbofFhJDwixBD32jF+GtAaS+7SPB4fBrfG1smSjBeq4LpEZClkuVx7
IpjjbIRROiDbq4Nthht3HFwxaW2S1Z9wjcBTmzjU35fs+Dnd1bcPqa72Up3WLjPd
RtcbMQnk9s80o/BQ+C53vtG6C/QQ+bE4j7DQf/GzzViEcHPePoSW2AYBWsfS3TFo
xQ9s+M6zTe8LH8aW8dgXfnpeWParVSgiar1V2GGoe/+oZ28WjC0AE1YnG7EgpiMY
7KVf95cVn3Q+zoG67L5zsym2LZXoneGiOqWOuNYJvj7NxVuqD7iZdgtWuvc+W9z+
9IN0Qk9k558VZ72I3qYdi42NWC33/R6X61IpJ40tcvfrmgQM1s2bGMrBERWRs1Uf
oIG5RHKE+UALpgPwboYFbCPmpAqX3dx+n+Ji1TpcvORy4c/MGcaP8729zWdi0Xq1
fJ65rC5fw81s+Zap5erYsrBtV+cNwmjpBB2VErp2oRldHfF5PdNwO67TqRfRjBL5
nDs1Gku+gStbW6V4JOksgYoUadMFJy6LVyDExGAXit8j/u8eAFrVX5XqQVRDBk+f
0U/xkg2otDnUh+mphKePmhRV6Q7A9dMoaxRg4fc6CcF5fq5QvnFdkoPYrLVZzcAr
WMJQ+qf2r4C3cxBObMF30QNMTbdOBH3z4j/TbqoK8XkLJtJlyipXeqVDo+njnr9l
IQvVgrsbGhn+rpyieRYYWDR1+dWlpGzLqFJrU5oIEpexAfjJdhKToqd8iXUJXK+y
CRRIfxaHiCoK+RUyTKhgTIDn96RDkqh9Y9lZfRXPUHYcBoKcDn2dz0I26jcSZimU
SqYH6DhjC1XqLyG18m0Lh/UahfurI/4CJhSXOtvOhXPiC5LSAwoUQlG2k9pRWXjL
dk3ZKYsvxaXBr0BWzOA5wwgK5RxbbsUb26aOBg1FvnYqJlG6g/TkICtj1zDLI2zt
jAmhw5+dSi+gCRB3b1HW59QuHa1fnu+R7b8jfZq8LYHN95s6lNkXlCByt+DpkrGh
2vQbVNyY/AWvCb3ueHHqa11pZvzwOgnvlJu7DOY8LdaFLWhS03v4LQoYokL2cG08
pcgg7zBU1AL/ZrR0/SUcl5xnQ7z2e3hi+6SR/15ONeejFhf6A8jCsJIuLEFip4iL
RKESBSh/ejLp5Q/1EcaB1ai6KQlpt+xao/cB9onIg/HhOnsjyAE1kngtSJP41WzC
K1RXEDGgM7WhJtMgElZ9D+rrUQaDKrGnW/Z+i/huA5ZAkEKICHH1DTVolxnyLsCP
uGikDVW83H1O7VLJrWjQ4pEMq04N0aEzffXWeqfENisEL3YAjOyKpuF5yEk68cqh
wPmU+seOC433qoYpBpRJMw1SgNu+kUDRmhdwEl5WlEZx75ImbPOJ/Jk4doe9Ctln
rH7aOiafNevQi8XDzfJaAyPWleG9hL87kRJMnjKUL8MOVgcuq452Q+/4gJ9V79gm
zUjK2dXqV+r2fFMpHvDXhywPVp60/NlvcaKd4BYLrKkNPiEpzDLX8ScJNhah5NyJ
DqzA/YFSbS8vAnFPRL+noOVirgHP+BncjykYFsx70ZKWI3PN5edLbFtniU99DBC2
YoqViMfyBsA5pWDrDkaa44drDRuPEs4HaGJItf3CaSir/mjBKQ0oD4yVi2bu4CnR
zgECVKQ06N3ZkFG4Naaeryrga2lItuIbBL3o94lL6zW7G7VA4KpjVC/lbcneL5Iv
++4cqkh+AluDGk6hNK82fQUknPkZjgD9kcK8BnLxCgc1nuBaBADcNXIQL83ZQbpM
eeqOmFokKrZbf0Y8PPvBiCNVWU+O3DnmWmdW4ekx0gwS9BstsKsP48Eu5mcnis0i
sdQJ4qCwZ2NynmmZwHiysnswjtNk1C6tQqdURsqABTwzXxKG8gXYq2j03iLrT9N0
1YgDHLje6CDFkcXyFMzwoRRl6htuoUkVmbJ2mnt0rizcLTJaFAt0ZLsHb6hhAgxn
1EhzxqHszAW3WYUAnr39xcNkyrweOMxlVcniuAGG2EgKjwV4gLgP4JLlid+s2jK/
WH5lycGBybsKdmu3Dl7YeHBcVzmHoTGXx10VfedmF1kIZP/suv3UBvKXhJ3HPxvU
dpttyRL1zZSBSiP4Q1bNRSYP28b3/IDfTqkBbqove9Eg21VgcsLfRplZi7vUdRgJ
rhKJS/V068dqCU6czTKH113TcIpx4dEBwLGHD3SaRTFerNUDWdNQuWZjRNPy3iw5
1GjEigsuqssZJya1psaeuiUsi0muZbQ+sDGyUXopw4+sSQsXcVVY0sC9NaNpVOZP
NPK5ZbOxLu8GPKX3sNqgBLUPy0pmLa2Z66a4Fl4am9n5QM1Q0aoEWQlbqAPlCf7A
WdExt85OpjPv94O4tgbKB6TKkPL3CSab9x/9KWJ2jrAdI/BUi5C7iSsk/bRbii5W
lrgWMU7Jf4eqDF1md6cClDcM2P58JBYTuQYXQNaOSUblzyAw0dRV3vc+Cv4xJ9Dh
2G9HNI1efzjo3vYiJv1D2J+/AG5jpxZtY24pBtv9zx838GNlBcNmv6Y6PoudFkLP
uZm5Zus1svvtYI7MBhEEGWPUj7L2hl0buQk22GjN1lN+cpcnugWOnUcE6R8puNsF
DkWNCOvsHlRdty6Gqk/PHlfjid8oJx+16aYKJpU4ztlSOR7A56swuBQBaOa5eQIR
HAGRi5E4d9s5JtqmRNFQvdFTloShFcoWjcGWkyS+SfrXmeDBrO2aR/QGqiCi79n0
ObL8+4OyUgqe0LHl47jRInhWwFUhH4NZQHvUcaRCU9AYZtmtOMBVdIoK+LVql5MY
CJauk9iiTSlszqsmN3dT/vFRkNDpTKXo5rBXfgoQmPiwSsjq65Qw3UVhr9ywdD+M
KVldIg/Z6sDlO09Ukr1UiU4MDDb2zsbwZdcZvB2TCDH2CMhunq/DFcd02NRE8D8O
tnNfXsnuyVj5M18KQmAlT4ad/ULAb++n/MtYJs49aVq70zdUh2MxQ61wgLTInF9Y
qK+mcdlCQhBW8QMafCwsQpV6zryMr7/ei6DJOua0NIkDZtuz9mGNjDC7sU6NeUb5
UwuEWDz0Z2VeNWtDJSyFAZubHBjzUY8thJvuCVBDFNwiPVayQYVwG6RcCO62hb9U
V6uEL8xKDuA4w3Qw1pBRdqCkYVNWh/mfx+lmdhG93fdW9o2CnZghicFjGjv+6XtQ
2d6sl1PCwAp5hdFZGgGCBtLBtg7ymVzBI26O7d1+D7xlmlkgDhkPdeBpPzs18hUu
LdkTYeeD55b8U2rnZhoOQG5ZhmFnqRgJDzLOJLhzrzfRUndQkNY6nEMTX5AKfnHh
Qarw9iWv7JkGmGfICik/hCyUq1nU9EG03bOaJPKP64ebkc4dNw7uIVWT25mot0f8
ZIEoyOHMTyhLewLERslumFx6aY56mjQDirOL5L6zIxGITann0lNOs+j4AxkPyxNy
9S7bK5yTQO/Ht6Ikd4fqgxQVo3sI3IaGb+5h8v2jfgmt9O5nTZqeeRaqMytnHW8u
KQt2aBByBrNFmYnI303B4+fkaWsra45FWI3hu8cdUKegDK1RC58FcapUJ4BmszlG
QHL4MFJ9vTQnCnlZJh/wiALICCTfFflilx9zKbK2W1RuYgzE9uxAQLfvKAA+/YXL
P8HxhWzHe2uG2R9flTtFU85LqLHGJ8n/D+FbqJe8XISrE8mZOfP0CZaRVV+S5Zgq
sQ5eHHQu+qNCOyHbWksNCAktocXV8U9UAnyL2MsNhqV1hBoQUGRhhGVcrsRAP7wL
X8cBMRyh+l618KJyqy7JrFzsp/I5X742mFWARAvz2gooQtsr9jodf3XnKz3yoXKU
F4y7akZ3LMZISoA6m6c/3/mOyxjELXjMlRSOqJli9kOhx5G9v7g+9Vd7FfnvxYCQ
14fFgWATLOUVmVUiu23uwjPRpEdJFbtrqUTR5ucj3tMMxJN03QY5hr/0RLZKYJoL
5KOjqON8BINtEdXuMuQyK5YxPPI9IbuW9lA7ljjiSknlbUI2vZEbSqw/4zfMQiB7
3A63F0g/YYVKzl4Sohf4CyUOZpB14TIV3DmqRyvHtoZzs7oCijSceAuH0OnGQSao
6hEOxkWP6japSqZBv1w3qrZ1DVe7VjAJJOmdbo5LVQNm+3GGqxK36X28hE25Bvsz
Ji4SpLex1Bmob67Y3xjqBgFfu7WRxNLzUA3GmEJvmmTuTmowIzHEqsGUGKLwUaJc
waxdl/Rm2dm6ZAsjf7d447HpzAT7yb2EDtH21PDOtXjyAG9wtOBtm9NUZ3+20MMi
Plf1c5rk8VDmcRa0V7dtIIsCofNZe4mIN8ZWVa3OOnWcIKJC2My8Hn3BhZofSimH
UkfBVO0BOAzpqT3Jvljem1w7kZujVsdsa75RSHPkn2/6Fy/waGOynBtERh8YmmLr
1MIVPt36+Hk4VF4oeVLNi9dZMqaukVIcouQcKslXPtb3/jzZ/qshhiz1VqBDFHDT
jmQOb/z8NB/aoT0OeXg7milojjRpfPPhMa/TVlug49HEPiKwc2HLXYh3iqHSAJDK
/MkpQPbuWsPqBw5fZB0xAWqSuPXXc6NtNMgKX2xjyz+xDv9DNSWXOdlYeosSJamR
ugg+f5kxzsyGEVqetKpwk2Oh3cF7aqCMfnwhxU2BpyPta0nwzbvOzWGXCLZhUtd6
IPw+mW/dQ6JO4rNmTcLYh2xeQTNdSMznLe8aCY7Lk+4LKL3EfhcFr5Flxkui8EJ7
YfUwcpkksZ44c3CI+rJ34f3/3hI7eFXmep8CPrin4WntprdWIBbDA/zbYkNuh8/7
x+bM6x+cMV4zblkvZ34E2yVp466ei2/ck7JnXVYxV0R+Bv+MtCKRidnBCHLNCCgZ
qV/6x3iIIvttlyDwUQ3/CfEMPR9WOKL3VEoZ/lrikEVFNcVIH/ZQJbzGrYoPuaGU
v/gzInsceytYsFyBzVbDq89v5Q/mRZShgBgTyPB3NcVBkasghopMe0TYNZLMTfpt
wktJmzgmnRXmLA8pTJMa8H8w7/BTr1HAUsiPkBetD28sT2CPfL/oAEVYYGlvm29x
PpADnBwg1HQE83h+SryPqsrENa1C3DcJUkcf3YqRUXyKijWLxBycupUaBOzOWi4I
uFxLK3+8dnIUrSue7vhWJflQZaEQ+2qWHlJnM2JmPeQs+aM9vlLpDpoVkiN+2urS
eeRwxmYPkl8ReUpU5EdVLzfM7D8I/LuCWjjd+N7E3v+bv9odmv5kDrtV350799Rl
SbGjy9tkefQAlAqKOdpA+pxmN45PFHUmF+L6XauTU7Vhn3tZyLk5hnwVWrxePv/n
eEkFJQJfX8CxWsMfed4/fbidmNgOhPcwYpkyWEgZ+5evzbVeW43ChdpVu04jkd0K
wxOx0NYTXKsVozc1X6JdnYU0lZmEUY+MsWAtdN4Vyo8TW6skTwqlcn8XzKi3zrBf
BFj41rTt2dIlQ1SLFOE+KUoK1deEQNzEjDcQdLBqLxqo96m8nlvHuLk9i6kWtdOB
3KLQWkxu/yTH+L5Tm2guBuxxavDbkP/+uVazO67R9d8k4ogE9jSfwJVXxjn9vymB
86ARnny1bxRqhhPC6npZ3LWHpb1YbIbgs9WMJsCHwvqmzrjY6Zsfs7VXgwUZw47l
7IvySLOxSUFOAmR+SdhYVXhFxE2jThviq4tjRnaqXfqWMJEEFa11Iq1lDOWOEBNc
O9gfWe/4GBatn5zIc5Ns+JuOjMr82QrzPx8T/GJ5vymdhLxfyaCe1HijoFOyRUWO
D9KNrc0mMzmBumoDFDcdAfWqbXXtTbSezH7n/u02GzEIP7OtxNCqwynY8ncNi6R4
og03OLOM36C0oZoNU+kRPc/11BY89TNdjhqOe5E6da4LWbiDL1JzzZCoG8FECOFs
1mH3F0WQojznykxr2IU5krPpCLFEVSnOuO7owdyUirYBPhYrtBV83fFQ4d5XNBtp
eSP7+UjCJI3wtJEhE42bceJGIchiDhWwB8Y4c2LB8q60y6nOsuLdQeBjPaWAytiM
T1nOYNnRZua5LTPG/8lgJYkAaMYYV3H2/0rdPRxhZQwLusW5To1MKBBKGawvb0Ck
fpQWeDq8UFmMEvNG0obrF2UEg4wHYDYgzADMWlVDYpy5IqlMNJoHchf7zUdLl/aa
yUvYPQAg2B9D9Ie4BGo7PctBvlBN2bbTl9q4CrLAd8vl+CETELER/8KKSQX7ZXez
WZ947hlxI4v8hyFNJfTXMmZ4w1BZGLt/ttA3jnMKbOjGZRrpbYxGy0dqfrEMySOH
B0tOwKh4XvQzeyyFFoJweYSZAcjyn5BRJNIQ3uk24DDSc1/ddV+XaeNKYtupWglQ
mK9vXXYdphpE+JKpDHUsJhgu0t4C/TWK8QyPpTpmIWT4Bb+0sqc+04UvSdCuQuBi
iS+R3Z6k+nEtrSUBney4ClVLMl1YHKo3wH8Cm/CChJ/Q5YaujKHXLTGfn035FQDK
Gq2ZvBDX6Z6V3e6WCgEUNnnv0eWgcoNHWWQXyVaEGZIAOyDhatNyrs9a0wuSLe3e
fBMIsclhQ8VQKIu4ET1JNAIknVsZuRJxR1UEiFAZYcpAqLYIyp1tg8aRSl4tD4tQ
S2NTxp0aET3y/0PerymusBTuqQ8gO+NUIp0/i45jaIS/D3XmDMEl3ddH6lYba8aG
jLl9Z//GxvIMEPemoje6BQySNjgtpGQvVi1gU+wcnKzv+FMyhzxm1cg0yyCZC2ga
jTtezmlmtbX6dv2jIshKcnEcczNJqMz+nSHHzrbl5IQANZfgaMc/JadG4g4MjtOc
AJUCOpjg4t391jJUxnImYExp5aRCRAXZbubFFXWhjPuZrIsmqbiIog+pGT9cZnuo
ENhA49GQayJzWvoYjP8r/Y6ZNrhAaRuZXCLUdoXjXQdmaUCzmcBq4RoE8RYsWvz2
BSawqRoTP19lgmBB3tBWGlPoeOfGrCVsUH8/KvcHOi6PXMX4E+S0T99e5YWh9T/z
ufsggxclWBayxRZExEp3MvRxXQQAAhtAWR+KDXZ3GP6mOdZ0z3zhU7iD15SQ2iP+
viuGCzHaP/JTHOaYLbWkMUqdOUE3bHiHv998BxF1KDhttHjApB2wpYbGwHXNaxM/
cT2mNpnVeRpZOCxUbJc4oItIemQ8AUeqN7KX2RGyYyx3Q1lhr3NcwjVq2YCxjqB/
4r+PmP2xX+2FTUy12XON+rmnLzaWOgj8X9hSYqLonCWr+QdjvvtFdn+bN2WF6mAL
h69hzGiiFphkgPKg8UHczJRK/sD1aRzHCJ5migr0qTKBXkv10AvL12bOU9Un5xXO
XGudaJyVtQLSLuZYhZvZjZV+hxfeKtJraT+RS/ghKe+moUF1D9JU/KauqjJ+aeL2
ZARQYyOYiqMnPQ3nZ4DLRPts7qyMTsDaNWhnEOl850PtUp2AhHMRKwMVlouhwsr9
i7ME+Q22e4h72uQrKlYMoK6Yh7lT30uovbmbkEZXEfR3JeCIdTTp6oxDB+Q5XYDT
EN27qkcdrCH6x090OksqZ3dtkEoqRJHrKospGDLrbHiU7KBfsekuHm/ikR/vdkjO
L1VetfVRDNxYyxnmFlrppQrC9f6OBlIZ4BMGWYqzK22Qes3OKjpYgeqxf/+QTvC1
9+irn0FKrhGRSEue4E3NklzOGW7RxqT+pGjm0jAKkesPbIcsALYYRuil4gDdSZag
Kxtgj5zV/Yf1fT+ATwVvXbGTpD8ShRDr0oH2ErWM9s50f0n+eMoBQqtl7xV/HbzV
7z+2CiYaOKtiDpGuU/t8U5jaJ3VpQu6AXdqVFj7ys/Ps0gwl7RXidbYJXtCajImx
17dVDKTSvGlOYNNpQ0d2iXArZ/08sxz7wO74jrVCb/VfBQej4BfRsKCszITScw9b
oR4WLiCPgyvpsu/50xSFbDxuWAIenloyyCdy+mFb0ytRAZENUTaCkjWF5JhIp4j2
ux8TLhYmsssOr1Je8Poy7CkBMwLBy+Un9nRxNBBSnKdq3brXr0V+pPg6WCcPkVeu
bE1TChOdGpPlvr7NaszoIC9+Oc2TYvaFT6arZUDyR9E6lu/wuq13/Cb35MnwLh+4
mGHIJnVPmV6YIvZqPcMUbxTOu1vQrWD3afed6Qh3srMneQAGq1vAe1+E2BZD78EH
sx9V/SJhqWJJwm8y0B56pI7pHIbR+2giZqGpDwjFTTcNcaNBhIcK5UUbVgGgHEI+
TS/zexn94mFSzuhQUih1I6HCqhbPWiq8jXUWIGxbPpuJVsMCflb00J3Rm2WrU73F
M7237MQ97iDPXniEzPcxwOTpdj/+enSJOT8Dxba7LpMAsNDyEwr3k9/RgNqIgOsh
D0pw+Pm5FeISuUJp2qC+kE1JAEu9bVDDUiuJEiZMCDo6b0GoOirCRxaggwZeVQyR
mHT1RRFzusMUlgfTt5uTyRCKP6XFVOR53t8AEigBZaVzbylkH6mvTloNTPhYMufw
QSkjRJP2dCPNwu+Xkz/PVYUCy/VzAIMV9siSZ/kbT+E6f5WgSVPkj8vTEUP9gtgb
+XIvOwesiHN+Dq3rfxo0QyJkPzttjuRUCsmAo/WwKYK/mZOWu1G9Q2qn+bJrEjBh
w439Ldze5o6I0+BQ1xZ9/6w8NLl3bdQVv6sV0gF0tEzQgzvTeFG2pXdX+/9gjc66
KfSuYbnVbmYgZl4y0LGAMhHZHAbhxSLzpQfHYMC/c6UpPLgE0mlZefBV5uPnWiFu
NwXiKpsOX3/aJaNnXGmrvIwrquLfkQhUIWroynjmYrSlobFyH6930TURg1V+hCbQ
w5UpjWHP5xH4S/fWb/eO/nX0n9NBjLx3KbQUtS6tIr4dJS9VmL8HtQ3cBZVNuDsU
xDGcW5kROGqn8wOzh1LUzAao1t6Du3r2NWAjpfv1Ms8b0dPD8htfzWgUAZlQ5JmV
yeii4QSwTB+gFUQFnjR/Qp9hACzxvJhLwwGM/FA2O66aDp6BTvIBc6+R/6gyh3cO
SffNfTSBJ93Ll8763skq08F8xvBcFf3B4lx9dMIBHWXNwKG6JSLjTiBf78HH/RUy
cnYS6m3OMZ6CDE9sP8ne3cOn2VB74wgn5+PYrnXUhisfFn8PbCVMoRLbSIU08cv5
Ppw6FLYyG8ozWOxp/c1DgFK+03vBujBBeKU3MQfJmQeXS7HbX9unKYPjuhFFIrxd
roO0JUK6ThtwoIUrvcv0azYKmuY3bTXM2iqrWQe2z7KGyAirgNJ/Ww650d9C4Dif
dgMZTOLqlfKldSupTQ67qVBRDA1/0fgH1HrNN2hNcIppinr1Id6uaNWn//WCshBD
cAt/a3fYaupeZteEJNTg9FAH/bfMEnSAmAcQ8f26oLKfwdwkATTnz+aTh/c8Kazk
IRkdK8jafE6M8zWjPj7wgNZDzbrJJ3uuZ0SSYgAJW22tSNjZkotIeHEVFImfhuya
7yfMigNNtZ/Z+uES05o7ta7wA6sBVslSDCYiMkcwfudHRipU+Jqgdab8i9ez2qyy
a+iDawAosDb2fW3fin4ptyDlFFUuN6QLv+ky0ybdiudUhZNhgLhj+qcS1PI7ixrs
FupoFCzPg0Ox3ScAdX/rVgcSpjku8452WL/3yDPDtdwIXJtZ87f09lTvBakfhbl1
SQrkLWqJ2GUCwJHjxD8IJ1M9uBj7mn3dW41MrBjUuFnuMOPPWK3OPZaGHIAHdJV0
6pi0pqsLl2gpyjJ95ng5zf4FBupSTCatZ01PI2IKwrJWpaJr1jE2yt35d5KWURut
p8vK0haa8hMG9WOGUAZrQoZ/jU2fcmnEdryqReFwZ8ZDAZ6vzSxQs+h9O5fFQB5u
ClKben47NtVugYGhQDGpB9xs5N0/mCsOFDN2Im2Ygyr90wP8UL435A2pCLam2lC/
AaTH9IlHcN3SKHdlNNAkuZH3GpktRpggzj5YNveqFmTHuJWF/Qtf8Yb28zB8yoAV
zCHcxxsvsihb8BBc2irs22orUKKeoydJDm1m78m6EZZb/m0CTYcrb/ry+Nb4KlSz
831LwHuCjVif61JHxh14pRc4Hmimjayr4PoEDIeUr0bx8OP23q0BVzpt7HLJUIHw
o4ojwhObg8ZULcGEjh3SkBDDEYKjezmfU4qFDRR8yUOEqZdMQ8buopMbTQ89iw+B
lyQHmBcDxxLA1SUS9LySxF83+5aL5gZvf3fJhVmw95YNho+HqDaj/MrZmthmD4Qh
N/j8g+yBnVB0JvOKhaJizgw+BuT9n9krZnUhB5wJFrBY1DTiXxAV2AzRCCWKpIrY
z5Y7jtxBkB96f4FGABXSMz5NWzuZFBrpuv1ESPsV4m66UtMoNPkQAzDtUsDxbsF2
YzChvtCid9p2eABLCGVXJNdYZ6pG7JSCVju4rpnMCzBfT9I4zkw8ESnR7QMVFMcE
HjNuqTSZw0IBZcrZcKqnqdxvNDpAfw76q/eZIevJtcdup2mmIUlijte6tFrHWzo4
54ULzWLrMnRQLrCn2+ekscgcXszQwb6CHdIT4PlX2V3CNPibRtOx6vm2zK0tl2r7
PanvplNd5emRpGgCFcGZ8zqcqAFxF8nOgcrV9QyxgncTJG+k7eQ+wJkDg+GMbymp
W7Y8fh+tVCYOir/I3EmI7aWBQ1zJPWkAhMGXuKVjuMH77bOCfOHFQP65b+ENekvJ
0oQXYErp4afadqfdqChjkyYr3PO3J4W2NSBWf+QkyWm0Rv/E0scsSvuQfrKjnREj
Oq+wEvia9lcp7cy6bNtCzsVZSEFKKLclAxRxPfrLPXUQK81jr7B0B+N8T3Jcka19
s2Q8LABN+1itw2LJQwguTe+NoHFK1Od2Dr9SYfBI5g1jUkGRlQLyigSfL2R2HTY0
Ty0lJBnotb0mx3F8fIZ485IjQmbN4VtwWpODCsAtFIshNT2GZJSOPQMWNarGADeC
tB1dHTsegtt3rXnoLqUu6v9nMz/iupf7FRPllz4eHxRZ6lTR6TYcfXM/82kjThGq
k3Uml3a4N3xGZwnE2JHbsmEcFekGJ/s2Aeg78bNt69jTfZyaF1ZR51fxiNo0i2VN
5zFO/qOEGI/HdoZckjF7TBOCYpulTzSd2CcoW2E53EltSUWD6M4X83d4FMBGqDYG
lt+HutU51PTtM/RgLyUzbfHuGed5GeNwqbsj7Rf32ZIt1inicffz8hqkF3XP92Ww
X2YCfbeu6rVNlvjLiWTmaw9GXKMjx/Ii3siXwyrEXrYGVjce2j7orpIvjqB/qvaq
fhfqGAe0E4hXDr2YZ0jYG7K+L9o/fVoi6ynXQLeThf+i+fpR3wfwV/QF+Kwt9dnp
Ib3EOi5geK4Kgwm/aS4rffCcJEepPYXXuOzQ2Lf8iG1Nc7rkX+ThuM6MTBuHJxB9
59JwRQ5V3UGCX1oA3fgeFKzjvrw5Sf4nhHPXG38wqmqu4f1LQJCTrP9JeQ3+gTmM
5Bv2WgYjZMI1GGeqcVQ3nyvkVaJu6ZGNNoZhT+M9r/V8L+fmmrzfegBqTSveb5UA
+e5dH/pibMdbKSvKhGGDhn8wjNeghh3Cd+A+l6bSn4b3CzVQlszpc30Q+qeH7qN8
RYdR8zuoK6d9uQahQ/eTYFzP/AHX9UH9Y1+zXT5+KQbs4+W8qr79FvJRa1E1KuKS
S7WkfRscqnzt2m08dMiQmpCLOWScH/V4ETgtGNppC0coE1M7GZEVsTkcCf9SA4Tf
aQ5Nd3RL4RFw6f9hOmo+Npt6CbKMX9KqMho4zPIakExylB9rObiYICTfzwolo8EV
UwDoy3axHCeAFSDAvND0bFazEZJk/wJOE01SyAru04NmrI81csiPKOJ7gbcLA714
LxBlZxiYotIJY0JzRzuw4JDUF80cU4RF37imqgljPveh/79iSQWcJRnvSp2oUVOn
Tt0SlYB5C70CJpnCuTVY0fpmtcxvPcTHYRlXY0Pdy8tZQAKyLnWzYBjXWkanbDp+
MuXVuge/FGPadARsi99BEJ+rnrGr57YE7+jUqE27i/1U6bhAb6I59h/HyaswP9CL
IQsgLxpnDwj7KascOQpd3y/tsvLfGlsDd9YEjjy4OP579VXU4X5ldGtiajAltT/2
Wo4+f24ztCgALDu9Us0oMkbFigraJMoif9Bq/iowmtsuc1/Co3EyWjLOjudzdFKh
HeTkmz3XnIum0+dRdFzmYmP/BV46f74o5gbw02auNtb+RUMeKDR76T9w4IboF2vu
tVsTxLFzLJTupZE5qjVsXVPF1C2FrFhxQk74EOLVqj0tzj+47G3V5b549Ff2buP/
8YR1kJIoDrKBlbgBry4nMkNZWXQ3LLK+hdE3W/fFxuM/PS2AT4LehnOKLGXL1UJj
anZbqUrlkXcXR0ioMLbCfYXYzDZ+feAkGrG/FwIiMDhUZyBjpQYe8gfx/TYagwAC
mSW0+Rh6iG9cVjvg/8ng1X5qOmck/u+5GyrtLp0D5IbfcbWONEVzY0o2zaE2h1/J
VXrdAZeDjSgv5ow9N51LzODJfeoyHSn6wEGn7EnsekgY/6/6nzv+GDmFdfx21NSI
eXF1je1ND6WyJT05cmllGD+To1xDsV/OcfxSfRksaFOGdhys0TOMlgR9SWJe11xd
qrqnoNBRW4XBUJH2TmAUfzwyhemmX6qoIICNJL9n6uHcaEGobjXcTKOdrTOvjsFa
J9YBA3cb6MXnipFx1NG1XKOLb9WQF3qlZOhZX/jxwazn10A5WP/qNawB7dsoWm85
DKCXxCAan2ih6oyVa9WNItGZPwacmCp8XWcxzRjr9lzb5Hti7vPG31eV+g5zn9sA
LrhGq/wxDrElYZU/p0fNnHdAGYu/1c6wHuTY3dCI/1NSe6w39LSkZeYb1X4F9dKt
NNcuz6IBvLfHtXGR9BR9WBLW41h2Evj+AErAl0EUEq2alEAziP8bHCAvMBWmVzac
zOXXxb4isRbOOPGJKiRZd3GhjfXMDlhhKo8nGgJGiYQHbMolPRzkGltSQu1tLdA/
TlJWvVbXgu2dM1xw7YFgNup3hQItFRgFLf1jhTtYqOMRnM/3kXSixwmiG1KwPJ24
87RLSpcVurz63zcPcAJnEnTmmsl1nZcKOhHqgW8L3E7pZkfOquLYRDyDfGmw5fMN
oqizATHdfR2c89312/68fBAHWHeXJoWRMqmuwq2NpYO+ZkmDQpJo37CBBzBsa+DE
8L6PsM34fCSmaiVQb2ULHYW5TpN8fY9HQzpyxmHT2wZSRx3ihg4tmag6kR6JJJUC
GZJa1WlfCYL40+uFJA0Pb4zhRhVfFTOOAs7snINuB3cVw/+lKLsP22vxbSHS6uoP
xkOO5NQ50Mn2CLsHFR9NpwM1EwqGjfy+2kZEG4KVJrU1h4UrIj2sjURksAJuloH2
mAon9/PBR67nabrm+bxOxjT9t4ebtvNb2ZfqTn8E9DetkwrIdD58lAgq5HeBovqd
kgFGdysXS2+CdeCb0wqf0agMXVN2fOi89+RnOyL/Go9qqhXIwXX/h33pONV1lLNS
dMBf8cGUdUmCN2Fq8euTJZiyI4DHGkYLqBJ9mRuUe5BZHP3mjXUhR7dZ93UPtweU
oDibPVIRhhC92wZZPZBppAEa71iqH5jFZfhDHeIi5K3YSz0eNLwemM/USJdt2sR+
veqCyDr+ZWLhS2HcDBXrkNT9CB3iSngVZRhdGUji3BOZdI1PMFKfbDAFblBtJAQp
bymcrI46Yjjuryjj9UHmDA==
--pragma protect end_data_block
--pragma protect digest_block
OP+5FSFaBmxKLGjERSw+j3iOVx8=
--pragma protect end_digest_block
--pragma protect end_protected
