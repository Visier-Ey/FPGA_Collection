-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
x/SeLyBDMHRpdLeTA3kGUsGNIdDB/6p8iDTNkErDSmZR0pUHm8BX7EQzIskyp4mVODG2SHWt4NZY
xBuwuiHEjOZV64nlQHh/G7+2Jpx54b2CHT65rlNJO2UelghdKzzVXEsYSeWEBfmy9XETUbBX3UMW
PUpPAlQFg0g6jHWhocyTrFsyCZf6uOAWEyZXwlCR0YukKarNy9RzpOSwNLz4rVz2CQJlfw7wk3pc
3TZujIIvuiNMfkCfydALScgACouvbpoI9DmdySIYW8v+X1uVQJlivqMzK0TKtD9/hu3wA4cSulUv
Ilc86R5fQ1+Uo4Cujd5aRYXk+4tAYVBa9TI3dw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8032)
`protect data_block
F9kUvII+k6Bv+E1lY7/0yXOCRnollqOWkzSBTDBTzcGSwWdCBhAZ2HqJSvmZ5rF/ylDHHwv+/MdH
XsjnQ0eGPlWKxexEaZNs4Q7jrOvKMMOsJ2BsAHsEkhAiBoEy9vB85Em1jBICA/mcBZb+Hqr/PjQE
Xmn1uQv35GYirJsdRfDD+jXpsOxVsxqDSLHsnzqo+mQ1tD6gORYUMubfZ/Vch94d7UiiePtWf+VG
dyPYQu8pDxi2AkQTVMzej75ntkFthU/CPtQlaPgOq4+Aj/LsSsKwZ4Pz+gicIX7kChuO784YBoQg
COHSbRlzcLpnNVb3vYUhpM7K3B5s8OVxAzT88Nt+krDb2UrY/AJtkodM6TA3nSXk4acyZU4szn+T
744Rt2dtymYbZbFC4i+3KPlpE0Qe5XXJnsVsIbRmQEPqd4uLHRIsxKrwMQN6TkB2W/ilEBo2BwLt
yKMGSNbD8l5JXZJpvMmwGGSZMuDaQRLps7vgPhFYRsLT3eqdtUXN7RoxLHMHp3buBnYRW6cj07wZ
/mKELZoEF2bwc1kUXisE4Qr7PIgYQY3/HHcallzCiaabtXkOSQzcVYGLpq6KVkzw13Gx3vzyhHGR
LwyUaA9MdjSFw20J24mnINFsxGve/uUEzmKfw3VbicpFg6I3P6R+RPjKi0AlDFciSODApfXoNGdR
K5UcB06OBjTaQ/CrQrmvjm/6Gd48KT8VuhL/ohLVO2ioG9Z94Mv+NH8FJ4uj19VmmUNFa8DRG1pT
fEr8QFNi3Z+wp6rglvkSOBvxWt9jDWVa5JR1Mw0Bu27JSMolj9gObAQfIiBVH6UT+wzdbm5ocGSf
UE9vR2qVW2pxCgl6xkUAy3zCzcASLxqgkOjs4pbn1F1YPZo0SwPapBqj/9zIdcsUWCv6qIrUYew0
Rb/aRsmMQscsrufhwgWbp6J3wyqAOWXivDjsslSdjWuqflqyT7memitQD2JIL4CSaybc0DXfGh6Q
ddD8mvNnCZEGZtsg7HvH0UPcVfSuDk4M6uvGlO06wL/K8bTgWsvqflKKvQ466Qsz0dQKdJi36Loc
M5gdDWgeGGt3kC96sy0vuaVo+V9HXprRv5modROqhz2Qkq88KRBaZ+C2hd+Rp+RCHlyPl1aqnv86
KEcjkH8VHQlidIQoUeoqyAbLu6dIuplrBaHv6Fa+2EDtNdQ79nt0F6rKHLGQB20a++JuMU98LtKr
O3iWtQXk5uV3lbPnQRO4RJhRwxZd5So6UssHaIWGaYJwpydpz4j2bKBFceuQtTexucz4OzY5FXgi
Xpd1vE2biQwRDPxKjAwDC0RXIaFidKhpNhNpjPNTX88T9+6nPbSKZxWZhB6SIUbws1EMWMr3Vo7z
++a/9ab1U27pU/dJf7bIgvxzvne9BK/7a2lvsY8Epy6GEcFc7BhpoZvLDwCtSdUDdqEw4oIOOlrn
MmC/+nmgjr/HNqMjnQn9mBYn2aoOt5m1UIsb+QIy+dqn00VrL/NzXHgXMMvgOwRkZ6FlR+INNM71
/C/kafC4GEGfZayoU5dkMj0onc+ji4qqlYo3y4d7olZ8B/hhB2e9I8pFIBQ9cQtSLlOT9Q8M/IQ0
dxJK3DpXvhpmBLhqWqRCJAGzmH85UGZ5Yt6YpafOvxv1hbtAv/XrWhcxZvo3DtezKIgJZ2f5bL3J
rz+Yv9gu1U5O/rxPAxQyi0jL9F8VY0XODf3tWPbWXsD2Yk7QqzTGcxvC3w7c4eW9Lm4VkMtfwtAj
dPtRDBTmEnxRu4HZCdBxHKA8A70H4fDCRg3ZwS3/zXULjwjfvKY7rfpysgmgcsEAjeT7cSum2Rph
s8nCAJsq5tBwS2BKUshtpFSH9bpm6IIdwDP4J5K1FALy6OCRXvPJ/f1Jq3EHW/YmqOf3ZFAGeSma
NSo/zn/JOPIKLOfDSv9mGzndsjfJK+FgugV3E+nqZkfCcdED75IsvvXQhcVMzvu/CKuaInMDHZ2S
EQViHusda61hjhfLLdLHCGpiZxWYw9HXnLjNW4FmOhpQ0h3ubArhbgNZaGRWLLJwMC0fTCq68o0p
bB3rs11UvRsU/XaDGINV+vXeCvxwhCOHWQLAgjsaciQfrQ5DaDtjUs8hUvn5kaFP5HzjoT6TimPD
W0bBKnNFND7HN4Bp/3wL9QMX1b+C0gDSM35jRXimRDrMskiAgQIYkMeZQbMhg1k+ZdIpNJngQvXc
+acm2QdItrarTXWFWlj67D0ijqEoD1ETIgENBDhLLvDudbm3gZmcfC0qBNn9J1gKBtu3/fzFJ+5c
gWrbbvJDlBEAN2EIjuztqJ4H7dQTd+yCWw3IVgnRq5JapEooh1+wkSNFvTcNPbhhYrRpD3MxDkSw
InPmB6/GousXqF0AZu7nbMpcTq28yyWJhXms+v6+y6OieeUHzg4pzj1Qu6zeuvocYvcuRJwiuJH5
lu71NSrhNeaDXYFqMIrsqLDbTv0up5ghq4sCcp3yPJjUxPqMcHRaynLMiJAO3V6ogHl1tw0EdNc7
Ddxb2Bb2K+LHKP75VaJ+97cYS7lnUFcLysClG4+geXhYckqTN4GYU4qNFXSLEGMV5tv2FdJs26FY
ai3z/WTxUwT1i2i4Nbe6sEFVbU0w6X/eO9VOdU2opQodZySS5u9Kk0qcwtSnK+D3w4H11LJQ/PW/
pj7z6W3zZwACv4ubI/DJCz1PzQqy7QvLQlRcHm8xhl2cEbGCnO+LofA/zevLq7X/ql9406m++jgQ
4ChC3iR66BMZQW+gheSNrLC2+GkrJt0nm9pAa5YMSEku4L3zDdn8om9M2wnWdYpBN1UE+QjKtMqu
CwOmvAD68G15glk73nZwV6/Bs/5i1NsDyb4uVmb6EUkAIcUrssdTneR+D4ErnD6LsLkX1Z6IU8iv
3GBnQg2DE+TQchpuoLZNiWtIJPXqsp7RrsHgH4sWuNMK/ZGohdilCUG/mXrwPvl4gAahzi5Ume3f
lfmeEWMgS1ZkpVLFBPnjZMd48QW5c2T7Fy6EqusbDOifwwfOmnYc0qIvoBUipXBnKIYx8OJz/9H5
MjCxgSwNPpdxLH4hEEk09F7Jp3MwMRVR9GRv6tGsLTGQoUW5n4eINQ5hJN/63uGRA7ofNxMDZmSq
k6+YufOKmxlJwk9TleYygofJxb+8Td4qgL3hHDZnTWE0InmkgddOcOHcVnrp7tOW7h0wdH6Q4Lvn
t0gHzpg8eSNNyMluOU8JjtcfoGDj14US5yFymdPhKuc9Sxo1/13keliKOtB1/c4yT0af42Du64fM
zguvTwjv9RkGZjO59R8MGmtt8TCZARp/e84pyqyde+8zCley2lF9yUqTqZMWNGCsA1GEeXK4ZNxJ
m5HTQq0dkG4Z11abQbyA6Cebg+7JDmuk4yzW2HMXy+cOTnWUxdVsN0w1xYPXJCR+R7r0xML2bXlP
4VxK3gxwkXNP1+YrxaOWNEJbVxlnWkSK/zxKg4SN3w7FxGS/WZHfFC7cL42gJsb8SD870+Ca0p/a
rGL68wcpSeBppoGt0KBzgY73t/gW+cuNVWoBgZZVoXQ9R5YlhV6qjAZvUp7VPKIVjegBW4PgSrNw
iNgMlbCeh9zg298n7i8+kW5y6eMdRBQ3HonpxNn8bOnPpJMJH/slIeIrkkR/efyg3kWLwhsE6iTP
NEBs9s3V9b2XdYTMe4R+vMYlFBhNN+H08vyyIpt33Bmq7Mj8jmTTlP7BKo9sBfDSUyCgXTt90F3v
ZG5cHZ04kpoKwOyUcf7g+Gw8CV3y5CV/3e/7yzvYna4UbbCS3Y3es9IPJ7K/FUgDnChp4Nct9uiI
iItSVn0Q7GTcOFE1H9Bh4tiWqAh/4Gg7J74CEpU3caxj2SOwNB5Zs5IGojXO2ijnDvsBnnPiXCDA
bk7jHNZ+JEO3wA+XGTRYenSGVupywRkry3RZtmA6i05Z6aK+PU3n0x4dJpaxCJ2JhPm7OBoZnUKm
FTzybdKFGFDnss9mKsQWqW6pY1ITAooWfPiuU0WGHfwZGLWbmdFBZzjw3pSPEtcl5ayF3j+PuXHK
ssIhxYvqY9gXKOJAM8CoXpgonnuzOo7h/WMhczxns4mKiGNQsaAeuuqJV6oANcoVDWz4DWQNPRLo
LQrMIyADNQHIgm6NcKKGS/Et8uPvZ8CaJpAuYyZyOFil+BzQDsZd9fOP4JnwTrbZJKkOjdEYSbQL
SOKEMo9wB9bxeeHjpVxQ9lzEkFmaWh7GITGq+0p0CMFUn+Y7AfD6byouyHDb56eZpyTlfiQj0ztq
0M++v1vrUDlyZIQmNmCYyPDALDxkiyo1ru9QMRRmSoPScVqW6QCZpNHnqlC24JbDpKrCNPiGZqfr
0Ieq7xaC1N+XjeP75M1T31vA+liiVd2Uu+8NfVs9vauy5p0BQysPh138F/Yx51BNhdIcdH7r/QHI
I4qJnscl2j3am/Hee7pNed21ejmbDCiJfhROzlK2zu2nkEIv5lsUcp8o7PXAn4nVeN4OKREnicYh
DvpWoq+pJ0LtTX9ygyRJpe/sCWlGgBbAbny+Q7/BAHJO8UUyBuDAEazI4v7SF2an1q2Me9yJkcdL
QedGUyQn+8FxzBZGSNU+HQnxsgB8kCPSe6rG+NVy6xXIVTwowTvcWNBRR1KSELxqINioLL0viV+b
ap2S60Ok3AREKVEmsT4tP5C+UfMmqCaAt5rugrbFKLYDvNCaylRo4qq6Xik2E2I95p2np9k7S1z5
N9U7te0bWxLbbJsrSXnPgDthSvtUQIDokwaMwfr3kYUepdTjddzr4gOKXQQ5j2IxuRTsTecGpQBJ
vbHBuQmjv3vP760B/SFFEyO92RzDSLJgoDhrv9il96smIexajraJnvk3MN21HjxxG/M4dijWESB0
QYmak44PU+jrk3bCMAO/zhzWhahE1ja+Y4SfcUEBP2aAD8NhNBxYoyXh1Ky3sSCz7LIAMM22P81Z
TyP7EMBWezO7ViToLEncnuUR2OzOZ1wVYsKlTHa/PkJEmCH5EE0TRCEwKrq/AjsLJGr3m7C3h5gz
BmHsonDlPsA0HkRA8vpr5OM9f6/wA7P6gq4Kth2adIt2CVgD1JHLIBErT/PEKUkQxSP02QoFx9OT
ppLJtyWZruNB5HwfTQcmR3rkB/0wTKe6QAD4qYG8AmDwyDkWz+Q1fPxwCFLZdL74DtpTXTmrCu5u
wZnRLzJ0egkA7IIx6pz8TEsGFGhsqU/UWUhMq5hF4Yp3jzTXAxQq7jz4FGMm0QUlKLHdYTN830XB
V8qmJ49qcqs1/LA5qUA5z25WOjVc/q0DXs8K+oKvzvT0gDLxNHQwJAEqvHU3Y5Lg+mq2++QVZd7+
Q9PEBBvydFuTWfo3L+ZDVfqJibK0JAB5NfupXvKy9sZR5LYh94nh0YNvye+HX83J5Z9jDVQf/oIK
/Tvrzv81rBgCsmlO4BSva2DsXrrehE1vznGJTCQmXYhBDcXH4foaIzmrT/AiTY/WEIERMKS3PPUj
qPobui0b9tGJJGO3QVWMl0/xOmBZmpN7BUgbNibZduEXclVQZs8BnVEc9jEemlCDYiWi+yPM0leM
GxpPaX8CzPNLCeSsM2bbA2ZqfzhZRVGACPXeYB0Y57S3SD1hmOQcFIvEgT07GKOvPSR0NNGghtLt
PEk3/MMH6wMeCAlbLV1GM64W1aeov2JcjYHZWOYYDxygBgZxAPceF23f8uLTtPhflUwlhCplfyyE
Mduw9wuOzLsLL3w+bfi92IUySCY2kaJHJ4xpehIAYooNiHGAg1V96StrD1aK/E76eqRkp0t3xgDq
RUKn0+5V1rrYC/1SE8j+1GnEpWZ6MlnaHtfgjPT0p0jRFzYqO1kqDHT5f7M+cnRJPIl2xfPrOXXV
BsNX8jeToeHy47k6eufb+LAG7/AC+4ec2god3BKay1hoLx/VWUfCh0PmhCLbk4C9ZSMPir7I6+HF
/N+TFnJR0xGKqu9Vck6GRR+uRY7rZfIUwMBN+cy2fP5QMsiYJpALZMQ1mn0PM0jHBsD81CjiX+13
GRCJk2EcCgHL31H9SL/FHN6xJdwBbi+oKsj0eZibvfoEttTsXdcz53/fBqjEkfXNuGULyofCD5Ab
PXB4gQwXNgLO1XVlN/8kFrGulVRY7pAN73srXUAerq7tvc6x7egSa4wlJDEbGkRfm9BpIdiCuDFB
lVua6Y1568tfh9R8XvTh9kvO3TM/Zuyb9aa9py0VEMy5SvOWARcv+IG9n6B3YeIYAQd8ighl26sn
rqNCMMAX4W7AS6CeWxPphdJoXxvoZrXR5FOoIKC9F9huVsdWn5qoYE6v9OvEj1qfJeP6o5pNxFcY
uYYzmWMfXq14Fq4seGe+YNbOQkaDo3fpkqW//7g0PHXNc/PWpCmL9fx57VNQCENNVzbnmOguSPHW
/w7Q/jDZX/wgwePSxwUYxEr/b4gVE3UGc2EreyPbGteW4BOlh9VkuxyDkGUFUznaSoHAf/wBL5w8
koX7zbfgrf71otIb2URNjUeoPn1sCPo0kVZENVsuzSfwf24S5WfV4zH+psCyK3rPAH8RYB1vhZMo
LEY+X1DM4PKSwxkJG8y6ewxnwU0FEmWUFT3kf+ZWq7X+jpijtroVC2GqQNkDbXz5QRIAl97zT9oc
vqimAHHRGlnkORecWn19OKYcH/l7a3kll2tdxIH6+8aDgWDQi+8YqkBQvQEKPEcF6CSyyv56khgf
9+k+2CEg0uXHhSoK5cUobLQVX2OxRJ3y5dVKtGHnbBd6wEkUU8R6c/6NtQEEewMNJ9z05XWh+1rX
UOOpMOYPnDi/wmFX5lDecEwUUqEckx/oTUq7UhyYJLcbmQPYcqXpIEs3ii+2utI/KPjdRt8NYQEf
RxN5e0kjIfD7P4WqCugUkXOdgp/eHZpui71L5uGuiK1wwLxq8w+Yl3Zdqy8eZUqgbInFDUY9A3OR
rpvKqeb70aMnsg2KyyTfeDEIzkLcEzIrRjLV+ymGYF/ad5vVYa5mYgezl1DLk2nyYpBK8LCSrdCc
0qnODEl/DfZY3ENPgAJbaF19ZidI4yapUP/KwaVfk5r0bxLWEpaoRwedxbzm9K4mn7dehLvxdjRc
5yl6XS1LvWPX0GJ1jKFuK4HgLpxLCxy4Ab6gOzUjGjtYLqbyl8Nfg6Js7wN8xcN+YiWoKebSMl6a
ogJs2NzFfcadoXRrVABu+bIQAm1h1Ncp2sziMyiLuaENWeB/OjB5DwulBwqESLJ/BwDrJcjBpAWG
62qnllFxw0mjwvCJyikSc9L+omhLJ6HTmLeBQCBk5icvmHR08TVCorqspUW6Q/0yR8gAZuMWL1jV
bW/W53pPHPxIZ1E1Jx3Sl7JwTY6TgfVfs1v8cfAxq0bmG+wFjeTeiXMBhZoI3ZzMjdsMC07F62Jd
cicVecDQGfyjrE9AIUFx9o/FyS3ujVUbPbeCducB5yByabhYk6hWqowlhhD/NnDLyyM+xnUk4M7r
Z4dJZCd6zrrNjavZrELXOsRMKYjyxkHYyRsKLGvWM4wzRqt97SL/87oSeQvbgio1r5EqX2y3nJMI
ZzkUHMrflvxyiA5TbcU9DaErboTw2MM2PLeuzndwi5NAkaSXF09ZLbTuEu3bTExz8eM70/mDuA4d
PHDCZ6KtKTOhyMpYYqzGWC5bWKITYrSoGcy0oZ+XdBBDKvbawALa4BY8rMKezJS7kx3E+MvQDD7Z
SA7sgoSxHX4n4dmUmkgGM+nuARx/nzgSV1pTmsOMe8fxM9f7IDa4EhBjm0F7H7BgRky6HhYY0I/5
7NbofNiKHz49otaMrLEKb3meiYQhjdGBuFPJl0LMJmuxUylCFaEoknupb65jmRoL63YsyDEA1Hug
/gabPmlVxeoghRWaTiUKUJc39U+32zkKbkzlZ4QV3CyVRZa5vKkzveGuRvUjIz0M1u7lya+Ld2Ck
ANERSZd/YBd0jiNnn6scyv519yAlh2NYcbIPtw4Z+Wm73Zv9rxlBkJurArmwvxSiMbyfRLqkJp72
Jy35BIozr57YBqOObV7gSEfHrTmG7vr0B3nWwF/69UGTKMybQZ8rdhZHnxbhnz9SfK5CXyZasPkd
xtuNQo+0lIfVE7nuXM4BltIHpHjHXjoJt1025cLUySe62GkUElouBxsRFrfFRbROdVuZyfIz/09c
SjOSEzXAs/BD4bkGo/c/OQB/YUC7nRPP0amyzkUVvJann9PCzKH0t5Xj117d+3KWAyBQZJM2+sGg
eb+flCMKjRTLa/jZCv/JPhzjHt8uXlTc1NaSdSsmiO3vYUOPN5EvJg49CSDJXj9/Z/+Odg02wVHx
KYvI6y63zgfnadesX2pX5lDD+XduGfgWXOu9fM4T/2kD2mB8xCZF7vqdOHatLbe8dUhvaedRAHg7
wglCDkIRxu1oB9/ce5YBdFNtFR7usV39Xgm4wKNTzrN5c/axnD43uP7zidyKgVQ6Iim2ACyOo5e/
Xpjxp9TeFiJwqp7om2SUabWHPDQVKQ1fyiOewM/lyXoutZ+Zc+5zVSOy8ZjiXoGIzkutMbvY6lBH
xJhJRnKtWqZaoK7v27X2vhV5PZwR2zINCLO+uUl8hCY7DGFBE/TCQrx5CYrgHuA0acN109y0Dt/d
VUZmzAAFmwY/eCLlNzBBj/7CtTbK5cHFC4umbjHOr90UdFBhu0PK8FeoSY+DLMw9mtusDOud44cV
3CWsih+uU/+j3xv5uJvWCvJ1BNETMtqQRc6+0HVgc6/cbv7HT8UOfAQEPbaUxOmyztD45QtGLyJL
iVmlFWgX59i49XsIsjvsMb30n+3g//+rsZoApMOXM1C3XsZz2TTigxLivssKhngCCAAZwZ/4KQN6
NmUVGUCPv2EV8dCFgE25/Ksgi1rzalOJUFW/lp8rmRH9xRHtObhnj3BsaC+TIBlnJkyLCHbWU5Ex
1Rtw8huHzH5IOfVWZCiCzTJyLWuAsjjxS97eYOcd1/MJtc3lx2lHryUTfAnriy7lC57MX2K8kDge
TFTzBBv43biYt/64wD3RE8qogblCyhaEk1U9zVrWmP6+QsdjzGhC6Q09JF7lNtKRb8v2Ds8V/ja/
fyft/NtPGbW5WtfKuD9BDrOVgv+uOMXA37LfM40HKzGWJfgfFsw0LhuyZHbedIQF3BXI/tszUyxY
4FWr+oqOtkl+CRdvuLxfALH+H55ySivaEpLcM3Pw3yicSGM3RyeBuPuAyXTybGLWGcFURl5dgd5b
TFhfli0KGW6D+yW2MQPUs6lUxMMoaTkza9KPSfMiBehVzF69c8kMNFr5vETXn2wo9mSeSIdXE8z3
Xm+tNnUP+lyLUIjyb2ITp+d40RfFnlOu51HBS8dmXEM3myAKcfHCE41HnrJgw5ICX3aP25cMH3kh
4uTI7k1+IQlRh1s08VEt4SUtH6KjzOdEEvwhGaYEeNKRRhscbFiyojT4ByPPPGPM/HtZ7lStmIq0
nOFIXbvw06W4lRrh6p5XG5ksyl48SHYlvi35yfkho2Oaj2ZXXeAn2pjOTiyzKROny+OgbcufwdJq
VHL7bweh/t+EInUrRtQu++ayShvPqAgrQQ3ZqAkqOZVbNT1frv8X9R8Ox3bUw6DEz2I+FJ+TRMbX
Imr5ulcmqLpyAYKIeG0Qlv5oWmWgC/rmlGaOlz3sY/9mmy/FVElgFVu75tdFtqvyb/snmMPZRJEd
UKnfsyPhx1VVQqtZzdni/C1D+HFFCJajuGszl4mvKp3+h8A0eO2hj6aUwF7j//yJW/S/jAxS3wSj
g9b7DRfHm5vHwk7v4Dqfmzjh2kXF0/48uQJ1H/+pMxDh00E5syL28xNSXeWp2+MS/sd+0wjvRFcw
UXYdzdO5wtkaYu4B32MFI4IOI6E/+RUOGQj1k7dpZmwjPOdLeD0lhZbII813hU8Z+v6n0rNtteTw
prlkhJ77iTLJBjGQR4BLEqSmSbr/RFxaDlJV5Dk/Oq/H+jCVsguvidvYSQMdh3UnHFFFNAi6yGd4
XFFyJfCDqlUlMudmdMBHLXRJ5A4WlxBs10badMkfni+7Mytq1VCwhTu7VCJERAm0pJDYCsarb7ZK
N84DbX1FT4r9eBzDnqUMSFNfVMoXaQCu9TZMy9ks+Frru4jigqh0nhaxJBLzTp8lZXouPXn7Si/H
3eeudMCnl8PjitWja5Xjvo2NVXOjXhqJ59U56I+Q1zXSDwLfb+GMloIaXkIQ4y5SAT4YD0Amf7zs
q8349jAoG3O8uMEm03a7pOZNSQr2L8Bm7Ha8K5VGWD2hvbD2sh2g0NvXTTGiH3BugXQbUqD+Cq8I
bKdSJKJp12ZTf31KsCqi4/uLmID2wM6dykO8o+wmEAiU2jSsLBnhcapQtwb+rD7LP7NNzjAjiubm
HZfhYm8vJ1EP3nk3ZY2PCD8voRfsSBc9hmZjtkmRnH8h4GhH3WTcFt0wu+NtKcOCjz6TZu5oyaZe
yiR0yyBNtm9zAo5VLoGSMsKI0yMkrkowqcP4l9XXlmce/y3obKm9U7afOV1YaftoaCVSx+GbuAOi
8DBr4R7Wb41N0e4Nexk7uzdabSIWdfzgSWlGkmVfVnup3kSpTJo8v1o/hSZQvL88W7g1WAzawu6U
Fsk9C+uwRTeBpZuVeqSg6J8iZXdoUkwMnpi8rUUIavDsJ8gZ/UyaNWu9mpfSfqzZUuiwROSmxMAy
xOMDMT/8Qu3Ao4MEO338vksE4mgk4TZU/3ByjlQSx42fIgtpwqt5RAh8VMb1vw9kjVdPTw==
`protect end_protected
