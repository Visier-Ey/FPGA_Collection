-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
INermEPFOheHNXKRRi5riWLkNNSuNZ6VeDtK8fP2lT6q2c+c3fAyFa8kNcuoEZoG
gIZPgMOaGQUkzgBg0htepRpoj0AllaSTXkBR/91B3WdRoE6gw2qWDr7ePClYNSP4
+/h67xWNpluuSnyJPulnoIxdrk437/BiayGS+AUksRU=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 7958)

`protect DATA_BLOCK
naYpkNJFvjnxrl7O5tZJH76Gm2TR1+ezTVA4f/OdvUKJyyBPo9/+Y5fbUnoNFd0C
wbFlpoEyrIyBE208wKihKkbb4ol8nh9fImbHIjFLeTkGeBPoI1Rg/Nf4Xh6nEgnI
R8f85CoZl8Q2BE7UsF2jgCtXDUSqpEtsXGWYY97xb+W2cqO8x/kVFgZuyryJHp3y
sEzk2pjN4Eh6AtS8ZCE/4sG31+vJNKiOPOM5l+vBOv0SX5cCAuAqlRJcAYpdnuvF
QQkapsxrpryLpRDaw/WXwuRvOvHQDTfaAYdkOenkwLkyxIlX4KbapN6+AhjV0Gzv
8YyQ7X+Mfj23bgdWPeF5jlnmq4IxzB78p47zkIwEXit9C0VWIY5xllwwfCYaXa20
ga7YxTHnF3LiMi6soNIBqTkedjVVgkI3QAvWxJNUlejALlVikf1O4RhgXUHK+4wn
27cwGdxuOYEXI5JgtdDbUPr6T/d+pVx4Ctu018UW77+BKbuKqSSbJ2yf1lNrSx7k
s85FsoVXumAsK1YDTdSHZu90xc6OLg/t8j4wFJlvtj0jkwhbvY5dO+v3a4BDsUFv
6piKMOtw7b/MiAN6Ef64TcG82/1unXYgbLsz4ONnKd4IPqdQ7X7D1czQTwlezV2i
HGgXwQ11nImJbqjSj8V41LFr7+oYoZLecLrv5Oei1UbE1pSkaRwNLuQvEBScRybN
iqcQhlBn1bZz5aLdJchHMdFcOx9udc7hhoql275QA1nd4oIcl26cWyTlfwrzJCQR
7XGkCyHQp4vmG8H3UzIfl8vyUJot4w2DZtkZIVZSAWBzJMiycquXdYbIef+OBA1u
MIjTvMZFn2NFZsNcc6cqek3XcfnwA7pxclZPxZUAypp4EHWNxcG6B9zRZFLUZXna
Vc8oAk3QkpAoFnnLXJyCf4mQvWMO+AFMqARNzsprFmerdw9aCXxomMpiwqdF4Wxj
9pJvoyJ7lQXixMeO9AExD5OTQnJfNYgmTpW8dhnQcOzUqFi2WeMwCGbDC0ZtRryM
YKVZrtEBSjQAdTbM48QI5xGvrdZuCGmrfAZJWkjqJLx06LfhkJPCIleRickMPMRj
dL+8KJdaDiY3QXqDJLJUWJomoGsjDXnU+xuerfWmYoIGEl87EOaq3NkzjIkr/NcA
e+AtOoMnyZ2X0Kn8rmJjdUcKA2yEV04QptYsQK6Q9fG/qpxQtcoBnfO95iuG1weF
pV/UdL0hbmBMhFQ+ltnYe69CYJGY63xV7eWCsaSioRlw8QYMfNX5XsiehFH1voUQ
aU+xUSPB99Nhjq6qMqR+QFu0OghHTMUcUS5756D/ul5eJLmb0fcrUTBBgHwiNcbN
hVPzz4OhEI5lo5TVak9BSQiMMmE1vSfZ7OA3XedROMr1mbSXfnQdyBXeiyOx+8VJ
VXNYOi96zz8gPh+up8+CvXr5iZZGgrTO/zGIDBIEfATsn1QCIdQ71o/pER7bNxHu
q7pomgM45t0EWBDzcYgWtZRo1fLu5jnVmDfIdqs05Rgs9evflVjGFmohViYCr9R7
ljHSETcYgqv0o0tzhyuEfbQM301DJjrozeSS5NwrqSko0jsUxyYqJU59H9GQAN5h
EuAKHbDE0nkuTHfemnakjuv/1GBeJvIFGKg7zc0hx9OBBDTW1iqXwgQM34WDQKM2
goBlztIF3ZOQtpyYpYCo8x2kg8FReHUHsTi1Pu0E7IHUbmzyiyIBwphfmmfeIHvE
znrYVSYQ+K9rznzboA88KhE3fAIqTplCN1fDWdwPXcA1vh3X2h4PtZRAvS7fgit9
V7xGyXhvV2b2FafXcrvtFwwGQf3SjaKv7F0rHn7XMVjGjrug3nA/aLrbm8exwOCu
rpycRf0MSQpLece74PsKHBvngbqUNHKaP0CUJkNIcUCpUBqY3glA5FkpYppjszRD
fBVmMHEIdlnntw9aR4fmJ5eGAJXEdm/RjFkyXC8EB43TTccFOCrS4jufPM/Bd0MN
noZ4GqwIG5cLhCGkPvtn43PneGThYUUM0Ek9+E9NPEzQAKDAo20krvPp17+VQZse
+wYWBNbM5M/6EpqdI9Q+RqWI1xnL6IqTKU/7GWbiFvCStRAvMnQkW05FxcZbxOUQ
zxv1bZrre4uIQ0lOtXIHZO0LrNkNuxjbHcPAsgeiUmlHQw1EK99mTUz/sQL2yLbd
POXiIMjJ4NyxCgpGPmsq3Okv60U8SDinRAInwIJdZ4NEysRaBnGJnIj1lTHA3keO
Ysy1AO2tUt0CR7k0l3KGK9QxoGB8zHr3Ca+b7O8PaHzRmVKVLlS+ZysRN9eAV4c+
rxMkT8NPLHOTGeNR0WFM03wbaqTnpCp7AoNgl7hwDVJLeEtztwkpWoyOw1L3r8Ji
0d9jrVvm8kCzMTDOxPR7PHosFsLsnuESatq67UKdJKvrq8HKRBurgrsnO9esZfuk
D3kh/M6NpINtpgHMtd3SUlI5vv8fpi7DoBkza6QUEvckyF/lv3zVPHyuKNiOq7tl
Jq44MGv3N9tZznglitCj2SE1PFzbWHK4LgxZlbXQKki4IuGCvVXCm+ToSlvPGEfJ
JWVBTUse3qB101zdHDSCXCTCQg9cM5OQmTYTErGsJCIKGp4Z8/hTl/205Lkg2vO0
Ofzv4XLs+eK7/NrnhmI9RurIBSE0mBpYb37x0ydb3VKfTBP4rVJqk4XfkOY34XVs
3DOoqvGyZwzbqCi+32GEjbF4R/6f/N3W16qLu0zdfc1LUJm3fTiQTNrn8DSB39Wj
T48tSFbLUr3wEwy3L9VH2foN02B/MKJyzyqyAzekFCPPPPMKYWk0A5XJgUUOiAy1
SJV1qmHG+abE6iSOx5VDEk335lXodysiC6IPIKAlidh8IcC6wJ9bOVEQEZDxTsqY
MHjZTXn8X/mifzmzNpQJBpc0jYuyovD2grOvtXYudTpkq1Cpo5G0yjSSY/zpPLrj
9we8uQIPnBsY7q93xx+GHQIXZyTVEE7z0Rh/IHzaThK36xYyGJGZ/e8khx5Uvm5p
7FdmOTqePQGq9sQk4qXEoDVLS3vabLLY+CD6IK9VlNBvXBor3bgHiBG88St/B/kE
SK9sDg5SNRtmqzraikOinO5aGI2hi6tXPhYDo+ZU+Fb+Xx2WNLsOwv0I1V/D6XOC
OcdrlMKjMOB4eVf5SiBm0JiIZmKBhdYB8hUoRaPffx8ovUrP4CnKh3kIl59RU1ti
NtZF2Ld511HlJ7AJgYpAbk8U469deRFSvx3DlhAygVKwF3HSC95l1hMfO9VxwTKN
iLnUYXTbsYkEf4qvCeLLJZNDC+UfY6UGYBoryt+kZUMO4KZiU7pIv93oRHDQUxp3
gfnQXuAbQLEUKee7Kla7HSxw8+63LZYk469pjjFiexf2++REEiJdxAJjXKh+K1sq
8CEXVRTOd74dtbu7ReW5+6QvWIjwqXXG7ilA2Fg6Sh8QbkBAiGX5tafa3oStxD/f
Ww6uM4AaWrte1phpA0EDVN+01BGrfKKgD9FQZfezsRItHj0YEu7yKFDXsUC0Ch84
qwbaIxaAP4NGwU+P5e105JTdIDwC/x159roocFw4BFxEZWWwsEMNosJl+rxaQHzn
rHU4gZKgKVSAWMHX+m1ZKQOSH1U8p3sgW2m2k59ApNlLIqMnxwmM1D8D1LnUTcfc
ChP8kbyv4Mx85qsuHFogwukZfFGvyBs8Fd8/glS9s6nJdQto4c94vbnFWUH2HNQV
UhCYQsZ1gaZmCiU2jKGzewNIL0Gy0DIo5f0CsTC02SblOfsNEBUkQzcF0YFVe5R1
2aZTcIWwbiIbR/qR20cAUDd8yBUTov4APEDpig+cKaK6q2X620kuisWd52rbpBAU
6lE1vS7UmVXfEhsQcW+L8kte1udeWJ6RUN9oyMHh+KUenr8M/SZzYEOdFjtkhO/J
Wg8QYSWYn86ZJQDMxqXeolpkKtgq/DR1q8Izml2Kma60NVRY+SQpk02Bxmx7tXxh
L5mSJOKFBY77La+nRaeSSG7RlKRC7AEuHO07P3Q8uBjbtG4Cgzpfe1WQsFu+60px
n2wtVEYiiZncqJSeqeqqZM7E/gu6voECU3tb4wLn0hf8LM5t66s+1GUZCvga2mHp
160O+vQv0qGdqngQN73Zs4esAgohiVc4cRwrUu0xzwlju5qYkVyUT4xBOsCcKnVC
DcMu/jQQU3CHH+udPpKIsaMIIcR7y+xZvMOWnRGhoQTogRRTE4TSr07zFKpgv8gw
FlNbEijrFsLXa4H5te3W4NPgzHLhIMK5omBGAewn4d5LfW09Ik3M5e8FplrdaT/Y
mknyaoWv2V85onRots4tuJqtlfNPmn68tShI3WHkT+TX4iwnUzFZ/ILDv0PV9k0Q
8f0rNume6XGxz5kSeQb2G2MAIPGRov/Jia3SIQJlH+YonFpYDup5+MuHs/XmQsPC
f5Iy4UeQrGUOvNZ8BtyZppG+KAesz/G9TcyxBTJODEnWKzJF50poK/O60oQHmTGK
V8OJU+zdKZPrPco/ZDF0293rdgK3hAm3EIxyNezGfA8fMrjygt6ScQrijHTVtvGT
Weo0v2b/vXi94nzVQXgwcCHaSOCR55vfqEETKB2K4y4BlTIrQ6VbzHW7t4VZQDte
EonZ5Hp155lb4sQL5DMaRG7QwaeEtOyVHF1WHK/aC9or1iHA156l4SKBYnn17FoE
RT3byLKZ2AYMFpv572oB15CUyqBoVar27Bla7U4wvLwpkhagVho1HOvZgpMVGjYT
6lkAH1cmu9mcrzcoiqO1oCCujwCL9cI11JWhGXUengc3UxgacaTdcD7pR2qZj3Pn
kswk2A5GujuuEPIrJFc6z33HhQNmg814+otHEaHkRQYuzPk64orT/BAw+Yg+m+rL
/04hiHCdoCVS5cp3UIceNn3kkdcU+smHyp1jvUprBGMuy3TFsCGlwj4bXP8uaNCG
NcHEMeznmQtjSa4ybxuYIZyY2lUjty7eKkwdYuo6kHCMxGfdLLrnt+LyMFLLlpVZ
Y8rAW0d8p9xv7YkUyOxkd73Zoi9xPMFKiV+qkx32Te9EPZfeaWRrF5DUqEfcv7vl
02TItXzmczSvoNirO5XZsb+DJek6HyAW+EOJFBE4ABWLDcGTwX+b9XhQ9YGAfmzG
ZDJeqYd/eJllIpsIav7rkth0QWm38A9F0HmmVsXgbXprfZ4tw1kbmUDXbS4gZR2E
WCJtC3jSWILdhEps++OiY+8vnargXXApIq5pSzpS1tluKFyRi7sDbpYmz70yskwA
HJqvKdCAT9eSjqTDANviHAhUU0YbQa+bcFuCJvBGJaqaivg0bqGcduCPmHRMexQU
zjk341txxkR96tCvf6G8u58iuRSgSiFpX/ofRXt+f/xTarVFPKKPfPZX951eInDV
drWoiM86z9HnhUA0tWJGHbdtMffT5hLqbOf4tQnCbMA9pMxNc8G05u6PdZS9nctw
8ENVMI1sQ7M4LbawJtvGKMF3tnKz+uOyjzDRoJxXRPkLKoZnBZy6zCGO/CQol3vj
Y8UcgAZruHsd9nT1lh9cXKdMWMlTmZa3FJe5AoT4RO2bvADBVdh9k9WpINyjSCpI
j60UOF8ZrIPBG4IHpk39Wn6L/iYBBF2xEUeG+oq6XiTetHBnE3BnQ8BI8hXy7b7d
LJu8YLmENnKiWogLhR2k13uBECiVnDGG0hNs2lo1lRd6UZ8wmWXnk+fb8hIDpLNc
7SLm8ucXH+G2LCLXOYqLFtf6ONtVmxRr+e68ue5sz0cbERZulPMpAa/hsdghgf7F
4zP3gQS4FcPGgzF4+5mPT7gkEeIw2z9AF2x9txZ8MpKZ7r/zwpXsyM3Zamx/2UM1
lR7uHlD+2TIfLbBRDPkD6kY7BTCZSCnrbXR+QxKdYNd5rtJLWfKvKSrNpQf0FnjG
1s0Ohs732FE3rCtvM73c9ChqCmsaTPDE/j4otvTVsXurCa7vNhHYEcxfskEaYVj2
juUUwf1r2W74F9xUY/dE3qo5ooSv3T2GyyCy1LaJnXbC/VGr49RfpVR1ovjul9JP
9CvHmF+D2O+HnisVY5/+Zl0U01gymQRshYYt9Zn+ToxEcCGQIIWkt02vx4Mng1Vm
KBQvQs0oq9g4JCfkkJUrSNJ8mxej633ByJSFrShbwNA80fbY5rFP44lsv1kpbqOT
BA4CkX+eyN8eNVpakJDI35qCMBOmz5LPoV0lRX6BdpyKrr+KpjX2c9P/HbHRCZ8E
HCmue8G/cU71YXQ4L7BIfmUrVjnJvs3JxFQZUtNN1RjdJ+l2P+XrwHLzPDiw1j6O
l1dT+YX5RyPMf/sFh3fE7IJfNHTIvpuEvY+KGDps7qGdoHI/+0NHHEAgCTNBly1r
kXzxC9NHhJvNL+zwxHhBbwdIV6xQbdzBfYnU88m9zwpbRT+e39T+ZSLmMd/Qz/I/
kbKzkApV+jZmZJOpUrs3HY9fWlKJ0CLEi8O0TORKdHTFOXFfCyQREfcy7Tud0gp6
06jjyLGtCf3O+Tzf9rERuys9YOnoh2a/VSUGgMCwpzMWzzKWan/sCGil204Rk1oT
bPAOYD9lUhzKvyKeR6at6OryvLykAoXA5r+fpznwygwvIwDLR0k9DXkc/RhgGD5p
WFMMjRSvNszIYjQhyC1m7CKfFpd5PqDViS4JKf8NZd8F9W6SXX7s91iqmfLEnv//
CO+ypj/VNywweaHGRZr0u8LuxNtJbf0jvBREJ+KXhbeIaDtIsnvycA1LoHEwyBOS
sCxfCQC+TcCSfHTc55gMzCbKSN3qkue/2LzMJscDRVnzksQmOo2GV+tQS5b/rvTv
mcLbTKMZHAkOioAK2v1+hEhh0Ui2J32xXFflfBF73zHiyqupXK8T9XDGvq2xCENq
1sn4XIRGCCnCjVdO0s0cNMLL3S2U6eg8iOwOdk0I4ahIvWPJcCgpLm8pMRg6+/71
IVDB8lf8Ii+NWhNc1scCzgNtSlJsJLZ1ZotQ/l18sUiyDcHllhUJnLSpcPXcySUf
uMxI0pgturVq0/RUG9gFutp8ZASLL4yPr+MegFTlCvssSyr+kLpZxG56wAsdMdU6
S1DceiczMem8qH9ZsdZqJntcZRxJ6Zuh4QPI/pEo3mNZQgVH1ZqGNX823rHce01x
9yYtf8XuM+h0upEbiqQcuvD1m5JOVErdO4bK0BipsyhZCvZjFck1OaJ2/7DytswY
eqd62nUhyO1t5xfgg+NC7CKSAEhBPZfqtTC3bZv0J5GAG/c7XwOcIvXlUOpg2iG4
KwhtBYl63Lj51KgYWQBfRSQISgUNFcTkHIY8fV0ZYruptXSIvaG8l+X1Fd3BGtel
KbTprbSdzsCvmIKC5D66h2xIH0tu95w1+85Y6SQSJiy5k4DIRHXmiJrjULXBw2EA
cLVM9LCu5o/7lvAyr1c+bvhFTlr1lSu2GCUFiUfyv0ZkjRfFKfuCEB8X/Xl3yDZL
NMbidvCPlDbgLxhwzmTpGRPaGchYph0CFlWZCQ/R/VGBvQvjnleV/EoSMbKJ1c1i
cnKOyFiI3gp1+W21NVHGGEUzonEpRA/qEou8zBY0Y6qhjblq/5+Ix1P0F8c6DuuS
OCzyB3AbwKjKoserQDxYPb1BosCwSQRJqdyAKX+jtw6La1Q4IWORyPio6J7xQk3S
bF+LX3DL1ny2A6QeAh404R8RcdDKwJD8g05Em7RkIz7MN4rQqTNB+qJEwhRaQwBP
1Mj2qtXyEc9b9NuP9HP0JlJ7Aqh8kDSZ0dFKqdsZVn0k7dU6Kvjw1XiSjhHO2/Wi
Wy7oNEux+b0OYGstLhMT0oqSr+4DxRtbBN+KDfQp8REagAdDfV5HRcraZlrjsZqu
E3m/CMUvFvl4eHjwnhrnXHC7gkp6A0bi0yIOfnLbeS5xdiFxzQ7yJslPFp/Euw+q
KPGGenYyxUbHodH/XA84UrbceuQHw9Dvfa1ajia0+nvs/csjGFwxh3CKQrdF2HdY
y7FmkW/wOmZfg5LhnWanQfxQfjOM+khTWz+HhN/WaKvAqGnUqKvhTWpUZGCV7fsY
+b7HTPa7m5MCNixeWU0OuZOxcFLs28plXMeNYEDjtXQAbYBXFWwLIMqIxoC0QtHy
lpuOGfzjCyT/JuQV3Gl455tB6vQnuWK/QPcBZL4OwqrLETwSfYTLyBt524L42WIm
hSe0EAzwb8dGUpEHws0WgjIcTetgZe95nONKW7XvngtxkrE0iGvDpLs3DkLPmtYQ
li/qTL9+RcdlqQCndOzJB6+2ZlW8AffhY8J3GTjnmeNquNLRNaiSFeAIFi21LL7j
pEP0kyfrxMsV3pqJTjKH0kB2d94jlHEv5/EcdbbOtutDxXXF1zymFyizPZqKGbrn
n4SYOY+WPLuzJn4IhmD4s4llvjlSKGxPSsHxTjoUo1BonqxAM7v5e8vVmGXTV2zl
sTdd6eybBd+4X1bIbvobs5HNy8TtxQJdiPUs6ugYD/RnSvWv4eSg/1S2+PhjEgg3
MhVbubJHbXiXD/EeaM2nPurS5GbjePruWb6d3z+wg2wBaCgunl2pO6+K81PlazmR
5CnSYu+dcPtYSPnZAb8jO5CQkFiwAhwC4g7R426eikQSf5FmesIZ9+tVJPateFSf
wFmh4VjwDxtnVnhuwZAPAQYmm+Si1KCRg9XFEHy+JsLK57oOaDdXVhu5SJHIRoBQ
fnE5JZ5O6KVn7Cys8bMrSDrSrOxF1B9t9L6Ek5/EnVEuOn7nMtZqtZHD9GK8jAQW
koNaRmfZ+LlFTe+uoIfM4JPxaMZogOrmnkZYC9n0HorNafllna5CkSAum03TmZmA
LOpCouXpWulgbuwor4WNkRsJQiVfWh1zOv99NiuuQI59hfAIkbWG+wcACtOkdUL8
HrAJR/mJo0UxPhRxJT8hD2bK8mp4sj9gxnmNheKQUUiyG9NqaoPK3cRrdwICX8NP
uVefEJV1NlorDiufKlXjaDYs6+LB2dG6tiupRhqSCfYJgRTQT4byXRuEzUfpoz2z
dEjb6FDz8PYzJNnQzYVcbOJTsRKDmr8blABPK03HW69khwp+inl97FlcH9a0a2Aw
nSjQe/fs/oEda7M0DimyOA9OfMOgFwS4cymjBTb/0x41vphc5ZhLccgjHaxxOVkt
khAbBKjk76yMgN+CJqzpPH5VfGdcecZOlOKcqlnfvmyDsHJQirgoX+tA1n+46v4g
3LiA1jm0QhsOb8PG+HqHdLc+DsfNICmlvHD12tDr+UdW+PAQ0iGSpMGZ1h4858bQ
nLeYnOG0I43Nu0aca30kO/3ljhC6QtX/xikMH02O/IMuAsjQNRwub/BFU3bO/rIK
JayfnBnQjfmZ56QvEjCDY14xlQj4GftDGaEkDvzFhtbWPm8IAcnzuebIiUPx0CQ7
ZoVPN/wR8REfk3TC4vk7xZaGN2nSOelleV4E+g1Utc4/poif7PAvbK+33vvY6ipg
7nMGOGm6nB8BaoKq06TFJGyDLIxUYttFPyddYnjaxkQAbolpP2c2/craRWFL3Y9A
nwUvg4pjOX1egkE6jmwMwUyU3wnS3wGsMiv93SRJ1az8RWqQgcn5PzWONaJfcms1
OWKEZK7SKPeVv7Iu/P64bsVucbVldVwFJRGU8K3/set+u8jzKiFffRkHkejcopGK
vPXb8d2+nG/ugUJbIVKcyiCj0vQZO2PjFyacOe/Oc9AGtp+FK01/HHf35TYtZbe8
rOg5uYhc3iUuK0G4UtEhS7Pp6wHt71rzkKBZkIK2JOwpxyJlIbdvKwcSOtmdpzic
DcD5+PCSeDwYsQSRqXZ4+AP0rbADmO9lGfRp5bVZBuLn0GJG6v5AwFTK1768g1uu
/fp4i+vJg8Myxq1qWoYIKB4mK+duIaYWxUMaHgTL68k1N84bhCwJJVzCM6+UTygA
GpoBgGwl3GxeNpfRGhPjXP6+bRLUr/PoQmKckO5YoNkt628H1T4WA0vLYaemCtNw
SSr+gvLMFmYTtBqi7Swi3h/o23Ueq64PFLwf8r7Otg+vFjPim483hkb9qF06qS0v
79OwGyP+FqMLOUZ4KipbDPOUiY7+iK3Lxai3vWd7l3JZkxy9criM9wpXEsqPTwHB
MCmPMn9fstOQB07aYXMozjW4T+1crWPC9JsLzz4qGh7Mja+u+VnVME2+xA0nWqqY
vRYa6g14GoSmOrIYytVfroiYJvyAz+cBrgr+f0PisT6yGmx2z/cWIhoM6lynHZl8
VESUUe11tSsNSE77bZ2U6E/z6AU6apmztC4w6ga6viroa0WRSFzgfjS496tG6TfJ
FLAlKOn1Np4/8pyDV4zvRr3xpWKJAvgeF1K3jCnS0lSGSDfYqfTBzYCB+F4wKkRO
hlH3xxuPPkMlzDWLGqOTPOAN4eclsJo+RgGp9rgMVVDD01TRVjc537+37GkoiOmj
S9/ICY694OPoC24MEqCRFP67ZayOit+z85tMu9OWEADUq2eruKecUd+pFxg7nhnj
RdE/YC5X9+5KDG+F47Vxk2hWU8y2ru21pezO92zRqSDzhAuKCawGWQ62c1IQIgn3
CHOOfITpbUGt0KLKJJ9Ne8GuSdvTSIZRXz1TWa8dzLxKehfWU6MWmnY/6gKOteDc
0CzQLYK4gzVW8nUed8R6lcNzWgRxLfPtfLQfwQUIwCBibWD4HI/vSqYMCfwolm6F
KYrpESRxWev8GqLJfpDeXA==
`protect END_PROTECTED