-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "N-2017.12-SP2-4 -- Oct 23, 2018"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
j7VgGe4fwVhi6TcrwPQQmlpuFJ++Y+Puq/7WUpTg+K39EOf6xDfcXH7QyHbyu07I
uGrpqZ5dbqgCCxxKt1zh2ucAEKjusCCdFh0J9PaVnArvW/012KvPOKWGbSHTMS7N
LzzhasYD7fRJdeinpJh4atwfqInmrgeFFlj2Ku6MK4I=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 22640)
`protect data_block
jQfxDYmEwgg3owNmGDv2wTvNM9cS6p8kZmnYihkEis3XA2WbCNG2xDAuhUDAa8mx
T9Qr+6cH/dOVXkfdNYsM/VtlhAXQZBFzpUvoeGlnSm2rufXjGuoJ0r7pKRKajOMg
ySqWyMJSUvEdnMbA5ok3WPMrbVWU9cLlAZvGNoYABMtwbXtrqauHpHkZ+pKclk0e
PrdXuIBBmSjLjZo2A7Ty2fKy+S27KpNnSH0WP87C2TmspVK+t+GUIagoLojELETB
FE3YJ+Sunju+8XzlUH/pkIHKka2lFdvBXhnatFSCG3V67qtuu8tZvyhmnPAoHr/S
DsdNXOE41f00P+8P7DSsIoabVQ8hoLBv5zF1Y0F+rWiL4j1dsLPg8/krZtir70iE
FuNEYo+TOXAkQutsmqOvco7IYqN1c9LQzBPdjf2cLpFeou4QPTBYSZN1envn9222
B0sOJWLU3B2Jehrby4dkWjISQfBZmH581+yfxARaq0Ov36KTNPPJ7x7RFzCWbwMz
U+DxkY6ch3rJStDE+PY1ZRAiOiGC3nft8TyGxD9zKLGgKyEggSJQOPx+wrzNEtWM
RZtqkINBzDemPpHS0YonaVTrUroO4fIshbzwnjJVqJinOxluEQ91AnvbYzuTHXd2
FHcvQVGKU/UnDw4cwbtkrhMDiA+rBB8aUx2ECt6HvUvd87zFcuoV5rxweq8I4Hmq
FW7EsLuwncwWTT0E9KMmCTUUahUbJ6o4/zkf2zuwOWkeheGUOzKR4xzyoddFvkzR
XHdeYBbuDxrBXcXKq15bsB/llkFEArk7+bhIxC9/5IW98OIQyfVmxyefWfLGJABP
zdMZrAL6+cg0CYwizZGFTtu285394BlNnkELkE76UPFylxF9ElzMYquqeykHFz7Q
8I3jTU6p+m7SEfW2wt+buuvOo3fvRMiH67IRKJ84d+mzDLY14G4JzPuYkL4V2l87
jzOsyIgCejub+PhvFhErlhio3osg3PS74MWana3HhhW/Ckqlzn7B2dncFd3PyeoY
E12ghWt/anfw0mpTjYORDo4O4RyGXPwZqWXcrDLj5+0rw3qxCgE9PsYptoOEenLt
3JqxQQcJEg/z4ftvBoA3SYaCxMGNglrFG3WLYUNYJ+H1EzFkRLQ7Ppk6Uru0qXyo
/mRkSoFZBGuaCJ4nqixmfiKu4cBE1z/WKuIu4GV8r7sY8zy7gNwfv+r4LjIoO23J
2tymaXJQwoP3n5virwgCAZ+fuwvf8PGQbv40OjGSUQycDr+EvWuYshR/5IAEtdD0
llIsBKJrhllKOAmUYu1umTgEvF4PvMZBpOGbtgoUJxYP1bgleY8Afe6F2qc1YOIs
qTOCFaMcIjM2E9YthEDazeUtoQ0mEGskNGC8CtQNR9dET1uqfWIV8u0Az8Uapohp
JTdFS4cq0Gws/npKRiRxBezTFDfL51Ux9RqkdxpEhiix2u9cOq5hKUrJgGzZ0r+V
rdjIe+fqvxp844YqzRkTg/m8kfvV42mlz5NOmaptmf1tTmt3aVB9as8TM0fCy6nF
9e19OFTSj0g7LGID4KCw1M/CPFGb7hMOiF/+Um4uEzfAp2BSfif6Iz2jupzdNcIR
h3IicsdwQoVnH30KXOcffy0B0vkC4ORQVBSWcQDKbgJZzvjd1zMz2dVIowLhJbvJ
73R6hY9rhEUvWBazj971BUVVwjn1lfs/ez6ynFMUapxhLvI5EoD1nHH01z1Bqn24
WwZXYd0zjnBYrNiC6vOgdF6zYcumsPyl5H7hAvR9xJBJA21PzcBlm4r0AINCIGuK
hCuHqY7xCPhczaFIh6zx1z3W1C2FAvTDqWnX87qcvxp37k9n3h2hvuqEWU0KqTMO
QfMkrsBCgBcLqy2eCaFJwmwAKnA28T/+vCWKq2fKN0LLIei3xgZuJB6hupxBss2o
WkhGG2pAgTJlDIiTMrL0Vv8060gBKGfAGvA5LTxoi5XUufg0Q+dyxPwU5LCUTdqC
xflkXA1Wlf3ObVpaqzgrWLIXWQD9KJ3EhkIqwKPumrmAAzeO8/TlI1K5kymsD1mo
w06mgglBr5WslOhztbgPf/TRC8TAGa+8uhjdGshhsHO6YQk0OGFASq6ug+yq6ShG
ar7eY5Xyo/+dx1N6HJ39hvA/Duhu7Kg5tzu1n4XJ0i/NkaZeRBo02hZBys/erhVt
0FdN9E/yFSh2D0xP66fPQ7k9isDj8pui1kDSHCc3r1nMqtOEL+xO5XT8HTyPxRqM
sBdAl8ARFsrRDe0EeXGHzm81KO7phS7pkOSuKtr3mGD7jfUoq/KIM6Bpk6AzvDHJ
jUFbK7fhpYUz9vY57hA9vyHXCWABTi3BesByfAIA0EYXiRkA7jKYcAa1G6H+gQN9
jRASJXjNwvuGN5kvB8//S8u11aSh9TDk0gdh3tRyVfAU97/sGz7Pvf5UzuZ8V+4L
00t2VLiQ6sVHt+TcglGYxpeaTnVpITCmTTReIQTv1WTgCy+RcVJVIQZRQrKwlo1A
1TlFGF25jVl6KS4Uzwu5zxkZ2+giBJb3vJvmAVvwvzccklj2CVFY3Q+xEWQVRoZf
qcHK+PtwVFvBYFwsHM211gIa5CbAm46/EOvrAfwx/Axe8O19i21iKEA9hGzeFYBu
HhZ9ARzgpDBm8Ue7uIx/WrHqG+OkHn/SsA3Sb/ldWrFPLNlSFLQp2R4dqo/NMZ0D
FnotXGxu/TywjRSiwets5sW2iEvaxGRIKOVoLU+VxkB1lYPKpzCAC9lhcRmOPCK9
ktxFSBi5oWa4Exse6HvTvHfdggmQvXNbbgOIGzPnHMzTpRR9OGZ2EgB8BNU2FtzX
+GC7bUJm5Ok7PQlkWaTEt8HelAXmkGBj/1me0lwr8PU5kOvY9k/gb0v2eWQyKs8l
+0xyZYrTbJx6RczFxnAc97sfuB/Y+ZU8XZd1eXfxDr76SKyqmf3YbaXEzkT9eW+s
8aR7dIgfzXcYYyDxVV2C71EWBL7lWJn+HAQD3iiUClk4nyP3frFKtqrm3zCb69O/
kygNXN2HOThMb+yDaLLZx2goFYbaLZ74tkznoZqldkuUwWHFmnoXgrUcGcQeSgeg
2/TPgez4ODmmlDAvZy5C8foc7en+nlMNRTl3Zvdt8IuQsFpEgtrChOr/h2bnoz8S
mjLYcjv+ALYW7gYSxwPGOHleu/03GNmiJL9EQRJh95vZoRHBgzJGQGdBRIpMab87
5BgmaCGOCTD4HeO2JqcKH/aFHluPV0UZkerrD7PExkLtwOl+MFfGczNzc/J9m/Q3
/jweZCy2eSZVpEmCZAz7UpuFlSyv8VfRypxv9ZeeGeA8w8NT5aOHUkp3SPqHdAkr
I+ZlU/w+rbhrCqEUlZsViSoMSPxgR2m1r9tfXIbBGVElg6QtTAlQiJjUoAtyNbgt
58V2WJKKsHRr1zg+qukCD3jbOyAnRrdBMMrXufD6RtdzukYJJ4n7K3Gck3URK/h5
3bMs2rEYtNzy8FjRSWUEm2oZJFgBejLKzAKk+fqFe/ZTu7bE0S5p6wHAj6kfD9Xw
eoOzyWSTCrRyjUrd0/fmftHK3NFZKwx4Q4fQ8BL4GBcQzrsEBB3o0B3b+X1buwK9
6vh9F90UZaL78GDES2zzR4iYTONf/kTA4ETHr6xPrj5Tv6HQizEhCVOncjYGLpVW
XQyV8B2DmPy9cKid4yLJKZZM0V4Gl/Sbt+NbGNVqwpHK2HUw8nBvrwaXqKHMOcY8
AJcLJIelY99H+dCVeBJVFNZG6REmhrVz1pcyKzUizul7EIZCIpcIp4ZQVdnXvcVj
oYeW0GflFjF0jNVhc7cRXfBC6SSckxxLdOkeFZMd8erURj7hB3YDzZyt62ZeR6KW
kR5qvJrU2T+M05pDYJ0MX6JBaJteY1d3cdGatlifG1rXekg1zBDUCfKGqtwObmK6
aHHdYYAAWp9r4NYFyXgofSALECes1/ZBFiuBMexbJr7gcCLeA8P9NWkQFxDUZ4G2
J0AswnMfEqaOg3/kag5cA8DvvVO9E5RTUsT7fNJrs9lImHYBnGaepUAPg/VJ1S//
/gXYDy3oL135wyTmYFIPaBufov0nIBjaQXlAMs5sJqY+7YLnLJry5afRZ2LPNa6a
3K7wRWZkTtmJ6FnzNu/keEZ4dIEHum/b+mHgLDcy0j8J3pN/qufPn5I8Gfom6OfN
ilIm91Z2WLZRSvj8OQ7PIX/5OklChkYDxqiIxEaQVUc8NTxqfuxJpsPGF+Np9q9c
JuojIUJz7wialIAbCNkCG7sGcNh6pXb1sb1E/SvMezK5KrWuizXqhoBghiB4Nn4V
SHCf6BmBnj3CiliDC9vxsJV+dO8zh2wwAXkbY0gysGRuXqq4tiNs+BunDjOKqYax
fFFG2yFIb44iBMqNrEMF/KewFX+gYlGlBad0oRlCYQkSjonaa3tXFOVMHV86XyR+
WNe1zRQo3L/isdDDURp6SjKmqHPuCFFT21lXwSaEYbtlhZwiUSo0Bj77SxLAGjcq
OSTYurgtE4qL3DGgXeFsjkLBwwxuhGjTMpcITwNYXqBuK9Tif7IPq60ZN1FHvBOS
Gly0JB9PeNzzG2UvqqvqeDvOuaiT82tgcRNSHtJK1ZTfBcxjNJqsnmBbJl7SK3Ms
Mbp0WrE+WtJoZwfPHnGvYqs7l8hCF+R//+7CX7cQtFWwpPLsSLDqC6BFdnN8BXGa
jC11gVT9nHIyxR8yBQGKfCUKhoHAWyq1JtSi+txncMZ+7pk0nel1WeYVpOH0lGJg
tfo8XA0fszw7eEwV/OetyqePi62/pTIpRmEjRYFZ7cm6PjrHyBq6YzexxROjyGZ7
Gej+WAeK9LEUzMbPLMqgzyAJ5zDS4E2zW7mP85PxCQq3X5REHLxukbjrTGNpp/Lx
CpFFmrL0W7I+iw/36emrcxP758WqUvGrCpyW05uUuQoToQJ09TLW1Aa9y8AIIvLl
cLLQycCzY+nHnAWIu40BipbpICvVYC5hshskfMuL3T9qQ6xqVt4SmWoKd+4shNTD
+VVnwRbDQRrcjg76GNYRVwj1oUDmf5GJ0EXgr2CIq2YWGNoHkcDqjs/RMqHWeE9i
bIYJylX7ZhNxXCWrCwDoILmiDmYZTdGS3+6DDLFeC1BxvsklrybRzB6OjfEUIUSO
A3AqeHEOFF9tUcSJCQ0UOIvqolk/ckjhZrQl09gF02utrVKM/46TuFM0Isr+FcxC
xWlJWqCwzyL+xngUp6ez0Nc13pFgTuD4NXEuvdryO6hYjVodCfrKE/t7vlsvLr1g
o+FCQzp4Wz6lM6TbT5eQYZ6AohoQuwry71Mw9nmxyIU1oZ3KRw7FP47HwCtITYt6
pzOoJcuBqeKSG1AncGd5tc4LmAxVnKe9j7A4xVNSQ9jgk1TfigIxr25v4fEPF4qk
iWFKeXzysGsdBgZ3SqY78qqOVjx4yUq1l1aDNT60VU9Kgt0K8icps1so6GjMmp/0
yTAIEikaURbN5FZqPc2LQW5JDS0pYNhBymofYBGmv1kBjPYZPmhhcKxL+EqQpvaZ
k00YYy46RRIlYj7p7VRhmJcZ3VvB5dLG10TvMU8NmT6wgy0YkwOGTQ57CUgmCasy
PZuf4YIoeb0nWjlEICY6urIM3Gt9jAN69qITABxpLRWG/joZRjoze9rrkilETeFK
fIA7X0GnIZALFBfyTsQYSu4Ow5ZO/wskMv6m+88yEFZ3ZbaKSTYbejXRIm5RFNPd
oC2E7Nn1TyFrigWl6JSQ8ywLIDt5/vlybp/Bmh89PwNNmv5Kni04HIUjUbWzs3Wg
COb9DWLGCtQX3lvsqJ8g9y+nLSOGCA/bUAqVW9TlyA1QI82Ajvlo6kkBCioztCUh
7AvzsRqxEFduy/GxhA6ReGfrZRdJvTyeN6CUqfEd/kSzx7oKLkEbOuiG+4DfEYLW
LqNugy3fgB3UMATJ+cF6kRTjwDgCr0I1UbdOLxz+9xUz/dK8U6M6s8BwZtuGt5VV
2kMx/p1oTHZvXYx7tzHyLhpNueUpWEQGMfx5Jg21p9yt2gTtFEFqAiQQUKVQGYXR
qLbK6He3+VKnACh5+A8mcWM/StjftCWEFpVtA/zyVDnhq0JroMyVDeyxDCMIbGbs
uOHRnAasQ7UZ9FHT6KBtQy3iqJcHJT92nFWiAFgpAwyYK4dNBXF6Oz1ZZSoKi/6c
WQw4vu3yKBkGtnlS0wDHLa0ivjiro6u3wetEEVdBoiQU899y2ezRUzrM5Y3mvCfL
hUbjVoaDrg3jq5LxDTApPRTNTsyECbkxnUU1GDHGAUL9VLPdZ3bbLQK7lT3fEbuh
dBCsG4ZDaj2QnSgX0Slm81e4IuRo8jb+D1xzlluCv+GTrdBsjcOm/fH7NqGghSkn
tpkm/H9DCakEEZ76+7R98uXl7PmIgFE2g2G48Ca4CAK7keWlQMMq+2QyyCQmTPXD
oidu2L47ENc4Puj8Px4e7ELNtVlbYi2UcxpNvvvkjfgblu5rtgCNhr3u6YPdFNH+
Tjrmd0LQXKcGxx/PqCTb2odkbJENtlbTsQZdddjU2iHWOawnhMnqxWjKAudwYIfT
n6eCVil9Rm6O3DMvzA+dGRYh3lkkfbd+RUGWPptkGF9KqTz992WpR5c9BjK0nIo+
CoJAqj/pLhiuzoLFHj6s6ARBTtqnUBoOcacaZWkA9R21f/qBCkBzmHOR8GHtc6VF
DPKW5q7bEXrb41S6+tXfMKfsR+BJa2Kn5EnzCGGIwQEGk2tfyYmA+wSO3MG20c4f
YHoA9zMXbL61SKxvMReb8Jib414it8LuszSW/vbExvZgPLY9F3Jz+vLqV9sHnxdr
WlO/eSn0EfPYz+Q9/duSP1dbYhFQXW/pdX4FvVVNzwvwj7/J7Nq9AXsQ70WdFEhJ
+0Fq5e5BCiQvsRaZrv3kBw//bfItJTehtiUVTaz+JJ25Nx2/8hrxmuV4Vp6ciyw+
X7jF3nn7p5jNQFLdrS6cruH9hxus8/Spoc2SRw1iqBMToJS91iU6LLvZWZx1+gaU
sfgBKVSvpi6Kja4Lif6jJJvK56nCeTG8elRClHPP85m7MT9yZ4i5Wnp+S7CXUOjU
odB+b0fHBIEnhJ6XhQtHFdLOTj+hKUq6eHiPP34r94TpeRDZfgZXLVx6yuCfuwLG
Ufjkz3785mkM59TxgaLE1k/r0Av+m4itCdlGA8Z7bA2x7wy+xHU6I/g/NOLRJSg1
DHRC77m5ABoq3WUEc37MeikzdnuV3YExOd6lmxeW1pvqPDiRounnuspnCLarvbaQ
KWFAbYOEq5RJ9w/wA1GUyjzL2+95yPh1VoLDybA9uH0hSF7KKdS5skoEZ/b/90nj
E3bnB1LQbDsJZfD6AnimBIlAmlh6mb1mhcTruJ7QE8fhriN5ZYOqE0LankjAwJQd
wkafZEO2O0vbLHAOh5KU8sj3cHjtdJpN5xTuvz93VXr1EsRIip4/Ia5jJqTx1mJx
UUD3MRQtR3Voef7EDT589YaJq4xkTzhVo4LbUlcNkUnwBXNSPFNRobEjiSZNTTHm
OF+52+EtuC71Jy6KxfaaAbuXJpN4WgcRJJzmjw1dq4NcFWffcME97FcioCxy9EnT
A9jiCt716NjZOzg+aooexxvpChDtrdIdaqKfrhZ0rj/Dl5YPUn6UGvVNmKwcMJoj
Cmd7Wn9fRNvejhzTRaTdPUjgRAvF3p78oAyZ0sbLMoCzfdwrqV9KSi6lafwu2zdk
HkgkhGD6yluMT7GDJFF888ZApuHgC/wDfeEsW5i3wr6vFSIe67/4sw6A5asTRGXf
mVBZ4TRCTeI6lnyDvKk+UJDiZl5yrKd3IBwRQzi7UP6z/eRy/xwi8dVy1EOzYqEp
+/v2xhGGS/THKMetXYIgp/xzSfJA6G18npFHy+r/6LeGjLHywwrEHPETvcEZUYIw
vLlZN0H9Y++OHYax+PEz9nS7HRYY00jWPUVGgR8MFuvxig8fr2hxiH+atr4CtUD8
wK5+1hq8XtRnSZEB2rZRSPqDZnmNtGdsxQhX4NKEz0UIWbDXhD230ReVtmmM8sTP
S2XUqbDaDPcdaGnGbAqE/R84OF4l8QfzrN1FE8XZAijwKI8dELqf+4PpclaGw8BA
rV+FIf+TkZ9x7byVaET8/5xwcAS8PTREgB4W+t+dGhDd52SwKKgjuJKDWHZtVdxr
uMttJ1okUUVc/aplQ5z2Vp8XfmEoYLUpI/6hiB3Ewmzo/YCI90IOVGjtwjgHzwWZ
RZx4d/T3fVFWai+jkpGYrySRKsHX+XGOfw0LBk0pGdVzzrxbuA37+/3cjP9rO9kL
Bun/XFHEjW3BW/ujg18K/vqndB1cX2BxQrIuh4m08xZh59cHWvyplVmXegPQEkNm
YcFxtuWOgH5wbPSGelCdSng2h5w7GzA1nB+rBcGYyUGHfeB2xnh3pz+dh+Uvqc9L
2vqowncct1sHEFHPALWtG7wZPWql/bX9xhSoWtXaLLX+GeZsjp93twMJRGFQC7n+
Vp4Abo/uSL6lQ589dDlRcQ192CNVC+aPjpc2+5B6YeEJtRP0YrmnG10ahyqUiHrA
/zYixJefOaAnEiK181st9S8YdqNA6SQNsKHdDh9NjVJWZCbpxaksq1hvvyUQMhiH
vSLTfY966IS1m2avc+SXSfGEX3XRYQ5LMztlvqrQZXo5RDh0cZVFgbIzYly24e04
fRDXXuHEqtclcgiFElhYMHHLHFaDnGJOGewcrw8ls5lrNnaSkzjtDS2w/xR+1ftz
3DplM9wJxvyQN2hmuezbP/xyvht6i3FaQJ6i5pcqKzGw938J0kUeV/zVjSoL2KuO
r8dh1MSs2b+q4RpcF/nVva8O/97cWdL/wP49rRV93W6+67ocA0JuDsjJZHDO3bFU
UgoikmlFpb4BJ9V77XJrOu8VKZ+Mwo8bwF06MU7wNR+2HBnUWov9gsgYlOLFbDak
ncBVoUpQHwNpUICneYjJycCfd9xwBexK8icrmE8fEgglXx7dAe2hoIbK0YpHaw6W
wJ+sEbCmoKwaPppg/zWXDAMZEvrDPbegqWcBXGsJ5xwVocu2K7dHrdxGwN3rLcd6
2keiu1BRxbFVtgv4vDIQ5aR74re20zIB7gc/jUrNFW1IOiLePj/egJSd38NSmCLZ
sXCo91Yrhqf+TLrmsy0nHEuqdv5OaapIxG8IryalcKemEGst1BH9aJK7usHM02c6
9Xrq7hYQyyd7qYz4vAr/s+j9TfLVXoAMKY5XtY2F1QXqAitMRFx/Ymvf6fxlUw68
O/Si+4luRqOppSYHoo5sfAn3lprK5xrJj65k3EDXtna4G2jP+SKvg8B3pk/nH8O7
YejRwap8cs2+BXEFG2Ic1qrZL9y9gksn8VzLCh0vsCIr8geogTIKdrAQpTydk7mq
MiAkuM3hQS7BGiAE53K9uQ7Jg/F5884nXZwJXk09kw13Iik6ajwJvwfVKgIEEE4R
+wqKB60LnhSyHr2Ix61cKrykysUkQO0xiD2dBEeJGUqvRwuwF4w1wiHuXKyy27Gq
kSojRIPgpCVcKXAWaaiTGaSAysn1OSl+NHU0yvETka4r4XT0YpdHsZJsN3aVnMAP
V1/E7yn/O7djRAcGMhS2gub/TBLUmCanhNumPL8i0paqdjZrQ1OsDIyUa6cPb2KZ
K12zILgwr8DCa+UTzMMP0iq+i93XcWEJ03+/scRUgWYjOC1g/n9HyAAa+W5ShBjk
+S4kaFlzHt4zLVuG5SU9aZAEhn6QxYi3vWJoVtDng/L96ZeqNsefgcWMZRqQrSPA
hXbKWFn6BxAs712VwyCt288c7UriBjGhYeNllxUZc0qxPD7pyXWaQT0btP8rV4of
tziuj+uVpFKkzBEb000SFFN/5WfnqeM7PKHJq1Eb4BbJkwLhwpBPQD8pIy7tBtz+
hI73gri/JTp1/NmfxW2NnDqyhbBmOLnCtB3f3pXkBQP2kTWFrZ1x2P93txwEWB7P
ADcdSUkbQj4pItpun8wLQ6sIw+CcFB6dylWQ5oEqNtkcjj130SnSm+cjBG0sqwfy
k1t3tkftyFFN9XPjJC1qgkV4Y3Xakx18zzyRhS5HooUfipSG5sZF6x4Qn3uQNu4i
7PWaRscYXvdh5G/RGOUL5BFo0XdnWl6LXMI1G23kJa/75Zx9f/mG+Yywa+euJ6ZO
qgMz+2G6rSke1psN/MDs9JuR10ITgqFc06BsenmDM6D1RMYpM5E0ZYw+AVZbFpNa
JdJ3slOsRf1Pfo7pSAFFJx1Za8OzT40B4E+bSssP4xWmq+pF835dAD69+fPIAniw
kZgmCu4mxXHurBSUpUO4Lpb6m/Z5DHm2Qy38S/jXj44LB6cZlJfJGXEEUYmJ4Wqv
F7cSSqrgvB0cd1PxPMq9pjIHihlRVM3xPBxTAchka0+sUQTfhChKagG9HTZxsz1i
cHFfuJbAvRtC1PHkr23+tXyvqovqzBeGfBWKqsWn1gIu6YyUh/SXqDMpnF9gNE1e
EXOxY4HhxcQl3D0QlJ5lJDAX1iHVmpPnTF90a4OAmBgCpe6oXJJpGe2evMEQguzX
wFq67Nz+BrwRtZuojJp9D+9BGRS8UO5xH2eUUfzecfwP7m5U1Hwmr+vWvv44TUzD
fhA7GiE0OZepnu9h0IFbnYi7+mvH0ZDQkdjB/lS6f4WryQLj3i7sjYUd/31wvacI
pIiDp4jXhLhOx5zn3XvKaONQzjY8szO8DfMyXtSnUtwEEvkKxslsQWEJOEqOxmF3
b/9gSPV0pf+Kx5BgP0kWTQtSSknrxwFarL65KCE3uBiCkZBwG2VcxFKpg8/eTq6W
Y87c/1aOfezBJoqIt3zD69S7yAgh1JCtWJZfTCM6kob9Kf8yNDVFCo2o+ze5yM+Z
6wsf9GxZcfW995S3amu6Eanj2jw4F/391+lWMUTlf/J6YMxeaex4j8WsK6duPvso
oYS7hdP3AdtnNMhc6cdRU/49Tvb21ecm9bR6TpGk66LBki9PhzCbwVN9ynIhEpsq
fULp/5xG+gW2RULKki5G3QZ/XuelP+SqLQPxFPrPh86Mwj/0lroXytSr8Pye8G/R
whwNo0R/+vq0fECaf3LdTEErMHTVqUGeIH+ql3m09LGEKYcRob3FhXxld6xjR/M6
2xz24yMlNdpfGAQOHNSi7GYtSV3s3/Ek8zoxUlfCsVuG2Kh+88zOyxrDQa9q1DgT
Uf6NWUY8CogGA81SPGCsdmSXzrXZqKd1enAJ/ayCfjvXTXUwZdaieo16szpRXsw6
3E1C1Y7FBLCICzb2jydssFuepDf+7KDXQIx5DfTBG4xvJuSlu/WpuIs3VuJbWnlF
48l5eeh1M81sTp4cz5ewoO6gG29YM2W7aQwgiD7xP8t8yEYsNRynaF4P43KM15wd
HX4zTl8ZHHGSyWYl6msiatRhhl79Jvmg/GE6qAC0KiZwPpXbWDoBL07knVeE3kFo
VxhYhlbaQUK9V53WyKE7NMMOi6+Q0p+3egVmSQwviUlsFOt3jj3mi6g3DND/dPRI
Ye3k+Zw6ol7FU+C3UI0oo9VOYMlzrnuaxvHtBAU3QzAPaAup0rnYNjQH4eZNeNYr
Ml5btvXouKrhM+rE6BD4ctB8UJUcOhYT6pXWuLxaJtYuZpV8IhQFuY4Fl2ExHqe0
QXEd5lDYbbGnM0Qx3UxbjnkfpRqsbm2U8kT+FuRIwfnwDst8Ca405ozosJgbZvLc
J7ZPV/YEbkVaSH+LeJRm8XNElZTzyqcclnRNVWlpRNocps3+5KQjZbIHx2fUZjIE
bTHguak0nJpWwHqQk328VwuvE7bmmQMLZupYRyAanakHOTEdEhFugFdZCDHLCmmx
g4IP+lzLldlUitB1bpHAXHlwLOgouteYDAuDpKD7fYoaqwG1QP6pQPCOUM3TAzZS
qm6nzQoQGRCa6ElBsC6nOdP6SSEx6o31QSb5lmsLSqrutIANtV4FgVNr1kapJFQ6
BAEusVBY9GwrLJwyQgjf+FmFOZ+sKtkI/+TrT0Kh+mdo2RNiX7z6En0piZSpTlgA
26Wf/U5qff0humn3OAQQgPJ5YQuO6WXpQUVTUOxrX/O0NEWYR414u+y3/5Cuc6Nj
C/p5z/L0R6lP5GDaoFsQ5w6ms8D07VFOXCPcuSHwyAGKmIoyzsW4VAOUuRxJsbW4
U8QXKqJ2BDfj9Y5KxlawDXKii6PIotaWr7GoxaqVGfJzIswevxaaMUue9r+vP4tc
i5qDRW9pnmam65j+/kit8iGMGiAJo/LaTyBZw1S0JTbXCiN0wS7FQPWStYJHfGTb
uMIi2TOUg8NsJR40D2OBoMsZv4C+bH/W5vHGk3xNXkFaKkjzmAptma4Nrg1Eg2ks
vR834eP5snJHbYd2/iRAXrISItG9WJBUuhoUarPR/hTtHHDOJ+SPEayzjldFNmWD
cl9tvDcjwSz1aJNHIR+VQWUjXZUO+pfPjFAUvmBdliU7Z7iowMs/9+lWGv1utZ30
A4cN5iFSvfQyW+cbxZme9U87lSXxMcIYJjUkTLkEUNhWJ2diFDj+v7CpzDZ3Q4Sr
r/1AZPbTPOhNITMtG6H4EeKhaGGZ1XDLAi12L8BJzPGWxPXmEZeINea8+7ufgL9r
OSsJqeaazfbJj68yzxzI2N6pd2AdlMwhyf3VOxMIZubFO+L9WtC77ZcczMRciOsv
eg9yeZhajmAP5jY+xmEfmlYUsC9KS4nDj3h68IDP2xy6F/DBlbDOxlPYA+PJlEPE
EvehND1sm1/Brn+kLBIey6WhnoSX2sGZJ7EMB+22e5zQ7sTm518Xg/nqfO55ejM6
Gphk6lXTJnYkZMqieEUQWb5Dxx7LOpmNxoTSu7NkC776OTdJOVNE0WedQqaGKBQ3
c9KyneZF93iurN+Cw5on2LrE0HxadjqQN/DmVh5K1wH7AzZrJoc6jiH7jWVHV0py
sebea6Sj1/N0z5b3wymQk+fQWahGfhUiLq9r/jBackVrgt3bbJzt4UQSBMfq54a0
bpPsnfzMP2Wo/pAK5yl12JJ7dUzleMegEW/SssRhI0UIwaARwJrcmJn4KAt5JdUd
By2j0IQ7N1vaxZSR0tSFI34SPbbW8lYgtp9roP5errbT6IvVdB83rLW9K6f/PG3d
FHUrjLKbAJab2OJGFsTGSQ0PFPz3ACc9EfXC12gep7QyQ7DrgP8d5SNQmikowYOi
VmNi2q2vJ+1EDV+0RBbQEUjBbZ0YFN+D1zFoBdwwCPpuzY7JbiWAQPr4Ughw85bc
1/fyaLgpQG2hfK7b2w+slsN2vTbnkZtRhLBDRhlkEYTS7oGksw7E3+UP5AaKn2II
5rtSXMLBfgBHEZhQtf5I8Oaf1YTEzKxsJyOqSJTwurP4rl76JeE8fDlmQ2hbVpLz
kjurzFiu/ejpNx3hX3eGzbKbFDkwWFE3WinYpYwOmucoHIDy4SeTkbVB0a8sBpC8
5mVnK4YWWhgs/IZU4WH+ZpFTR/f6BI+CxnDtVO/iNIXwcjgMJHjZiqjVwwa13MGM
hy77aVvf+BMGLSsmvds+l27Uk9Cv89X1/jRbtcTlmaPnMWn2DJmOdONs1WKkcWAR
LaopsQ1Rtq7iQEE/KUvpQp5yEeut/Knw30uhX4L94nB/+kXEpITalzZojgjdSs0a
xz+taqhZ9KJrSu6yvxAdUMirpYF5ny/8uc9N8ft7kabCedZw7PhzNxruplS2k5m3
SgHl0pa/p2ANLm0pttIsW7ky4XG5jAVTro+mzapvCtxQaJr0LYxrVH11aj8jUj/f
TRS+qVGYsfuUG9agv8H/NeKTdoXv6f92dGvdwI24QZ2O9HjY59QPaQJkv8odvQAR
pmjkxLAhP1WzV8F1tYRcDkxH+/l5EcbsgoVG9ojmiCFNOg7QL3K8PpUTtOD8Tl1V
pC62M54R/Pe1KcE6Bwk8wa0i9uiVMTtNeUrHeXjVt1G0YhlxjrUSxR4d0DUc8bJX
7bJYrWAevQsDq01hFsrSVtB+8U/Hf6hjHnDa0fFUbAWOpUBf5fdQTeQvxp96A0YP
5GFD/f1d5dWn6yWDEFj4m+MQZaqdaWBTOMqSpdCAya3B+4ywxuyEwE9g33UtK070
Qv5wvS/P1QlwGsB1Tw/nYG0+OdTzMiqi5WpOECp2/RDS0JjOALPviZatC6UwpIWs
mzGDtBW0tFR6yOmt7d7SYzHEy0zXkSTC8cluncOvt7TmSWlG4Xx92plp6mYoF0O6
yFVIo6u9uRONiDdmfVzb9IAgG5poe1hMSTCtWQ6ilp7eRRghvSWObDQKMhm7D16E
+IphgDd5y+0YOwkohgeKf8erKxVcncleoeJCbm2mcB4IgqBu53gXZbZlq2c0c3uh
T/Tai4jzIRcYmc0xl5D5oPYTBl5eY41fB3rbK1zC5VQZqB76FS1HbjCWKTZzyX2j
qNJzzXmu1wndcIttjWNqaXVimSBuGe2hqULI/VbWoNW5i9Yvd4qDUS9ER9yW92AQ
GzfctJouGIsspXvt/G/bMBGRJ+cyLE9p12qZvhP5CM+bAXg1DQqwCA5e6Nnx5WD3
fkIytX903RFvmtEgqliborREWM6wOnEGPJV/Nu0b1IUSV9RyaINU7PQWLJ1XGHID
ubrOpQMjXBZtRMt8JbdNWdQR+kZBcIxVF8hYWa3WaZwcliqAaiQUKyqaYqpZZ7ND
QClglvfTIekL5NHRtuRa/XHZKB0kCs9X8gkrm+cfjdubP65hfVhosd9U8LTM7oDp
6nYyDipddlZlP4LHU+EABaGxfMHDlCEQC8dSkqbSv+SOADIwyYMSxZsHfHtYUgLk
1+x0M3c7+RrvuQcHfLhdyQKbBEyj9rQzPolX4/F49kodmUgxppltgxZUHhqXmAQ9
0hXJfY/jP4m5oRSSXjiERh7j+tB29kPcxULrH+M3HdRO+zoQpvs4BF6ApSLViLLR
5XPM4fJwPjGaIQfUwyC7LrtQm7VI+NLyBGcrNWgSnWy/G2EODwWx6IbSGD54R02w
pjaX4eCYwKBO8DLR2ddfMi6nsoLkqbgQ4rgyMxSKbf8lRFiElmJTvE0jjk4jOrIp
NG7YGfAHQuqGCpHuhbtn0Z6ANIKSpZV+Ehdyi0Rs1atjjEmYWsq1HllaCRH/a2yr
ri6JDbo/99CKsAm9lqZl5my6XuhIsAQkbZERQ/EF4i3/hoaxQVgTzrLRv7ijqHiU
r3j9mnzwUN7UIHXeSpa9cW8dB8wpVDqdTw8nK8FJwfAUumLpT3H/hTXlNsuKvnJ6
4f7YB+g/YcWERW7JLTpiYp6hl+trQyLbmOx3wwPP5t4bj4P1zQywKMrQWW/pqhJf
Soz+nkvppDu1t1rim/lD43OQpS4UIXrpo3KhyIib3u4/Mmgz8ijUuWrMwWWeSQkW
iQC79HE5NEugYhMSir0IyUVd4RCugL78YSoDJm3DsdZgNPzB5FqN/jA5ytllDf6O
+NRXM4pqsL+QAmcNGUv9UwOlTFXFG8faVxXwjv7Nio2kCy8gv4NfugGx40Jfg1Ks
72D+EGcIULWVNr0EpF0VS3LILQLk5lcM/0ybHBsvBc63CW0Se7XBVCKb11VnNSzs
QSFcpQB6dTwil3X+NwGl4/ggT7wEl/D/gr5PckhZM/1An0K2p2RtmvZu1fYrpLYI
OszWHCpKJfb1fUAsuW/ySPw98QS9KjdwV4hl4RrLXhh+9CzVoN0LeUBFYvcQeYD1
JsFr2vtjqS6dLgIsRc4/hTmFTJdwawtYZEV06M/qNBucHhG2KpoTmVrrRhH0xXip
iWn5GI29nlb9coqD28Pig6DLzHgJKCUoSp19k9mfMPvbMkewvoFePk9Wr6bQvYJ9
erGw47tFGvOh6vrwhLrrquvV2OfjBFOQZqsfSkhc1+Ufx9cOWvedxo29JEz7urDR
70f8qWRin+lxZzHk5DrFzOTUoYxhXdkHKJypBXbwo0JgjSBFp3Evq+yzCHfTf/JX
kp3FFPzCYEBOAmyiffbhQdr0L+dX57eHEd/Wd1aDplcAMn6Kluk+p/SyUTgLUfYE
5D92B1vXYwUZknjGstZ+NJmj12cDZC8pyAoY4Or7umRPO1A+yOROIo/ajAlWKUJF
NEyqtKt1tZI+lBN4OhZ4Amy0ULnKbk0Bra0LWAXjO95tqvKqjpaX/w8sdwhRRVey
IUdFQFgNSWlgSC+elGb89oZfcDOoyFTc7sbbormSMEgMH3zcPLlwmN65m83As02U
gAwIvETq1ZSkH08h2J8DnlB6Dwu6fBQY0mvDUxRZAYc6OdoqV+VSqyTmPogXw4Xc
Pn7wI8eMGobFtLcUwqCzWlYLRNIXxDUFBqUDhVzB/HtPjn8CT7V1gHQBjLObTcz/
GLFmyARatASGVJYuGvSqvprxAr7kqmTwvAIRsube5Au+7uHOZW/rAa0hIIKIpkSu
iEjLSxXZt2oEDAULnTov3q3MIG1Sq/EOb69sm4G9zEFJh2P9TCkpXsd4z44IaFiq
zKExvWlmeP5jDR9JQgxkopj5wRLJNMbu3bjDq02h+Nt9Zo52KE1bFAtuqjM99iQi
wKcVlTgaxbFJ0m/ZOuWJSulc0ZdHCLgMQmDGsc70F6JMOGZLGyQq1ERRAi/+HMJH
eF9j5BOoluBwo4hW8A4bAK4EB+wrb2irIAM7qL7QvVhvEqJsiOK1nQzkBVuzzSGe
Eb5c1JpaQVa0MlwY7PpEYycBnu//C4yQ29aIBlFUDo3095ELdusoHR0ymJq5tSLH
wVpJQANSQQCl61spIrwJN7oaeGQG5MubgZq7WhdIyYG+6fdMSQ8qQb9HSEiTzc/T
KL387K6AkCJ+cs0qmeshI7Wpf29XlPh428Fbgxm6lJhY2WAPUqp0Cx5WC12CDiIN
cVtg3pr86wIJS0klKX0BLcc3kK5jrOpgIxIo1AGuSBlPGiT0UstFLe67ZS8xuAGG
oc1z3pSK0ZAFNp2RkcSy4PeK9NREPypP5LIVV0VyqTPZ+MH8XGKvTZK0k/cjVlLA
Z+v7IRaA5anqyft3JSPN+cgS3OAtIaoyJEZAgMC4FPygqBQOdLO5yEQ5zDapLiMr
Z2QWAr1X0Iu27jKKHYNkTNKRHOF4QegY1edMTgrOSZrAcUaiZQCKbh5WnGAFVRM0
wIk78Gg+p1g6CGsKxYQyy9Cq2d7ETxy5aEM1dyG1tbGV3A+hh31xCiC0NSgMKkri
N8x9P4NWovT0/g48k5kXiKQvHRgzhOew4POMwEBASBkg1hqlbH3mFJAUJ+fWrsp1
Z0UuYgaumiUSVsSKCfrBBN2/LQtazHHiBUOtWq1YZ/Yg6m/1iFonJEtaMKxG5TOv
eHl+hPLCml/I7ttTVvKGNGC1dzJlbbjIw7oL4QCHMzQNpWsdYUxmky/kJgzGCZ56
LxRqCvNaRBwANHv2SLzcr5oRSamGcDjcYwnfdKPo9ysYyI7q7zQYaprR751z1TBM
D7gRU1GEKCcV8eJu7K9xdjC6t9mr9xAG+jRhni4vSkkLAgJOe26uVCwX7jSvPzFP
FDEhFOkAoG5wLQnDmuCGquROrL3XSdAOj9YMKmGrXDY6q2AAIsLGQNy3pPp0dGHI
t2ZpAsDfnoFqHzLeibyLuctC09lURWzNL+8cRo4AYb9ktPK9awYW/oo43YL73XCC
VC8Z+BpUagwvhJffgPhaOAyK0y2dTX/wEWzXyZQXVRntoCJcqiu+NiYVlb1AdNB6
IreImopij+wV2xzC/rYJCl3HOXJS64nWF/LaihXmbzKn3yV690La9zJqBTbtqK7f
gP0ns66NaSTLed3JxXp2GItRVgyPffCRgarldH2Ld7mNsO7aRfnetKcaudLP2iy9
D4A2k8HhEvArxZs0mLXRC0Erl6L7YQt4HRhgcMxsJIHMtL+WB22WJXzs0SQcmcNO
OfsiH7gX7o3FKw+A/Xe/eOOVQIZ2HE7C38XHgv9SWzIq1xDHgW3kt4bnk24qZyPq
6GcADbpJrxOR/jaFk7EOnjYA6hOpXA/PNOLiv+X0dWVUjviU7X2W0bHZn6S18ody
aEwkXCe7Z4SpMu2pJOSmf4g90QuyKWJcjOfeNHgGnX3H66DM5nFkwu3JNLPzo0IP
k10c3e4pGQ6zugyVC9AIyaLgkdj9RqqB2BZJNdGpqGd0PvEkKypBO0mQu9Ig7F/r
fuGQ82chtD4dC5LIoqX3ei/IFvxlJyj3caf4kRHCXxV4DBfUCd/3CNSeITY4Ge1J
1xWNbUYROFn+OEiwBP7AEJ2DL3yIgcafCqbMaJG5GLUoA4yzfYhogrpM3dbX411n
cDpQJLWtAYGCz4kLWjnvSe50MqXvDNXRAbm3htiMvbv8pouvBbwT29dbVQl1ODzK
AcVSPIKAMoYhQn5dE1h3JHn4TW2SMvv4aOgYqeUVDG82dIrqR9fDQ/kgred1Qx4C
5+Bg0d73mLw8L64czFegYXKrkF8tH6Z1Gq0ESDiauBWQissUi1tflva3TjTSIGsQ
rjO207DcnAE4aEkaoZ2rjLnuy2khJxe4SujkIeDMXQxY6PwabkImcLYz+CxBS7p1
v/DNr/hlxENj0jV9ULnXjQliUsSf+zNxxH3oR+fslHJ4fd+nfhvo+nZQtFMvIKBC
JNwGuFqsYUP6xwNzEsdO0HSHMm7zhFC2h9C5Qq1r3bJaRivh/xpN4zonyMtktqJZ
mVKO14BDFFyaRUB6OQjhOYLZau49t0EH4Pt4L4ghrPXNUIxRgaDscIVS5R1vz9FM
BhheXbOCQmUz80q975I9qzQ15aZpdZn5yM++kKZHhGgZtCCUyw4Roo/l0g2WhiQ8
R1x5N7212yRhCDkeM2hRKEwxj6aJ0sVFsHrBa2wJFjTRrO2UJjsee4ESxrdVSv2T
8HE+0T4KWn5wrAM+xD64UPkkDhAmcfXGBt22GKRkME44fwgZZjw19c3ruVXewXPE
ki8TnZAQ0XCxCLc7cJizmpdNMdTTD5zPQ+8lj+lpNFytXLe6fPVdSKbHzqD2EGTV
6UeP1dlodUqJdasNpRZB3a7iilv8tHjGiOFB3RIukMCRxlogWozkc+tWfMlHvpY9
nQ9i2mr7jT2yvUwwJKcCyjrTG6osZvkEQhyYOdOGuMzlDofF5xZQXCtGXzd+M7SP
gYkDrGxkQiVd7cX3PcGi2fSAjeTBX5jwDdvBJEJ/tefwzUvLsxiduAZ0/RW+e2zx
f58+bxnaRx/XGstBot0e5dzsrWYvUJIVf7r39EdmIyk+z5CULgWD+dECJS0YKKce
KEmB94d7BQo6YmQq9aIa11NM06u/YL6cAhqWimUrW+0QW1U33orkzZv6/tY58IMM
iRAS/hbKjQ76nwhYP6/QaGPKELJg95vc15caKCwMM/ENFe86/jcucGQWqyS6qsTa
r5mRuZj3A6JE/KrrJs8EFgZMMc5GKfUc5QYyXm2CjUvxBosYMBBH5BGXqow9UM7Q
/3eWkIBdXlIVlTbFjy5O6XX0vUzN8OZG3+KSSP8e6h0J2r+Yr2maw4kdDjeGc+k6
0xkkuhXdkL+epdxfS7aFylYDBHb5TPw5gC80lm2qFORD2aEI0IPpz788s2xinf3N
Wc/abCb2kW0nD/JnWz/fo7bzBtz2B+bMd++LPxvMAYY4dGwdLx0y97H0rYNKU6R8
mU4A+RKG/HOv0Sfhy/gI07ZUKV8AuBasCUX7n+uQSpv5gT5HoXzB1/6zhi127krI
+2nKXENM0p1ww2cMT+wJW0QGyvRNFAXhdTRKF/lqxWcRpNqrmZUbOA9OIpfl9lLm
X23EsjYtpWSwxUZVdzlV1eRJfAZ8vhESquooB566QfsJUjUMeyLKnOwmZVRfynnz
qkthtz7OLfQ/hNME2Y9Hy8quXx3jWYr+RO5POrg9yb8zphxvanW0xLXnrQfjiMB9
+EPktz5oJe4uqOoFZXQ4wnyqgvV1elzwxMn7ixgGsa8FUtLCh4tM4llQYHL29zbl
/bsuDLkX/dER3PdEPpToX2dJM+AlH8h/fp9vktaJUVd+uzR5Hp3nXFfQvMZL4eXD
0G7RkvP+vZ6BKze1XMfAtqKou/VE3IL5GFpq9ZPkgzGOL+sQCXle+de/nnutZp3z
1dTOfSUBs6pMyISxjFME/6wZViGJIGisapHXnrPZn/HGeZZGfISMH1bP4V2GObzl
Lo1Acj3dI8jwhrElMXj2zv72zJhP6B3gCcT/nZJKVSrGHpDFycapbTBLzcw1SBwx
fcmHLUBY/C6uVxVp0Ij6uhc6yPHCwA0raBQgg5KDcFVxpxSXmIEhjBwM1x3vS6ZO
taALQN7RTBe9+jHdew45jhH8bZhVJ73kjV5n/jVZo0LAYYW7Rhv8EDGiY87JiU6F
e+gWkPJV0UnFlnumYglO1AR5jlxqVD9xgmf0y58czxkUQ3BqCRZCkPZaJ9wHwy25
9MSj0dQIWJFD17xnZsxeIAQd/hnzO2Ys3BnkCGtttBtseSfd3rRA/etxvqzkNotZ
UbsSLTCweG4wRx7GaoJA76NWbhfYG4Nwc3P6+SMIXMmnBhLJ23+4JCLoga3ZLBqd
1fCATgCk8q7Y5KAOPu9ScXFJU7UpEXNB3DrCmVOrMfO2yB6+W0JYZcOyf5+zjL4p
1715oPApxTtVSyXxvwagFKg/kbZs1fqJ2nKIvkWW7aAb0gfCKCoWdvkp7hkDOyHl
+KNTQ+nUW/Y1HN3dA06UPtPEFzGBdYpRHeueHJH7PW6sj/BXWHynwx6hcUKTVgLA
LvJYbhcy9v4XApkJr4wXajM3aJ4JoGvIPdqfgyIGF4np4zHpDsN+1VaVXwOT+vfX
io6G/+pbuAuvSCHbnIlq/YeCrjXnVLpvvvs3p7JgEZOFpYBmQ+7unEJc/EiJKIWB
BnJHPYE+zD8fH4znpi01Uztwm7nxQEvj26qpAH79ZbgiKNwkeHlTP/hw0cQ7ufU/
CigzPDoaCVkjRM/CXya102lQP04tQP4PlBHOPzBCBfYSAtcYJQv1/KqvsLMedUEz
kgMygui6nmmWs0s3dK0jBekV2rEkK7YeyzPUAxWeZ2Fzip7FqQ2+PGW8/btwBLky
l9Y3J9XTkfpWQdXeWswSNQkNc6UpzE/xmy2BiLKVaVdUXndSINf5l0iKOStfgVDT
VYnlVJov9CPnTc2zObrknaEn2TBTWnoexC6kqjB4IPAtqHLWFYpBDRmRUfSCA1P9
yZfDEgw/fxZs8TKe7Hg9Gs0VZ3/2QjpeUPWurnXNe0zcgrrHslyM3ztmo94qUaQr
vUIISvli015ZvJtB6XbEjNbFZ4LYtcwe64JZEMnZfvG5D+To19d3EQhesSCYO0D9
qBcnTDVQhdvVd/+cVYfzmhficAHivUI2eoKQDpJ/xgLZINBStKFe2/BK/esgf5VL
X2QiGsxQoLuBE83gom1LUl6fZvpX5mGph2BsTdqD8WEXUe0FtfwLU39xLOwO9M0G
UYZNpnf125SWcEp9iTc2G/4nyVePS/5isnLUbDbmlNA5+8SIiVCqJzgr3KJp44w0
fL1HwvCHcwF1r+I7Z2x0O9slIBmk9/F6MkUhOx+vdh3fm7DQ6gRoSnNzpxNp9Gwt
FOT17SqUDPd52ZaSJpGc609qsftx8Q8vJXqY7bjEY/TtmWi1zUy2bUI3p7P6BsOq
MA0eTe/LXB+mwyBgF5nGvMdCXeL02RCIisK8K2liW6pWDvWcO91xM7mUjLi4PQId
nW8gGC+wnDmPyD74rCasih6o/W208UYatBzo57dvm4hqBVs7RZSSJzXS1QiIRtRy
s2PC+vsj34mslVRfhu5X5MhzpvXtB9m9bs87cid/1i5rU99MBv92jvxrgGxztHa9
LTGOZpCrXPmha6BP4ANYYOukzwmObSaptYltWjuApeccqeQj3ouL/AV7Y59WJIHH
jQ6Htk6lXIgtPUZPOtkgoB1TBjfe50KbwiHqSu5VHzQX4LPalg198Rzrf2Lg/hnH
4JK8Njlokn0EyMjLrMJSbNkmZrfKdi7R08WIG7FiQZBZiEebrHPTLoidRrmVI9WN
sAQR6mFFXw1DMG5Lt+6n3d4TZTGWo6npBEhRrmEHlBVrDNtwNBHw7Ymj9dd79uAP
teEVXmMaZO8np8gNSohgyiVkHSbKNgRy8rwLDCrbYjdoi9yDt891ngGYLVffcJCh
+Khrf7Nk4JDUHok7wR+j7owUQYxsmbDQucpddEgnaQnOmuHKO/dApev4I6TOLewV
oZ4tAT4QujSIvn1MVMRwPlKLuCMXrncCD7ixVgCjRlpQ0zKpgpx/UWFmLVZCmSFL
TcPpM8VeaGA2AX8fYXfb6ucEOLcDY4H14com1Pe2VTiLbFYvyw8RrUcngzAln4Ch
P1qnKuS/OoEgKw9+gcieGAI/cbzWjI6XeAPLDuj+C04axs5BdJ2LFUJWw7oekZp1
X5yOkAk5LgKVa5maDrT1Oh8HpWBPoc1AQC4Uc0Q3pVBY9gd8NivwNzypqczTLWf1
EfPAOUfr05wH/S470jgg2Bk3yuiqD3dSCf//iPLVuOiIEwvbw7Ck/lbuGxh59djb
bgv1OM1FgsyHbQP8z1YdicwbIZwPawIgaXL1eHoQpa6fpvl3u0S6VxQBH6QU5jEF
PNnzk6gJPA1xRYTG5uc4Da9BmXsOBae3LNbO+W+pNYIa5QEX1V8rLVJbn6jIEPLU
ibJhTUVSe8nnbb4VR389s9Zn9ZxBgjqhiNsGARdPkUScpVmcw+ymBPslhB7ZPbZf
4nw+hNms8bNps/4U2MKOmd0uayL+JcOP3OCEd3xb3cl8hwUPlVfaHrkF5mVHR78C
ZZtUVXuuwXjpWThabM3nurL+DOG0f47pFhsS5qvdZt4+QXLF/O69JsM2w2KgVjV4
0O0Dl4kTZvL8ykweLMuBTPNBjFdRCN5MmM2XLXhcN+3m9Gwf+HFakd2Jmfx0zJna
JHoeFqCqT62Pt8lT9TPISK3uK+F66bugl5IBaVUWWJef702Ft8rLB5bE3Iq1r3YY
bzarcbDPkPoirohV0W2Q9wXBXwYM7I7w2WQa4plR8QoMEbooVpunM1grrP4Acr9b
uY3q1+YGl6pTIqkQkm4nFH7RTDt4mPPeWrI9BtozGwI7opBNWrpMBSQ/FXU5REra
6rXVJFKSkOsclLbz1mM9jdCyHjHPaA5RslvXEUQdqEPtrqLfFkROW1PA2RO8eveG
F/P3kLEcAEgUuk1ax5BznD6TA31yuYhW5hcaGrU1c5pJVcjlCj2ni6ynkfjJLys2
E8ytz/nmq7Smg9idpeD0nvYtGwWcd15H9ATZX1kkEB690mM7UrqVACnXNEaghQcL
SvoEj9ko4Vz/D4LW9mh8Bo38O6qv9jwAYltXztFFqItVcgOPyRjoo7Eu2ZtHhBNe
Ig2N3v+3QeP58A2YImHmTn5DL0gE9IE8nstUPACfWq5/dLDo4ybx4JHBvLbyznpq
2z9TvyPwsBHkmbZ/pYPphQ0L/Z8xdvag+WvnPAcbNzx2NRks3/BxRQgnKv0gSu2R
oYOamk60vYZRinB76coz28nxPNY3ZD6wqWg11hriD3kd4/7SoOjwJenHAH6ZqSFT
lm4pbXXjck8/Lgv8LkS9n8XtCmeBxn8nCVoJ2vDRYsxSXpgamXNI53EjdUGJw25G
KOkPoAOkMCC/GCru17tstu7G9O+kE7aHCqk4bHvcKnZBuOjepmGSY1MPNMFjSc8R
npdlz+VWIrigRp5OmA8MRqI49pTGU+xlDugDkhcbWNlpIb2gryB5xcv/APgZGkJj
JS0feEwOVAx+WwLomjegrUifv3ZXmTPxz1chFAkGjRTgjqyHRNXoFFKklWf2mwPo
xOxsSt+OU6GARO6+rq0gZTac9Xx+wBGu1e/boGhOFw9MqGtNuCu+3vGyVtxp2doz
f7IuPLPe5INW098S1Q+70lk1OED/VFL1b0iWFRTnHlxiArT1Pjlf23cTxWsWw5+H
4uuxnZ5A2JffhHFx+WnMhnXKCgfZVMS5DCDDSD9B52Spa+hDwWYWgcblTxM46c+C
qOE566Trq2g0hOtDdyujGbdAGgKfvRm9pw3R8GTqcbysF6A9IdBs2G7I6AndYObN
BDaB3I8omYyvO0OQ5jJbiOkT0yM/DUFfK+lPXW6/ExjPfuzO9tsvEkoacckk1ioP
Ezfs6B+9QkjIxNV4gUl9VJOj9U+HU5rl+FOtzQWy83byHzZlJxYSNJI0sUP4CRtG
6U3ZYlQuiBRqzUvW/+ekMhBaceHZpywG7DQQ9JLLuQsrf/XC7b4go8BD23FYivyS
29tL8V+WGQp7wN14UBfdFVD8R9Z4bzfl5hJQRq7O8iticb15NwTi7v63lMRGPi3+
aSJz34OvnaRtuIpchJPCbNa8QNGn9cW0Ojuy9VqQ3FYV11VMb9wPyWjjX9SZntRA
2MvQmyFy+d21N2A14aZeklgaKjh233Bhdh7g5mMxZ0t4tDd1Fg5dFjznkjGM3x0z
08DXfUmzk0SDzif3uQOqGhU2VmZOiOjrzMSs4mvm4eyLZK2ugsnguzL7nQaJs6YE
g5Nq2UPovt2SIHmUqrfMtAjkVsrkAlGgQM2woeDDXgCTDAOIAGWCqHbUVvyRaKut
vrX3mdrf5TGpVo+5P6KNfdD6ZvXvpJAAPO7wTo55DE7cV4R5yk+xqh3xZmghWUke
xxsMmtv4V4tf9T+CykD08QTZo/yY0v67Q/Kbgli1UjJVTvWVa7D1VUnJTPmJOVIQ
k65IwdMv3r1idazc69JZcS+ndaI9evWXbRZKJNzZ1JMR/o1Db+JT5Y4THcjw3SCb
C+BkMCdIOoJnULpvSQFbuGkxN1W7VALx8uy5ffNYmz7+ALotc6TPbeysEuBbPPPu
qM/4MLqOvJWxcTlKES1xCrgHtJB97l8klbJD/YTFHJrmFdElTtnmdESsywkQOARz
o01K2fyHca71ZKEHyoqalfG1dZyrP1sb1J7/3xrELC+ZVCEuW40r9jwMMcQ0no8M
ixF0Q4YWogCac2KA0gH+3UB/OVrxzLpcQPyEgIvS6wId+Wl0f7mO7CsIQcKADHS/
fA0gNxJMYo+rowmDa9Te5wEPaDFLA8EcJqhHzpvj0k9Fra0z5RipJJQQU/Pa6vv+
l2Uqfh9YMmEhMSF+GyG/NvLX1TuJK9rdIDjWXO2ueQPzWbNG5uZAwnC18EwDj/qA
ADfIeDMyRymZeSTRSunpkYvr+dMnq178QU7NxTqvwcbZFEJv6Haue6GKJrl+W4Yl
I4f+BXCJURP7v1ZiXwz0GZXu1bdjeO2cil6AumyXmq/eoQ+gf7YxBw5NJdq+QdJx
olQ2Z9vhZ2EcCIqvsTTx85Lk4LLnUJ2hxXSGtu3xOzPajrD0CVZSog6+Viju2kUh
49Q23eGb+t5vRiroMYXA9mef7wzJMRSpDFEL/BXbZpxPq8mqNpgumPSfyWveZvGn
h/udrBllFSRKlbfwr5AbYgPjlPoD09tnspO+JUFo09iuH1L8fkUY3Qz3OTTP50xA
z0v9a1IlLmo4lFK63R2/4TIkbzABy8XTdZh4cL9rIpzCt5mFbQMCZHadNvFDnH3s
zUw0biAhj6qSh+YjhMggT3bEZIDj2tG6HAgMqerAzIqwnMyMyduxFjFc5Hu+l64+
9wxlfiExZdalKBfXJIbvZnnggzF7j9B08U2HmM/Fw6qMDEZTHJMXIXVA5zz3iBxl
YZ5a274PzHmrusbZQp5J0ne446vLPRmfV8nmAhBlBSmiTR52/7X7th2JW5Np+Ru3
cBxLBbSpK8oZV+5O4DeWG3fLwwG4bpA3UmJ/wmknDe9dGA94H5FkLdRBEPgURqNo
Obtfva7sFqm4xhSPzZourBBYmo2HBaQiNrrFndvpduK+kK3ZBZmaBpwGFHmIvEWQ
2cemuy7V932jBWZPN2xJkEPcX4FiiMInq5YYe1tiwOMyC501waH94+XeSFwP4ISa
BCDX/vwVrPp+MgOpL4KPRWjoEsetYZydfsmQPOE/mIDj+Ks+bdSG6Arg3DUsFIw+
KfQgkwOBAbV30MRB8i6pwbV3k1YuprPD0RQ8WFzAjyYKnVFdsQhJqyXrd+D5xNn0
LUX+OPfVL7oEH5IvfA3auPqTZVRj+3CSXzAIj7USGl8lqU/p8EugN4I6hcG8KXig
pZv+VTcfom9+ZrMt00xt7Mxsn7Z0GQ66LfnteRM8xhcFM0G7r+88AKg/tzCLKyLs
Yq4LhOe5727Wn8S3se48zYInqlmHqAj5P9uvByYSLqCKfs9E0AZl6ry0YpmzSnwa
TL/UJ1eK83SPqVjOzhtPsHAQ8p/ULEhq4mDjrn0q5tkowv2aEH/JLBzMJLcsA522
T25EMp4oICUpfW1iaw1SzJrThxzeJsEU2GG1z9e6jdyzqcnR2NOboeyad7I/0muh
MGBV3GC6in17hyk1pliX496AvK8l9LlZrcnLSg8/Ur5NyEi/O4L2rAELy+a41H3L
MmJJq7tZbENZxKBcPiKmgmd+p09EB2PhNCt2QIOwBO75+D6sRrAlT1kDG3sW9nhM
fUb18VJ/MkBoNUwemJgHfaJWuXgpiCAAbVxaN0XEt1fVb5b7poRWmpd/YoNjM6gZ
V/4nlTBTn6ZR5r8Vc2yQcW7LsK/GVoip4EylCheUxBmKFZbVv3nrTmCXJiwdpyQh
BSqumjPs1+RPyI4u5A7H8bzBmEPUWll7RRBQJzCt/LPho2X5gyfbNs71457tzP3R
C3OMB3EI/w8LUdwEC0NO6qQf96vUSaCCt+jwMNEeKQM3T+RV/+Xcgmaikq49oazs
v7p5FD7Xo1lsimc8zuoXR3Vo7u+8KIxtwNEFSY8DTPt6efOlXWkBnVPjXdgqH4qc
TfvAlnI4a8WxxSRoD4oGS8JG+T3CIL5nuTnxHvnoZk42VZAn/NUq6tqsLNlyjivM
Wy53nAYt6MuozIkPH7dtvmCdjSoQlmIeChfyjQpQnD6me4CSYgXdSDgQ9GFUrvcB
U/20p/pAE5wA8hOfnwgKxJpgn5/+tzlGwFfgrAN9tA9OkYvT9Tu9q2dyF0NPU2im
EQbMasEfRk3itrdNSNHBQ3LLJVltXD3dup9q92O1gCmpD3XEoFe28UL0FQYyckoh
Hc1EABepx/cYJlzTWPu7fbDztLl2wMl1/HU6Ukv5qOZnM5S5vCMhBgINt2Y8uPBK
hRI5GKeIYgmd+s5xP8+uLbpj0EDM5CXLGYmjH8PlF+K6ZbWzIUclEh2fR5kZRJbi
yRqeVeJhz+EGBJieIPRFMhoapuhAshFKq66wloNfwwP0WIzA050LH8kajMe/AvgR
gQiIYGbIQIyI2faDjJ/XKKpHnFTBuHHEJWYFdXCmVj2/RaVvPvnPhqyMl1pqFXs9
28gUAv/fDW3Fz04cTwfPk+cgwh98YWv+eXGw43i4UisKFdyJJiLFFJRNykA7tfbm
+rgcj971TOAaCJ1wALKkyk0aFh3aD4KfW2GK+ohrOxB2mZpwsqBSDqrNCq627Qd3
ine5/rc6DVxcvTpdf42B/Z2Zls6xFMi8hsxW7nmlxu/mNE8a+GhFzpZJXHiaVFcG
YQid0vMAlXxCDZuMKBqNb4TtK2XCvCaeOPd7YE5q8VSxvf+BqFJe2UedzmvSDmp6
/DWmJoM9dBhnabAWJr/MNAl7iCiYjioTOAR8SsOK45ViPd1Nqc/sdf/R9wmlfkcv
tjryqGNGeXITdmWGeWuqB9KXq072yPN6nAqgEFyhRksnO+NBtoHa8m3ippMf+33x
+kLIjyxHHVXlCoypj8NYPUlw9yTepL54BsntLiL9aEFPMo4kyrBSep2978A4j70c
CLt1mjMMnvpDguxDs0ZmpzQDHrDwSeSUzpmPdZ2Bx9HNGpTZUGqeZcDPk2jfIMz2
87mCmhxgryGplx60tx2AucRv9WDZFlzxINAJMwTDahF/E6fM1lWZ8WVFMpYYd7zG
4XbyVDvT1iwzn5k7sW511QJQKgQnkQxNNRlLEDNFpkTusl9qqqECLULouS31mVq6
r8ZU06jc7fi3gCQk/nikdwRWklv9LprnMVIbHvBm5Gt2J43YEoNYeDcjB9CHiMII
wlj75ODxjeJR9BbnHMJJ/atv7SAJGwfaXM7LNL8voVivNH28dj0S2XwkXOlUdeuo
Eu8tJmluaF54swqqege7F6/Sw7TtdQYKoNDQlZvM3Da8AkXh3A7Rt5BcFNk3ZpwA
uqsU0c2kWl5PZRMCKn3hUGi9gmBu3FbI4YD4ZQ2vrk01WdQ29MOv4OzSwGpiakFZ
K4196R5DH9L2Z8TdpPaqEYumGpmMGhArwkbscuz2rykCRMHWVJUk5Ww+oQJ85lKH
9+sEJfaeemSj5bTDev8+WfX0zpVmXIotSDBvEWNq19nYUWQztiA5CWioSNFR3kOZ
9H3vHpFjAr0T93clnPBWWnhJYmZAheDELsqtkEJfU0vKsYNE9Vl8lv7KMUFy19Vl
3JhBZ+3nZkHKS6fRP5at+dF/Z9WGTCXn36neJSCuuUo36yWSGnm+QFgVzHjGvt5H
LrMFdIjZUPbEN09F7oyV/8VgHLb7mfWsZjbm+Ix4SXXuSNJf2Rs3tbr0KxsSu+TI
EmLwbKykr3iwar1a0Y9FSGZ8j75IQktDzxN729lxn81QLVdiLy60uOinUWr22avS
jaHWC1TgBbz8FMI2APIfV7l4WTkr5Qe1kJitpgCuVy9ud5v/+mrJPlll5NUu9/HS
UFFLK5aMzsjhg/p9LeUzZVTvaY5hV7OGZehiTWwOmeDkv23EUvnBE/XCgJRkC/fy
0iOUluDmcwccORBawOFtiUnPuRmV/fnXJ4wE1PHIkrJGNCVJbDDuaRAzSMNcPJKz
w9v9Mv2S6AJNf/3LT18q/Ncf1G8iWUrkdWtjMF3DnFuMe+zRNKV5ggBknE6Wv4t2
1cbNP+qP9aMn7amGyrm5gZGcY2/NW82KaqwRmFk7ueOqtBxOGFLpQ8bctK+4R3O9
89AY/HEA9qqyjcXbI0ivH6eKrAqYUPnF4DR9MKbLYoC9+5NhK2OPBd722u7WEy0i
9f+91JRi7JPfgKEp4M8N3LlSrHngwfMhTgToGM11+h8Cg0wH/tAMT0thDXtNCmYC
gHIJwp8uRZMaJ3lNK7od0eagEsHJiLU1PwVncQKPedWmbLXasu/8ZpHxkeZT7mYN
XqxFdP8Eh/havTcD208Ab6EHWTfGiOnpoNgNWrN2iOGe5477OBZFJr+zCCfuEWf9
/LsImgyuCuLeJQTdfrAcGiIV2jt0w6l6xDVvEkRBKGv+r3JLIDaAkmgmh9DKtZpM
29L0RgtGhCGtt4GH5JsEPzFkbpAtvq+ZdUj174UAx3R1LSFfYDLvPlacpNc0FCN0
T/jOis54crSz1igEWAEX9if/zOsjQyS9P4dGO0K86E0+1M/rLWMCuc5JGCuhoTiN
fwwWDNaxNbcRdrmmNe6aOeC0rU6fQhVDhzmyeqEO9sMp9duoHqxuq13cSqJ/3bq8
TvhqyQ6q9kFg+68h13A7vkdzqwEHsyUrKniS90FG/T4SN40fIN8TGpBHHXIFjjA2
ObBh3EO6RCZYHoOl09u+xIBBOJQrMyL9cZgSbFUvq9JAxODF+N7dodFqC4nN/Kyd
WZBzZAS8y7I4Fc0k+cNcNlp8wWwWZIydoRb1rMv/pF1Ie041TjUj5gKbZ/JzJEgG
bDfUMAYDytfyWDl0bphZh7TNW3WhqCXcxjXgf0i0VOtjoMbco/KbM8Z8DLXLq6nV
Gqr4YBrs4Zo6Afkf0hc43+RxbA9O3prigS8SF6NPfghf7Ga44UiHo+Rdup1hzVxJ
Juc+6B5HFmG2fr1F4aPBQuxU4kYc97Hup+TmQcqeEXZNQAJhrUT5jUxgbXp3S9Ks
vrNwnFFF0Q/UcqxqtVi+734Ba96kTEv5ppfmGoGLr9rbc/mWM1JyMJmLz3iop0ff
/ZsengMz220HGm9fHCour6GBdPrH8mPd9LNAIU4p05eHCPKOZJamfj9EWySfMfe+
DTyixyiSoSMZNI95nVzLwEjAYVub9j9xvLIlxBW/7dNVyK4la58IsSlXl34pvi//
HmYrZe6Hi9doxp6gHAidxSE0ytCW4z/di9QZ7qmHR2BRa8an3KMiYH7M8ST/rpFT
QBfE3Z4cz8uLSHBcYbS4in/ZMkU3WB27wotUn8sPGTrLQNfMUeYRnoiiX1qijWhe
NJCf0rFaea23PNoDo0szOTvj7UVp2u79tPVrj9WRMsxvS799wIKvwxwe6d9G8bhS
HRbqHoViNY1C1G6MBK5AykmvPnzb1AIUnTmYAnf/qTzu89lL3X4a8USA5/UI/lzY
g2X7iSzwzxpVga3/lrPAik2r/+YFC1ZlRmyDPXMvq+4=
`protect end_protected
