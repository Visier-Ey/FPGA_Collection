-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "N-2017.12-SP2-4 -- Oct 23, 2018"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
GW1KM+eHPCWjVOOAwrnFey3mxQaR7s1MpWcMJeTODSe2PsmyyTYPOGE/QvamXIZ9
Zn2ywx8l76jWRYuBjqaJDH3izEvY3ni1Qthpcwc+LVGfuOvqPknZg2+Uqwyn1ewz
NJM9sNBLGMoyl5uZaL4gPUGiugtSjERsweZRhbGdgUw=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 7712)
`protect data_block
B8cDTdyMZ3G567WcqgL/iXvoI6TxWeATF2iiiEB85mkp+N1kNB687n1zY5qsdUoy
YNV3AWI5dX5K3PBjaw1rtaLmstcXfEJ0po3MIiH9pNvmSRJshVO975XCw2YlgQYD
MvXPfuwLemld7s7WH0NcHO21zRjzq/+gvIPdxH9d6fZfQlf6cr7kBWqLmMaxjOSc
LE70Xlln49wSj/Nh0QJWBszBOK6HGT7gbrTlHAiT0+T42M+0mCMvDNd0jYMhw9YA
nuC8a0DRxT9kg/y5cKI1Dyo2pEZ1iMASxLnEk5JH77QZMKfexJ+i3DhWXdc88X6S
iCtZW6qg4nyYATLNyebDzCxZkh+KAaSadUyiZ+/8UF/fOVLVWbWz/Tehn8tGKoEC
rD32bhIvYdEsT3Cjly0+pllbBrhaegiV19oSF39x+FB9BHgGqYRQ/z9jnR4Oamme
ksE+thc6X5uyo4RFJ4Lp2VxOTALm1lqtlntWaId9Jec6wU6h098cPkyU0nt51YBt
+2O3ZioD+2rWql+ILZfeV+VMtkryVCIEeZjl+Qi+3cZYcyRjVsYYyzSefIDK17Kl
sqacH1dSXfu+cGj6R2e3UongzBTfWAkQwh+qLCF5XvDUb42V+XXTAR6zR/30EzZ9
ofoA8Thlw8Xo71aA9/AmrWkx2tyKPVNA6Q7WaPic47s1LmvsHSRHS7bndk5kqz6h
c4xGryH0eXLmjDNWYSMtosk/nrUKxu3UpydYXCaPxjYDi/jJLKF2SK+hxDMY/ou6
u3kAlGTtJ6g+DSB3nVPfaB8i3spzvMQuZb+czZrmkC3Txr5yNacL4zBgaLG10GFd
h8uEDXUq8vuXqHgcH2WonAErD2nQcIHxDafJGRIseF/H5qqx9fGKcklZdZbtlIAX
Ci8IutbwZiONQNDjbA+ZGNFkphCZoV4dCkQdZZlr4jYBJxh6uhB9h6dJ1DaaFKGu
h1VPzlZJEOR7NAqRUnnqPTvBEl5PXX3/VPCgWDB25TTMQSxaMIHD8yUFigEBTzCd
W1vOMfl+8qANYFciXpuigTtUyu3+E/Jf6FxHmjqELIu+9uf0TgLYSYxHCHaJM+DB
FfgA0tBXpcoTI2Y/lQ0Wo3wBEixtnQV6KqHfkMHwguMSl1ifKyFqUmXcEterzbj0
yNzrIUxBT6YwGQeuXtfdlE7o5WCqdBRSGgV6cszdG4XsH40u9hubTBeic77WmKcK
3v0pCNlVS7OMqALMG8yGV6hEB54DTtvWeA53I5SuiUB0frPzRDnBbS3CnDpsA5sO
DMUnTWWyjqonA2f0twlcvISmID+Uoxur3kZYOZlMNXdmjQvxVwRiXwFb+sKGXARM
R+icG/pi90vQr+pgSmgl9faKwugPzPGL0/LwTEIu/LiK0bxCtStN39fzCH5vk7Pa
se5QnPk4FiHN1zIDgncnganWqGBcuma6YywS2Mh+iKGWRxtysJhXXPZFcEiYhgnD
SdTEAc/2P2IHGrnnfTYqhy5mc2ae/fOn9QsewX2/WwuXWgBSISj36FQ5q8UAEyNY
Dcx/Hcbmq0hzSyJIcX2a/6ikG6NVi0DXCdDoWlRD2VoO2LRVPCNpeeO0nAQE1WdD
0BOuyfkSvgW3YYV2RilQuKKC29IsfJqMwoQL4fQApcqz8OEBpePfA7s4cL3e6P07
0oUxY0A6b05UTs6dTmf5KbOYJkgfIbK5pdJ+QoQjOjzH/ode5I65hOFRdHGK4yoR
A3+oEOX5SSTQLZWylF9KkgEci7fkVS0WvMPXw3+i/JRnun+Via+SwOJedKm/JYfZ
ZgcmlSoCNl0PI3eT9RUqxEHzoJj0SmjldCBaeVehKPGoxkHPSEVhrX3S4nTIPrCm
Zbv6y/kb4oS5i+8+t+u94TWofEAp2gXxrUd2+xH/dtTguP2c3W968j5EnM2Wki9u
LvOxnmGLZQadAQMHDE0LIKwjw7Aiz2CntFr8T3eS1WPurXaFQMldNTTQrKDDie1f
nJxjjp6s6fNu2hfR5kf1kWo+Q1L7WJoQdZwHfFzs6H0Mtzqw1+ux2wZr4NkJJ5KZ
FyMwjoYQyq7O3xYzgu2aroZYVm/PpYUVSpuqgSE5brov8Lp8TZPbDdnlECJsbZsI
kYjBvyBlS1N2OPmzEbzeHxGriCU7rRF0hoWS4qoHUExU0dKVR5WyrhgCKQIg2fpy
0PcH9VMkZrAI5dhLNKapnEPCxb3QCywv21PwYJodL19qWfH0SowwGELVjHAtKTBF
GHgzw7IPBZud7l6fVKQ3o/2POegn2nIuHBQpwIud1bgoGLm0MR54OoYpxLBqK3Lr
g5gMI+zPQ8YOwILrwwx+Bxdxp/VFcb9sSDhZgeAB4/3T7nshiuUGffLsHHtAttBm
O1pomJ/DfznAMr0HSjBAGPjDTe7hor4+eX9IoidIjp5grCrrvLavmtL4s3U6v6JD
1hGyu+KlMRyCwgrmDnMxxA05tTHCWMddWCxRzQgdShGPDwE+xemgiherunefUrq0
Kjztfg8fY1mNRa7FIeRb9WaQX/MzMuTuFo6DzjHm4KoCCThTQ0hdX4TzCcTA/H7h
BC6o9isEUq1S1bJp7HQv0crsFytectFmKMcP8E3NO2Tl78AAJ8JuUIhgnkmtCFF8
R/SUj5Sx7FvJquPT8xYyAaBlVOU2nxG8glpi+lw2/0Z2AjWg0iOry2c91m61es+J
SfynZTjUwgblcDq6LGiO3px07YzBU9zmiccUGZKtstTjVUfkyqTW7GIdimAVQdXK
E0sLLew2w4rVe9vw4FMlLm7GWGUjVwZh92WjBN7eTgEV4cbGq3wZIye2EbK+Ja3m
529dB3V5kU9Rory9v9AN+XpZ8/Cm0AnREvvE9XJIYHX9ea5DjX9E/EMBdAP9On7A
gwjlOikWMDVgidwVc2IaRItP9L3q7GSDEjX2OyUWjhKpZCLXMTSFQ7R8x9U/kMhm
DfL4HszQPtvB7Q8lz5j12n8/p9NIDUyMccEEYySs1ggCZUEMLXV+ryirt006Gh2v
ujzqydbIBn8UDD+Kyj8iSket8fdALOWbjAxap93mrGSf0I4L331xitlurZDYEmuh
bGofr1napk0NmZoWN2WusLEnHG4hBhiZevCSouT4DpjJ4v6dH5m1GG9nB/kMpRdl
/kEtzLF6VYcaTHsgH5kMek1ch/PYQmdFP3MfOfoqqVPUAVMvYfklGfjJNJd5FqbM
ueJRyE01TjYdQezP78B6wHFWFzLgdrCLAn99B5CmF/EFgDokSkME0aOieg3GseS/
SGxNlX6jfC+gCLYIGjemiRp1aGHnyDJ5Mb4Ipc8fK/la5UrrIwk3Ev8OdO7oN1G+
hgYBTwnP6tKrLBrhhmaZFrrt7hv4oCBC7WG3h0Hz32Up04IYjRynNAg/kM5V/Ot9
W2+Zu5OWw/CY/71Rs1utKBWxZEU5iTR0FMFkKJGHpPRMEkOAWEEmsJXI+59cDy18
R73mzhIhxMl+662BLLvjgjHQGPx/W1qUWlT36T0/9x3NFk4B2ppFgX/psLwKUjER
2PZhK16CBqODZY2ZQ9NNTuNRl2LQec1OkEfjydKPBOH6bBJ/B+994e1LwUWEtOcK
ad8cR2wI0XQ2lBuXW21+FmLyJYPGymBLunCIpYDo/3rojtjJGhMNpupJOYEr8g5Y
7kjqHKKB6asRVPE82nIwro6U/95w8qpUnpTliYA28kyf5M+E+UU8tA8jzc3j0Thk
O81mGqS2kjg5d38zdcRPl/fPeT/pk4+GpBst1DHCkuRU05WYWHs0PBiSGIvdrrEE
E6P6ZrBl1oDnW/rHS4DU4ZKwAE1h0LyeA6CcAU9kpVvaDWuYjGx8Yd3L555SYWQJ
ZlTt9GSlFBIC3pUExRUekgOtmsEbMkIYzZyUNRzU1/c+/xgvJEeJOQlg4HKmWvib
Tp13MQT6m8mE+EbGptw+kjc6YnYCnPRZnqaWWdzf2QK/D7HNRoyJh94SSOn5q0nA
KSQ0AK93c7/FA5QST7rlMn64fs8uoYWRXHmlDM98O20ZyBRKIEZN18aXfDX16CpK
YiyFGS/9CU0bcSUR6vOI6arsRq0mxP7Faxb86ZvPgAZ2wNEycz8Zgj8/bz/Ck1Jz
jzAFWqxyelpT3uw0HMpvndudZuezKlfH/nU6gaN7RrSGSFBPkmVt/l5Lc+xSqohM
WDXgFSEhLxqwX59p+NjWpMvRSZFCbDufUeIc/N7Jk597Z0ZTIPOZ1S+QfMfzy4us
aZGeWfHTuIfu2J1HbDSMrelcqhyJO7ncuqgFqsDIpnHCW5Hjp6+voXrusavHBzP0
K6vRNFlBYMG4CGshRJC6yTEk4wlbZySwtqgwYBrsSxCOZCd6pZCqFCPbclTZYmta
HrXywncf1axHtxSGCK1oEWYwrtVYDnuEyfX5eOos4FCS5zA3WYG0Eow0c+bBU6vA
d50XdG7hjO9wL8uSjyGDHZthsDbA412UzuRpiCtoWv7U1EviGoVWjKRtm++aFp/E
Y3qS22yRl0cjgZNzGSTIv2oAniwP2wkGSKDTp6CW+oOYnersItf9257QaSZPxrHI
GGPvrqv671+BS9qIPahEn+m/kr4ZWwpAo99xNSIpN/olnwKdI9eIUGDZlCdYSQ98
GtgFEQ+onwLDK7HZD4aoy8KMZ/wDKX4zUKR4w29wrCm6FGp3x1T0gWJ9Vi58a5Uu
Typ+xuYpzGoOLuBfVT/IEOO2bbS0RGckbboIhdzvEPZJn379e2MtGy2N1t+gEgMw
biG+k3tdMOF9wk7Hxba4og1U7xKq1NY+dw3ma5/PE1ggUYpTlKvjGU1mlJlXBlcw
+zUydBrw13zXqKPs4qhisPpE2A9yFg30vdStxE4sd6YP8jqtdhC4CAbp9mVJHw/n
OkLSbEWjwYyT3ubWA5X6vp6nE/i07fxQnz2e4+naPEJ+QzVq5XEJSxrfzDZ1SVWH
NbiaNVieuTqGYg8Cr1/P5YWT+IOgSm7NgQQU3tG848QMUjO8bcxPCx1F9gtBOpjU
NlIdOqzAo6czz7iIIPiu5azVYHKLdUtAjSeY/GE5idStQv/0UqArHxDeJCDXAAoU
boDiu8Y/0Xz+M0giPdZ4T/P26KXjNGU0hXK0EIowY31sHyXOOHT53pgJIO6mZfSY
KW/Yed/e/Bt989/9RrxWfsofi6w5Yc5GAstyeWxC30VR7x3njhnwdeBWL2daK2pM
DN6ZBFLkKoIBPXAb5c1YuPXCVnED2u44LnMUKqrmZvcv8G4RFoJFRhtTsy6E7uO3
5tkHjHGAoQLPf3tzGXe0Fo2UGOrTPtfZdZeM39Qubod4Vj6WesyBQwocgXG8vcnC
oAuxsCR6qrUdtLpo7aj/qPFvmW/jESQ0Ep1y41AnnpFKVJkZmynzf25crGYkhH7R
rWlUqGD1Nh9lOj92m/dJF9oxOWCEfyNpOWt/kefJEiJuEjL498KgDmReq9QTTpIn
XLAQVh5IAqrc7oDybohdtOp8c1ZSVUsWqIuVJ9PSbbnhLbM7iK17Udr+rLtVlBEW
ks89JOrU726SQ5QDO3uopw1CBlNYiLgTK0yHO/HbFtNlhpxkzZWnAb1uojIcJBRA
Yd0bInrDfu6dAv3Ez09fEcIh2BIqQCd13OlVpJwyUwkX4q0pmsrtRgxVhg7dbuww
0onIGvdlgWAOqkkGf1pDLeqdVIcWyKjUIXO2ffI7nY8eJrcd8BHrMVvjQU66rP0e
6N0hme4nu/TdhjmxXJHhtuzaaqUdnOfN2jrfXVHDKD+C18MZHC0s1L73mFuIcm7+
vul+Y1LyUyTpw6ht485t8ZbrtquEua2xBExUVGfltNbInIPxVjD/Z05xMtQEoaT9
zYYMfFxK/lz91AwfWfAPBYVNcQL77UUSzr7p6+QBd9SQUgu4CtwgEIw8N7tMLlnT
acUH2FAdY3XzaWXVTfBOL74I+DnITXst5c65a7+PheK74HZmKnpqQEGGQBI4slxh
UvTdUFv+r/U+uGEB4kLRY0kKCKVRvZ4+DQYmicx9DJu+sSiiI9Bo5Wb1oMaD7lp6
UOFXw+IXYDji2HidE679xhdgt0L3kVEOT5MwnqfhMCg4OD4KcGBoQGmznWP5F5Yj
6XQVCNb1j/6l9sGkBAvN28f2c8uRvMRf47yH6OL93jcCkEoOFXUO0XT6F7YOSU6x
LZ4ey+5HiRMvd/pjkIimrryiedvt4Wa7Qy/AJ8DtKwniKvxNSvhYHkN/O8YSm5TG
QzD7HiqtpPNSKQFD86JNzp9epeZC6+2mPT7i1CDdkHgfZBmEJLXJ5KrwaecyMz52
k5it82pCKqYKdtUfURbU9Bav9X1AAWC5+A8+SUiUkF3pL9Qnw9IRJW9zA9IP1ven
1n6z9Xr/2499gpDLNtv+uoOpzcfBxmHC2RKAhzmjPhHg3PpEtT+7pBZ2mo+PQhb4
Ih2uhesPi/hgDggPVJdsFeFZW5W9gYKSgdYFJZCtulq2RJ17SY4roXdaUEtJcygB
/Lbaq0Kl1/9A4FPKTFwND8d9SjqYhd4cxQEPQCHyqtL7WTpL0Xcmu4GqGf2w1Ph1
GD6/p/bB+aNoS9BKb3+vCGFpd3B6Xe0N9XD2YfSB0hwCCG5QXSqwQmHVZWqSsIYK
8noRSRe1Ud+u6zTTKjXGtG0MpkGe1GRPu9Q9BKUKd31nC49EhkKO2rVbCVCWXhdC
nDZX+E58hs60Z8vPY5j2VHZYET6yHF7Qi1wzynUclY29DzGprSnaMBHMJPIVG38B
na/XPktm51cD0HQjr6BZAGZ4JrUWn0P6w7TtSLRQ+HvIE4lyZdyr4fQX98j/jNfj
jg8woL1EoxpiFuBX3rsh7WhhaSzbTbWP0BxTV1sCinG3Z8mGNmHl9wlefYFrZyav
9cYf0SwXfioQdm5okPiXeRKyUy4YMgCLKB2vPYLLillNSD5stWYhKnvoFBFUKAkK
2dODMWpGBHCmmiV//dozRly3VLyTB42qiSzSEUGo7sO3RNIJE+1eMhHvgjsC06Y3
g5OO3aILKJ+1/JdrNx0GasiHM+3E4b3EEfsYpnPtz26UUVTSzaQ0zYn5c9207xcE
ciuDLnu77zjHnof3WcLOjDbGa4tLvG6GQFueZsVQNy8u3OAAOp8Wf27WJkyYBaww
j5u4XOK4JmpqbXJc5ziorjYKCBmUGFPbo5Aa07+B7ZHmsWOhSo0Fmb/uqGKCjZ5e
5dIYkCNF9WJlhtgKufWdbspZUXw84KjgyTgQpR2IiCnDxM7GeEHro64Nl25OR3Sq
B9T4VDS3fK9wrRyxQIQ+AW6X6Z6Mb3QLlle4eWBTapeoHeOpRFLYE+0H9Mm0t8EE
3LuC0zgM3Sfk32PY8wmfG9MYy9l85PpK38myA4NOpXdzI8f93iOX4cyYFFYU0+jQ
ag02PxTl1lJybAf1l+D7o5dCy5iEnGqB44dO2b4LlcKMq4BE8Vy9ZGpQsP1F3Gzw
Fmw8Ibnx6V2UB1fet277dSmza4YfxXwwCmvxw89fqwTCsgHN0wzX/f0yelXRwr8m
aUgh4lISYmGLXrz7wnp7KcQYbeWCP+uzfgPlALK3FkROJjIjCaPIDc+H3HMPU3qd
0Z+Acln6mQm0pdkUdNPfEoHQ/jycjkVO9wNIGtYyzqy4s3ZeH7RscNMFAGar/xmC
gw7vgkZU7Yll1McsIeVaaLo40i+d+NUZ3YykxzEQbXt8XmDqxNu75aq7tu47e+4M
Pd83kjID4vWzArS61EY17+o+PYUkWPgacF9SL1b3Ci2Ml15wQHz+f1L/CV2v6Jim
L5NznCeyNzRH4ggNvf4HLL5X3SBRzZJUk1o49RR05G3XHwRtqZRwVk7fxZkM3KI8
e1xFJHsLKf41GM+nk+NdHVF8YiK59OB4XNnus+vrLIW50iY8lWdSz8FHPGzy/XpU
1biXN1vaikiiUKZXkCH5p82oQic6DNPfo4cdOIP7osStRsIWfzq+8Kz4BtRMUBs4
3zg6TKLxYEpN+Y2Oab4839PaRjpdxUG4KN4aK75o9tX3g7ggIOGXAQZZchFfpd0N
jatyFJX/6hAbgPPIHkBtqkG6bOWiVXeNBDasHnXwOTtbWnnV+Z3MiY+ASbydtOgn
FZd9wFFJTC1W3tnF6Eo2KRBydSL4LEW5m8usGfpMOb3UFYaJvpcAPu4IRmb9jMeJ
2xfk90t6jhg41iFssVPduu08JD5lewZtV64rNcey55xBFdxbYLrMHWobG/ZxXf8S
x8kfhCRrLkFjS8ebB1Oz0ps6sJBWmW7/n86zlA0r2DviIbTk+MEROXnyQYzgskIx
CDzkDsfsj7/VHcTjE8k2K20YWaxLF88jXcjG/CtFVJXvj2iMqcokjUbexw2LMrGr
PE0WyZ8xSQu22S3t9urTdURxHEg0VBZxiO1KrPfjonT8g23Z5C9VLlCkK2fsqRaq
tEkbYFby5AjfB2XxeMXnzy3aRmZeqwOvY2nkd6GAK64+leYZvVJMgk9NuGQdzpSE
+fim63TvcPobKmLUVMod14oB+RKHsGTNRsM9lhYnm3mgLslDQaHmAbsW41ZRKJQr
XLqBGvL7N7Rjphf9Kfdy4s5Jk0xhYm6FNq5OKfKMOTVNlC3aid0INPQMUsTSwYUG
Tn4YW6U81wIGEwHtgZtB0ZGNet/dOENsDpoxcUXrib4iIq3ZUSvcc/ivUUEdEIsT
cceFAKR4Ja8T4KNbtAm8BkmPAIkEHzAw4Os5tes+YYIrrcnax3r7Owdee6HO8lQK
t51NMjzBT2hRO6CnW0+FE3ZrXxXh1dLvpDRMZQ/ZDVfpMFF0xDLYwbnBPC93KVbw
pgzqnKpYTRfiEzZVTgurs9h+pnDaL12Wr6a4k5fy/lJqky4v4gcFY/1Y6sSdxnm3
nkip6dK1YQ/j+04Aq/F80SXcTP0ANglSMamb5xuG7s7Luv9LIimU9j7+hxBma0wP
n88kZ27+NU1E24KSV7Fdd4wDib7S/UybGpBbN3UjWYvv2dkYOJbX1PrfuFa8PWhu
44nReUWX8HuJk3wqdjs7m//6dMGBUDrQp9AZuU8jo1mi6jlldnP+PkYozlLoJZa/
68UZNpVpNI9Nbr1sZtuaN24a9UwrLminlTmgpGs61IFPHxDKzElxOeTgfnZrpa28
d9st47kNsN3Y0+zWoZ83eA7Qtl/oH4Ny6MbjCjXKiAui2u5ioGeA4YA8UPZl/+1l
+iHC4IDFSjQUGFySHFPi+oQuhmmIFqhJ5aGGaUrjw0p4U4+Ro+HzgLJkU726JWF2
atNahSDtkPp6UK6GndzbVKkoBb4TvxbhiXkY8eytVOZuU99pyar8qdS8NGT/3HIT
EkJ6pMxXd6GxKcf2gB6gwT+zqisR0x/NnUbj3RyyVRZwzBrL58bjp+gpYH3jR+EX
NFYS4eo7KQas8YKj1ysctmg2FFM1Hn5B2vTg7/g8Fl9Jo75GKzqDQ5a+5hJoR08N
1qUICbM3XazdK3RH36EwFA8CzxuYZFT7KtlcNSGc8fgLM+xHEqZoSjAbryKIKi8G
X8grpD0zhTO9CCyGvnnnvIbK3ZErWX7P3Op0zyp/CHuwQxFJ8a8r17bX2A68htY/
kQ/zEuiM6RU6aqdYxgTeltBK+QbwixyX74F/DCpzmzdKRzb/egBXQwk2RIfNp5/+
5xqs6lmapRm7oDHJ+XM0pUdjgYTXNk1D7LYoGkH488e8SbrvthFBW4oIE7mmC3as
b8AeyHGCkyMekgHolZbnUt90r5u86FPLrvvZsBguv72uTibXHPoE23qjMLgmuRPo
yDHzC92fRCg3vramQ+BlNE2OIOT/BMdC5T/AyVIQ0mCv2Rnv0OXR3G7rEyuFQizN
xjXkbLke+Vh1F17A694dfkXfFmgeTDTCkiNeE/dJlPNn96qmzu0X4uN0FY7qaG3P
C0HLEcI5jM8AibwoxdWAGp7hCrAJmBPANRFKb1F0YQsHfTD2aRAA2mTcOX+Uq2g3
a93T6+VQEQM3hbubMTVAkCbSbFZMK0AinfvRekVfeXwJOV1mEo9twpLSM0reUyud
0zKQOUEV03zya1ThmHMKEe32Cg3KBX9X7RqSHm/+vjmXjVGCX10WDXEoqUBM0jh0
0R+4STeNs2KgYo37HJ13VZtiswZyeGaWV6AhXi7GVF/1viXUZfnQHxnGjoElcGR4
2y7kD8MwqFMyTr1XP8EAr+0sNc0gUIo3H0R1AQjx4XcPdTNnV7C4nYxhWP8e2n3e
1CX+iy3uF+xr7k57DcKxHyB7hU/kh3GUkcZ2ZgbQgDZGV6kQZ6PN7N7yYv5Pq9Td
En6j5fTiidulj01ZIR21MmW3gNzdGI6D8ZwZsZ8W044=
`protect end_protected
