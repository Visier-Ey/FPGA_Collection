-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
--pragma protect begin_protected
--pragma protect encrypt_agent="NCPROTECT"
--pragma protect encrypt_agent_info="Encrypted using API"
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
--pragma protect key_method=RSA
--pragma protect key_block
kduzwcYG6ACDDjw8h6ojLM+n5yeMCWaNjjJ7tgmaAoUNP8NrrDZ4ngUqa2fRFZRK
9/6J8BC8Jv/bsWL1jWIy1jVORcXEQ+RZq1fy0jaZ2QfqkzgwDj+qroLiGLMe4WfS
wxjH5Sy0S+vhRLbUn1XmNRy0L/k3u1/vs+dQDGMWPiKUz0NSODjI0aH4biQv6t4r
lOI0iesiKr0TquV7tSIjnbo0WzGWMZKVD3QWt94SOott/I7qgZRV8ejCbnCvTY7d
QynvZKhRkGKMNMk3oyul9UF35BcKVom+iKhqVHNtwXApY2I5tuzoPXliJn8U7X0c
fzzeVt+rrqCIh7SMimimAQ==
--pragma protect end_key_block
--pragma protect digest_block
FGaYvGbZzn/qpvNFn0IlSsWCaTk=
--pragma protect end_digest_block
--pragma protect data_block
+jk3FXX7JAYEc8N1HeDB4b63rgDZKEoeFkkJwbgUJy+seUh/VRWXh7N7Fyycu6aG
+swSwEFu6VcgwPJGb0nPUO38gJ4pxdcgBHk1WX8EedNPhft2R95A3/JTTLBR2RNr
mCt9H4hZyuONbmLLN3vrS2bw3gGChK5x0BjJDaLWDo81bFwzT9901UrA2c0L/e0a
LwfdBl9wpH4RpaLt9ulET2ZLEhzweFVVLF0O5piQnmQb4znBXYSZb/Nw7i5TwH9q
JnZxQl2hLslWUqtjCe7K1P4iKszi+51TlB9varoHH/+SWDP5HbMvrMWv6Wz2QFhr
LmjdPrjYKTLdOSrI3h1n2s9MccrZz5fnNwKEFbuFVje4dKP7psTpyPo5CpIHgUj2
JZl0eb5rG1Poz1OlBVuhk0NuU3w4ZenEhuID8a80fNkFBnrwYZV4YbBQIBqmWniS
bsWmYxlwb1iZy+1/7UtowirgiIoUXCnxe/rMCLFbXgwYGCT/yIAjqcvEbCbcPL2A
7v8EiF/eHPGH0bOoNeg/zK5A6+UW1GSNVhgJB2wCh+UPtivnAhH6b1HMkGhaMNTV
5kmhipOzLCrAMwg3mPlIVKULwDWtRubBnrQ9kibIQDQTVW6V7p0zrwhBKep3+xvf
aJWpepMdnAiKG8kfzAgLtfEEGFENJ11dG6+pkr4Y/SqVY/05KUJrO5wXyW1jmA1O
H80/kpOXMJ+gZ+xewHMH+Yw55Bln4LMjrnfpOp4eMy6nQhjuszzYjWcTLLznyOmX
gqbftxTVcaiTNMQqohOJVs6oxdKWQszexbYp4hDcO8bq29UHb8RFrlFtJUDiHh/V
g83E8o//eA1tKm/CPClkp8VMdvNTaYoZ7wTcJIWTj/S2tOn4IbiCJgHlpNDUqGE0
MBAc8slCarpGnkRuSwUj74q3+9irar1/w1SLNWZCaL0CFDfySalTy8k1AgdDDCJy
tviucf4Z9Tt0Z0As81k+Vvaw3wHYCNhs+G+AwRuGnvcWqPVP08k/EUpIDaxJ+Cym
CZN8cAKNbJlBsG03fC5ozwbJoNP5nCVWVtu0fN3PDIcMmRjT6oQWO1NETlf5T+0M
VzKuySl9MPwzF+N1xmEVY1ZPSYodvIHpppSuDk4JNuJQeLKi57FZd/gmlv7byrWe
qRRjmNY46tEdgqILoaZG2IkqdsNA9ZN47Jyaoa91EC8se1p01KMbzKniUY7yTSJG
tr0SWROgaMKfh7TsFf/6TeCeTA3iKZ25qFQxTpudkPtsXQi+dKY+mc2IY2d69rw9
So+yQTymIAthB95sgHFj0hBENmjLacZhLvklluzaYN1hZth4k/zH8zmbOrIfriE0
i+6s90L73WLSE55I5rojOPxvfQnXArxOiY7zZdC6UsZCyY7qmqFO3p8KXq7TAS6r
LIAFmZTKY9NyEndUbf/NbKRLMlvABQDCRleVGNZh04DgmDdXD/8/n509D6odgzRD
J3OW4Lst5iHZ/r0scFTTHOHEa66FW6Ckc5fbxdJMHewc5GSRcFl3vhVupHviKbMV
D/CoeC6mk0gcfYtnZFtLiqDpZFI63mLv2zgIS4wfBshS3pCFcXe7PyT9RXBjA0Dm
V+Em8YTVBc+Avf/WJLyZ83AvUx7snoadqHivEUFHVGAEpwkS3/YM25ijNUOdhaO9
9G1ocB64xWi1rKPlrj7rUoUfosy4NRxtx4wny2h3AcM9Qey5LTWwe8aZRU5r7g50
iEbiZTfSR/VCLpyPnsA6WlyTcPzBKJ6wmZQ7QWGrhQEOuYdLiDSGVtzXG/R7PRCR
so9Iuf0USfIioBiEFRGMMTIqq2tR6Npw6/J6dJWAt2pWw/cPpyRlsWK+qPpVI9bM
yFgMqdwLtrQA0uDnaB2/KjVs4SI9P2Lf8EX7+mvCH3XUD3gw6y2+LzuxsCZiE6cC
mYEkql1qX6XHaJtNVqolbZoMkNOMttriQued6VPTD3QolxFojdjCOd31SmPHeone
poL3ZH8LF4O5BA1Ej34EqSaSs6867enWvNkK6PFbp0hBHMCUh9JyZ/eHLGYMTkdx
o2q2px0qwJYs/GqkXOj/bxHCmWmlgJevnKl7/L1oWOlOISZHYXr8q+tEZ1Md4rkG
WizQA+KU1N7PMD8b+9VPJ3olNqwj2Z51g+GEOfEmf+EkPVLZ6KFY4nNdiRAereiI
HCTGomJa5I1XkmdR5/AXEi3GLxhzpwlPHTL0MS2ffUYy0DEloCP8jByhJNywvFME
MWkcPjMMMD2kUJ6MIdYe3p8Rk4WA1MiKjFRgmob++GTIL9yECmYxYIhnBX129wJM
XHMzpebUwSTtrPOUCB3aa/5/sITPOoHQnk5C8PGnFfv6nWTHzEYlAbjVoDep/Tyt
79b1HDnVgqDu15PhLdEb53cjy9m+lNemlX0qbGTxfi/harX2jtJmjyrpn2GeUbK/
MZclA9HkgZDR0N2DDTW64kc4VgSeM6Kp/eDugHKoh3A4zxgiryxyrTOK7t7ELvsb
xn9Z4Eh3qjW8/H6AGHaRY6IbEy+lvkhSGSnjfV1c75hsWFIehYItgHuqD7qQvvta
iboOhwCAfYl3SjeImZ61kPOavS2QoBoq+BI02990UYiyr3XfbRWwHbOCEiAmeJQ6
NfPSxxJkm8C+6zfoVYQgCphheGs1kVJRQfVBWCbmXDoJQXiLIrmCSoEkvsqBYtf3
ULMUn8nIibi3CT+GvT79JOqadDW9O2jzZZo9AKWIzzkVf6gJpKz2Kfv6IU/tbgUR
4AFW0TzGLpWVWYcuJIsyU0IK2BFhwJBOozsZPDa1tNbNhR/O9nvvq1ADu6Q5ORo4
Pm2AMyauDUkbS41yAF+lS5Hul+NRqlHKQutdU3Ff1gu0UQDmlig/WVxmq4HZHvw2
5bspB1ja6BeA5N4Od8uwwZ5d2B6aaF/WdsFncp8gjBK3jSr8db7cv3YcZHNaBVSS
Cd5nZ3hzE+GXKvlJTrFxcE3i2t8ArN6AKAQdxi7RW8o+lFqT5s/Ejpg0372NsQuh
VdQGoOPlAzle8YpTyePKyFuuXLe8a72jMmeerxPE0XQ8eX503Xx0mwakDOGL9Fig
GjIeq3/UBcJD6kahf7aKQazMV//MOPlYwXTznTPgmrPGI/OerN+R86bNY+Hg9arD
XR6hrKxRmHEtXsDpxGUDmSrTeEFYbUF8lZL3EnDlcMwCEh8TxDZ2+W3b4btOvlN2
5PCe5NZKUEyb/16JqI8pf05yzFzWvhez1FCesuY0qu+ojgcVzZg3xuCYbERrlScz
WkUJWYeITozbSQf/zKdSXzrLvbiHrNdN5EPPB2lZzMK9Q718z8zxdixdD7QFwBM8
qlBgzn5zovUX8K1A2lqAdT0F3sQIz+JTNnbv5p/WQosmDq/pD+YSgBCYrsLPZmAT
q6EWVcrV5gtuOhaFbVqsLiCg0FqHeGRa8S0q4Yvv0H7NJkonuzkyP1XGTvSmBZ6P
IrCovSLNK52068Tk6ejh+13aZrKTJzRPMPb6/9Pu68/Fh213PpD1xgGSzYA6xCio
B3Msz8Ezqun14QZVuhBjJkO0+diuwGHWScF3dyRhvmQq5xkHSFj+4A6tYEzR0prG
v+gGOKr92pvOyGPxVF/N6s68MVcYZMcfbcNXUUgXEIsYLSBk8jyk1aMKHjLDlW2U
rHgMyXp8owKn6Zee8+F1CK3GnNgjXhkq7Y72c81MPpVmm5MaVasVsU4uU09XOBin
cXB5TSpen7xsUdngoSSOPAznoImxlwIcXSpLoZo76kswzcEC5WgZgiPk0GYvtOr6
BWf8WITfResFd8DwMOvQi4OMhx4h+C4K1jKxAob0m2gylkPUq10bePFHohCaDOO8
CIguxRtKYXju4cPPl6FcNMiheX4cxg/H4X6cy80lE8iaSfKFL2RFBRz6sEQuhQtH
98Un6G9NjF5UuHI7o6DmFIV9kK7JqRiUJ9Nz+jMK/FHxo0XUUAlPPAWdl5lYfhkJ
cd9XsFM+NzFAUV1+KN5Gaf5BSlxO2Nea89Cm+Bhl4HkrzQXGxfJYVLdjg35PGX0x
rGWCmwEoCoV6Prj0kFYk3EMJ786rRBM4BbI9Cxn5ghjFmJOUszGTrm4ZY89Xe9Yl
FCbHlU1IU2NJBuUusnP6dwMtSJ1d10QfH4QuHnZrSjkgy3aLYClGLMyb4sCRkFvt
kvgsfxnXHiIEpe5XxfDNz437u3z1PhCkIkFqCf90gwt4A29Wx08qIosQdGn2jQOA
FHpvbTEKwLt6iuOYShoBKKfW+rczrr5fRq/J9Boe80KwpSteiOPWgU2IIFl3qsxd
O3OrVQ0Zgc3W1fFpVXA6ws60u9FT8JajyQG1VlERMZmVtIy/hw34G0whlHeHEpjw
fskbbX6U3/SFP9dAgLWk3d6ywUkSiac8QblGAMtLhFp1yj339XqIGHM57sT9LcC6
eyJ656N7a44PCvo06QgtgoHf+4ZUmIkaCUzuwT4BIQv5zi6PRthaGXniZY+qzEbO
5rdToTKbVc6D4/F9Z2SxSoQpDFSD2p6hjdZ72edz+In9a+ZtyEUe3oWJENA1KDgv
/YRoVnpfMpKJ20eN7JynQbsgiNNHRUj9HKNlrcJUB8YF/Lox0So5t2WU33uHEWpS
JY4eeA0T//FhX5rfW+owoL30txLBrCPFYl5HVY+n5CNaBiKScWDm+81doIf5hUqE
pWsZcOkchHVGWrzLdquXgF6soELaIT7b44vF+RFTOhIkb/cWmkruMhKLEYLTLhxH
sfcB/45LkI04fwi1W9NDshwLdV4FUu5G+L2MTXmMLrLvNcxrrZ5jgTdURpGCQukL
Zpc5Ol+O6Sy+xxU4+pZO/wIawqhhLmClXdmWpCxMTfJVvNoYnSiwFoOLP85KJAH0
ZErbc0iRKjWxp4UIofJpfD+/jh0HPNiLuSEVlZ5CWlEr3QjDUl5befLwdNNzA40h
9p2TwFNv6wEzUvKSAHYex7WazjHVR6Vu+Cwwh8ONjO5zQQhBsi6bTwRG9ytAs0FF
KEqeCdUPQulW3D8Mf4dGuD6T4a17eY9yRnyZxNuKltvddaob1agX6LiKmZTgu2gV
L85QtKrVhKDiUUzzL4b1L8jTimWakTqOaLp0MUAYjWkX+zLQfZkijFQAWv0qvTuN
wHtzgNj1Fkc4Ji4VsNUW1lOe0z9tJl5BZ0BiOhMy/0v8mrt54Jsr2b6+E4tUtWlr
vYtX6yeHqZ4UdHz48M0SCXN7H8PqxPX6y4phlqQmgmWg5XkBlAvxlNhTYXsi3zY0
km1u+an1kc5brBmpqzNi3STmEe89AKRh4ZFqGqeMhZ4JLIH06mWHJO1aPHVsh9e9
6BFI4Jh8MMpZr6qfyocuzLr8NvEkjcJqHxpTQ9VBaH9t/CsHC14E9EVgZIVGbgI1
CdNPUgm5ZkSiRWpLn8YX3xs59PQK7/53kOYerxksru1UpD1FPlZwvcL1NYfSsq2F
Tn3PQcx3xe3FAizhvK9Ja7k4RLJEaHpiK6io3mbtutshvISgQl7SX+SQnZB722t8
gP8X1s49IKnxkKW1e7ed5LwrNxUFqG5UF8Zh5w/iTCax4CeQXMDXw47gc3dr4QYO
0suAaoJz+E9uopiXcvbHaz54fUrBa2qJI2ZBCXzRBIbPRiO6eVH8UhMWrRLpBhJT
ViTzX0efX75poiAPFXbBrhkh/QC0RROUG1kIzaacCatiEZK3tA+5YCVJCQMd6x24
NqRd3VLvqYXShtFlyCszCG77+beaMbOVzJnbyEm5cWyS+BsnF90NmdVAR8kBnI1T
TNXDRW98xFTam9hasUC26ZcBEQbhhKJiPIShkfNY7UKP35Aecu/uCNjdCHkDbzsR
Z75hhig3tivdkvzfBnLAfqEDAmUJgYG6iB/Rm9ckMCHEafsomLlv/wvFyheJMWtI
gW7w40xxbP2QtDR1OA45fgufnpTV4TnqJ2D37ODuqmSrWBxcE6RW8sxiaZfiljW/
SN7e5QTXMxH3x4MckbABPePBdggXCXj+Wk+GycRD3hqh0NRsqwukpr/fLzUs8W9t
XWcIcNlsnRRN7zoqNA3/jyOVKL38tOy6MKWRazwpK3L2RXOTIXw2FHj4vgHxC1/U
mhgnIQHRyePMAMUoavhi9DOL4yPaxt5ti1/+Dfi3XY/c4HtCpIB0mZN5wijnAQVx
uL2yoZbpAvG12K86kN9hFEr2LriZYorNlW6dFpplkhoBGBDMHz3LQd6RONYh2sOP
dm9pXBvkOftBAFJrNid/tKa/UPOfh/FKe3fUdiepRQExCM2GuzcnHQy4aiFC1zDY
hgoZPHLLWJX6EL0V8ls77O+nwJdXkPb3NAKstWXLO7C50AXEQE8yPQzb6+roVr0i
QAWzWAqmoP8sW7s3sDUKZ0ew/qHeneVUS+Sd2SgUHDYQSEXAi4GYRTe4z+sZlPXc
fRBsNQ8nJeAj3gXF48103LxmrjIWWt/+J9P/A5XAFF8m3ZOiDKbaGcqRbiEi9NGD
WkJ7yTSIMj7OngxfDcvzLkNzWqcd3e6ASg74dKcazAvxuoUB3RAx9z+hgyfqpRNN
aAOIwxDpRoD+4Bje5cSjVFiFKZtrDkh9kNbGzXu0nodvxZpC67eKrXhczwmOgEh7
EGO8xGi2g2nvgirx/cVRTDZEmUxiD1Ec2wdR8rXjnQM+6FwPh9QkGnHzZbKU6gfK
y3a1hOofyNEyV6VIlwT0Sm7qSvJlIpcCj1tJGAr6ec9v4Gak1VKvAXhwK8OwA9Q7
WNczz4NIPcFAfVWK7b6sEl8L+xk6kMEgpLICWjBZ5nVOehT768ceipZOkeGkqS8R
YfnAILH/mrhIHxrh9WgqKtsH/DtB/+yO2YLyGtgL/qZyQU3YfqbFvsJljME+4roX
YOPIaRctfJTvTxANnfB3zhBLicNIbIWZY/wCSsgR7GeeW3Xy14vuXE9wJMYC/GL9
gjksb8vo3QJJ2MDxHzUyHxsJ5MnRzeyuvzbySDv//o+9RdfYsscpuLz+26r2TM5e
V7cRuX394aDtHGcj9TzEvdXKl0JiVVJb2dBBxlvXPqWINXET1e/9iZ1X2UzfIMlD
wmN2uoZ+t/tyhqx/g9ln1xyXZQDL+u3B2+TFcd8yV1k7vqp4w9rCCjcy5GLeWqpz
BfUhHGu8wBTusrUYJKMuf6rfK+5BdZFBrGJDqMDQovA/fpFkdgYOgGDfb4UbeMX0
pQz3Px4e38B7R/Qde6KzywSsMQ9E9xIj5QRAGmkSsgmFeHdlsnEW0UtiE4G1WquO
ps1gh4mCNJgN0r3zuxUIWbdIi3CiYyxv+k7zWqfNkStiyB5a9gpQ3SADWsdIDnTr
LCq+4RuTxVLNPwXgoJh2ieLV+CkdsYrHbs2MWm7t4fs4515kYAtFAFizTEShKoX+
l64N9BPrukZUf2alPLUdyIYWxmFeZD81LIWlLfIzK06L15VTPsPgOX/6x21u+fsf
tURr8rFhLytO4AA5xkyva3EM+/Qto1DBsrPV8yhCulvEge/+vT+Vl4TRTYFiThxm
DkaaFIj/691rAe8ukost80ym/M4yJKavuIf5USn+Kjv45/qSSmPxDHcTlbKfkNem
2OMWwlK3hvtY5u4g4YEfRYswIvKTZcjhoqHHeBJZwZ9DjSzXdvaZ2Y/2Vc/xamt/
pUYBfpzgXfWJt/Ir7r3v1LF71O6K9zSjvMf/Qo0/EFSrUFAR9qTvG8rPT78Rckp2
NZpVlbixtuiJNz/w1ydIK2Pt52AR+7XaemA/KWtHQ7K9WkW4Q6T7KLlCyIVFjpLz
f2joMB4wUu9uriK3OVXifJyflA9+u6LRI53DfkcGqkp3EilAxFgfijpkY5SbwlZt
TOgQ6FNAc6EiZDr+SmLnexFQuUWP0uSzovcHZKzqCVpLaqOhzuBqr/13EwkNGpJS
M9Q1S+6uvpYPhwynowv1lCFEIsOr4kuckSMN2tHOz0neYLz/IFqnMZ1ayhO2iVN/
wTzLHxJY8GpFbrFRBR0gXzX6zkdHMRVg6J1PbyqETQwW+zg290JhS/M4PWw5dJTO
CZOj4ginVk52iB4ZgJ3WnvRn6ns2i1hDzR9vUHfdKd+apeCDNTs04AF9NXbyRtgr
yR/bzu4cnwQIbIZDXR0qxbBN1ITM9nLLFiXMdxw5tGZe8mZaUZmPRtdGR0eDew2K
9Vkk7BT/pYLCidEdwpD5RGeK7/glXl9UI4Fop+jAn9jbcdSag42VBFlhy5ndxpRr
65BRKe1JAfU57aRFMLlSfyCtNFKLLvd10A0w4XK/5of0cdIcDK/1q3M3oGs4RUMu
euxHczMJ0z7JgK75wMJrrKp5IC8tEMe6iPVtRa/N+ihZX8OdFnJxGbUY1jEkegA0
M74JrQrUbiPM7mFSGeugJLJd4zrIVH8g67lo5gTA6JeGh+Ufk8XJvMLEIvHXBtPE
Aih4scfBrIGm9hBeXDxmJc2wT0sbrSl6FUN3eaRldnlWqof9mNYFzPAt5eQHiBU9
rCMafrctufOiOxly3MtJQlvvoKYqf4pNqnPBDAKjwkiS37BzXz8JlRq2GPoCFkdz
VIpxzbh2CV0b4J5S7Qk/cPYX/LxzVkbOfsYi585/rt8JSvo/3vb1sPjikyAqHf1x
7HDFLy+twqTSo/vRzEJ5shEoCCcI6BzsUD9DC3ePxI25YmEAfbm6OrYP2zf87uZO
rqnV1e+GmG+Tb4N7mtLxkTFAsT7G/CqhDHMGIHk8ON2ZMJSpYsRMLZRxtv8JhbI5
XASEYDjrhharbAF0nEiZKt8ZjQ65Hj6GhEgoj5D3MAHC3m40UUjyL9uFLLJagitu
DIQzwY9CZG7y3WigYBKMn1ZR5xouDeahNsf19yQ9zjxUelt1YdOs4oQJwXnhx7vp
SCzI+C1UTbZodtlqEHZzta8sIs4Uo3K7ell6WPiaDo7GtzhfnYA4VdsUd0/Hofqi
saSAdLONGPgTt0qoM1nFR7xZx3l92gZ0UbH3kQI4be1/xh30oHZAPCt9YV3wjk3J
mHBn1OF31+uqwi9Ljn9icZw/0JzJe9o/D+mkZO9Xq4/ypMx9WHDRjvY+t7RVvg/O
2ln9EciXPRExLvimjwrF63lIZ83THjL3XPWTDzcTQ9aOGzNklIwpqWA2djGeGJIq
Rc+NBLSadvsrNCR0H4LJU1u4VcmUq5FxUwuDMcz4/bLNNvA4EbZ9pkwcxgBPJd7Q
qWc+TMxxVcSTl5tzv/VMbezty69y8U/eAeGiaJpRLMW/Zf/nzj7m3+KsbJFdCDVS
uMT7KjAvLIaEUE9Mf7z2adoi8npY8+8f2aEFeCAWXntrboni6c4L0ECRCt7DjXeM
KPCFdcWNRvR74xun2mxEHlZiMb3lioltnJ87GmhFq0IAXSJe293qSm4XNcXuTjWV
tDDSkz0UiwHaaalNyfJexV0DKmP1DMi5KtzwJqDcqkkSCQzJK8/TgYOzJghC5MF5
5NjAhO4NIn35JnONmygLH/0UqbnKZGSQ2LGMKr38XdjKfy8bTJWyRaiDdS18EUod
VkQSxQhhnu6Eo3p+LGGzPnSDWTOCaCwdouWF381h8Sc3PX5FEN6mVXHmNtBKuQgI
gQGW2lTdYz2lWql085GVovGKEEeA4ELQ1HJZmvt2/MHBbIfEXCoaMWYBUAkhgWmu
HByCxxZJGnOr1FdLpXGZpLbaBJjgvMGLyT/c5k3iNv5sybVFwlO/vOB+LaOYlilt
Qwy1HLvvRitfNjgXQ1pGXHObSttq42LTksUFXBOk981+5CCcgE1KAT76jiykFAz9
GqHzClGKiKfuxnS/1q7YDefS88+ef9L6r5KJq5VofbSU+GOkXTNwKljqpKo1IPh1
sYvRdDBsA1IySv60Ug67+UUc3ALj14eeiHxLimY/o6pEObEKGGusvxhY6DRJrWeQ
wmn4r4HTZSuyaauwbNcf6RGEG7Zbpic6JYKDIbqEQfqPt5QKTeHa4PPLFPlLD8gz
NSdonjTkghmtUUyLSYAOnjE2tLM9hpXA1sotxj5wkdwVcuiFGDhKOKWlczrFDtgc
tnsm8ia3S8XGg5BXMKo6CsuKmemnTEeEYA3wUtIC2uMojs8/n9c9thiGbdvA8GFH
On0CMm5y1Mwmq01nBWbPGg9aNn087pi9nZ9UhYZSAkLKCl+I/vYQKyDPyrCuNzsM
tVfISc71J8uKhWQG6xbO5KfjP54XZrn+1ngdFoMfeu8BTwn6d/G7LcfMklkiI+cO
K9wzHWBTyVut+o2EUM3N/uQs712Z8hoX2v6pWBjQrfXF/5RKW1HdmCi97qWLMo3T
pqVruonT1VZpV7WKAse93h13wXkvluXYJixhBWz6ObhenjtDdJgbeL3bS3qytFuS
lMd9KNgJiBEIhMcg0sToShVrgQaqAJ5rZ7MS1KEy068zxNYAbjLdAdt69s7mXrlD
M4/3ZlfHviMI1UeYHFx0rEnZjAqtgfU/SYunwbaozWw2v/pQHPPiwBJ+oI2+dARJ
LgXxat/EV+J2B0WFWhKtQIu8cQOlyDEvbFjv3VQCYb7HX1fQImVxitkll7fljONc
C8FPoLYb2bzSmeJ2Jzkf4I/nJ2FxFTiJ8UKZKUrvdq/rCWKdZEE6ReuaPlXEVcAa
KXO2UOr/iQno5bPzlY/ieM27UWTV2cIqxJidvAsikOPDUKpUbe5lV6H0enny3AdX
C3sBz5asgBjOg1QXcg79CXH+gI+E8JTZC5cwbsIv55LXzCGa1/FTMJNCEZZfpEpx
HmylbG4IArHqd0TbuKHeGTtgiQbHD4ORKkHIe28f7SOUAVMDphBddInD8od1K2di
wduRURZSnCTxbiDPff9LRJ2hp4JngViszMkyOhx8mnrWc2i2iKLbLbCyMQMugQIq
2T4arUHNwUClIwRmRomD71O217C3O2jTjEnBFEQpl1fDSIu6KiL4JrDKAiIBYfpx
3l1Dk1/PT6zUW74cuX2BZR4gZhqZhKQwlc7S3NAo8osUoea+3LXIeHnCtTjbe6q4
FznNYFap1qcznH17mbKuvde77TRljDYz/Dw0oTIfsf0W8oSF/rZde6hUveIumKjY
49Fa9ssJjULDD8NFd2+7tqswDzuTpAxnlfA7S5DB82JSZX68AK5/o0UZE09DPz2C
J6Z6EAZQJJgZbb9BLsmvhbVtnfV83ZLLlOd/2YMXfb76Y7GPZKXFPUMW9Hu6VmP8
v6Kw9yV+wxArQg4mKjI9oqP7SY/wKoDpUviyDzzK4ZV8psFgA58ALZa1pVOYeUSr
dhs/eKZrcK7JDNKbrOrzBUTj2snczkgYEwDlbIlwG/vfPxOQtDogr2bRXFJJl/5a
ass2UsAy/xDBy95Jb3emTDRx1LKp6vp+0qHsgiuKZuAjL4qOzUbp0QqSf5APPdS1
ctg+E7/pLcJx9Dvdaaz/amnSq9SDEIqBKwoMyBg7IooQG1eYqTsJnOP2xvCXR3k3
5N80A6Of0RGfJ/MM1c/+YO2ji0OilF2Z7yqB4HdtrYTJcR8hXva2uKvxLXIzptQB
fkYhtlrvbnmeOpFXr4qJgck+99i2c3+WPTp2N1MLjf6FNtvna81A/y4oUOpGk7qc
IdOtuObQ6IE9ClzLjdkcWYB9jA1HQd6oy3ZYBpJbZDoUu1JjX2m7w/mFJf1v9QeV
0FVsVRYnKuRVJGnNXlJvw/8LpO2A4e/2JGMP0GgNlGfq5q0pNjLffpWh4NQNuiiZ
m1B0ICZk4gt7jQOYyJ4IWaX5TQ8uqPJK5xyFiBEYSY8qplq2p6xqlKAqhNjFTAkS
mM4Pj343161cbuh3xEq6F/S3xRJNSiqYFvvzFdjeeHXCcihMhgg1tHRI7BVeWQQq
E5AZl6FnWAKUSNYgmb88+8C2q4cn+9OrhIHSr6HGkUKURltzbpJAhHfSJZGWlPKN
o+SAkHQoSvpd96oiEcsHr5DVLh0XppcqLBW0sG8yrN+Z9Mao15Dd4SUYzrSBQhu/
eKrggNOUU2McPMMnyC0CSm1d/FGfbAperWA/w4jwuxoblC5k2r8SZTJpDbvnemoX
3QZnb784Xe0fV9Eyqj5zUH689xuPSvPsnqSvYwUaFrkOqskSC2Q646rXoUu6zUHn
EMLH7HGjLPpBhWB/hqXSODciTRlb8kNW04vy7jYZdcbW5d9P9/9n1MAiLZpeYEfk
3fckhYHDp1YWJYjkTEQcQJozjhTHsnUfzKQ91fQ9D4VNgD09hdtGukfMRrX8iM1J
id7e6vv3F8ksHvC4QfjVWNOKLoeoDavDYf5QIVZ96R7zTcC2qtsme4RRAJIexPUG
wb9+6zmgUGls82LIr6CHYx9feuqmG7RIyRXZ4QM5p/oW2TY5dGhf3V+O7MewoTil
4tVYphyoA0P2d4jQsS+BcDornOQK53kHUEWDCyeL07guMAkSdrrhgXW107PoraPZ
PN2uwXhyRDQSFUkhZu+6yxz0C4ZCH8fViR0aCKND1Bhe29b04WUkLIKWCr8PBW1r
4o6Z/FtcbXxFzYyyKRyuwaoo81Yrx6EzeIm7MDF7rk3/i2OpFdgk8Ke0HArlEZe9
dmk9EyJ+d6E9FX879E3ENF3fNfPMxiYUSuuExPTGmbT2wzi0TUuRRPFBLE4OLCtI
GsQxxMURLJWvNH+mnTcHMCpVvy3gdpskR67HWiRDBqb0S6eA+O+xXH2+Ne/DV1Cs
c6LY/ApVqqeBkKmgkcgyD+JfEBUT19ge5+Zigu/C/2qtExUqu/TcPb7kz6RLSwlv
b/X00uR+KNNRCaoXgvHsOFnpCnTPZYsQd4HbxzJ7EZyuBo7bGDQaPYlOWmG3c1+V
RHTwkpNfIfsQzNZUDJLSZ96AfFsemSBWlyPanxQ2TQZH/3mC3dHVw6uEreaLaJvl
mbgNArX7HrHGnXGDm9pCrlw6aDpX/bQWa4/U3aPYh9Nag7RbrGE+EmZRlzxT3zef
rkQ1GERRIJ9gsUCL5OMn/C8jHtPbEU7dGamMupUhsz4s2HGk6HQj0hC7m6UrB2lj
SiQ4SaqVLcaLfBjWPRUYNt9vZBU+/0ne5M8EGD4ENgrspbcG19ScN1+4H8QdeVFv
2ThzZy8JjjbfheEf4NUDetVS03ICWUvy8Ahl7DL59r62/QQFkAx9m/L4sRfU7CyT
NI83vW9ZsqSwcH/hC6WnNPdSES0AYjxE5o5Kb3zqFBAkfLtCQe7uxx8JoSPqP6Ft
0UbCgdyoVjr7Zyub/9xcDXEQ+5THpQL7KLpxGyOvCtyI3W0aSs1BzHxCPxtiZ2fo
lSzTQRwRfDUqzCAYptIeH10fEHrzrQSYz/+JPe5Vr4GnGLw/LPtrA2iCltT2MR3+
PTLhFwX1uB/iy/g4d6MRwbY9rTEM/Ir4N68MF6MQJ+JDlxWWBQ21DQlBVVDNdpzE
/Lp/CoMEqjKNLBLMwdc1IaXD+NJoiqL6JfCFzFLNPSbzIvSfVbsHyKCBgawuSUzh
OcMoPM3bVjN2pWVXdT0Olj7DJ75l/693ntpYBLBwWTfHKMz2wmu9CMUnnbyKZ9FA
NzHKzwlIexWpTJ2PNta38Rohqfvu25Bfff7SnkIDmoPWbIFDCqYBtN9rqZhOygka
8ls2zlsKsG0h8Dp5O5f3ufOJYskzvf7dXK/s3lF5hJpp56c8uUDLK4xxdgNQTFXx
+Y11Sz3hOAMeCkS5tduFMhHFM+9jYflUb38kurxIteQ2v6o5SMwqYEwumPQgurZx
y1bC6S6LB07B4lumaAxs4qd5ewz8HraCJKHmNjHhZRK2gZGIEij+c9aYaprrNXYk
zUKSrIRRDFOyEIBx0eU/CCmQ/9ImVuJj7xh0eNE0LpV9yBy9eOchm0hlXN6GzDzG
XP61Ogm1hRN/fCvsHmo6jgTzF6GsVZewQWErCPFcaLdodK146wUjfHQ0ie0PdR0y
7kYiwhyo70WHpMa8Px4YHZ2q20tf4qIY0CZTXnKYWIsbbD87quPgkBGMX5Pcv/PK
6SFs38yCyYfH5XaIZJQ2kZ6JBT1Ltlz2DkZthq/cIHNWxU+kBIv62i72RXuWPTL4
JjffN0mCVZg9ofVMyIefF45qDs6etFJ0LIhGPTLvEuQB7klmyHWreHUdzNTr+WoJ
8NG0RAirQ4Wmra16XB3wtLIvcATdIV0nrNjHnIjk81M9CK9Nh2/ABuo5eHsTt5UW
Lo4/sHLVRmk5M6O+meVVDg6T+XGgRuc/4bTZnPixoP725q22yGoqtRjRCpzugDis
moCOmwFVWf+VUea1A5u7xAwCcw6j07u/4/risbeApliPq2ejdv7Gdpi2ENVnQM5Y
XGdjFRvX4ZZBAYIh8M04xTDs8NY7mxnHow1EUvZ2R8QKKopfvGytTW1maGMrz9st
HYtV6RatN8jr5c6JZgFNA1ig4GWUCJunAlvUY/FtKzAmV/9jUcl0mpSqFQvi6JRr
/FujhNSph12GO3eqCG/svo1rojLY/llVyWR8jxPwN1EYJugYdccxUKkTXEJLqfjh
f1BOCSWcO3NmFLHX1c41jrtqrRV+hKYbXLxGVEJqXiaGwpJm6Xnfe7d1l44eRFWu
JPwDA8ib9LEDXdoI7b/oT2F8qwYBPMTFiZJvBqkkVuFtNip/wi3NKtmxg478FY3Y
I6v9qzwLr/3PD5CfD4Op5S0p3A2HWV8XmJsYzU4KYnxCNObbyMayKmL1a1o0AUcY
8hLw9rcgLXDsz3rc4+bDipxJDooSDryUIOB0ZmuYH9ri1VTa77ttngVitnxWomb/
FqIgYwrVCoWIdXphP4Y/Kg5RQKYP0/HsQsCxddgEgBzht9FT17R99cQkGO521ZID
4Swwr8A6pjQG5sKCgAP96qd0+SZSn+/6D//2r07RlVyLfz1jLPhKJ+kHjZEdMjiI
NBaASznDHliVh9EiNc/rRAdkT3a7zmvsp3eqQBgNRPbL9pWE6mifTqszx+7tHQF/
yBjGWDMmFRDFDBgXBsYV4ZOoMapE5uaCTcPA8p3w/q4nTQz0rJ0grKupsbucUUdD
JNKMlroJWAnPG2uoNNmWmVYtuIxLDApbsOEsTUoxR3+QbKAaokDNvobeKLPsCqHf
ehnz41ntR9LtK4bpNlpmDPdau0ISir1BObXjFSdat0DszHCO2GW3Lg19RB1vBTEd
3s3QAqA4Jj+vNPweUvKnPgCJ6nt6DrdrL3HJqWBx/izsy9NEPizm3FZOa6bTC5NE
ttvtX3I2FxwrtArph+jLwHrMi2G9Q/9Yp+djphq87q3zerLMDh/r7muRwxyHtseP
qBUJuOgj1Em9ZeJz5OUJzp0iVVeGpj/rW05pxGK/ANDQFqfF38tUKwSEwWoFIsGs
xt9Gry2/qT+h2MUMLTNqGd/2WN2ag94agxYh/GKVs97mn0MG6kK1PlS3rnVUljeO
4X3jJjGGW1WMZHvzoUqUwPuuu9JhlyuF2oSyyZaNPG7GuVgL70AyDtGEP1XKx3TG
YuLGGpfk9kEdbUGPmKd2sm0+Hp0jLCIq8GSVo/eMW0x9r/CkhWJOODvLrFeb2Gkf
BJoAI5hoYRwQxKG5wvTVkapsHzPQgUuVFC0PRjDKcZ4vYrIrm147sH/Q3kHXQJT4
2F3wTrHPORWcbtWe2a/tXQNwe9Lz5WeFwMGH7rxvv4+fwkKA08+0kqQWNZO1Tl9E
abUhiJMY/HP6sH0nVSKAf55O/6t8Z9FUK+hybrg5ph/bNYpbSBmuoNF445pwgckg
Vs1yjzEHqZZY5UEhTPcPGJeH1uxabZnn4vgdupoycR7L+dtk6ObEl7CEJw4CyjwD
Ec7aPas3kAZDaQDZhMsp2W7Cpcyflds3W/sIQtDIlfEjhkOtL4QZUIgdmIi9URJt
wSJGqeQrN2wNsqmDWRQ+AaM38RYU8qY0oNdLiSO+AHRMeisFoTcZkTG4Lb1mGIkv
iWFlrap6lTcsw5yKnsoIbAMhyZgYUKS1VC6yRocbhYPGTYEvsHouj4yUqNGWeroC
nz57CaPCNf9wFp8PSiU6RSdQR0JlGm1oE3ekorgF9Jr4lCfgkUN2a4+CAPkOeWoo
pRs79HLdoibKDiVlkU3y0/5U8Kquxkj/lWqXX2Kysy7EzCiyE145HIeOdrCzlmrP
wI8d29G5ZmBOfqav9XXAGuZmzih3lQFHsXvWbLYvOzodHimEE2Pe7hFcoRD/eqUc
C2F782OQOFBj8RJD/dX8ebnA7HKa7mzkd7mBSZfeL0VZSNMzD6ec4Gk0iBJqj+e2
MmToW6Aw9scukNQSfD6vZg64joa8dtmCBQS4gbc5pb4qtUAOcyYatRfQ0jENVZIx
bex87IRbI4if6nbxxLp+nBGMe3gabRramRfhVc1M2oWT7X78J35aEGrCUPiqaX9r
swFdQ8mbdozEgbYlQ+v2qpoJnOe/nOGQDAYz5U9wzCv+lbJl/+8DyOc7VnE0qqlm
vs2G/tbVgAhrNkcRDXhl0IaTTEG7AEgrSHHaeOCm2+l6rUdz4gvZ+U4mKiCpGT2i
OxoeWj1lzlJcb4dotH8WkKAtcInBwgLLaYDDopDoKMoawktuGWqEsoGzM3pbpHyp
pMUj4nPsX0EcK3Gr+a1EPc+91CTw9lr4CCacJQf+wMSXyfAgawLHCWWbe9tOmwfD
Z5Ju/susaLvwu7v7n2wBoX+80FAulASxYjHRw3GG31w3AdeBwtBmrN2rOGBklKUP
CCYuEUxxQzBM5tPMz7UoCuoMlOmTUFeHpznMfK3B03tPxcwnMYUfriyrkdsf9paX
ey9WRoQxhb3ATbyf+LDSUZ6l9Ctafam1xLZAZdeoBBR0WK1hX5PWBWisztL7XqEX
w/U2C5Mi0k+V2vj+fT7IZe7vbwSjqxmD3/EJjOZV52VGbyP7I6CIJRoxjIQ8EghB
gbis/2kQHxq3dTvIl6BL30EMmwyAxV+XfQg01BtCfTHJe+QCKBhil81MKBswVZvB
GlJjnuD71/k1urCiBg3qSCAHzlPQOxf2R5hfGd0ev+Nuw8VNVtMFtEThppVXX+Ld
EGV1l0KLIGqjXq6Dv3Z+FGat+DMCneYlV41pdlXFUwTk1HdRd0qolRvgGHNg9E3a
NSd9tvb6ylkBadOnGrCfFAGFIUYo2faGmX7O50fQBVE7IPGZOK75lWXa4XhhCaW/
93Nmg3GlYqdD+YUNUPXDosAPMu8NaFjXDV6jKBsKpWTGx/8D0hNqlTRPCdm8b3gV
uXCoTTRpJCMTv9iOVVylNR7GSMi9YW87luo6ImnxjA1vrtqDY52iTG+ICPpMJ1sj
XOdj4/3RGRVdXhmK+GySRZhKpkRxd9A/5TPRx0Ga6ua601pyWRLd9h/42fiHk88j
OyqZgPkHzFfGTcnuPtQIbANwTrr/uWbZfiWSCLzoUnUw8YXRA61t7XzrF7PjVAqX
7nT4y8nu0LcFP2nq9uy0kU4BPlbPOjCeBLsdQyPTZL1CQoXDKkxMkRfVBXVtR0G9
LaBWjUIOr3QCIihpTJczgvEoaEhUz30NCu6vWOzXPu2K+9uxrMD6QTVOX6p7ll0q
wIfzlMtttF4Pp6ZG8IuhPvMH+f8ZA+qcnt5KnwSTFhWQ7IDwKfiZZNL2x/1oI8IT
V0aPRNOKBLBWr0RNp1O7PEqNr33Jf1GmFUEMFssvd2sBJLoly/Ad7lvDlg86wDvc
GTeJcTiNWw+f6pzTxyXJNzEoFNcKIAWdWTBBRf4d8fZ9BHIAzWWHCNjzHwJJs/Nr
2Fs2Hn9LWQRuYmaqdkbueHHAWVGpq/ls+GqlV6pQatX+7xEWdbCvutyL/GFnVes2
ZZQBxWomZlw8DEvXBsfWotTBylrzwd3u5p2g/znGumlLC3ZHztN+nZ1V6+gpKJdE
UJjoosf0Lj2oLoXsNnaKZS7C5oaFSBgloDa8vozfocUR/jdDn0ttqhJCV1b1Xv8r
O5z/lJJ3gxFnMyU9MhSDjE6+J1Pqk2BXD+WqGFRmjqGoHfIqOY71NGMeQ7rr1dJx
yP7oSEgnkXppr1+hERv4c23dSxoRgIYEZUFfrFvfoVGwx2f7s+f4/QSH+yJD7rAk
3wtrcKaIYtxQGDVGPjbGn5QMG5wdxM/zRxyexNNFBtI7opG77/w/UG/BAeHo4CCS
FDt0DMsLQZ82yyzOqOH9beQ4am3ZcWoKhcY2e5YfFuOlMsWvIDcJxPGJ81xDNRa3
K8GFa9I9h7yh5/wvt8reiTwU4gcR4lJ2TWbj5n6gtS6FOZ9DRtXIie39OUMAko5P
einNMEtfGJNX9/40noYe0woWT+uwRtTjF99rrPKlvgigzdPNB/9PyE54hgAy1+cd
nnndNL84McDqi8x3riH3Zb7c0o+4nIZWb30Fr7y5WWPCkklHwCZhZ4uKM6oVzncV
EC0a2wFBmDkuT9RGK5mN3mkRyDB5VbdFNFpx3TcOst8qe81Mfv+ygjuQgIiXZ4xT
ktqlu3kVLpEWfkcBLP5v+pd5Y9rtxgKPyNNhEcFcS/yG4DylSsQA4NxuHuMMtEyX
jw67I9moOor9GPQMz3cXT4MM5gq5y/Gsgtn+Kkch7uZNUmhh342KOti9+9hNwt2A
HVRfrRYvXar5LNeHzHA6dGtw5fRjbLhcrVUsHsU6DSzB36i29Lb/7qvUEqkcAQ+X
bcpg43nNLE9QHqzXSchbSyGDi/uLkQH2AJVa5MhD/nWcwlnzUv7N4y0PKMxcOwPv
PeD5UdkOIw0uDQhCw0XPraL2cF/tCTr1OixHaPq8GyyPwCYnh4oipHGPNFWDo2M5
22q4O2qo06EZHsc2km9Nzi+YW5fWwB9r4TcOHAfzN/pzEALchjspSIav8cBsSChL
idEHw9c68LPlE6FDnZwgCt4AhSCSrfOOWt+hysfcxDdBLL/a/ATLo7sRAYKkwoyI
OruuqG03Ga8EvxyDNiRw3yAfncuBRKTkjt4NcWeqhhxwPPE7u1HKlFUq1se3N+gv
3GtRsMFrTXA7jwE9mFQBjr3bhWpN2P+j5b4++7rSbgHoA4myJm6b1G9ryAIEH0w6
WD4GdXi+5KkRrdu+CcdeCsZCWKL3EO4W0OmpmR8ammzUhgiOzqqLgoDzkt1N10Lp
Bm9uJ7khjRaxCZ+P/hgPxasO5ugGTdiUIurguKJyytKwjLZIvpLRRgDGE6IXplSP
JHc4SkBemkByM97JGLDI7pO2Do/8N4AmyPFvEkasYkpjX4STWPieGuQJLO4NgQ+f
vXN6Ijihl93sJ/d2cUmaxcji/YLxpsPVd9CwtlqxvjimGJ6Kj9uvG5QNx94GLRsx
1gf4Pgjro9OsGFE5RDP90DFPmG5Oa+paxwcNzyln7RDY5UYdpUspQ1N3kkHjZ8Hi
+d+0Jwv4keqU8vj+VpDOQ3PNRUdHGper+ch9GXh0n44FvU825SzwmS7XCKAHyadP
bDqb2T0WyoCbMgs/FLwhLjyfH8qRwfV1VmlZ04nPCkPqCONKSMJ1gNWsDzQw0y9f
rApB6MIHxAtv2OUVxqRyAFwtFRrBXAjKkl5JPV0BoVeYr28xfYZ4Def9nRwxn/VZ
v/Et47DJqotyDOLUQQ3W0CW6cN3170s6HA9dldWltBTvRlJpujLOAW0u+vARPI1W
KfcVnYWFPnDG5k19/QxCam5Z4Zle0GX//pYh5A7X+xtnc9m7nQCe4lWUJ7xz4HM9
LeH6vDDOXluloN19ccnFssYOOQib9HQjrPwv8zpshVfczubaoe4CAtNajnyGF6iK
zZmy8BhT4KIKFy8SWSO2wqY+K6B4AR1Tem4ebhvVwhjgdmDu9pPP31wIHOOm3n94
Qi7ugEnNJqqnMEHFz9jL+D6gQlEaDPmrTeiCkzLxF/YYqPLxOUu7810DjiO+pzAQ
4nK5yho1Jf5K+/p1IxWspa5MgzzNtLfRr5XdPDuCFm6PAzvwzIsBR2tHTPZyUX0h
voeCDn+R2PYrcZ8L+R0Wa9OKUbN8aDbzwMT+Vqr6chJabYYh06ORjTk9dRnd0NEx
i3VhReyL4BILe7x5P49O1Q5dRX+A+MKevN2FZij4CXQBJsIGtonqBy+9IPiNfRdF
uVUBiQcC8IDTo+dio7I+JDp+FM8GhPHWPviPd9CGvQKsOX/3S0kWzPh2AphSULzF
gKvO7mZZxNcZ2nRhO+GzH0T5H2l9jX6suXvKDkA/lRp/fTAehDqRGqxcDgMRlUHg
U2nmz+mS2Oh/mVCDIRuqNM28/aDmS3f6yDZ+g0NPbx7nj/aKSIv9J5lTzxbnwPVY
BbEiejMUaNGLdGc3tsEEplWhLpyXmkgye+OQaLa3TE+y54IoZpiJjalFahwEMKv2
IAUzlXAmjchSoEVv2Qf+GPwcEitxHyp/bwuF87S7niMoRkavClJpxtognK6kYOuk
Dr1872X117eW3Guc+q5IbX5pxydDLpPTv1aAVJi1sqqIEYj6GTMCheoKw06VR8t5
1RZgCLaCy6dO00mb7nk2zXWAs/hixNxQkdnelwN5/LVfLEQ5Dw4DEQ0cvFlstS+Z
yZB7T5GkZInWyS33HjKFVa8CsdXs9hGgXTa2hYSu/AQ2kJ7jakdVX+2X2yqDuefn
WjPel2abvz90ND3lw29oCJfhyYnr4ekyIaZzB/QV2a0sNgs86UZ3zP3MdvbVO9/N
uPJLmBMaqUAEp+SBQHqIt2Arb1iErsfxf4/MnG/1ic1HMKjalA64l9e9AGE+l7gq
D2mKZgTeSwH3OuUDfwScXros/54ah2xpoGIHyDs8GmIwfRE5AvDJBsGn5Fm9DPqw
hDALrh6f9wOL5a5p2vSWyipB2d3DOYRTEX3GvqSiPYd3nDhVg7Khn3rMuKdBaBfK
47l4JXbpYAnnLBitXaJ7nv/clKu0ETuoqv4639jBtdHoQPoazYBm3HgxfCbPD++u
lzWCTK/74xkj1wdZ1c+q+TJq7W3p6udw+TcNAQBYpz3zsb9g1ZvYTxt0HJFDTPzq
BjNTDz/f/iUjSiJ8ctDEUFCD8BYB7QDe0HPbc286yO46j8TavaoVrpx7mKNcFAiW
1rShmP05ftVwNEZUkWMYC93xr5xNCHS3oPoPg9QYNot2xX+ICvKejsljSqDA9BHq
Qr266hV0ZEwBEAy+0DiKJzBOoyRIeMXBcr63SL42/e5FHdZyG1z2w0VS0gELXUva
iaSQhz2Y5SP/AEjXT3p+PQXMYWD3AFDKvCKsxDVeNa2sXuXzj+3/kui4a3ZrB95g
xGb+BFx1a5SvKfpFnKzA7QxQmSIf+Ray7TlQfc7zZZh6O5owCqrn4kd/+c4P9v+0
lNSS08XtmV9n1AA/WeYlvxdFWeKhCNjiFw9x97IIMxyAX3XMMIyOGR/z280dg6tm
SSi7TBfBm+obtnhvZD13DYYPbaqPQD+vGkOlM6oiy7yV+tHF/SW59SO5bXj5dEhv
CMK6yBR0beagSamUfLFxzFKhXeaciXuKtu50ojjBqrhP1LhRGKYTtoebururNrEX
RHMBqY5yxwaoI7pgUwD3AGfONZAOaRx76K298xFTHRIRbUxr4q7UOgUp3dLSbT7R
/6ar5KaciNbugb0IpmrR2JqW3YZlM3jqv6Hdo/MfSF2uWUwT5QEtWtMVCnYzw8Pl
G1xM8lTqT/j9Rb01iH4SkwJXvcWnuHsGOhpkXpyh0sKUoS7/zo5lBkFa8Y2PsqM/
x42NSQVuyYt5pgdgHDERp9hiIViumUcwe3YQjRmHhe8F/GKxbyTVKYi/PjSs+Wdv
xJoftNycsabdwhROthi/H7YN6jjBNbaPoMLsf5b66oaGSverv7Ylu3Qt18wJW0s1
sIz1BQC4bgsk+sM1pzxAl1Y5kzebo234hQ//mf4iVUivQQIwcG3j6LksAgzH0rDO
05JzZJqWBBLdMd5Ul0MPN2PrIn1cnCRahENo0YASVayma/RFAhNkKXZi+jW9eV99
NiM5r9MhEFRpV7ja4kZ9k16Jn0RYXgU9l47fZEAvW5g9crN69RVT62pFpSn/GZd6
nCes5XAFqzK8Jiz1A7/Ta8Tn11w0CRCsDUApadO0EMkbicRgrpyj+yE4GJtEK3Rd
JAjYimXQX0YjPAp+hTBl9gFb0tx4MdAyVLeVGWQnMRHpuArYMD1yTfUQ3uwCFiwO
GRx8Z6g3dnprq8KJiQTBpZzJrapTvAmwvoNJjdMZn62LWSWDzeYKWnDby+oYdC16
Avq6IZVRqUPUN92RWd2i5zJ0I/1jdoshZ910kuaOl5j+gm5uzmMFC+es1R25/3kw
m8J5u8m69+1H2zfUmVbqwsMVNOYQOQMTd9UhIK/YpSONZne12tCgd0sm8qGiVKKA
BVlZlg71+uAdunYmbGKjZQtHg86nL88Sf3Vuuxqf6uCeMy4vBYja6P+KqHiGnd6/
7vFJKguiW8W7WHwkIjF4+Z95YGDbTuoVh0LDyCDYrXJSt4X96Z8QPkz8ZNw2G7wr
NXi8bSKnZgpGOjEWUhXFnkKhsKbufpqZhQQu/lBNbE3MqR+nB3hjcfjz7qUNhWvW
UWUAuLfCbJdMAJLbkULiPQ==
--pragma protect end_data_block
--pragma protect digest_block
u2ivtuaGou4F7evmvlulloXVCIA=
--pragma protect end_digest_block
--pragma protect end_protected
