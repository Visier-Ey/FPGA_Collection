-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
--pragma protect begin_protected
--pragma protect encrypt_agent="NCPROTECT"
--pragma protect encrypt_agent_info="Encrypted using API"
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
--pragma protect key_method=RSA
--pragma protect key_block
pTaOmfGkAvXXee2FV7PxmLopJZ6ls4G//GnIHP2idBUBKob76OsTu85Ix2SOvsOL
mpR7LOcpKZdE9z+OewnCQYdzbWPCevEIvHQw5i3Y6djdlgoowN3RVX6+HxR7ttvk
zAnhg3czdNCLQFH2716xz+OuGSx1ycbSXCNWGz9MBRP84gDPBRXaMZxQ98k82hIj
ri7EQhG/1Tr9qwgCFvsguu/iJU/9acRetIJedG1IbQ0W2LcFbGkjKazBYDPPg70q
zCsZRm+dPHWKSMEMeixbRBX3eR7zJK9XCxW3XDOzMZ41d42CqTxDAY3oHjeu0U7b
D7xVszx/ZhgTZOylyBrAUw==
--pragma protect end_key_block
--pragma protect digest_block
RCRNSv4AS4ki3B3PlBV+mGAS9H0=
--pragma protect end_digest_block
--pragma protect data_block
sVTG6GoRnqPysqIdg2VVrQbgFshq5FnDtogZ1ViUAzxPqjqUS7FHMnMLVyWUbecZ
bjpJfeZpmnfuvM/KPKFtU8ygbMB8FS3eM1yK+UK7C1U7v/uFgV1PIPJ1UneAuVzT
ZNjSiyOpWUBtkCF5Sv1BUUDVIPpEknkUykWWXHXCu+T9nv/PHnUGk3iX0vD+rKnz
GIm/BBqZEjm1Y6f/uGrITraa6TyQw77pnigZvSXLnW8HHhhkIBO4KDc06S3KXRHx
00cv71xTYeew7DWPvYBUO1oqFHRnHOmSgI3fCa/3y0/yi99SNJ+OgDdaBwWeAWEO
C+oGunJxrAX6ud7NmO622M/neUwJEVWhv8C6pIfeZBdG9vi2MX+odH9ShjWjB2mY
PQZZhYrGYcbrmHHti9uNOgcdoagMuvdZoA2PDiy4YcaFh0WCcUweoNwAgAMIWCs8
06CPD+z/VFIGPEOEZjcQcfogONcVM4FNvyOUC/gHMMShZPef5ozwTafff+iwfiRX
swKBAbEtqRG8AdICEZ+OlwNgXuGcoGa4nQlnWeETZFiZ1N6nja64PB5hZaazTXqV
DixZgUqRanwRpvCTo20+mvDkVtx4KfNc+DD0o9nRhG9SH0LVrH0hgKCtlc4aJy70
s4DI5tnFlvlmQ7MRrLSDupA56vtkkUqW3MTXULh/kM3+k5ygASCZlBPv9G/o9kbf
vZXkpOcOsZZm4LKEG7mQmkgan/HcELLGYmpRKESq+eyjV5pFkDLcS6Yk5ndJOZc8
Jxe6cJuHkzIjiCeznFJAJk+3KkmJxRollJL/961sfrMziUsq2cTZH2IKtAqBRmLN
dL0YIVA45+P9tsSL2hw2L3z22/RI896JnnZyid220Cv7KR+ozUFP5fwXS84gj/L+
VJrngeMCRbBh4O1YKxsxb+crwv2teSAGT1hPY0gXj6wFbJdR7FcRjzuRAgyRTGwh
6oKQJxLYuYpzOoUJOFgLRWI+Sz4h8MWrDW0JXL1qj8jF31F8AcW/FRCFoEkE8N52
bwA4CR4Rixb5zxJH3D3cRNIEpHprLc96Wx/IrP/dnskeunL65njc59mSfRbtyyKl
NlOuuCKMjIT/HdxDDmhrpCFx5CZsMBCs+rZp4nh0aSgfGKpptn2ntE+1k+B1C4vs
ETamR45Y4q2CEqahhmZUd+lo3tm5kEtNyiW8it0F9skHZq+rfYPklJVxzzXR7lph
Nkthj6K8gqHbFu15f1yc2ZW7fIqM++r9Wgv8SgQif8VV0pJVHu3WUClD55Nb9SQe
l/NlX7hTsNhkmhF2E10c1zj6fAmUurfWy5C85oQ8Pm3kPVssLgYxbiPuX6kHf4Aq
AvhCd2YrNghR7cxntV+5kIgrmch+qhmWU7HlotTCbhwcuL3bMUS7PK37W4GuCA1F
T+2ppKJi9/TJCkGq1jry8M4GSWwU9qUtTaEDCw+TwDSDJfV3M5XNZ3zXDU1Gyt61
OzwQCvo6eTWwUTmTKLN/lX4jUqXZJi0peFBmQdB+VuY21YT0R2WcHYdFPjwH4rE9
TZbYAp63TtbB0ucb3995P8pDinGbS6UVWM0MyAI/tyDKALHI/6k1Fjqhoul+Wj8/
dffRxSkva1LX6AGziUj09l8OtBbgy0i4OUeT4kd82lOih1aPiZYqQL/q7EvA/JrV
tCFYGJFZJeHlxJWzWguq8IGHgZnT7EFKFRGC+1oEgkapqQGMuZy94yg70Ipx2/Ea
2zB+QjOSX0mzPI6P5Uvx7BH/kraB5QwSPjXYM3GF3Zns8kBuj/UaspCMRkTky515
yDRa+qbteimxF84nBZ8oJVsQ9buBmjw3hA3MlL5jEqIwzWbp8UOH4dViAgmMD2Zz
Ie2buvv+MiLTfFw2f0SBBGzOMxI1nhgudJ4mCBwQvkiM3rjQN34CRZ/lc/u6kceI
iK//futPGnhmsHKlSPArHlpa0gfNy3AqiDpMPKQ1zIiCxjyMV+0IJZk0p+78gzqL
TR//wGdZb22BHt0ZqvfU9I4mMgNG3MJ990TwhDW/UXw1keivrrDDQnlvbG6Yei71
H/rNlZ1nQeExDz90Ynu4xC1W0HN6v1lZ9pxBxUtLWS+11OUBKUy0Lw6EkK1o0o80
tmaTB5wUB+6z8ljeykRVCfJSJ8ldk+8Eq61tA3HBSV7PjLX9bCF0+hEaKWvXQNaw
6ttbl9+0s1oWHX1AqUVkmDkhIHrwqAGVK5I7eMkWRO1X5qqO6xRrhFy1XZxrVYk9
Z5qJwIbVih7Eg8q4QFuDeBanwQ6G90nKsJRdyoR6k9sPpcq0kjjvbBtN4fxMv2Rx
/0IkCQgAfzhv3T5RCEWCVwsnA3w1AZuZYx6/c7VX30rFbJI+VmqCPVVJ+tTF3qjO
UJp6BG6zUJRcPFRD2dC7tHwmVrp7h8xbf4/pbXGp6Z49ZKolyrjuNvaSvaGWKfMB
43TIPf5Jv7l1UnWlgrKL+9oS44lE09LrqBF6gN1IB1rP9jAj5RN+WUlJmqeoSBTA
Jn1lEhcWSnVb6ZGrEgHgz1ov37t2HwEF2zxJ80dQ8NakQx/QzCO6UKgVOUKblijM
TMPlME6EAnG31u0frx3+SA7EP0N3aTK4C0D8//okDmmhzZQ2GkRRcIYI0yehufUm
2zhFDFhmSsUhZ/E//5Q5VBA5gGYItv4I/BXB1APCHnEmUJgNhS8JfCiHHDJyPynf
OTCppgGZCnS1r/Vg+lLvW6KUUJGxvIXkodY3nbnKIxPvcA+bT0VGM/m7GheYmXf9
4OuonlEHcMtzp4rThk393UnkdIU15zGhXGgtl0MVs6gEEjBFMkxACMB+JcevoGzx
7v+417eCsQ9E8DEeEDXvdC9lmOT3Hn+EVF0yIhsmI82NYX2wEwyDnpb2ti9kGNmB
GWBhtxYeJowjTay7baZ8xb3WVy3k+xyIapN+q1VAT0ioR4/PNau14triTI/WLdsv
KBZgT7dZTVdzJVdKIkjdofNonzYpEeiRyP2s6dx+h+L+8YpuGTXlcDEAjRX2TUtj
sPeVZUU1D+J+f4uS8SHHwGdkApy+M/KTk9fO0dL0DHZurizRFrJKxs8y6t+SAhaf
QabRwwkRB+HBSm77ZnoUL/V1onqUL1kYcDbMSBMfrt8FuLZPKdjJT0xdi/33VVMK
uwEgydYecMv2kVkNerJgYCZssU0o06MtjLnhAY+pKFs1R3toy2XUmm8FEgiTPo26
BitMNPUTpwuhAZNaHqFOEVf4doPVv5Wz8KIHXTOfVI0LyjgdYqMMOXsUvCif9Km3
nA0e3PiuuPH+SgKw1beHb63sW6XOC+QvfjHhJYHoheLW8mkERTk0rrsXEJXRjw1v
B52CiaRgojdwtg48OGPqO6M4q3IgpvleyO+UWTi6d6gFr89Pdqn4wdvuysgxoaQj
M0riMbHYcjG+54B4XTXjrFJhQxRFEWdNKDpiD81lCbiy0VQuu/Azi7c/1LCUBuE3
hTGI7fPvUyM8vcmiNJOCZQaKzKQDO7DFnAcUpKQRg02YmMF0fBucRN5YVip8jqWm
0BOEmQCR921ARklwklIHoIV6I4a3cPSTkUtqDL4D2x0YfvBfCnQYTebXQUawLuH0
JsPDYjrqsbUIePv5HdXcpXWfTX1IsNo2/cXfSsLOCBDEy/WNpxCOghg0jqOuzyl6
rxkrZavY04lLWyRYIlRg4fBFJe70KizPqO12bUq1TkdcUtshXHele72P1M5MIvo0
4aB6iKKaJbq7ooNeblbRWSGTFYGiJVqInQNko1R4d/OdbAcY/hEbvIq8lBwWsNWr
TIlLqmiGpxB4omWoO+GLpNEE+kdQj4SXe35SccsOK2Bd2+CX9JJQK3hsZBGCEm7I
UtDHoigiV6JawDAsurPwIQ7fISWi4CDRBr42Qnc2GN7s2ypps489QiEn+V+tpJDZ
BxOzO3psx5TYNyM2QxHFDXq2swF6B/xZ4o01ycF+iRM02/kFFX/nRFTXBrToqp/4
7IkseoyRdSpneCLKsXXtPZCQz2kqGNfriub5deRkstzZlzreLxjAdrT6xdvGvnN/
TcePn4NwGMfxyYXqOFbzZpaLgVrrvfHubgK2R0u1MjriBpJCfo+Na59iwGrYlHSP
6KBgzlixq5TFD51tzq5z87F430iGqoHw+WzA4z0zFUb7JBBAjKgivJ6DRh0MQtbG
EoBWYKtWYdSlmYamU156t2awhCN9kvWw8rbwNCZV86MrfrypaDPbEZgAzuxrJyXy
RavaNb9zDa+xcJkoPGrpc2XeZcNVYOp4xCRHfDhWVAgOV0mShoguIW5uBrYjapVL
WCCleWuVexlgBSmXtCDx0Jgc5BbXHNG7w43aPVCxlAILfFwZpqngCuPBrVRCAak3
TZIN3L8qiEvnWdE1fS53hfLdHIOz68k/zIju7xLc82BuzRYDF9Ui7I/fjgW+ckU5
y7/PX/12DSTmEcLwpb562zs3qbszdLJnrz7KA9UdeQ+GYRsokvkzPINKaGgKzZXX
n4mKuLJ6xRjPFoIaah89A++OtsdktlRg/jlzn7XUJaWE8zXc5ms5KN0r+JF2VD6R
jxV7Ukz9qFY3gWdNCcgl/Lf8D1XojJHhcHDlBSHigdXoc9bX37VFSQPlnuGeosuq
QR0mKIcAd6pgwbVHJ0Cwsi77c05DKxOglZecz1F1bq+xg+ay+HaY51ui5pf1R8OP
TjX7dLSns4ExZnGnjUSVAT25CTLUkdumbA3OmaXwOVY2ZJoGsj6wGn0r0rvulTXT
2K8c3ByelBuWZmCDGmCZPYTYJgW6MgtDSCSwqYxO0/ZsZeZoScu8017HxKjZhxQH
juldVhwGBYNsUKvM/wMSNRYQLO61MOFB8PjbHSM4AibFzH2l6kYpxIvk+rxOyQSU
rBDw8AnwMpV8f9jDRD1gLbg65mRtnfOxVFtA8YMewtZsGPwuPJW3R9gTmfVru1bV
GaAhqabUFxfnSniVhVaP0nqhw/xWRn/XuW8rqxLUYr/WIYaqpbrjZSoCL2ahysKt
gnCNOzj5OFjDrCHT7Eh9mxotznzvV/u33F6KQm3AN9tmuOX+L0KbLk9HfcxXNvgg
SYbRD6VyykuE0eHvMUQfTV4eVKnEV5TjFwVXozfQxDopF3yhOdfmld7fqjhiZjea
d+k6mmzmt4Xi5kTQtgJGjTFFbxtvXIzwR7cTGU9VHmbqfvCUNl3LkgC6j4o91toH
x3VVT3cIqjzANgQmnjKc2GNiWD9wraYPr5OYfoNcv25gjsHWxqRORDuW8dCfuMtf
O8Inwem+ukB/WAGIdM+ly6kokZxmleNxjmtlXoWlxWM/BkOtYR91pKBYU5ZPPrBq
/W6mlc3Zzn2NB8gd6tSjFIzWe2S1kNp1MEK69389o7wbj9sUg+RWCbtWZvUijtDu
a+KgLj8Vl1hnOgpZicPlKH0Yi49PEQWjdRYFm31mZ11IVXIXauLhfTEN8UWSWRrq
8WI3Pd7m7n/JcZCNeJWvkIioTAjRQjto80uYMh1mXSbiQMzUouD5iMHwkreRzsSz
b9kz6e1mB6k92c7fVc67Ny7mTWEdqMYrjlTwKubdsGgavAla4AUgjDMrnflnlm+V
QBelJF8qSwLl76b31kiYQWUKlmbl0ya4sB4wbpsyXFC1ugqRQGhAAPGM8I4igJyj
w9RuvDr4jDjrYctgF1nS1c7rcV8mlP2c8YgvhMbwWoESBUiPlVk4t7tHr+GvgsJy
1O3SHy6lg2M2RtIckb2n2kbt/pxOgLrBbA6mp+xIx418iuzfwkG+fH8yCgo7MTSz
p8AR+KJOmcICY3RayEGDA2os8/nhpAfSmKMjpIr0pqXVM6aTPf9it8v50J6HKhTv
/AdvxrXDGfOeJiH3NVqsfRLIcBVFxuA+PjK2DLE/pvNqMdS20nN913RZtk/jOzNQ
AZiFExTXfMaiFzJMGgguW9JOomK9L+7ydFIXonAEP+H/hJC1Rw3IrsrinSxRLAGy
/byRp8QNDBXkuT2cxTT+aGLJX18SFzaIWtB11lPL/YFogIgOCDhaaKyjUmYlY0Yk
yuq6k/qiSiUbemA1xxij2Evr49BEbfKQmh118e2WlDkT+lS2FjjeDLBm8jSf7+0L
6DMe2twSRzuN19L0Q9Y7fmz1imFUbaAeK4DdLu/QHTjj5hVbnh0ArQhyiRZ2JQlX
HaxHAC2u+j3ssNrzFMPC/OEFWF0V7Cr3mCLvU7PbpViLDWrhPo611WFPE1iG1Rtn
Kz0hG3vZKatL8xwIb57OEcWO5jbIFmtT8mv4QZHiUf82ezxloBrNRCfJ3EQX5tPJ
8Z3G/xgfcogzS1GfSdsY7Z79k5d4CKOBx6DYjSv68i5ewSYR8pRWMxK8QV2OxBST
UQ+dhtt46FuL8WNYSp1iXjF8J1q3rQXRgh32c7gV4zk91hcnfAl3MgM2+fn/tNG0
TozhPiv+bQRBBk9zSr8yX3vdPSW0qcclp9E9Qkp5Bp4Ska0t2PeYwM2FE83LQ8p4
rTRizkDPNV+e54j8l325VC3EsB7tVel1ekVkL7g3uFCyLW99o1kjVyVX9UMP7OsH
LdUIMTK34qAaTKu3nf2I/ENyx1KsPv5N4QALSORg1HsJs1LPpz5BkD49itoK1kL3
OnHOMB3kheLk/JvOeEBRn1gcFENg9b/Zf8fjdcfNnn+VHry4dakXsGJzaJ/D+2Jz
P81OtSPhQLKbVT/QRJ4/93Jbn9vvtKU5SWIWIySryKJCCcagVPKSgyZUCp+XPiQP
kBzm1+qLSvIA9ZlZx0giWdZo94nSqpYJQ5ww2nMCp7RwyseSOMYsd1Bwe3YMtpkY
pfW4cu6we1u1QGo/obQgvHBrdSaJUmkKYfJi7GPutb27QIHvfzpx1Rbqjva1QTR+
VbXnTRfLzA7QiAG1UlkSewol4MIlbsaP4bl73zUNEumHGqqD9l1TuNWzVDxMtin/
W4g3SKgv092wlg9rbaHHiliyA7C3w3ZAfIOZbRKBQf6bf4csfsvzmhoj+ka3rG9a
JngpYUwqFkS/wPhDJhSm4oerwBddmU4D2ezqtpgVJLw/rhim+jdv4wOSCgPxTtjg
zFHVRPP10QvHjwwtQ5WNfcoklDJ2xYnZmpAfTr4UylAP/Cz4yo9TdcEcnCNQFFLE
CFjV8/+SL+BJu2cPD4aNqE3n3zEr9bFhF5jR4G5ftyC1bzg50EMZ9DzoyDPqP6la
Q24teMKH/wqH2MKCvHCL6kbV3TgzCf2ZbgnNQJJu9TQDMapEpI53oLymvY3NXJah
SFdBuc5M1Hm0OW2sjQubHY9dIiMpWBIicYvOp1emRfTNAILIW916pwuOeQfZQr1l
vkOQCVzjTZEf77LGHkJVH92SnYgGmkWDO74rVEpb3N0F8sha8fdPvZFGUqLUQ2tu
dNICInluWBVQvYbhq+J9IisC2blMY5E6spU4V14a5bXgqATNNLvGc1FeBC0l7ik7
iFxTU4qC7IInERdg+WYHZhS4vWbdb0RBBPOtVCJ28hVSkCnHJXogEbpRy9Ssr6oe
ch25MvNm+q+ZKPmsybi36GHCI+eeA5H7Uhcm20OtMc4C3qjLKBRED3PGG7rVu6aN
KoWWaOkfU75YMMT6flIqrkPFr72Bc7MbbVbeVFkJBQ6szdHjWO8xT2PzMoW7l4nJ
9YeATsqMuo9hBC2agnh9VS65X9v8OSCM7WCAdzAzNtxl6iBXIv+Yrd3PgX3bxaEA
yXv6oxblyRdGoJLt/Ow+JFYLBUiyKQ/qRlG69PKVSlPUNhZtOTqjeSbmvebxa9Pa
qAL/NMqnU5JXTZWtkSXVvy3Fgwj8ODEDZLhGfMFqV5XGbeSDteoVdJpVizRD/zWy
yzmo0p9vjnFw7FBG1IBzCXg5EyKrh8iyKg+qxNnUcDM+PembCJ9B5kKKLNWx6bVS
hBJrEOWfuwJLM7balYA1mgswgX617hRuIdfC7sNxtHxFPPlVsqVNGEAEVg5/mUeB
w51x0IN5a/VsZdmgA9zbcL5CiRXInbisAI9WTg8fQA3GVIsczwpoLsTubxFVmeB4
caW1AIWXUFl/HmWWfUl5XNLheXcEvxeFXG9unUTzABVLggGDiJel5zZiKOMWdS94
6h0a4VbBNYeqdzUJZNZ15Y9wjUEOUJOL6FUzN3aDFtkuLw4KPxounrfu6k7jyTj6
VDeDA56YvHMgDx82hOZyyPHg4+8nCH8lZ/g+Ex9CO7yUFFCP6nCmElyUiKWatpG6
EUG7FryPjvQqvLLKP/jOqiYdJCukWbGBC68olkEataLZxVXD3a4EOXn3rOIP19iP
zUqOK1/qEYLCwisUp3PzKdnSTJGTyHgouF/iNCYfg7CHqWp1lTWhFIrEfQGKRjV2
gimQc0u5up3O+WxSprq8U0xwKs+xGit1g8uQgJWvLjf7gGIbAinG7+FRcTGxsgbZ
J/suvSjD0m3Oo/ykwEZIXtALMznPQWUPTdkJgLIsJrZNceVXpXmI+BWs/8Yo9Hr8
W2pLmRGH3UtoR72ISMuVPjniMFOhIOiesyWSw17RIKNFy7UhMJ/Xvj03OT95w513
g19a3Rl22OOBsDsbBK1WvrvJW87PjphJI4RYYi8dINActRQLn0zB0Ey7pstipahR
Fw9HjJhkoxmJJIWgnG8xE5DvidOkwxMO5UM2Mt9NJUuPX7P7uLZzJ1iktmWXNto+
WlOvHIHFFtTLY8DpOVfUkijsdh9YawPec1hapB+uhIE2Kl0cR1zxJpTB6I6b32+C
9Eu7XOeB4cyWWmsFIcC3AfQgq5KdNHE5syU976OdQpU6zly2hQOPIPK6B+6A7wsY
C/nhaHxg2FncK3Qv1MipgYyyJ9sulliI/lxDii8L5wY4yW62D+dLKxiqA2mCiQ7k
+vIHAZqrkYpoySbmb3NyyopaJ8w5+tOJ6LYVpNDspzXHGrg4r0aPBM1eUx1zjzrd
Ga7fXCPqywaAtfHq5MlXmCozCHeKkQYHv6Q9bOx+swmE5QrYeCbNecpIq4Z7fTuQ
eefWNcyrcwwa0V6mZc3bPTM/2UQ1CbEGk8efai1jFeQhcsRmEXMcCBKehoUg4PKS
HnG6705M2vqtrc/PgbgBMe768qwrd9FnI0jh9nbWRNdSwueJqa2nFyI47R/2s+aW
Nv4iI6fohbu3dtCsmlYNkWEGay6G0osreqw8yYyfMVYx3r/T28Kyz2i3Km+dipht
rHpDQ2LFnCINojECac+axlVBcndmnhGkkYF7bMFUg7+kOliahJJxP6/klIH9+pmz
D/7jSJ2OaDSm3M9b4WR8k6TNYo5BDdwLUqUvn2oipWfWSF4VA2ly6hMC2wXslDm4
BSY2eWwGw9QBuvOh5GRyz4O2yI65oRv0yeLw9XdUs1oYrExw/zQwX1cGzk+4WKex
3rT4ABLaqi/EHdV7f5zqRGB36jKxSfM3QXCjT0bLzsidQ6UZ9OzOLdnfafi4tHOj
oEVNa6akfW+T+Ehc4H/+EFEIwmK5as/Ov6gyKM7pknMCKgJtZiv184G1IQkKpsqv
wTpnl1y9GqMuJAAzRRMNEjpo5uGA0jdP3ccCE8uQIsJDkKtsdc2mRznxeAjM8QpZ
QAlfBu0YPu4QVNmpTTmZmlOkmiAp01ndGViE7H9cC+uFEoVQlm31IkTpDajSA8Bg
MVdi7SIKXLvs9PaMnyXuWaAj7HSn4+A4/MBKns7UgKF7KF+Xo+lHpxf3z3QwFwiP
c7Q1oUvBQLMg/O4oqN9RTYl6JBG2FOpcSrwZxxliJoEZ2dVVoIFs29x9dY8uRx8V
W8t7N8SZLEUAbNZgKaLLUqvpAsiWY+MMJvEFXnYIpefPMor/GUcz4K0klntuQ6Q0
FRWTRHUk8lwlHL92JLf1Y3fkxpzXAr2Fs9cHiMHCkuUhR2TFzGE9cICfCyN2/p0/
lA5E+cPfdRvAWsFqkhREvYAc5SKVfq6MZ2sMW/Zu1tLhfGgGA45E3ts9X+BGTy9/
20eNIAteScWOLZ5pp+dr6Jw3qYPTFY5mM0Yam2MzObiicK1k61UEitCbBV8dGclq
A1E63DawkVoB7aIwXk/77UnYlmxqCcHCs3mqUCzzdy0A2Lm4L8nn/DdmvhxyGc+4
1YxV/xEuuWoegKEXATY3aPdTZSSdY3lrN05xllvnEvjR2a6ePUKLzM89mn9v0WPs
7v/Qsy2mWWnooZcyQ2ruH2tLGs3yruN7SEEzeQ/39YFw05VqRN5HJsENDJi7VZpt
I3fZNvJPPTP388zadq1DGd+k6Oj2m82nAG62ktDVimwKXG3y5WyHkOSks0DBI6X/
uEsIIe92IoH1FVxB5+NfH0tWWlWlAa7GGaEnReSCAO/hz6Gn5mSsoprIbTN3ZStN
EZS7yQrYKKWCwPxFdWsalW8Iyc86Dtk7Ziwc53ObYWj7OQnpeGH0RZJc+0uTRXLz
ZbC4ktGmqxsQ0FH84EThkg4UoF+oNiDa1vEgoWGVk7cdS/rGrkNrBy+gq4k22fcR
TJDItUycX9F+7bKQqknGKtPAivsbTB7n+A49qkBqx/oBYHLld+5wrZTblxheY1LY
kVr7XaFJ7rOkXcGIASBhp9btm1nnGPVz4f81whX01oQnl7mwJiuyvsIkFFYR6sN8
M6OkYNSYNXKCG3dpyqs0s02WC5L1f0RIELGb3Dq7SfYdMS2TDXGG6USOpjVWy+Ry
vcZdrd1RiUuApz2P/vMs/4q5/ShW4j9Mk7g8ETW4Zml/KZcaTehkJRAx7wMauo33
1j7KS06v3JTwcu02fKDehqJBIoo9i0L+YU7TGYG674iMT1EJvbzGLgV7ZIpnF/vl
2VNqblHoHEUmS3H8pgyspoFXDTrd74O7NPTT75p2GtxOg2R5IYTvv3WezYApi6yu
7phr84uau+U0V1puV2HpRM4Cz3ku3uySOzmfBEe+3IFGU3yO7hH6ivLdvocQpRxF
66scY3fhDN/5eM7BC9YgNdoZuzMu37XIvQtAVv2oVzaf84v5so0uUU3oNGVz3mdS
EKHhCbRx2rlK8t12BWBL/CVpXSlK2Mfhx/NM9qyeIYmrHHFd7x//z610GVhrr1rE
t/OyMLjLYtY4Z8g9tl5l0U3oMIBf8aHgTE9vt/+dvjEw9sQtrt5Fsf5ttBG12lLt
Kh/iDxBEFT+bhGAmimKHXM61v+zqIA0kPntQ0tdW9zqsQhMksxwC5kqYb0LDUeT4
O3veIpMdwu6ypPoQF3AfWhCJ62IPHDUIK2Fw1Hw0dJRATOMc8CkoE4wtL+p4MEyT
o6IJkmh/X8YyMgRhugxxom4QF3Qifuov45llV7u5hlLrU82sp8NMmJQxnmKkyMoM
6K9gwkhHLVZjRs9dDvxKDpYW3sQYw0AAWxRp/1wUlqPFOdqUtzQ46Zp3HVPH1XQ1
jOFMkSxjYdyMssEiQSO48vLakqsIxO58oKXDj4JwH3dkbay/gdJeuFqFhbYXXgnW
3KxpB+xJwpJJPyBT3RKuMByIJxQ0V8H6WxIumNXwOygK/dnbB6LSaW+V0wqEoN1y
RURgifA1FUsowVNIaqOf9rbcswbf303K8acvLEEr4rtsTOIy7U45aDovixnG3qrj
oyPXw6su1VcyF3Xq/NWciTEFBQyliYEE/a522S4ZvnJZa0tGKJBSkix0KWi9vpum
kdB3pBwNuOFCQxqc4D5sA7O05a34ZL6clKFRJChXigaXP3muQWO9DlII2Cr+vfK+
KPwnk3Tza2k0f/bTH6Z6l2ZFNaDDiD1RNhvpUa0Ezyq59iir473gpzjuJXTB2GVP
xIzMXxJazHKQNGPh06IoedrxsUwxhqWMkzsiv5hDbNSW9fkYRIiNwRLWch7vUjEZ
w2lHXNhqOKUh+N7E+JTXdc66rWIdynCk1FIAxTGKrsShCq6JdVF9slEJ+1RI9swo
4kImwGWg9r9DpHOS3kAWnvXHc17TDyBem3nyjmfeSDIs8jisv5gI5DGeEbaN/A2X
eFaU7SCJCgVXnAKMpJm53Bmkkw/VakTNLHXFmmX7o5pX+l/pGmzOrPeEOluzK2mU
1e+tNDX9PWoP3BCqrzryyi2m5OYXv6jK+rzrxFb7Ylur2i6/TfQVh+pQ3a4En8NJ
xYJd7ViO45pxh0ubIT2sUJ3cL4FdsU/xaszHwn+ihskluxLTK8g7NK9pv1G4FRLT
bd72bOcd7JMp02kmhP830WgMW0cRGlIktuLsA73FVli/d7n/f2wmU1sw2iSXE1+i
kBwPlBYVWdRwwBf0xzxJ1A45aXzYo5RzkeFHg22BvpANh2EWt95ys0bBsLeOfl3q
8nTJU+sesxflYoeph5peeEVaBJ2pBnCshRwPnIA1eYlm83wFiJVhjJLWA9Zu7vzt
xpuvsRV/HCw4lDftWk3EAohv6Td8yA4s5jjeT3UjZpmQa5P9J3063AR1DQwPy3TT
XyswUNtjEsaT1e9zl496X94stZdupcwK9vh8JvPVbQQSkTUy0WBWolzRwauiOifh
d6oIqFfyDs6D2UP3mAeHj45BZPdTEspYY4iuh058WOrsxADpQcPRBGR/pdz3Sd9C
gCqfr4HjzmZBAfPwMS0r4z6e3Z6xmR8LmtH1xY8B2RR8kI316LA9sUwkFNV2Q3Ox
NRO1azXUcbh4lae+SL+bEWYS/Tuq/SeLkqvsAwdfW3Z1+Bin7bLiDDXok/veOpS7
wfkQt0Xvu8TTtSZoNnSD+ClR9xjUK9JaA9S5o2kBIdTtEmhtCcyfNdA5XDnHdHuN
ZLwbViGeQUTLOCxZ5MlxAMOyI2FS99YWrirO+hEyEKN+HeuMAjZFHZMXdTugPlWy
h8bhxps+FC8HR0XE8td/3DR8qQLy4h4ZFhfns7VMqQxsYNrtAbDALWvhtmqtY4w8
bwN2q0KA776Has3lhxSNL9S7Hn7yEKWCs/BTgly67yLxGD/8W9Z9BuEb9ySBwpaW
qW3Myqw0vzwpCaAf/lx42FUILHKEXxoyK+0QAyuamiNefEiHZ2nwJdLROXOnnlkc
D4Frhrht7dCqX1aYqHu9mlB63mqeHOY9w5DaqO9gEIUOXtvmD5TwkGB+KGZ2CLs/
gY/4k2JFdarJJmJsgG/3BMJsQF/ZSGj8ECUV9f+yecwAf5LHnxAcGRFkFXcOAU8L
w9BcSQIV9c5EGFFN8erLyg0bKso0565UT1mwNyf6pwS9W9Me/XuseXPFWCVlCthZ
XSY7bYKLZ9pthK+YQ3BN+O1/w15Z/LMKU3QvzTabLMwnLwwt8TBtRG1TfMCvKVZp
bW6YL/KyPHolr0TlOLiPRcTLMi69mNgBs5eUdcO2CrHB/MV3bfddW3hWMRQBxJ71
3b5v92lF2g7A59nNZvt3W/Tyz0RoUGykO0R5sHm6WIq3yLrP0NK0chdZEaKd3lSQ
4auTh0ctKI+XEgLT8mMpqHvgAMci7Zc4W0uJywLef/fjnsMLf12lxHeqskls+4MW
sOXNMYv0u8PvNQ676raw5xA/VQrWGwtKQpgRmzIIUA5YJry7GFSIjdp9JntqJMTr
08SwoD7iIq47Hoca/FKiW2kOTX0GeSqcnmtdUKG2hZ6TGwi7GW06rH4P2zlYLoWi
8h7CsNw0x/SGB3Z9kviSuScaDRh936s91WGB6cZnFeHSFIsBim10AUkAP1bQYTLn
FTnC6Opst6XM9pEm+5Vwwnd48q34AFWSMJOnMYmCDL8AWUGlPh8wMLFpqdiXgeDd
JEfJv+Hpsiq55mFhyi7nYs8iwyVfoWN3EOxGj9Mylp9f7WfuVnkiwpsVjIbmnlOp
z6swZWOEwlUlNlGEUenAj/7tGDsnLy9XMC7dAgXkniwW5ihMyaMkEjMFO4sv2Iz3
/YgfYpOvMwoAPs2knLsbTVCZkaPhbLAf0N6RCvd8TcoSFjWVB7sv9vW4a4xeKrEG
jD0Qd7g0mc+twF996czWs1rTeBbtxKLpmBv9FjPoSle9tR2WIrGb1wR0L24RKRKi
5kIw5pL1ayDu+zYzntQlgWtqQ5dIbTFvdyXUjGxbCu/+os6H8jyUxlUBF8tU91oC
gdjdE3m4GDqx8fk9IuSCsHqRjPS+SInLDj4j17k5beya+mXLjZivoOOfrJxbesCg
C6S3IgVdr8f2mV9YEjiwVQeXVwHRYJMjLbXsUipAUyysQ9bVHvLlqk/y+w64a1a5
BMkOtScqUeTzykZAzaMPks64RSF4v6nTfCgGqcRhNi646NOppJqvR85a+9DVHoiL
mQH4DpA1nWuf64oEOzD4hj1nKXmU5+8S/wFfQ1NdkGsHyDVbbv92shFaPqSohmyU
ZelBQHjkZ6SK1KoXQvmADnRPI2MBcmFCe/xFkoThjUUviR7n5ACQDR44sKOIE4Bg
bscLnTjZ2qF7fWYTiNjKxtyjpiFNc0jiYM1VLGK6/+bU77zCOV6uuqLdCEkoW46G
UcljcHQ8zdd/20lEnmOIEG2GLqKvdNCpyPa2QjBurgLfxfP9rrQsVtLEf7xvOjv3
4fGyDW8eIO87r5y2Sc/VEvEG6s+KicYc0tefjouRH2JuQ1c1JoApRmyfm1vgZ0Ap
cBQYl6KOCNPoTBxG6IZHnbNKahxvFIrMYgffU9WnR90ZSqE43K8lGn3faujv6IEf
rVX/p06ox1+zST1Iuz0dI/TUnJAtEl7bgjMT2QRKGwAXcu2I2JA3FVSKkZPmMKnS
KLdDrvb2Im4zoQmcxb9MW1CIZmcOlxk+Av65BIpQL+o+hBfgvBfF19qWvF794ziw
Ijg8XVhMmWh0vgqCJX7sxk/9kPJ+UrdxkyPLX6i/Uh6BZbQ+Y352cwzGRkixV9zP
iBkslJOsD093HpRoeJcsUhws9tXyRxlFjjvmu2xhM/ye5mhyEbONRhy6NReK8wOM
Cn7Zcd573SUPG4Q1qsfmIl4ANwtRMrXCpafIFYY9U37bSuAkW0Zr2BeIt3CoNgcL
/0m2Xu0xZYEjUxrfWReuQdlzJCIm5INq4Yz/pqOmmpk1HTzd7v3as924RaS73mP8
Xt16XftS0ojI9G7ItS3rFnCaohdEmDFz6H8ad/BK7zR1C5AQfTN/6YDljC1juHZS
iB+1LGJ+V9PENi8h/qWUXUWUXY9nneabefSDwojQl6ZasKKAxA+pvTs/4+nkc4+o
NFldk20CMeAvMbJo/1px36SoqdUgxPeiyxSOhf4UzFdjEQ8F4uR6pwhDKN8tlTck
KTOAee5nvIJ79oNqzdDUwngAE92KWeV0/VeWEl8/ajA8ZqlKpz29wc93T8ZVRSji
N4kknjmDW2gZ4KT+YAhs0XHk5sAOh4s8KKCmMXwGxXxvCPf6pniSLdJcNLneU41q
q4ques0sSBwx4xAjMUaKtblqQbvhS0pW94aTUZTNNJTpWaPpJcLfnTpJyS4IjwGE
/ldVIzg9iE4yhQfXiC3hYGIYM5K2DBPYeBhZuUl62/d47L7S466MhXjWniKeX2nK
MdW/sqEOV5xwt7+uqK0gRNoA+1VbrThBr5PFGepUHJWG9gkpf+gbOZvD5aQnRBhx
9k8gBqU7rEUadwgX0snNSfQd8jzELlbJksh0CUeiEaoo8iqBgSRp4yRRaYE+jXWz
zsc/4JKzIhbqW0DcWyVXGm46v1i2SOz8Ishre+UjffDVT+/h2jWQAF0STcP8+uyf
2Zcgpwq3Qm0HiEPxZjR4aueyndKidDISH3RGspkf7CCDp7z9Y4M2zJt5mu6U/Fm3
26Itpqmt92PLzTFvbNUuZpYbokMnYZjfG4+eWdmyZsz7jsq1Egh2eHqfbMR8OR3G
HtS0GB1sLKArlyFjhbIF571wcybmfFs6Pn9dH9qpMCZ+isv9cHkfvqh1eBN+tpJC
rOR6ReXC8gN8qmY7zn6yJ4GwSb2ukI40Tydaaqbp/12dhtFAyJ7YaW0WXCbuQ1Ty
IMGF5LWLnJJbahJX9nppWwnjNSbxFiTqONv2+MRecW/BLZPlVZKq7a2lyV/g2q13
S6KSJysYO7MeYB8v5QBHW8tbd7A9B6Xg37Ul72nr8IRzT2JaoO4pbWmVxR+dKuzV
T0Zb/4BfYKhTFROT6KheSwe9Shgng/RWXJc02/XWb0sKrjIYLxqT0wXZIBYKrW5m
uRCWMR5iIAd5FrFEeX0dUn50N955GKpuJRFDpnmYR1lKZeo95KfKvg61azMW4Arl
zFK0PfDdFWN0bI5rpdDqicKww6FLPx2YB7JhQCYXKXGZGB9FRQkHKxepAGnGT5tQ
2aXytto4YFuWcLb9ERPAhRxXZDpp7J3Rdf1gokRFea0cNJb82eiSlZ5h5OvUSf1x
L9krEWr6jD7XG0ETVYD73JPB7tamBXJa3FSQZdHYOVUHjX5Dyl4Ap/BbITaCyYQn
7OKQiKWBGGpeCZ8q683JHWXjK9Tkklde+gUjEP3K02ZBFxdUw56TL3+DGQYydPRA
zbKFMqqQ+vYCRp12bSWhuKgjtYZ8szq5hCUs/6UcJX/+N1VIP58erAfnCjVxleDt
ePUHzYTjetU4rTkRQFn4kQMaggwny8WUk+PePLqJnn8GmOEx+rdSS4jpK43VcmPl
EYVAwkFoqFPyneIGSDYCXGuPAR/uywVBaCCnmGrngHhx6oFF16jFvXq6j4Fy5k85
Y2/n51zSZsTvHnl1OimUE4hcbkRqCjxXSrURZmb+TGv060Vk1KsFx+0lIr28ZPqJ
2icbgnEZCj1wjv70+13XfgzkxVj0fiWWWoGHe/Mkc22YXli5sEcfeN2eJHEsHHN4
o4RVf4WayykoZs+w5hAlqpaeM8xMp2ieF5TZlhGiYCl502AfBI0AVcA7CgQ3SEMD
l1ZPlCS7kS6sQHJcLXzHXMqW0ZkkOUfe+e6sOE0E4/K9Ml5IrHCPR/QKXci2XAqK
BoWPfmJbVjRlLTd6m4OcnvPwGarluiNLB9cPjYonfT+yrorEceN8RAL47yVzfsoY
txfVOVqQXP6swi9Jx70nfp2RbIrCU16aBr/3IkI8WYEXukvPwH6kYT5KLp2xhrby
bzwkXZcotw37vnyq/P3DeTWrOZGoCHuaKbrwAc6D5MxuzEMdhuTrDPlVWx2iuZBA
RBvef+BZahZUth/nXba7KdeZm7jZ/gO9MLLQiqUVUG4IW7MRRWp3x+7usiB2IqUJ
BKNjY4pJWZTb14JolTBbiAnatcO/Op7lYJJNAb18hXrGIbA6FhP2I071bSJdtTev
HuzfRO7BwN5pC6LJYnilDDBjB8oSvSCJ1Q5a+E686DKoF+uP1Z/C92i4iyYb1SEF
yfXBYCj4cjrBQovZGAhnIWaAj+reBwrAp6kh4vph2DT1zZ7YNSBkUWg6HLpTQQsC
AcASHE9Ut6UHmVnTeBKtu+CQKYFVpqBeh1f3BTqIs/+Qp5us+u96G98TzdHRNmoZ
rDVw5GdwTDUr4h1gyIcYOkbLkWwxZcRHVOYfIqlvLawl1xpfmSAKfRDEnUQiG3hj
wqvZg8DF9iCNNtGAygEn01CGrJ2oLbefLWA38gieF5uDnUGJgn9UA9HTdzn3IU8T
rdvfqmW6ACRI0K5dvgahfH1wp+k2i/cJZBIjEuGFKJmj8Zx850msr5t519Ud/hHL
sj9oh65CJqdE+bRdFPNuMtR5I2cz/Vnk/Ehc+oYR4IoonEATYcoVewdb3c31HNf9
c2INz7CIhO2BltFvqANrz8ju8FXdalpyTytvmLtycTo+gt/2TfjBNOdlQ/18srZE
PH1LcQLe+rStiOtQS3UBczutkbgSO9+lqDljltsEdN+0qnHNIqXnjCxlJkCaFteO
mj/NuNFb7hR0M7GAz8udsns13k7lc7c/teaBERpB5zxkxWGNpvjNht8pCz2X2pHs
i0xYPTNFb3W0xbnps5gFGVrDkgbveepv2XyLLchH7tl3pqj33mPG9iWJ/dEl+TfO
HZqhq6vrEO2jiCJUZ2N2dcZp0F8GWh+R10+dkE4EDHjgrspFItD2eFJKqFwsrjzd
7f3UEQcD6KSP0QJmldfQlBYayv6Y3CbN+Rd8y8LD4WeQ1ezH+EzZvjvp4/A6CZCc
Ht8a/WSNRBpqkRm6d5sifWy7sKxkQ34BmOKhmVwatAiJsu1BA1WtBhS/ycravMu2
m7aL+qZfLZn2Qut7awyK6/cBHASTEeE4aonaAai5ksrBzqt7j2HhGY50Wjk5ZRnr
18215w9l+XiAPgpO1hcpd10zdXVvNGtu0QzfgDSLxdKide3WGXeuMQHUUl2arPS6
XiCzf0s8/mBLh535iPwza3YOVmZaH096HDdJazXulQuAfXifU1GYYT4+x2Ns5Len
iJIfUFVjO0Dm0w2crGPHTd82ms/cfKpLyk2/MW7gEX/5vH/l2gVegEEdkhYtcIpu
s7mrEu65kO9E0cw410qlyuFcbFUcAcgVEvJnlM53maN5E52326yr/cm/iqJcb2Hq
EMWysVOJStEIOBZ5MhuA69BtDYhMc28A/9609gXO09l7RDFXdHQhdxbL4Wcw8j/C
fLNw9ijC+YKwLuiKhRi32+knvf+kzQbXhKGIvpjk55HgODT6Uqh/VnPHV47Wi/wg
XvAliW7AphqCgE2MgEtB6tg5xxNJ82knfvBsksFZq2h1dY0aIQxNeGy9pvqj/MDg
olMqcJvOpiJfRUoPTVRkezYnSKvJOXtQPl7d+strPYdz6dEVrGCORuPmNACgrigy
YTOrXPO08jc/lhQVgDVtT6y1OdlWDDfZUbTj9JvaI6pD2QUb7M9F+nEkgGpYZXsu
Ak8//gGv+vCm7D094SqeTjtX37JGvWA4xGVuDqupbrQnCseMZRP8zzxlNc//qbVd
dDr4ivcifHvm2PitVpOlPUcNjG/ocRbk/Pwkd7IFwPTlgA2sHxPYQVc9+OhJtU8T
XjYCjFEUBXwAFlutxfqXtA3Yjf7fvsLwh+PAKnOdaUnYe+Yt4Bu/t/k9iki4GkM2
mGSdQ4tkHq0r5/bgyv0BF9F/E9YrxNrnshTImLN8aGwlWwC7BWXAMwVOW9NMompM
vDTcl3+t6nGGYKSoYyKNfAh0FtbEd7mOZ1GDuMXELyxZXEmqPxYWWG3e0Wj+vfQt
xEwS+dF+ZpuObK7nLIVD8cPXGu01rVITSnD2fQa2tWiAYBxsfCaIyXTIJiRUsx+j
/hWjPs40vMJGkAt5bcitEiMNEBylJgogM8M5aeBMjoZ/6uWIC4Mm6Y6OKomIiqUx
fHdoqbJMODANsb4sFfvGzGVjGyVtvJFUyyg0jpdBpxSFdGj9AGkesUp9C6Xo/z7m
rlSt1rk611cBVjKUjINFOXscwyGNLTl0/65WpbBbSNS7i3gotaUfXuv9GKOv12pG
AbM/1IJ+ADCPrMFNtXi96hToybb+gEJl0pLdPhzDAPccttZfr8ogpSrzfiLOs/M+
nLgXbU3feT+07kOr/bQ8QqBm5tQyxWodMP/Nhdn/0UTcNQKxplcHd0LIk8zNJIxZ
IllqwNgX9MOw2wPXWbHIXrCWOOUak6hLs28WNJbpXhA17fzGEMDoMgMerTrXZU2t
iz0s5/opfZQGPW8W2CLyK+wWcUqPoUE0K5UL0ojdhhXczqnSJSW1SbcVAmLEY8rS
yLA3odgGPOlDJInhSvZDYkbEu7yoOKcQ7m8Gplm21v5TQ/B0aOfsl5Bce47rqxDi
VOV6vBfygG1KQ3jXscviSJvAsFp6/iVNjoxisIiN3XSQiVy6LUu8FNt6nHuGpQ+1
IUgyKN6Wh0EnFTyWDZKdzfH3IR5BZ7bzIYRnznOtCySV2Z5guO7ZKqFNN8D3knNA
VVQkSxJ0c3MmFoqr661u8mLNoq0pGsNKOkcpsMFY8pb2STm16my1q9yHZ80125x3
/ACf6fwLb1wiZn/X33t1sJAWNfDryVa2A/y/tw1gvQMSMJ6IVh9ytEusT6U/1lel
NzmOTe0e1Pr5RFE+Xa0JFFzXaQRl/g2lT59ee7rwQ2UpbgpH/1/pAH+/gdmoRcRe
I7cnjomIWH2+3w1Phkcdl+4asWSI1mFOEn9s7GNxDlBPyVuSca2GnNM2sOL+Gw7Z
GiFiE25sq8zd3vcmSMlDXUgTJCx3Bztx/NYRlhC3YG8NYC0lOKWrpIG/CZWJLmjs
cRgS7jkl8zec6Y4b8Cy2zmm38dxaGJQGnZTTUW3B2gV25ahRBYLZy+bzRcvbmeKZ
UcK7sSd4iiB+OBWtmH7jNPVoC6vO2qhWbKeatg7o+Rs5IqLH8AZvZVQw3GGtzPJ4
+NF5JilwLn50TIGbbkFviBXI6iczGfGPhjxdyj5LWbvvZ56HVLnFq8klckgLnJn3
zRjwJ7yOAA9/LWip23AnvZGM0wrBaWjkDutC7hVuuG5XuuwHev4WJOzx8x6LRXLT
cScm3ow8dPiTQ1kjMKmkFLlvNIdGSZKdyelWSY/RbtQl/Fjohw4sFyCyW9DGpyJA
7cPX019F0zkG0kgb7/BGM86aNfpBsxCsH/KL1SysX5Y3oEL29s+upfX6CH61ILvG
7WOChg2I1heyK72UZQhRX/gRYCH+vx+JFfLZEcPdYMnqOnGl3R4d6/yy7lzq2PB+
cWqOlxxDKjb16ZTs9Z8cEReTcCrLseHTYxK9YXmQNpjSGNwXtRcWy7gQj3C3sRA/
TWW8/5fCPbgCBUBSEhQWIUcvgU10VQ/ToT6N6uAKlgo08zsLZ+1UumSBX+k82w6j
FxTc/8N/U0JS//3kmCJRb6B4w1UrEaq380xuchOD4i9qWpYVFu6gXG85NIAejOQx
FePHG9NfXc3UDFVsQ6WCkUGBMV0Uil+3z4+Rvy27xMch/IU8ACZ2IbOi/I85jvEm
TbsjMspdeSHZvKJvZolE7VxhSsCks/8TZb+rZh4vntWpVBqEKiId02MG7E0olWho
Yt0aM+scspckbb4K3F4I2OzI/6pWeuTKM3uqmiPltAQySubRaxnqewIeWcoLGzBU
0LSPSZRoBGzIiLAHeq1PswxJlB8VQSsT8N3+UL49AFGc4GOycODH18P6lQNFt1vY
njehsnQOy9d+cgQkpVZjGoaymnR0nD3PRUtvxa364JGSoILo0wpkXLwWKfRvawXc
f/hApjHVmNtxjFsslbhomT31tVzjEcBAv2V8j3Rjyx6Efqae9ALB5ZMqPRMvVOzY
XL6gO6Fiz3gmwf7h0T9vrLzmzlNH6zXZMiDZ6wA4n+FJtb77BJV+YufaAYhnfQNp
N7DjrTRowiRMqgxuxO9z00rYuFSKFW2EhJuOk0V61y78iDJW+IAt9AfNTu73ncc2
UD3oInkdfObdxpudYUXTXPnEv3NRgSjWNRbL2lU8RYxsCiJSl6RQ1oFnYNAEnTvE
zGnUd0VZ/o8ZZitsC6GOagWy895XrAwTtQW0viUfbUSlH+kg4vsq0JGWEmo95OvX
4+mFSr5Ua2m/F/h1k5Vr6WVvpYuiDSFNshwr5dVf8kidk2F7P6mx3t6MRR0LynFp
/RS8B++C0KqYm/3a13SCHwUW/N7+bBalTXHGZ2RlD0D11Sjkz/JsVYVQzLglbbua
VRX8Qbvlq6zgO9EQLg3kZj1LAY8aiQ9G7uv9GHqgiJfLa8OLTwzUSbkaWs7C/bqk
GL7+58jXB4vDayTQGa1Awd5gFn8kbQR3ZoMcaQQBVeg9fI7eM6VsB/wwSNvJgRKw
R2P0E8y8Dx1yNz2aIxLaVf8e9YqvEcXAyAVNN8MHW9MwkMhi09JFDBQTJSZc7WKN
yF07HZ6ms1wnatgyGLFQr0gzlMHOm86aaMofBY50/aHjO0UZHtTV1pO1b9Z+NP5c
ijv7YMXZXOgt8S+zRTI/529VmLCqnORCNf7p16OtOYxX7kEPnRWIKkaSKo75E3a2
QOgdS7XIOA0Q5LJFxlY36bkF2oBM4iWG7ukHkkfZnFdZ+pFUIYv579clvvG0CIrn
Oun4zM9iUHQCSf07upw2BXXWea/xREQgSjalVnEVyb4PRsQo08qeDMYlE6w2gN0Q
9Gfh8tc9/OHKBIL83JoqnmIZRDcv5/Mpq/2UtK9vwujh4XskM/kkjbvIs37RTrdT
GYlVls0KerylgrgLzVUoTtsF2tIAwbmdsy2JqfrAJWh8cF+uF1inHDQxT22dUiSk
aBm2fV/VxsACiY/0xj1QIjj3bRdwB6cTOj4LqLATcQdRaQMSESeYhhgNKKS16mwE
R6aKSiOeCXoXcvzXnLvMpHW9UbvVj7N6lLr3aGDwKE7qfWA+w8DIyK+sqyJ1pFd7
eZqhJgTFJ5R+odzFaBMGYTKVAHopsxk+XdWllRrS8d877wDCRP7M8eZc540EkkP4
sqdELFFeQ3pHEUQ5ObzEtetwTzfuHRqLlx+xgIMDD3JNYNop22UQhhzHml7otkHw
kZj6hslKD+AvWeBxsygAWCsZCpqCC7hpE9mwfwB4M4ny0kTP0b+B1rDPiMp2qiUj
6ghiG4X5oXU82tFJMyVXEWYTRFFLj2Rq6vE05aNfsyCbKxDBaztfdoAA8Z6SJOs9
+ZJmoSHRriUoLyEgFK1c+5awXdeniMLbfA4vS7WQuUsQj7FTjSqiQnqJ1/c7nIgR
FctU//fvPw0nmT2Gxmpb8YUK0ffLQVpa4Kr+sQqLTy/Os0D/kvdLEp1sBSGSZbXc
NOjmveeT6Q+2igxxCKVzFexPZ6A19+Pa3Wyj6cs2/ra0r1UJksnBj3JADDfZ+HUZ
ujCLTsd0DfeH/eusxg6w/5o9pRkQwKmTBCbG0n+fzK1arYb4BDUoWuziVlsFHs9x
m32N4ufmEC5c+bqpOZ7M4EtewmV3SwHU49oPbIqGvfqDk3Li7hrzO69/55TAmmJn
VbGIbTh2EcyVnKc/928h4jTiklgN+RsRnWoXv+HyL65ZPYBx3GDX0bS6Qxg/hXtk
JjcarZLlMsJKyEIyN9tmG+dI9h/XXXoNl4+7L0tV4GqHsk6N6ScpIZhnGLmp3oTi
HNEfz1s0LpeLMWmejJcTBMaYidbXZyxkIAKwvyteCZBrESVnmyAHDPpsqwYP5H2K
JlridAiB/b/Rm7xofqUgswU7O6gIopsZystOJvtweknJx/40zjM9nGZoYGnPOv25
6idaZb8g8ISCt8XAiDZHkfU0enhXztFh/EDD3vkRASVw/Ynrt+dCsTFSPK+FiK1L
pXeaLsv2vKr2QEbh2/GRn4n+nIevlwPvm/F72Sy6mdIKGmjCL56oZXYsIrH/BqeP
WMF9tNNjeypPQi2b3v5JicWq35dRdKu/6siL6YFvlXJqL/mfiMBqhtqZRQQDBwbr
Rp59FS3o1JMuq+f8qnug0nervwCSbajnL7HNeqUHnEMSUnO0ZLVa9Mw/Ccg+tE0U
5TPpsubrrlBGn4J/yZI5yiSEctxWSTGjXtFqRBodUQpjnq6S1MG7LzZhYuT4KT1r
nQwsaFD10VgOpAOO/1T5RRFhRcx3AvheNPXLVBcW1xpMeHu52qoJhZbDQ57p9yzm
Lh3DAk3IP4oU8KqLa1/iLiyhD7z8XFkN49tYDTwSL/FafdYlEcauzG4K7Dydolh/
Mcbo8zOZWlRiJsVeuzNWVZ3p4YTPAIAeeE0IuwGrJI+Rgxq3Bzs8B7Z1TYgnP7Zk
wf95hzFde15kT6E8u+o1dd3ay2m9R1INvIUN6ONTIQbqPWX1y0JRlBKNzLSTu/Oe
2NQinwlz+fJXwFr/WaRJkymuqwqsromCND/kEBi8hsPcrDZfmHvid/Nfgv3DydsW
jNrL6RVbq28PKR51z8uCY41lQRIVsWykRIlSO0cRUs43hZ/tbKUayt0o41IhBTdG
aHtjQtIsYZY/jtHKUqllV4tsUhfOF/Aa3rH5n5P0Vtnm4H/XVWXSTMi+bOe9MWCz
4ta/S1CbFQu0oEn9YVblmUFtx8WSH34+WfmKLSGSSmvyt38rlT8SjX5hjHqWEV4U
facKfGyoHsDFnhpZ8NyYv6Ms4NJhGjbDJudymgsR41qDPTtlxzcvpOjMsAum23i5
x7+YeRDI15LZzIPm8xgoh+1FnJtYgISKBWdiq3lXQywfbC+ZKRqXF9LBng9U6j9c
RNDpnK9trDvTyepV1se3HbKxA3fc3ONjgTGT15Tiehtq5F0yx5+NAWfoc5oEvsu/
DbkbJHSi1yIdPAptuRznvuLEr4tLTyaOJD3tGvUYeDVodCyDPZ92fmOqJU4bJle9
0r6I/iUZedgeuVAx2ypl6bAL+ceiAKwmB35eNa0w0LWSeWalcCkMk/Tei+kb1VWn
vcvOHqSMChUBDafAUuxXWm9zSFPUWysf3M67gWLgtubHOOnrYfw6xQfGG1j9n/1R
p3zCLkLu8geHyf9M0rkZKXsWx7dutq7aTFGE7eAezcQLQC0NvSFaepm33+1sm1oJ
umWEJea+sfN9CidCEFRNVCQicHoCkE96TFlhsTdSheoGDIjP4hrwcbVkVWGC5kML
L243WuikpIwTN1BG2sd0R24hflNCFFjBLxpzDM4yVAfqgiwOZ4sX71EdotXYaIw4
cSo/V8uYnHlh/1qP/M9EVrMZ+4vJiEwx6hlcmpF5Qz6k2TrcIPzaMAzIJRmldZvr
wJW85jXzfTcIWsoIGLfUvcemTGKi5obaaoYv/toN7HOjuBFc5MyCLGEJjspHXVQc
Q6flT1De6dc5IWXM7OkOiCiOwhMXtS7JfuVXT3KqrRnXaJkVfjhYenYnmr48IJL2
C54XupIOixRWP7AyZdrsPO2I/7g9aigMiq3O+tIAf6aUzJRR86MdMKbZXmdW6lI7
0fERuCAEI7SzIvj5YB5Rj/t1JK8D31JuRNIuObaNJm2KNUkJSkaul9OuHEVrNJv9
e2p37/KpE4PSJFuC7JCmNN3j4UTZ03D9zUwmq0J19RtjCmJDygsVWWxdZDOljl9Q
MpOHz1HRAY7ohz+3o9xATKnyfizrO7/PSV69OXMh6JUa8ii0A+fVzKY++bT3j8Gl
FiQ0XtX1DYTJDJzDVhzW3D6nO783ZAEEN7CDGxBTxon5mOBJt1Ns/y4N+0RFxANS
lWOE3hpFQDq9LQ+n2Bb3Q1EOavvbJ2uT3grukD+YiBuPgevwA7E5tZvyb58NRHQp
VJbpjcmg+kSKst11bBwRARxH7bMOK8kk8cpyoJpeyr9B3wZ8dvVntkCRQj+4tkOK
LdBcfsLGwz61K0thkWR/aIwfMgzJlLjviUdKxmTu3a5aLXzSwY3WReEaMEAWOMLA
ZhVRR6hU4QEw29NBQdSrQKdi7FGBIn2ydynFSq+JAcK/3hYX3Mzm+HgMIA4T6CId
6Wqp1eCRiUjiXzy0XQVDg4QzmzdIIL5AHphwCQA3GcmwRsHEoEAjOWXSVefXLB7j
/uzztKA4tQ5gb7EaWhHWPodA5LZ6Gk//1h2rvXxTBXC1uXaC5CVJ98FBs576lVXu
zyt7vaOTDlWNSpTF9SpJ/8ct3EUbfrEZgAQOu42zwni0QEUe8IGIot88kd7/4ec6
oPsLU58G/noSYo5GCrqNwhy0d/66LYAHfWCNxrQo0rN5mZAUB8MNuKF+Hlr22O+q
duqBx080ntR2aYCtZ0eVdHwmnib698Wr6WqDKImjspA2glSoX8nXhA84DKkYwTl8
Q8aQQZ1Rp0UrBz0d3ScKgTL/ybltXLEIrsxo3DytBhzWDLmBKlMdfg4Q0J2EZLFT
za8wH8B+4mOyRy/FXfgnN7pYD8EivgPx9vYhNOWFpVNegg644coJVlXqMrBio3hL
Yo3R1qGvDaZ8YWC/dGBLDyxhQwaNGr8YmL1ZeNY6h0bvKfxi3xjPFpuWozujou62
IHnXjEuDFmEQXo2WOohXqcbJIhXErYQxf6Zn1dokGFLw7kewx+qCpFyv8rwASwys
eDITf4nyT2qn0WdZWu9yyJdEPqYMeLzaLbbot7lDmKGBOcGeC1MMEw/JmrbKsIHs
RsSSf01OiUE2AI1x7hv/sU8EBbDwvLEpX8VuQehH1NGEs6AfrpSvc4lQ1NwJ1T0i
8xeuWHk5xP0aCyxbbdX9qpH6orazCanHkWNKh8rfcLvZ2pidBpPaE9MCg9FeyRpr
FC4sAZiMU7QwqQG0oiY5DhUMgue6z6h59RS3qDZlEzm4Gr7TQIaAKD0QiZqRFyL0
okIKwPkbm97QcJW+WizsgOu4as2Q3MPcc0hmm1fEMSHzPSk1rUxcoo1mDUwSK7Bb
eYE4H2ouUX/Jfk5y0ihZsKSgC82nNXVnSIRopnB0aBJIJytOqG3SzJu60hY8+20j
672RMBvbcGNt0hO3B5+VLu+yzqHz0ucBI11KAlLMXIwIhAMT4jpLr+cXRaPYPfpQ
rfWbTiPOI84Co/R3QojopzMT2oZGmrzh9SDd2i84qab42NlDa41PqDtddiizQq8I
Py4SM8RgEnVaVxWL3F6RUswqWTCeiq3cBdrJNBFt6U07ZUuct7TGklxbmCODzILn
206tWPQctCJ9ire/7L0lRlK7KGh8aLlWK1hPPgI+GHuMyWy8r4/5vUC88cbg3KTE
RZqvkV2HFGVJ64S0ecj39ubF5zcrTWCosaEF1b9guCXbffwwWo2YjMQuJZQNjgBi
1/bwjVTMod/WBhkHdyM8xILKYKR0wCl6foRQu0XRlpqAZxNeSsRIIqpXUePElzvz
X8lrHMi+j8tvI/ESOJm0gjJfVpvje9ustiliD7Adb8X431FFFpOof76c34yXf3Nh
WZi7Wc6U/FBkkTexm6SWsVzMWOft/yVfeZuZu0GZUPLYaiIcPe+GF38oVQfdODBi
Cds2dx/zVCeX6TH7RrYAnBZ2N0NM+c8RFMGcHdZ/1fwYyAl192QEvFhmGQNmhwtM
hTq6fU2Dfvv3562arwLByql3D+nuu8fAnyQ+5adDt7Zuxkg3Vzdk1Kw17bOjn14U
mqGDg0Met5gcvtlCVH/YfTJWFmpfAk4sfKAqWj/MBR1vm0VinALJhj3Q3kf4i/OI
dr5/5Y1K+ZFf0SisGHviTu5aqul05PEMECucplAqvP4Sq4lDwfo3tNW469cERQcj
ETzRi6eQfS0qWfv/vWq1fBIjyak2SYsCbL9U7dz6OEtC2Qc7u/0b2H9qqpXXQqLP
5v9Z8dDEBwLvJgVO19JodWQmSJOtq5j8B8zpT9blqQxyBvKRE0vpTiLZFNFtgxha
gDRmGts5B2zz/Uw+q3PaD73sdXQyrJxx8gpUXKj4hecwfx6ZmPO2KvTSfWT+E62P
3T/3oJNBRCNgr51VJ5XKrHXZWE6mZ8snEiGsWIWYfghQLLol2Mqo//4Qf81iZJGh
/C3wLrVTx48RkDTA06u+NhvP9Px62fy63c9MqBg7zyLZ79VWWtCnVSToPOmTBwGX
SOQD1GW2bfOXh8NajblYi7p4CzEBvJDgaJE8wOefEnjK+9MxXiOuhdUNLtdsNPqg
wmVUeg/ey8cX0LPx+cQuNFoCVXO/CvBpxDtmI2nqnk3eaoLXzzk9eWPcRhp4SlMi
eoIXZBJkZq0DJNCgkxm1QeZyOx7j6BT9wtnklv+7PUBpUgEzvqNFz4dGlKjqnEsb
cOck2iwo38nPMne32JTLk5Q4uVqolL7vuuXuHBRbdxqqAilUUe0fR+tKncQoEfTY
in5hfNx52iukQK/hkef3n07V8hPleMejQ07oee1PfK2zIELAO+9X6MYdlFwllcIw
NH6MqYmD/WuNnuAopYoUUF3nnKls40grlV6mwxxpF5qcXw1hXvDYOzjZ2ImlxvDB
ZA2CD02Khs1ZysSxuZPqL+Jx7OUgsoSwkq2LdA15V5nae4pXc6yLrfxhwy2qCjqn
b3EIFsFVnnCP5LhXqOxh8yQq/9vh8i6EFtB865L8H5vXRY7p5wc1YUw0ajuTDZWW
aULCAJgIoFOA0xdYBuWNn2A1SwiuZE3GbY1a2XpTHWgLdI+077wDdy3juwuGFex7
mLbK6blGgJ9XGc2zgq9SC9h3/aZclhlG0Hbwetu551IgC8i459ua6CjR08u1jchV
krpGDH6C8DPaDSVMEmvbNV07m3M0Cq64E276HEJZDgy0Blu9IrRbrAOfHNTFfKvD
TCmliFYclNeBsHH7/5+W41v/2b6MzveL1I+oCXJFX0MR+EDPfi17EwDeYr0gnIXp
yowkZE1GWjwJ6F7r16RgRsc3lm7ZXOvnTPv/LsSGc9CXVaMBzQfTxMyc4KUPRQIX
VF7045A0YDmmcY7QAry2dHhE0EVaClbjkaPU7LM0lSt8w7bUIS2BIoKCLmCkCMr0
ifKsOtTN567x1P/8EFB2TPVpFGlUyXiM4gPof8TfNIO1o1UY2K+s6LL+tDylMlZK
zbls6i8/W7x0Ysd8YPvwkH2OOGw28BA24rbJJYmZ7a0mIrJ85TuDmM3/3HT1+qBh
D4TqvT2scvMbC56Z2AL2X9o0wP/6jn3oO0sMcjokG7vhbwLFsnU1/DCTzO5yfgK5
tGu7oelTmjJZ4Qbbd2IYKT4BWctCyoiu0enYl5mUCQYZamSzmL95FBJvOJ41eqPL
zJ3fb13p9K3JLdYbc591ytfTpvj9C7zSSejBU+kzGuIfGeDkzrFqKKAfswUrBteJ
8dToqH2cnLelbUHCMjLlqRLBoJdJQ0WNt7LBB6tjJpdYN5oPMODfaR2VhMoCIsOQ
RjH1puZ/5VCaLD16L9kea1398KhYetmc46kA42OEPtH/iOkjKnBQ5sgYi52/Vs3Z
FtQnAPfj08zWEWj4oH9GzPiqoF7txUy55X+TwijlTIC0A+ge669mGTGk0YbIOZ8W
qeKxBrwiLRN87eR4BJSpQg1Rb9X5OMng9Lh+H6wT9WWuhCowbsZxUWhS92dN/+A3
QMghlCZTdITFmY/PfU6VaxTA6q5dPCQi3bGDUZKAjjeqXSGFy1z638DPZDjjDB08
oypR5tCcz4PMuCKxHWRQva+uz1vGgWaxSs+hH7Ast/f2+hv+UQCAAM+Ezhzbvnj6
ynl+MG6NqX1we3O7w8p+5H1Gw2EZVBZysp1VFnnCZxxPJ77lHUZGeNwvmWovonhx
iMJ0VMuu2nXOJU+1v9iZ2BigA1JXMaMWh49FWXGXj2zURJewie33nciLDCUc3GhG
k5H62HyZDQ6gL2wi7ZavtbrcA3PQzZHgLOBhJg7fRAivjCpfsLv6KWLRZfdc/qCi
NKWgIDwbtQX4KkcCUgJaOmB+G9s1gLuKXmRHWHth0zIrl4LLy8bTDoVEnqlrwoPu
PXy4ul6VqI27QLiQOxfU3ZkEhmrudBbNBF5Pwlp8xBLBN9+yh+i/hfeGqYmOEvVv
iv/hb7i+qkoZ5POEa9CNUMZyoxNtQJkmzmbMKgfMELt2s8T2LdLR8vebexR+XI6G
HmDk8Co1VZdQXH23m8OqLNs16xKkrTyg42Rp1EABWrHRxYeu1Un2JKuI2LRnb2EX
YyqLRP3kpDyAQNyaW5LWs2jzuStOwEaQ/iFFLfcqsjQCraGIqlv4D02IUFSl1RPa
zNwXktdR/yDga4ig2nCU5Acs2pu8+W9Ce8rEM3ubNk9upeiOEl2opoNEbF5IzVLe
au/yOZBg/EqUsYmDXJySw521di4LaQLJyNH0uWbLtnHlfOrhaDIy7eTzTzIGJfqk
pVCCV58PX/wBTsYWHa50mg9F3hb5e4Pub9oQVNkjhajwO4rsWZSXoaEIMroKIZ/8
B4n2PL4Ibx7zT3PbnvHhoWsvABpI/MgJ0CQ4vNbe7Savfun8OyAOAabEk8Cg7Us1
Z69P32rWA5Jz0acszN6oMkSoambB3FRoagX+s/walCTH1wZarjO0a6gUxeU/3Z9J
Bj3ytzDct7B0I/zpBWpUiDuu4nxnDLxSGocGTW+Sv/hlWa4v221slFudpE8ALsYc
xJ8C9BFSLlOtgDsXDRptZD06TsltBbUVg23tak1LT83pfPPE1hc/UpKLdVay2+vc
eRnDVi3XuvJNhRPJ9R9tLk0gEKQKuufPHBdxWhzQVGi3e1TRjmDhlIlxUrhn6989
Pe9h3ushqxzICXX0ao43wj7UnZJ13CvUx216GnUJ5faf/Uq47S90PCJwzrNRLqkV
Z/rXo+0p7CaDOlfYO3KyHFJLtmtfh1MNCXx5ixymdETef4teZKeqQheZkKfT50zu
9tAsQyzGY1dXqL/aQOQTjnPxqp+4oOG0h8Q8vFclZm+d4TRnTATezvRoW7wFb6s/
YY1NtOBOTeQbGb3X8OmWZlUNmZQsrE/E1cDtYmvRsPwLEZodunmtLl9CqbmLLKPM
s119Z+oc3w0sjZFxWEwDdqfQFhwC/bF15tNpNBXH0X7EohY4N6/Cjh5XnvnlJQEM
fhdRbBSwJlMAQ9Q19bgVLp4do7TFiABaEui5tE/knCQ+eVOt9CEvpk5mbocygJdq
q0NBvQLL2PqbrPwIJyvGFTmmwkoexDfSVs3+tsD7MZrKpPiJ8Yuzd7UnmEYRXlBq
pPPEDA8rXti6v8f2WVl6CUHcLAsTs6CKZrHEnQXisQ/kynSCFudmj2778vQ/PkWy
vcuSsMIA1RKged0zJYUcbdrROmcs3FoIdiasJuXxAbKH871X1rE3zb2myhBHeTVX
pM48tOHccVTl6m7jyZyb1HK1M5URtQB76rBzD4vVOWAhm/XrfkSdhyxjOFi/RhAW
ay/t3YV2S1HS7oPfd2Ful7nfvyBrQ927R//lRURdvJPmp4m6fSk88RL2Gr3UINbF
YKeBhl5pBaH/qbdGEyukNKk9TLdbwx6rwZLAURmKLzs=
--pragma protect end_data_block
--pragma protect digest_block
RMTtW6Zj8zgVgjLXFOoYrfDKpvw=
--pragma protect end_digest_block
--pragma protect end_protected
