-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "N-2017.12-SP2-4 -- Oct 23, 2018"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
K87jqmDOpojgpVvXFiBw6dVad/qoav6s3Glm6iq9ligvnGj5esCmuckRa1XVTq2h
XDTm/w+IbM51oNa6dCUEX43RRSPR0PQBCO4YfWreoK/hHKYCvqrEBhzAf+JyqU7q
nnZh8/MdELn3H0+WEKfSmJXYtg0N3pnGabmsKJUCXko=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 8032)
`protect data_block
PMQQYJ/GAiz8BPGVqFTeFeRCJtkGl9wJf/vSwHKg/eBFubdyxBv0iVL8aKnx7fKd
7PTXPNQZ9CaINq5NFzBVkPqTKX6WWoYXv8jHUgouEM8ISV3++2ywM8v+yuiGSWN8
WT1sMAiEwSE/7Z5oHgXOFvZAZsaUbNDv4NdIVy23IRAtUphpuYS1EnfmMSHezQRV
hOCgYF8hEPmQZUIPff9/Gpl5Mlz8zMWd1jALKg4nvjzJZGNrbnuogqwhe7JK/l9m
LnJT/Y/UF0FRo5kvXOz7Tcj0lX10vQ7sMIyHAjF59tKA5QG/NeRtkvddpV3jbYxZ
EErXnHQ2P/6+QOnCX7ivfdyg21jx+cj5iEbV8VeWaVd7SAU6Kfuvp0wELg99EblW
zdxsJuTCRRaN1q35rfj13Sh1MKCDjoq2XDcAySiSJGGwZnAtkDrb1q5O4kHh5ZlL
7Juri8+tlyyS2uAcSaS5hsnw5hoeeA9CC0E6xsLvxXZK1nUksDwtCIdZbJljMzrH
YUTj2+aynYExWQPTOLf5DgaE+iIlZHWXwwqvxE66DNqJ6yo9H5+388MhYycm4BIy
kYL55ZU9r2N3FgJuvZdYTvs+cr/9x4HM7H1qqro+0ARoX+BLRxMbmsUBOePzDhGo
1IWWT8VpXsLUWAdzq1JZN8c2nOLuRQQuIRt6mo02+4QurBA0UMvv01wRDPITd3/f
ochzF65g/W/Ju7Wfpbiy5liAbjFb5iEYkuAf9MSSHWvg72WJz126o5VBcz7x97wo
WDNASJpKr3G4XGWkR4fJ+UsHVQrZm8fbM82jNc7naEKyeVypMDLfCrCXmlPVkF05
ib4J0ghmNY65JcZ2d37w5GkcooaSG3XbIYgQ/XZhjCpfeIM9JejtuNckE7UrUtuz
CVGzA83CimHfUTsjRRUbaUr1/NK1mjQhqOeJLimf3a4ek0if4tnMzFiJD8SOz5zP
CGbl7kbcIGU1Prhmd+0GN7rIT66MFh6491wMruw6FZz6zd4rqK0vkMMGdVxwAmPi
7pehG4fkS/1yrM8biZC6Br1DnMSDDXbriiTSXZdVlFrEgKVD3hM/84xsxdoQ2kcu
UlirLm9NKXOlvKc/8/RqXJFN+Ghd31MQTqYxpAblP490kSURFc1/JQD36Kx8t+BO
AK6xWyVlsVM8abu0eEgvtJOIlS7KmrK8cqZ+1P5Q3ri/DKtSQEAHk3r0ktjjKPwC
jVAQkVuipSuiIUqFlhyw1kK1IHDpWbCyiQGSjIMiDuEXGZEQA3ODE9tFFFwn391A
aN6Tt9T6Bj9AcalSeLN3ryQwN0wdkQMVoi51V0yaBL2cNlF2rhlTdi2aeNZkqwx6
KEDA+jb7H5E0OiA8eTsNCXNPbzHBVS+vyKFZkdaxbvMagoBs6jmCjN7uLWjOXLsZ
egytokA7yVIWRgkbCxfneqYn/iNKP8i2JLf+lmSWmcb2uac8lb9DcABgaAcx2vXO
2MqTTgtLVZJjW8XBAiEiB1Vq4lwVwe8U203IOrr3DDgxxkumslbMi40SIWk2lMjG
WOhemWPnSBmhatGqlKCEbl/vDq+VR9g/jufuBLqFtOxEtZgvmvYn5UWH6zI/HZ3C
Lee71uWBmXTn39ywycxksxWK2VEZQEO78Y6ah82hGFsGAVEVpYWK11BmtguHwTw4
qtzXnfgbLUt33T05sWwUDGomIDtFRVjN8i+/zT4NijQThviLgTZcQ+lp3jc233dQ
jlunTtaPvFsJq++ONzi8nvA+ayTSV35/QKilMfVF7UKqJ+vZ8TMqufFD3ClANkhH
gWDCy8/JjkG3KHWlMP501GQfAlUV73t0b5nnGKUK24Iva9R2MKYnocgyfDgjnr5n
b800YHFco/4bVv9B4VG8uL5bAYzJ5fMpGg+DYqARimOROEFvxI86jB2Gs9FvKOL4
MkPOMsbOI/UOvP3MviMjMhYoj4gcIODCa57RbnR3/hY51iUHrYSMHIyg/Qd6MjqP
rIJyhTzvvONxGNqiVsjqVJFxto8fqCIY36NzKBA4et1ZjB7UVYODySBJGN/e3SyA
uybRWliGQemqnPgujyQ5YDH1toZ1BjhAIX7woh9ZUTYFS7uPXwF8zuEi0H3Q/TKd
W3LCs4W9XJvCh0+T+2hlychQE81OH+ANvGb8WGYraXQoXXy1khebQGkcUn1/WpZA
RW5MCPSMnhqliTst0KUeEbPwswM1HcAzfESkloINqo4kxDH8m2KSUhL27rIElHmY
x8619nhpOG7bOGQkvqknrmdgu35kMvb//2s9EfBkwTOq3tLem0//zBmVMgXJLaeG
8OYCwq/6qhMQFeEhd6W5gzhv4Y3EmCW60AiCCZxrC8YQudeo+ImeZw+5wn06JlQe
e9fQLoCob394f7/VSdgxS/J9Kvf0gXUoZ3W9Bt5w5tDAHMUd4BFkR+ZXPx1hsA7m
dQ77U3Ixs5lRaY8GXW+f/trTIcjxwXeNbBJs49vP3f+roWS5j0nmz/tSbfv1Fwzq
4LlIlqhDEOIITX8fK1HPNrlfBoO/sRKIzLCXAL6e4Yfhhy+ptNEEB+KKAdOu44hA
zT3NbKegccdLv71cBeLwHM209324MoLv2d6WFlkmfbme/fZ25nkT4uAl2d/KUmcX
tncW/vDp4joSwzfx2EAkswoo7jYaPAfzsryKpWiK5dIl4FzoiAY2CRsOBGVOvv2I
3ofcwp7RcLzXTTW+fkI3N1HH2lzYZJQaTUPrGEcVhZBT20ruj0y5eYmp4EjgPmfA
sVhnGO1m7EtwZgJHGf7zUWcisNdseBoIEqkUo5Eh36la3XoFToEZOV3n8VL1h1WB
mXBBv40B7XA00F7AWjxn/a9Z1mZ4nnF4u6zKcrIsgodcCGlwwvSi/gFdqMquv8xM
bbMvjOdOqhdw63BkLDYqTjB4pYkPn2vz/2DQ7Mk8/KA9EL5/1zA7vQD7/te49mkU
m/yKcVPnyv1vSa8PI0BfEAWHItDvCxP/KwzU38PmFqcT7/2d6/g8gEJ3UNTBS0oH
AZstCdI2Mhi8o4uMOGUUw68C05N72v4OQfFCwZzyNgCRqH8nqeREle8xBebUeWk5
07dYHQDDLdc08N2emjvZ1jqjghbzRGLWThZ5hK6wvHaKfb1h39NLlXvGLBFZ2Rl1
m8OsEO+70dh3POiouI4pRO2Gtpj5Zj3D1hk4huhtubQ0rXwSpEXMQ0fP5tqrTUcc
pgXOV1EH/ZG5kxyJ1awRK8MPKZPepksKk7PbLtMHS7RaK/F/DQ3OFANTuf+2Bo9Z
B4BFsnUJ0sipuiseYX8+dZgdptYAM1Dkj3wmfa1p7LkGDdaOB4iY7xCcWXM59u60
/q/J3WzvbZbZEXQLiL8/DVQi6T6gxBBSOoCjXiP/WqFgKuuIu0PxcIw3Kn/Nrz9x
p/cjTI3Fif9pLe24nzTtls2hl4X1sdVILa4dNlBSQ6oVSpGdNjtjCa6DF98MQaYA
XEE2DMxjgrNa+zWgOISb9qgFBvTi7DpL3buMoo1S7suBluvA3Z6sPdT454HWVUp6
6nVEzWuyFl5O+38kcFt8cW/0PSY4qQr04IbrHVjyDVON1z5neUr5DQmbXfv9/ciV
VHjhP5uXAgZiaaN+N4Pd3o/nGqCu9Q/sXw0swtZtzYPkaQs7fti++jtl/D0ra0Sx
e7zho4RASLIeGpsIOCEoZWYQeR9V5lZfsMDX5jhBxRKWAk5C1UThD1p4ISvFNH6r
OypcFFUDjG/nPphoL4nFAX+NQ+x0juB69SUFoadl+hTcEP0hb+lxmOCcLwBh/Bsu
ysz/AB0gpRTaqu3j3oQr8gEyhpXG8alONjpcf2/jrk0LnEEZDBcPPlGyMWsj2Jdm
1IZRUKbvlEgxZFIu6WFXF3GyP308ykL/CcB8baMxLN71gc73HcSr0EQdqohE915n
ChLVqfGLzpFS5nT2GeAyrqJtc3UzJYof8NlPtO3GpmWPxgmLnKtGkfOJK6ZDLiJc
Mfmeg2ytYm/8VcB7iaE44K3dX/Qr65i5+LCb5PgAaMuKsAG1i0e8u1Yn03atdaNO
FXMAOSFfuCdfXv49w3XaIa/pqoX88cZhQjU4Ig1VyHLbx3LHRljkS+ToixCluYaF
P2oCMRefLzedwtfijB59sx1nnA+7INejQtJSbGRB5pJDRdb8Y2XePiz/xtndZIRY
5NvHEM7V9CFpX5GVP6GiIpEWqKfqWXiigi/glGTNhRDzR0y7sumK+H/u1rTnSR2M
+k0Lq71lVAR5LYXi+BpWmyyY87QIKkLk6j17tIwumkLKSR3r2GsywUArovNPfT8G
P9lEhhiGozezsx5s5MRwLOWkskr1xY3p6/OX3gV0xb5qHytecU4DRefhCdxGJ3fL
BXIkSsMXwR0ZiGCS6CRphGYFYHpB5W11d+rg4/O5Tuebv2oClMF9+7XeDIpsqc+f
Hi5Z7KpMDfNMCV7e3yE4vCxmnJXYiiJXvvNSTEn1SPp4QigALuRAZNeq8nYSQPlL
GZBYw71fn92lKGlW6v+WxnmoqXsfL8Nh5AGExWKoNxFhDAdmLEm/Tfmh0Xp2E4q4
6k8Uqplwo8MEl4bPRBJW68CPRgK59NB59Q98mEXJGD0IS9D/uD2NautTeNWgHf7e
IkSTI2yG1f9w30tAu5hg4T8HUkdqdemS/yCcibRsqhMn/O77yIrJfm/qYQTlhsJd
ZrJxo7EEsHt8on9iUIcnsZFZllNh1l1bibBvEYO3zlboC9rkv8IdbVOWT9q3UrWJ
64Zs0As54MJDfPSPOXdziNjkMrnlohUiUq1yQplAw+3YG/FC/n2NeYQqAHbi7IyA
PXyxJrMc5tNwtorEsv5NsYP1ALhJXJ9tS8H66/RPAbxuRBGmfy9WGhSNz3OZ8S39
cm0vXdUGko6dCD2if6xScaSyhg8rQWhKMABgR79LBkeUSyWz0BfnE9Ji7H+uFR7I
rHgJarpm2TMGOupL2ILFdpliLf76veTJxohLx5fCKmFJ3wLAkG77MaGokbvhuYrC
vd5XPuUe8s6o0KJlbswRgw1drYHbTS72v2wYmXPPou43K0tDEXS5qpj4Mwjib3Um
yGe/X13txfP90LtvGnyfjnc11CmGGbjODhfAyTpwvklI38KCsSe0B2yv5g9HYB67
Fw3JQjVOU8N1IISlBBNFrSinxS7nK4UkfG4IZej7tHXzGAKbnpjRaIlUT6rb/ib4
g6ogtofqPeem50Eg/Vru71tXc3bOyIEftuTCBlRKP0+quSh1OEUOumux7GWAGMAU
bgm0nTicQ3JTCIo8hzR/+9PCnIxe6eju1n5u+Pjxes9YOCJaI6OfetVuraW9pzdh
vmmr3VIX2V+mbLQ6Jnr4MMSDywwxCNQnl35893YIeNHm5paldC3/rn6KQGmEPbCI
qu7r0qxW/tqxXW1S/RTyxGefImgDNTAEDeiwYlc4zkRj0VWG/BriEHn7s3Cy0VmP
tD0aTxreagWP1huFcvAhy25Wt3HMxQO357h2NQCs0LmOYxE+fmpwgA0w80wDBp38
+Sf7VOIXqaLmD6JAHR3weo0mzpBTL62ydTanBqUPolHb5cRIuJEeFUEV0q0ZDOMz
ptQffCSNNonqECVKQWmZLq3H5VQwL+SIPzuP2UGo245iYpBOK6RNvrIt07icFlZO
nOuZ/y/8s24+c0RtRwmeJ7VtQfoftSvQT1QA0iH4cgpGHdLnazK1AZqz6o4MVDA4
67yT2c+Ge3ejTzptCfmpb72dp4NffwXu07ZyDD7PECclOFe0iuH/X/rqFMfvGrD8
NfM0nKoa5RITh6GUx4EYXoFaqOD6fM7tzc2OSOqcrLh3RkY/m6d9cNGbGsOp4IUX
IN1OgE69YDaBKNKveHMiRAMuoqYXALf35iOSlYzwreQKXs06BjjjSHda8SVbduUP
SSc3n3sT/VZEWCQOh8fUqYDXr9cbULqgQAPUHvISmqP1TY3Ve+xG1v98g72jBKgA
GPKngYVhgnSZP3xQfF7vz4ZPS5PHrakBcXLf+HA6XYSImqMo+3WmvDDnwIrIDUmX
cuNjYO38PQ7FuKeQnQIFDx3VwockHiM/R7SplvRuRuERSAwW3MCoYDQ0qd0h6RGP
HvieKc/6STKgRl4lTVXcDjqLhtBeepWGK8Cpleun1tB7+0A/WrMvlKUHLrVkZPv9
ygQrSX2MhgorP26lm7YZ8m3ZAjDz8uPehOMvShf1hSvcw952iDsWPJYtSG6RfSZ7
JZmb0H/SifSNlHiVBiU1hBYq3ZSbo7PKaB4ZXV+kwfg2zZfbqq/3srAKaYCbbPC/
YImyh4JoA/ycxh8/qVu8xtiSR2toc5pgRSXCm0Bia3ofCrJ0qCD8kt8KsHMZgo0h
fuFskTEtxJ4lsx+fqWSU5JrxkrBP9afO6XvQ3iChBQdua/1LYqBv6l9LzIhd8hJw
unULYwu3buY+ZrfsHSxTCRX3so4KoiSgq7WuxMZJT6z4iKhrogAvRPD/RE3Rwv4D
8XoIbgjXK0ut1kQrZti3rIftShbi13dRTUsXa/Bi4+4oJK/fvv6lMwuUF02qsCFM
UCRqoifHE8fk11h7ucxfA4Us//nlxVNVTbPhp5hXQVdQuZyCIhO/5l065N7c0PBK
iEo80sO4kOjc5bPMK8s+JCqeaRRMAbLa4eFu0ntP6D9a3RguIoO6dxQeJCGFzEQQ
0f98HO22jFqSdR3M+QnM8v4mGoBOkeFZLEi1XT9o8IlYbmpt5EWQwhPTAKjlgkJO
JZYqkUBuQLJ+iMDHH4T5nIwt5huKm1Ci/nk+A/mPDh+EZ28wAAPBRtGFcdo1NdT3
zuyTPC3XE6czh4+P6qcbkatVOkiMC2QCbwQHYwUjBcU9Op/muxr8h2yY78j6KYQV
ouFpdEPac/+3gTq04K5iKbIdo+NF9EpIy0jw7GYiNokym5zpdCipERm+RTvIgqUl
Az2D43XcuQ3sWTnZtFg48QLaoy8qpbzFO3b0wSPgeo4BMH+qwRU51odk0BJgInzb
HpRFVDgF5To9pybwktkmX89O2j41JHUAazjYatjvGDr2kka/uYNcb7JJc4i0nMRB
4u0DaUnDtFCO0u/ZKZPbL1lXXYW/7VRVDDFIk5mJodM4K5jX8qGXdoFILE9CsyKu
9yWcQiVwA0rtvyExSI4+CZmw8UpItsyeCfmKCGQXi5djKnXkZJEnvCh+JRizww65
1x/lAgRTiUKvrb6Zp2y3qKJ4QZbPPjaBbL4BeE4N79VKJ+BhswpW/hyAATohuGmc
8ly0TVWmZkdy8vlrOyEhsMhBxD8XO2ab6Ov3TgiFVXrmHBNGJtp8RYvmSJrl8i0L
7G1pZ66WeJSRCxHOj8QMiYZ/9jLWW2jb13D8gYDn43t5E2VpUFQDKdTbWjLac37U
Dwom2r/1VPoe7wnuUXldHVUFt8FXqmpRBpcoWmP2Ef1QJaAAYGLwPZZewwsNAmtz
ppxeEaOok5dnTiVCYF1Qf0H6mKBWEWSH1Dq205BWBsHzqMuC7zIXwo6EVs/mFlkU
kcQ/p7NFLa5Bki86o3ZRPeUMlfxFG8ztOKdgQzsSlmjemvooHmKgWVfoc3rOSgMp
VwXOYK9WPXD0u5BJz8uWOM/RLLFpnPFDpBpscFQkC2Ay8DNnTevECOJZOwkR+yn7
HMg0LVDia4PkOlZOC1ZWEQjx+jlPeXqYqCQfxWTmsn7ddejCcG+5O7AbNlF9vbj6
ConPIKMQsiI9o33dxkdtPOdxYKiiKJhHTCrIVd395bP18ADR8e6fqiYNemafKUZB
i+vLDviXKFgABSboDHPNlrw+johpfRdXqp4U9bmzEryDfFQLuyIlMn2VOPROFjKs
wtaQ2b03rdj5PcygulbA+E/15Q1WkGPcOnsZNh2CWlwjpMiNvMINDSL8rCX3VuE2
ixH+fKaMJ7TDUdfT0HTeAh07ocVoa0KZuztoU5bRfTZg9QZLP4U9HFziNWnQuFYT
xKqu13xq4dY1e8oFVaO2W/OvlTLh39McXH46WZquTnPdmRH7mze+axz5kRr2AN6Y
IQTejJpkdneRQTIhP988duaTnNn/o+IscUS+ERP2DrHhU2F6fLiwyYWautKDw9hz
pEqWgXpnWiMG5rQlXxa4fxtQ/A8zGkQn0RsPVniVHeGDdBjRlXbUVQS00VzlNh1l
24SYEmGeL/CkuaPfsZ5XRz1F3kfyUHPsXkjd6RJr0xEpXvSXtHKK5B4RjfF7qKlj
nOVd8VhJ6xsBMhehVUNiX3e0GUZGLacB0K1TortyYlTeNsekVHtU4ZZpIJYpp69f
cS73m8Z3lDBKztcYhmq4ZEV3HrKYKBt9WFDrwdjC6R+k3oP9CldfCf/6bccXmI/u
7R9FPC6NHwl7HUcz5D/KVCPf63ZrO82CphUe3ifEvHHcqald42S/DdWERXZrQFPN
j5FG2yYexbK2bsoctienvBmExAZCaFa3ZUViuwkoNt0aWE1HMwM5p+qFctxGpCUB
WEe/7Qh4q9DYaMFeidL9odw9Nt4C3fC/gAOiAcp8Yh9wtsrTHmJgySZmAjjS3V/t
aPxQ788EoY13fdS/WlL47ZNmMG84qkRw0f1mPp+g37TkG1T8Ket4a5QLdc/aacHt
9MXfB/NUk0LSu8GqcQ6D4oa0Z9ShuBw3BGofUV0PkYEsBQGdSGJ5fdnK2qWISQFg
WvuHyKaODQnVz5DtbMTZ8JaIyHYzVBWFHt+3vnmXsxrPlHXXKn2vI+HNyPdBxgkn
+fKASV2M8O15W35vHNW8CORoeAcZm8hQbJjZ68bw+tBwj/3zWonqqKAl1JKeAdLg
piybPE4oTVLyja98jIljRpCvIKaXkrCCMgaDNhQwIVgvpZ1mAjRaAX6o+s2w14n4
b5S2i3vUXzkfGXFZbVwQgZwE756mplKCzIl+tCLUrFZKu+Ls9+iLwQ8L1Q7DJZAM
iM9dKbQ7OF/T4xh14P9TTLLZsu8rfTpfFT5kAYx1Ka7r7ODjR+TEzNk+GuKkVp7+
TgIuE7gHwnEfEUnotqt2pmycg1RjBZKXtdim2j+WZ8q6CB9Lgyi+RQ2XPuw3OYjB
d16acwlvcIybX8wP+rsIOClL6WQbM7vMIKvtNp63j27Qqo6ebpe6iKlHTIzS1nHu
wMd1TrNklSrMeJleIcK4jgXJc4MBid+Z9VSsl8hJ1dPHwS/PUG4Pm4tnSRMNVc3i
Hw+deUFc/mSQgfxsHML+FTAPUDGqFsTE0c25ya4CJVKG078DDw1cF1+CeEvwXgEk
+703PlynKNTuf3UR4mpt1U7GzFRitIKEqv9OYSUVP3dlHxAIRfqdRNcngtcnkIlZ
1YrCUKd5B46JXim7lrHrCwCKTS4Qr2/TB9p7Q36N2VVP9a4y4C4JnpThU1zwFxB6
PA2aJabpH+wzJRigcaNTTf8ICThGZT/FTS2IwIff1kw+HEKSKfgd8Z0uc52y2Bnc
E9gpjLt2xlTimI3mx1eZxD6RvG7gmbVP7gvPLVtQfbpe0XD7BLEWskyibnw3OZmJ
95tPEAbjbX5VMW0PZrfy+ClQtpwwozD3jukXaJtSyni+7uGoGIDNlZnqcy1jqzXj
WcoIUOMc946S/lxYo0LO6BFuMYYErYyfZcJ0pd3x/VLxerL5j4iaSx0qwWWZDWdU
DpHiLq4n3+QbeLilBeyRT79VWaFeqOhGCZGNRuXNBl6ZP83GhdQenby1kVQTIZxz
bOqkvq3vYvP3GRmlK9rgUK4IAlCQfDbjsqRD6xQsFRa14cYuxkC+wM80b9QaPpDE
Q05eEIQY3fDZZFYc9nTOQfih5h1/SkKiCcbQtv763pKkkViBhEHx5rz7Uc2QsC/7
3vW/TeHtajpFjp6cbXw2i2satZEV4qMayITh+qjie79QYsavCwgoxsF5XeuVXv8u
idVh8xfolN5M6yKidrM413Nb+i+wGJk5RSBY6Nh9sZbytzX+qzdwrWbrROxrbpp0
ZocMTlO4untRaz1PgEm9vc7EbobK7W4zzijgRm3+aPuHAtyu0OXYhAo7amFsCAG0
9zf2uXbyFa087vvva8xkYF9fjW8RkL6EMu38eoDK6sPEMPOGsoTfHlR0cTgaMj98
YdsdRe1cSH5zo5tlo2f9nRGuAkSp6gm+8Q/X7i5oGNX/nn9hpDOS+lpAHN7efmM3
kQZ16ysuXh5tK0rDgGx8jDOaTmiMcNFrY4gtxcFrnIjy89J2z1lJ9czY4EnFnWLC
c0vZ4JfNsRamEfeSQbojopS519Ee4Vub7Pkj8i3r1aijcSf9YWiOw8H4kcD+PSo4
eelpkSIpm3oitl5SiWdW/m2obcyipOlJL5oChMWLOQnNvAtY+AbVgDiAP4Adb1se
s7tfZolnSSnKZ6Cg0cuPH/w9l7A/NzD5EhcmI1p1PxzoR/wpE8UYVoDZG/Rwd03T
s1Fl9+787+z6CycR5f92rtqWwMXgFJERqEMrRfatFHQaGoQREzjOQL69IuWxreuT
eVrNpGKg4iSIZFjELU77uxZ/G+fXOjyh11Eb0Npa8xEvJyJrfRA1eNVzCpZhIC+u
sWFEfPUtGe+FKwfwxEOeD1dAbtG9mWWZGcJWdSial/ijI+b2AtV/9bUY1JzppskF
tf+nYCPcDAZa9XWN1BZlRXRJTdbzgdH91h1q50Ct48ujPzn7CU6LX8L6ZLh13npl
cXg7rOSUuJ1nJ85yHdJXWBfuguR1KMQaSa+tNs/Jg8pnqSGEwn/v0mNiY7Lk2ZCf
Z+IEYux6v7ta3E5sqAhUyA==
`protect end_protected
