-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "N-2017.12-SP2-4 -- Oct 23, 2018"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
KvcJJFw1pJ/FH6OTHccIqDyApJH+NMz/DBGmLqyfs/ggYqULL6UpjwSqeeisWS4z
4h7vvsTSobohbCeNhNTCDeBmAz0hu8qofp/2HYx7nAOHvWWxvxktXO41lz3qcctr
rQVY7upYxPEURS3ssmHL06vHZKZvJEQ1Jr7yd+sYhxg=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 28016)
`protect data_block
e1zZqy6GDQzYG3hdawhQ/ociSpavfGH8wSZCy+mES/rrLX9dm2YhZOHkBE7KrKf5
fHkCWPkY76hxQEp5KQhjQ/8QGCNH0gSahg1L+PTFLJ0duivwNbshKsph++nIh+Go
SqjrWf8LBiP9Vy/dtz3HT0EKO24PtxVGlnzQNvhZr6HAVPG4mBfUDlvq5dTVYddC
B04mxhnOiJ1+xE7IMkAXZ94bUUGJPS5/WPDorm4cvKvQiYu4mSKO0KG20pD3QYMe
BH6yaoDFXGD/FA19MHUNyJt+AR+qppBevAm5zHJUW93MuARSTgY7ywUZ4qqaYoO6
BVgO/ABDLW5NcEeOBNLcg8EBDEXjfY/K6DXZxPWXUL0x8/oPW5wU/tExeicYIbkO
JIMPh82Jcfv7oobvc92XmKaxpVhkrNYR3rJGVFSevOR/LHk4U+dFeDehc96VJF21
fiGkCc7Ppt1/QtahqCY5Z8uigKp2/H3PN7EHITQIGeMegVdUnwe6vQjyhG1CqzVw
DbY0oA9HNAdSi99dSThImPBbdnvRasd48kAZxUnVAJ3rXSSRFf1BVr4HLnWl/x+q
vQpvnThUzJVESsfQdws8Z1xye5trb5uv1mxC2/OzfxnNQVDk+IpuragkIeFEYwan
rSAqsvIWRRajlY/aIPk/egJmhYrZ64/c6BSwRNn1QnXdchP159x5peN/fthHzIrU
M6COCRm42oLhJ5Judg5GY0iySleoWwirdC08eKnzj/BWBEJ2PVdCtaUQGFTGb24F
7deLhTlKAs8TGL6RyWf3Q3My4lXbj076sWwlrwU9IcZWdyjN4IDacRHdbpzgB+Pb
91p7tR3BgmUQBFUN9nnA0ba/K6Q5/IG0Bxqe/vh1TxrXMeGNkOjuy0fCE+R2ChSx
7gUV8x7RwMDA+hvTuBVzuPqnGoSegFI2llZuWu63SOHeHLIszu4Xu1nKoUP6Bq/e
j8CYwwJBzN3vUB6dBg4vr12Ecz0EvpQvVDxP9U8cNztcw/yRmjufFmPsNG9dAJtl
k+f4KYIYIjZhiW+vYApNuj+9/UxgMFHnywKK8dr9A+Fyhi6+uWndZ5Gj7d62z5Ys
0YGpQSuVwZGQyPJow/7iHxsk9f/ZbCYJoDBfC3zkejxVlRQEVkeRibjhowtq8Ius
G7wR5HafohyKZ2mo5X7cQxLpOlWkGOWtZ0bX9uvLmTmYc6w3UWErtfVentvZ/XQZ
YZqn2A21JXXpYAVfzCPY2vIrhkvcFhQRpaaxzSokatvbtQfaILRl7UpfDwDYQK/D
DIHieaBf+Zjqh4yjHqONWHVjTvdMQf51vCPO86rR7bX7Us76Ay3iaiGoeJfunF3b
P2XSnP5whmHP8jNr3m7ex5ISxUqSKpJrOcVVe9mqv0SguBwos9RnokaJNehLgReq
SwQQ+inhwKgeIoL1+q0q3wBmyJs7RgGRUY+kOL3ImM2q/RikjoShLbDsdPaY/wHj
BoFeoQEOZ82k7UuWo/a75+pe9MEJd0Gi5TGBfFs7/ecaNfgJZBS8FDwZ0FSnuhT1
wd3wcT6j4OmpUb7ezsQcpUb2V2Y7fGpR9TphlNT/VANKaBtaJ2vc4sLwotLzzFS6
9PibR+Lg3owFf6O0YYD0Nu8marSOmIOAOiPGZFoEa+vBX+aUcFVpQW1qfw7oFTjx
4FX6qdx+BEShnL0NQKHk5rVNKJxNjIQ1Np2YTBxPbw0/A63uXLcxFtN5PKHf0uZk
t2a1GpAMyVsHmyO6ulKcUq2tnpEgeOdaGhsPu51Oee5bl2yZ8qyrixZOuX5ZKmcc
o5e4ZMD06Ba6t1G7f1ks3sE060fWt9NalLjqoaErBII8AD8sNLK/SG3+E2b3fJ40
hf0YddX+/Kd/lkUsU6Se58ELOiK61FjAcX4oHs6GwTItTZ/prw/2XUg1bBkKJMjX
Cy2kjpFD6FtZxiFHUIEaHQAGUHt2OdgEV8gdEim6KOif5qh73PbCSDs9FtiwxbiJ
PnCgQDoiraBaCy58Jl/d+r9XVVhMJ8qXSIj3Fs1QEqUHWppvXCEtvUpbu62qTrLC
LXODmpxw14tFIiqoNsp3sOdEP7DJA9/DXlwHs5eBlZQPtpko6yZCaei2NqZWzhbR
TEEXFpHq3pTDwt7Y8OyykJCAsxhTF5hHMuK9XPtcXO/JvCmAqKsSxaN7WuYUEhfu
5VDX3rp4DKydamnRu1HIYXxqJS4LVXtPIc0AQLQB4yJfOJZ5naiVl+BL8gcwPmxr
ex8Eky9bMxc7n+YMKOKXE5kvClFjJxCErSbev0fVntwnBTM8F3PMjVyTp5d5IeIl
vP46atsbXhx6tLaWEfnKW6fpV4iyyycr+MpWgtCUnFyg1fenSRax6cN1tFlWcBeU
0C4VGy4Xuf3d3P37WM68aFUBzdD3Ivl9wqYbsZWKkhXNB6jjDtp4pkVLHoU8Xfnq
DNHbalxZXh2KpsxmqiUGIzvp1STNlnh03llmQB1hEQRI5E+ZIS0SVUHC8oOtSoim
s1EkPGfh1rAXGQugkqQXubrU8nBa/JdVvQIsR2EBfXh6VP7WO2hZvt4ALqzg+jCc
HxqeVDQgBFR+qAt88nZX59saWMfExYWtI3dBORE6kdL9CdD5n2cC4OJrGjZKFtie
CdIToolxh0Vu/o626p2jT0iaEZ7vrd0fKPvC9fXjez/gCWaduTjVxmYJFuFL0HfG
7KfAeiVqxZK4ZTs+htGzGtNbS8CICb+k6fRC20L/YJWOK48n2zchfWTVeZbEQvfA
oWWW2XEVEA2+kwjtGwGCaPIn5N90UgQ0YEHtiP0eBhKuNZHwO8uBukghr5qyQsTM
3uyzhKEpl+W93WnJi8GKLXVsqWx0MqxfhxQRBbJqqweL/ZRV3FthDUKIQewSXeH7
U6Sh5dXVavx2kS4OWsLFTkLPNUqCQrbA6mS5AUZCtA/qLbXpHerS7c9tYOzKjfi9
j+V1kFrivIyQoiQFWEvzF/JUjF2LNNCtEVJk++Q22t7SMSXmArqDuBKyuLL60HkE
yfDe+AaSgmjs8/3BgxIMjQpzKS0A0Oss0QQVstyG88zKwEpyZRvh1pmRp8fhnbpp
Mq9ZbDO513UVfeGBOYw1nL6o8ILzVB6m/jJYhjDkVMqwaymYkSqzZW4FYiy5f10o
lcUkjuf/y+aLus7ttBGtjEjYx1igUBt6zwcQ30fDZSEpV85DbiAYrkdAD81t3Tic
wlUHVpvj2WVTTb7ynrMk+IDeiy3BRTpDSN7AqypJ7oDYAvxnSTPMzYa95emqxHTy
5DxcAehiq8Z/yvZoqSOXUl5vOH6KtKHCuu93B9/JYJjXMJIF0E0S3yJkBR4xjFTh
vK+gAI2is9zjjcntZM22MMIGtSHkfa3QPev2fXsbvKUucWF8JXMCBnb/jtw+tjtV
rVuD4UDui/NUyt9OdQ66WUpwkAiK2OMKYMMxKc5MZw1lveM7fvY7X+RASvURIn2g
ccglC6t5SVx/DPqisgkrh5kwrE4d13DuZ1qRQKFScuANyQYpuwJwJBEjqbKXSAXr
tv65QWFrBjGAuE3Z6n4aOboyDSrvmbEH6dOlYzGQuaZeMJq2qnqrDRlfy+jKNaJN
ciorIZafijucqcpYJKuxuXlaZp3uc3SF+Ben9TibGCqFIk1TWKwi8fe62QP6Fyxm
xB5CWkOdwbsbTf2uzQUvol24HgYeAYviRzCWS4sPDvfU1g5hATD4xvT9HqpRvIfM
ZNAkH56teeTQi6vpvHn7bChqKO3/KV4387I967uW0rhkkfoU3/Y9VIDJHt6wHRay
3ZababXYLioa4NEwBXO1+bnj/1DEQrVRQDAxb8fBlM6g+y96WMUtfLnS+4UhxaM3
B3XJjEefrLh+JfmZ8BPi1UPxaZPSa/AxeNVFJAE+0NVZUnydQLXs4//3HnIYSQUy
Kr8CKMhZCcaq4X3s5C+u7zacGGHgRcpMmdiGCm+QEPyG0r9Y5ghXaip57nrRVycO
T13fPsTC2h4sgaQkSIkcfpv7G1sbje52EgPCfrLvY8tDRLQaL9VCuTH2M2p8K7Oy
NQfqIMaYAnifurNNrlAmCkZqzdph6JmJQqFWr5H0dPtwXjVHFNH+H7rvwVdZ55sC
eMHbjl6P/RKIoVv4gKdmu6STqVZboJO5ong14QQaSk99UloJNoEXvrjno7LwFRUr
62eIxAbIUBenYmtd4G1BOqOu6L9K+ZT9EB3H0cm3pupA/W+3wULO+eflXDz25LRU
AVbB0OtoF4zdEmIjNqI/wanjspxgolYmTS4al7mYsFf1Jav++9UopQqpYRjQAhA6
8O7FbGZRcxQOH1Jbrd2HmWM8wNilzmMaGn4vZQhqSGuBDuKVyV5hiTckoco/4Bwk
sOQO9180noyLDeVvWMypWaJ+te1/g3/hDFMizsbMLM+tYKiEeKCTQSSTWZoowWYD
3gqBJyGKkQ6aYdjIEPh4VxggbV5/gp/g3S01ynwcI5xdbUIxlxSOAia+MTzwO0+y
CPrqk/N0aME+hTFmMHryS7RiYAatzDdyGlWt0TVVVJbEkT9eWVbapWNO8vmkNN7Q
TrqI/G7cJszRvRXwhHoReNMnxcdcrWw8ZvEsX/p85hZOqQnJmnMcCO7HEvr6OXWy
gRMDrIRtnyxWrIvOI4mgv0n8BXE2hJHOtbm4KW/mdcDS8ztd/YLLZRvZe2+BS+XI
xcDcWJZzenLsUYztzunMuqh6OvnscTLJg8UEexPhpun7n3gNdykUjNVvreq8qFI+
LOHQrMCoGO50i7ExeTHTOHVQQBjQkwT1ITk4fdfiIzsawUMll6tUqMofN6lIUNx2
v4hxgBiKsfZkqJdOON6Ad+SNKDaxDGHIavbReC6n+GomFHHXibndoosU+txxQdPQ
S4EpGKKkEdsZ57pbSj2qtLN5hpO4Lxb9ldytr/l6N332ETuB3zSbMUqnAUeSl84D
IyZ7NhvjqioBjMPsf9diRwHTkyWAMm2o24LRAHkJiIHEo3QAbVN+Sid9qeZ7Sy0z
whiKszROG+93RUWWE1vsLgHqNFhYql12tDjwaOKDs6ye1skS1i4p1yFamkNil7hL
hYoSpa28aom9s1JyO+ZgrtSQfuE5HQ4G+W4Dqjz5qyWbVtOI5EunIwhL/S0hWPop
P02iILkivCdMmPOnK5u+Q4inQL3jiaERL+E985HghMavZzWL5siU9zRHaETzM8xK
fnPb19VTrFAg7w3jKU2zUY1xFQo7a2wPUKqNlP7AJevcvhKFrw6VNLmaxpoxP0Vw
Apjg18ZChG44K/R9ihV4ROCPbZFihgTFdkgEV9POSL05gvhODb0bctUk5+SeO7Dg
kTcs6F7ZWejOUgWzts1K/0peFuhGNdAENBs8hLxW3SRPO8kHKWwSNlJC9zPUm/gU
xHxiculOK3O3OJbjBp+LNEbRFvzKMU7Lu4zmD1CnAT2RDHoJWn+l4y/mOfQhsWBW
AtHacu/kK6RwXIE16AbcCvYLsm58gBNrFasfUMDZMFuVHe/xq5HWAx2OQJzPFen2
/hLFZ4Ic2fYVAGNXieLRkJY6A0oljh9wK/UmHPXA+fQttirbfvgtOoxMZ4di6IxE
fRVTRrTXAzkgHImksW8HYIcfLsKaDoGAnLGAWw4lavt8LgZolNIaKj4WS/JSZiYq
jgZYYC3i5EwglJSSolvPRs7H+vjRjOfupeo2Hd11zn1FHyKQHusM75dN/86QrUKV
shbbe/0/kx5qYqAMZu0htMLTAgl24sgW20yc+IXDAKxFDMtV6ZrcKINUE/AUraX7
w3x/8hqrPIl590QvOfdHBlXEsACY/12kIuY9W3XCY/MqRX7L+MroIPP/Yf4/1M7j
WNWTxDjv8AE16T0O3dHn2krUGfh+f2v47UJ1YqrefHTwCoamNNfMVifVNbAIOOAh
dCYQe4ZrYHWE5GYYJZnSR6OeUOoOy5VJtORG+0YuO0OJakdjj/UIL64CX5j8n5vv
1rVVjbHYvVcaVkx1DGC1uiyxAhsyZeb776cm7jvSB4max0cVPqead67q+YTvKlUk
ZE0J6JoOdO+iPF3LwGLwoEYsA3Hh1onhNElnfAh10VwPCMVIciLPvDWU3SlUex6T
MaTfMG9jO7NsX/PUUOidwYvkIOD770xNJ6Du8bk/xi+2alVtEAT4kC4Vsp/Y8p9O
HRsRFIxY4vhLj8mHHy1ZZil9+RrbFqJePzeGvyVNEgDg8lE7aGbBo5+LLyH8xd7J
8/tfNUxH0so28OMxce7nz1Pz6UJ1uIIPpo2SxBpmg4rs2H3AMnFI/3yBpA9ks/Vr
SrtDm84prr83f1gefL0EuPuAougLnUYfzpOGiG7bNS1vaa7IU0rdGcduYoK5pwwN
WjomoiEIyZWfbpApPrpE5IUscNQrfRcgkAIulT5DO5TYGSb70FJhJ0mJfBtIjqUx
vf4+G8RXF2MThNefIOCcr2QT4qug0BAQCby+OOqg9uV3ehylmL6nZ+mQ7LhJHODy
ZikZpRXAT3/JDEuKY3grNmxs4xE6t5GGcpeoKNT3H4vcAf+zY1kBdOal9NDt2Uaw
vMP5x80HIv20NZVEOEOmi2XGy3zUsYoUSkyii4a1Y5I3cFx4S9eKNoTADkXb4fqo
Vp/NxhtYaQAQsYIvPuzT9ArRiGZzQ+GLCVcW01FE0kBeNWT38zVOAxbyz8joW4t1
iyWk4b5hf1Tfh9OhWTOEOKyVk0xXkJqKTFIApQlLmWyGNtuX5t/nVI/AJ2nAv5Fs
I6Ed9QyMiUh9ScaZeBDQBG2NsDtceLPFeeYSxkI0VZuVd6zAyHwJBq9GMj48dsA5
EiR2QlVjouRklEIDg6Kq0wXxYKCgyAe7ZRsY8h1RnVEVUql+EIZv5XQF9+tHN+dq
5TrO01b231W+nONhxPLFoBS5t4/xMitNIWpNHy1x31ZA/ieGLoM25bfwxfukxGnm
w/iTM07/INw2xB/aRxFvI7r1kMhJBnIzpmHDTGQNmMtfSwZ8yl+juibwJFw8jmxp
v4ol5z41mVSDRNa2SDBZYGiQgXKywbsWBrAakYkSXYr+hA/frw9fx62vATetcCaH
V0mZQepD7dGxtctSTUJr4LKZDWlNAQTk6KEEvLgOT4RrkhClzw7gqLmhfZURnR49
Ef01hNW7rS7beP/ixoMQfAHJwBNUX0jxr3WVLWtfU4yDtTYSJmHS8EY/o10CgOAh
J7XCzSGIN9CxoXd/l1IBczAGyQ/rGt6TECGSGKmEVzcIOE28Z9oL2oTPc7WyvtMs
t0F42sihmoEpprMF4ZdoSC9LpVXDb0Ujh19ed9bX1khB0qkhCmJo1ArQnE4hlmPs
/AVSpuQ+Q3yoMW7mICsB6Ua371n5WLReugcmKrAUYGpcV9wSNwwkjKOGFSR9E89m
X24a+R1X8hBtGCI+5C2nsagc4pMuMozJZai1N2E5Cp4V7rO40SANQVOl0cS6hUAt
mbLLS8l8GA8rm/pXaZMibWpLl7CO9oWQy8nwwqttH9aCw/F6zSAoCUp9lQbygO1L
LPNxO6kk0b5AOkezcpoLj+6Dm6roVd494WkEhi/uhb6zIbRqJoLw++DEQeaSFQ9t
ugbz+NgueCwaG/K7DjEQwfOwEl0hpaaXE/cMowusyGoSNzDSz5qBuaFy4LEeEBnL
XtzjaYPRzgQx7Qn+4TqiAjA70MaQC+fAJl2RlU3L0q8tsa0vS59NjYqKm228Q7jo
Z4E1TfvqVk6JsI1d2h8z4Pm17/vDglgyFPYrpYm4oXAUPPYQVEnrra3YUJzKa1Ul
b1Xzt5dTk1W+zWoHmOz6Wb5G2Ib/1DGfQ6FTcvpHY43AY4wSCxcrfuBB6JEb/Cj1
dEuM2tRGKZY+aohyfZE0pwzsv31LQXpoOLkkq5vXk5CAmQVbBOvwbWNreBYC4pU0
yBLK5LYxev7e5eHYTIMfYxu2g6wOdVOHXTBQRTWAhX64AAjOjrBZNFWfmd6Kao1E
sOl/3G2bFLHGQSKNCQgRhq4/U0iM5KZVYuSp53/tOVjBJKAgU4lzKzKFRKdzUy9r
UM4a11s2JO8+EzljqIRjahcD6xvX15ge+VUoTixBb4gUWJ4+zsa7thKD6r938tZ0
svzyexTUfaJhdfEornjj5XXeYM6b4AqoyCRtc0JVv+ec4tLGFXokFl3f8Ttfg+PK
CoELMvgQ3ycxvxcuYKO/Oxr94k1YpMEJoiQ6f20pblkZi9bJyAyItcpyRfEH4ScJ
g7lxR+xSYAMAO2YjmevCodb8y0qZuSkUvC78YJCRWkNW6bTf9JFTVOi7tYSUBuWz
7u0CZpWvgM1mAvEVtSAffOVG+8M6kKAe30Dotvvx/f3Lu3SNW25SKgRKR7rENX3g
iWloyEQJEYU7IjdIfEtpwYfud8tM2g+Mgett7ILs4r8ondZYlkVcEz6m5R8frJJb
RmxcB5rot2Tazeuq9aZ7q3o3/VCwUu2Z6Q04s5xVEfLTE20JBOsFFUfqqwGGN1TU
ihfizNXIF9DMnsxb0iQxjsy1ON4XtMpfpSw95Cf/YGCVkB+MNwzmZgZEErcB7ojK
Vaowad+khyF1wxnXZMndfYHjdJrsI6wrFIzs9IArEAWF2mGAGqFyTRtv4rKSpaX/
2qdXvk65r33Ebnni9gKew6v4ZYxdoNGyHDLt+PZUKZaQK9PV1Htunt2JmY4aB4fv
Rs8rCH+lxb2yEQqJNP+DbBJ+XZx+6NMGmvjXxzpodX/tr7dqDIQIxkA8jDct4Pjk
GHFsTG5MhbGJdCcgvaLH3uuclvCwze6t33HqMF1Ehs+494DaEGG8s+Dv6BYV9O2j
DvZ8kNANJ8X7HcgFcMAlKIBfgx+q8FO67UuBCR63puRAVgrEPYiai3NB9OAX5qAs
LjVWCSOMNAng8NKNOufR2uBAXTFup29IWVdS/H0bJ9x/3jLm0htZUySogLOn1+79
VQMpyjILS+gnYi7jMyMitksIL7slqCkkPY2bRqEv0m01H1IWxQ3RSbAlEKl+j0ZI
yOLZdEEw+J15mdKaP9d2OFc0VvGszQEDR8eXpJXbRA1fhJM7+vRFaUnKVkqMi3Za
A4MmYnicuH6EmW6+QaVuyZWOhwizXhftCrLKVYq+MhLU+qd3wUYq+RhlZeLzLof4
E6QWxjVzofnXRQPe5nTAwN2DaB27ZIaVY+BF574yDAuU8cLIUtB3BE0AT9orLp4P
3BqMKutiurHTHpwhHIolts2JLS4cvBVhVK3tCMAnkkfueSL96lHse7r8sfL5Chhe
xW/lXPjpRTmQaPqfxapZ4LudPKwnsfkWSGebgoGkPB55oVBVRfiWgPp/7WDKqgta
TlYuZEG6JXIAHkwYoKjTlnr+PHtEA2Zn73qQXP/I/FD5w22Tzp4Q9vrX17uFfc/1
LLwlEh8Hrm6Rjr8iu1CrdhnZwRz2i/QezsJWGpKZW95VEfYQg9aLVeNLvyLQlsFI
VR2S7DBHyzF5t4SbfdSNOMtIxMrTVM8Ilxaarx2BU8Rw/DGsiL3gpWcvbAF1bXU4
zl1aiXszl473Nx4fdoB/6rNe3O1Sl/wIaDg1FYRGTHAI+4hj5gYUblY4BBRDGVq1
V3fQ7BVKM+xu1LusYF3M3ycWj9o1paT442jdQ6EEUHje0lefdTs6Pkn62VlF5WOV
GTcaA13IU8M5zWz181IXQdrnSos0dh4wv+g/SG1p6cn8gdK25PfAwNgx/z3DS6dX
rz3xuOlaB0UUBfxxkbxm0Tev/uCGNOCJnGpImKdc1oyTLrZJzLS4wLArprVLwJTF
PFkKwkn6BG6um9UhQJU7zw3Qa52hivkeUo5I+qrp0m1zse+p68AYzLnC3haFXH+i
SZMLS7IW1tiZo+VjEDmwmCd1TYC73hli2Drq8rw7Lq1mo0m46+L23aOknmRTbvD5
kYGnkTXuFinTOZrM3Zd18H7zPp46o3lWtQUgrxZu1qQ/fJnlEC7jTVJTEabHjf3m
WV1d6Dyd/KaG/MDg2nyK9VQoVBO7pZzf2tJ7b3CCFC6+wxpgU51q5jAK6sJtTVkI
Jh/RPEI4DNOsP9klyybu+WLU00kbN6vG29FsJrxEhv+B/fK0hcIU7BS5Eh7K/5sb
hbRAtyA09Ujmqb2F2z/teP6l0yicD59vz39s15O1+aJNt6SkUkYOXyw1aZH7dfnA
n0xPETbShaQG9b7aVbPBudK0sLeZ994yWdiXUGm0bU5GgMw7kNLDlg3M78m6wOEA
IgG6dOPjBU3Mh1fsR0oaAq0pvXR7S+DGOq7MHzofthqO/OS5U4TFwVOzObjH7xgX
4z3cqhm7bMzV5J6kI8IIKvXdplueJ+48jaO21f0h24VbPypRZRDR2PNkd0zH1I3z
jTv+egdkhVpiAU5DNmhpp2WPd7x/zziD4eRoTY3JqDCVe+DRtGciW1AkujSmVBjA
+8ZyJW/NOjJjwQ6zWnAAEAPNNPSXmcLOF0uJSnZ9oVOlLq1X1/rWtx3jmrpCG0oJ
CsGDotnelRcMkT6pAwRcXCFMvA8zjFe3taCu7QVFGoX8gBLerhTtEey2/5AA6Aha
tOE7xVAdD8bRR0s38d9p5MBoCAmT5LyeIPLTluGGd3Zd+owQh7S/b43BPgoIaK1q
rVVqqygMxl+b/EkqdOIVtJhLx0a2LPBGQfzWY7OpyFL76VZ44ezK4h+KNKizryPV
FDynxG/eTQh/i934tJMRuArW9WtZjXfW+yZMvvYV/sCncImeLYuj49cQ7oSeE75O
E7Ai3t1JLL7fPA41s+s2B4xRl0O6s1S9GthFm5nQRwDreK1au9Muou8LsujEthrl
T8S54Pu7UkEssKY00LR1vl6JWFa5OVzVzNytj5SXWk9JXbg0/fg0iCM9XxfIdYZQ
agiobFPOgESWFWgBA902OC15XFbs7eDkOxyBIskwDiK1gdSfhuEtu0E6hKeaJNJr
OnqEIXdgGPqSDSRCFzdnVjDQgwPbRCp4OryG8Qz7nGgzxJZrl1RNKRqzS43KjbHS
c7uUTbgFIxQkRMP6dNMjO6mHqrVcTNrZW4f9dYqbI4TS5vA3OY8oSZPGtEXOexOR
RISUePlS8jBBDeYkhKfH3soWKDwecDGJlIgBNYXLUpIQS4N/kfSWaX4yuVDayNBQ
SeO/X4Lp4i/bPBqeNJxdR4i7YZE7zex2AiwfDAzRQAV3o/0VmjxoD5jos7Qamwh4
YloCmBQqhhdwz8rI6sJXF2Q4fPB6pO9xZI6HIrOFnLYoGAG8isb03Z/QDRyM7/C8
GEa2qYZ6c/E5T/5sCqMW4V+tGw4rfC9Lr/2sB6dm4vPvxCIeg42sPgtz3lFMlffg
dZse1vNh7SABiZCkcNDxOlpTfeOhnpGMQLYYHNFVTnmgo0z3p/TdCBlqoGP20Oob
l1yWySC0a1xVVfBKIeU9o5FkWmOOLr5BQqynx9HTNrI1eY4bGXRo+vVERfR8Ip/g
Nn6siCr8biqsNKdYERr0owon0YOiuGrSRzGM6m682H16u20aCv40A8P+Q32zh/EF
NWV03/0YYfXhv1Qke2cryy29YamS6V2lnttCRqZ37uw1zehZyD6QcC/q/VTPIpqE
2yI+haWOXdXIL3xeZmWybtOC44SFrMghiYjD8Do5BrUoWCl4SmGdvcjx6vUzKZnv
8kKeWtTpfhmxWbt2jr3K4b+oGhYH5BqPeJERp3pJWhVTp+4Gi1/kiMWW/P9LM+ud
fpJxhUhf6DQGl2MGQ/FIH1adL0vyzcG6a3IiqTpozfinCqzjgTw0m2Hw2RoKZzD8
HK0GaVcvmK1zyCQTrLEl84wL6FXZWb6ZYykMSJTuC2wm/LpGOiRstmJosDmumVW+
sYkIgrOou5tpcLd3J/P51WYYdef8wK1sITV/RBaa6B5fGdsf41YUwg9/lwfoJx0G
sdSRJtGQMQBlSpQacj33lh2mv7j57FQ73uqK86NrKx0oH2BBAGjyVjF0VehFiTO8
vSFLgBgVcZkqPAWDaAFXOjv8YWPFXfT/CV1KTyR4EoWc0MEGibsDbvJsPRcPkSC4
bFp23QmKuYkh0Q1D9RGykKO3fzWswLV0F1nqEEooiIDXCWx+gb5BZvnF10haxN9k
ZWKIxy52aIPITTU+RfN4f2qv1cMaJnuvM+qAZf5Sfhx4PM7ZHibEG/y9qcUv/koW
xwFFWBsV8PF7hauQALbGIuMLoy4APtawgmwP7O6xT15HWIr+rLzS51I5SfNWysWr
DjsFk5NKofQHHgLqanIVndFZbeMr1/8tQK/NUxQeovXIz/EIFIgJkTbEh6NrDe+b
B03UF+Mlmd0NAo1LwLjN/WICpUD43pXGVTNMPysnS3URhSBDS+S8LZNSDTA9Kdem
qERbQXTYyCedEvrq0vzuU4TzFFUSSp5WXzBdoBrouRCUaD3ww7IEtopQGBJfgGi2
LFa4oIOSUVrZ3nAXEKzub/I9psb6PNHH5dg6NfvRHHbIcDkViPmK4Uv6OWyUyoyu
+KVVL6F/OzRAqpz8g0FANS9Xw2aS64csaD1+W/BNvn6KhDSwgkLeFl5QUuAcnuTR
/gPci6GLftXHX2vxZedJ+L608RC/58Byn67blGjNtiQwmLYXFkemy0qGdpTS8hAz
6WM7mkbscmjFOsPdar3CHRwFLOeadHjHyLtNXEzBqkoIa9lBlzESp6JLZd0hr+WA
Z6wqoVptScaSDyG97EcZRlmhBiT9HWy4QY8lKrhexOxEYoJIPieiallI8wU0X5fT
l5Xc+iP4BmYM4iKVxvsuCOeJTMz6ZKC+9b9zF6FhHLIqMJWiJ8fQjS8vEgD7kniL
I1RfI9P+xW0AZbQaOkb4nSglE0/FY33J1hvfk/aR60Lw0W9ovilMwzYr/0pbl3U6
nXRe7/FKxEFwS5z6hTqhioiFw++VM4+wqNtYuwjGNq3Tm1mayqOCT3wMD0B31HLy
6aa2gIkl7m6i8Q+Gaj1PvAI4uAExz05SviQ0mRChD3ioyUjtPan7Q4cFqtxXIsmc
DF5Ats5eV8XlQig5tDsvFR3wQTNHGuQCjN8iCML58vFovv/WmylTtR/n3DaRK2Th
DsBnoDaEteNuojarsxl3Kr6ChPGKnr1Um8xjRwvt1+gApJs+rdgxA6KVMn5KCjWd
WOrQZBcM0zcb1eYjHLjWmGZKw/o9imAE2DQFz4siqLteBLrrYc0Q9WunF5sMDROp
Hu2D6gsydqE9zViH7sWJmDIMNcQICY+1ZkKTQP1Rey7+R4nXCoMMLVflCCqjubYT
nKLDpwQUq+n42mL/na5VSyo6FjNP9asduSb8RBo4bP1jp9U2QU5w1ZQ0b/glUrR2
WfnnOy1tDwP/frcXyFF/5t/rzlMQFP5B3IEqdWuDGjXX9LcM4oDCROOV79bZwxKD
fSJLqvr+hXx7u/dnUmv8ixZNLsVtY/okqLCcsAyJOIJD+9sYCQZASxnIhZKyb8Ha
6vdl6SqP4Xi0htPjzXnwgE/pOyToMq3yfSxZS3mtlbA59gwUrRJzGcHD67bzufMz
ris8Fv0nq2ZOwIsNXodi7l8pupYO7YaXnfYRBL6HuY6fhQXSmMc8mv8mR1jWAayK
Dfpkln0kBuhmZ6QCTTq2Yp6oRu+V0z1BP74eDq1aHBJcBp58W5oT+Z3qQbprOWvi
edvSkBPJ3Vcxz80uqggNNE+nk8H6Fs1p95YORx3da5vgLn0Z1mhMctbCPqDbAezi
A2CuEgp/5P15um5NOfrFyeTosBMUCqN93YB7a5TORcLXW0OiZJeebVFXqHieYr/S
p19HYBCxyQT+b29aMnj83B4rZ1Ov8FQbF4DMuthyTKCI6JbuNNLHBEayapbsO2K3
QDeMpfBEgrIxishIpW4KbEpRTe1jAPzgyUNB1M8x7SPOyhlRPbfNdBt2b/v2oPmW
NNxfdLa5yCO09U7zmI4xCiupSnQKMQQO0lOZ+6rXdlXUPtJCps8Vmt9KVCw0mpPG
HNMWqIKIMgtdKm39C6nZZCLdVivxwJH1TCHS5bNIxdPy6XkbcUhVoZpk/kblNbUM
YJixywaQdDEac0PIt/Z2xLze00FZ50cmmf5KQIWoKLuaa9Hp88sNjH7mVOCtc48D
DAnDWDGTqf8V00SDbAdJJi4Qb5qTSrsULQYk15yoGS9zPHe4N/QDul6/5oG11cjY
jcyvLWn0TEw7qABqUdpIYhMhqV/vT5n5E8kN/FjcTavFHhlrr1MrCmVs9lFMnq6W
u9D+1NITWjSN3BeOBW3eWz1KB5F7SdVeayyvfFfEvtNXwn3NQQ7DkhTJ2TxJT8Fp
WNiVh9lO0gypb71t1rNwKlpunmKq1vl/Zz15IYH1knKDt1umZ+JFTivg074oyDM1
LMQz3JmmiIqVxb4KltcUYmNrEYOO5S3A8mbki6+Zqd9dKlY/kSRlKFdgi6AcMB06
OmzB/CRV5dVRwvsu1t4hJkDDjghgOh0GUGRe7m3ClWvhRC1p3EDmvoPdyM5F0016
7GF38kBltANEPawhHod1F0ZXPyopCwUMMkPQyo1obp/3Cbmssh5uo7ft0VHg3y9j
LiO99/AxAsy+f9ZoLnxonYENLqrlOEnRTyAFipS/CToxUZ8xHZJUw4JtE/PXn9Zz
S7Y/6ZArPnRr+IMo0x4Y4gos0eqosW+2NXir9ChUDpzt5wih9faGnLc2rUQQ4nGY
tz3+2H6DYVSdieAlD7YMwkzOZuCDiPW+VK+qDV5h/VOaw1cdGuMmzXyjBZ/Nefxj
Z/ebswLiXy/4pyysAtAARNbmheYtvnCjbHhntzfBhEJ+HFPs5bmdy+EFmzMoc/H1
XqYwaBYokyhXE2j2JARLPE4NhcZoTRS/xWOiJSsa2ZJI4x6EyQQj5wC/n8dqBnE8
i2W1evhARCTI7Q3GmAPoq9dmtgfLTPdGW9xuvUJMMwTNqO2ACrOEFKZAeyX4n5aq
84ZXI6oNzGEseKZ0BU8brMqY97J99qQ8PNI5ROuY4kBQbDWq7f5aTJ9Pq6/35IGi
TZAyNpYjgGevmTh1G/l2RIt/QZXOlJoDZU2+pW9Lv5Ql8/MYEzOPO1BulfL1t0Ei
LMntHkUbEJsovm+eEAa+nsqPk0k8HvXX2qlw8ijRWsh4ygBmJzIDrlAokEkDAW3s
XgFKSLrZ/VuN+8je61ehU8fTfGc001hV9mDxzNnYYczm8A40xtKmMUZDJBAvTRjd
ABHyWKE0m/mfPiAgQXWc5uKlZjJZMsd8Y0O2IdIEhnMzp8fQGOQSy3DHD1690QTY
HhpDspkwibp9CxB7dOl8HJ7Uw7wBLtgo7i7deQx2mvgf8bhs0p4xSwCFZ8mIOY/f
IDyi/xkhvjR2+YAsOMvJMaoGuXoWA1r753hYWwXW4EU3ROAJRjD/C1g1rgj9iQL8
Ps6HjnPoNY1VKoKw9v3GV8F4paLmh1JOUbkb7jSMKUGtWM65+TJGcKN/zf7mW2D0
fk6YggdUPWldOrXGisF+lKVZ7bJM2iRN57ebWXfjhNiW9j4wm/ldUoVV+PeqHN6O
RjDki9VV5TLZN7Yrgqo+HTRdx5zvMw33lpSw25Ck0ROF7HZ7WyAuecSPQBR59JjD
Ur6oOJSI05s8yqnsq0xEfKRt7C1xIYET/OWz+4g5i6SSwjkMAr6nOUadoqbnmzhS
C2kBpu5L2Sx8ao/O3W04kCaIYHkMD4Ywx7jocxmU6n7pvlzHmZuL4Pi3KHOS96+D
AgPDKXF4WIHRoI6QI1cWCLD5SVwKmppVMaUCQiTR94vRWvJVkeXpYFiYvSuh9qOf
07ezwj4B8BR12m8gwABJvbpdKjsQb0WBY4F5DtpFtcqd9OcjTH1/NB1Kg6GgRgPc
dDj3+hwN8lK0Ve4WlBXCQm26EtiQmC9kS97XkSENwtACxLttBlqah9nnkqZ4Z5so
FUJwjR9K+PkDTCLeIiEGx8CWuE6n3f1/7zyrGjDm1t1LnxlbRQGOtFc8S1R1vKf2
i+IXOkApe1M8wGlpbnUejyJiIxyqsKpJBREYKpli10YgB+8qWCQ+3XB5YE1zT+jH
xNYD95ExDLirdMa5EUHrtmQUXozxbToMdl0hU/8rcyXKQs3qxqzUbeHn34AXul2y
xuMCWTgioOTc6U5t7C2jEIRf9ofQrklSWJE1C02e1wGg6llTP7TCfHxvtVkAjkd+
tg/0DXpXI/wd9ru9Tp74BGNKv7QxNRfP9lahfW615A/lv3OE2XuoQosqh8MkxYEU
zp1seiFkUbP70ryE3KQQUnnS4NK0L4YDiXKQrdpx+AKTNWDurmUS8dbva38sZxOv
8osWFoQUc54qOQvQnzPE1OC8qTayUVBnXeRw3M0+lR2gL4uttUADOWRmLoLzXDFq
SH0EI6iKDat+i9jtH0mAoa4IXCBRwZQeeklS9Qk8d0j3XjrEF1eQ3nkooksZMn0q
xujWESxK4GCwesn45LdeIFaUnov1BJv59qlPcBLeu+pXkIZCvVMKBtMMycjGUSgm
5ML0c+WGlUWD1HbhRoRQGyCpM6c5uuWeirOclvfEKOe/e5TsV7VuTCvVlE8kqwFy
eHf+IhXsl8mSbjwAOVDT1jFHQzBVo4CStLeg1QK8otc0PedhUR42x+143Nvs830F
1mjUR7QpwQqqpIgjb1YuY6PCyWmr/WO8WYN6jrEHvd2sil25shMpp4ssy1ylzbYv
lu06tf0yYEneKlUhPvjMuP4+ydN7pMZxJUcGaSzofVEsugaVuwbPz0L+PtilUli+
AqnpT/4eUhd2b5kQueGpl8XbSqXB6unveLpwOtFCONIQ3LaE44onNrqNgYqQVznu
68oyR+s1bJ8+UlTGPpZ4SHgLr5Ckc6RPhMZmPGfO2sma/AGIZHdBaFScTjZiy2gf
7UPbitkOysUBornjouT2pmTbZo+0rWUsIRgCVBr2JuYZ5x2RbCwEf3TdAhpWmLyj
BkbVQcMvJ8CwiLtirQ1QNGauqRJkMrnk6E25N0mRa0fHep1mA2zvPsjZzKER5Ekw
Uh2BGARrv10cjpCvskdRZcSsG7CRE/z/cqtmzWdHx7RHFCNvUPfDgVsFnuG1G/mW
g5vhueGqT84cvppymo7+PbrhuhXRjbpCi5WehY5oJWQ3NsUjMmhZnBXsR3IefYkD
YwL0wGe0qifg8ka6wAdVGN43Pc8BhscYe0GUUZQg25vvcyADMkLpB7oxE++dtodJ
TUV+oZSNMJMwRE/Hh1BVTnMDCFvVpprNH+mDDbE76NPxPLxFLQU5X+Du/isX8wct
1skQQoWq20Coesk8MKMxuI2z7T4DFOFomlzXdDiTAHw5rMyk3wK4AkYP0FqqU+W9
sT9XqFXNNAWd2YCM7COGfTAKerFuKnAnplTjhjNHzao9nPjDb6Au+0u54Vyd4TzU
r1ca0kCMxq3Ie0u0qGp6dXA4snRWJKa6XMNgfsaeli42U4ylxRGGbE/aYTYX4JtE
DDYQkO9wsx6PjRd+g1C5fFvKnDX46VZxcVadh4aHpAmU0tR3c6IbrN5v2n/rcoxR
nITN9Cm3y75cJmZx1OPUm6M11c00uPtf+BbEcQGAY6c/AVjGMJ1KHH1Aj1/k1K1q
sBPeKXhiDccl3E/45B6cgx015HpKB5xyjuJoU4WlytjOEm79QqKJ/lysFrhAQGof
gf2QbXPBmUpU5gkSA/PY8rQbvkmgzBf6OwJSv5Eo5EGZchA8uBqi2nNn5IM9JdTa
6mEDq630h8MgOH3kVnxKH3fiKIJSwQZBPtmoqbMeaCyXA7Ud5U1O25KAY/K0X77X
DI55vZS2SmLnJD7GPEaHA6QD7fABEdBevYfostRjytxtaxNwYSor2B8MP/uOdEvv
NxpBAfncLldol2sDkUHur/C4e4XBgvbPBDE67GPsTg8kXliAZqRZTl3P7YIDK5xt
Ysf6OEkmli5TYt1aFBIMESue6oY6yg4DLLbsHnFlzi8XP1+eXSCECdKBp3IPHd7G
4X/HmnuJjJr9DqOCwlAwjXjlL2aEMT3bb9pqHFH72bDyDV/GL7iKiiMaWZvdh4vC
J+zSLDiGYTlQmReHwWLL4xH+ckebquMzotV8q2YvdxzYkZH9jLNIifqRC39+jNl8
kTZ01Ll1KyTEJNeDQf+IKoUjnzjulW1wPGFby8x+zKdwVp1aYdUbf1l8clTCek2l
qokIXlxZ356njdZ3IMvdeJcOuimoe+oBwlJzqovRa2sOKC/qSsHFhDfuJtxmiN7I
bE+KnHYSHf4VvOjaZFakdm/oDFF9BcZlRdPzHfzRJV7kcuIcq5UU+iSPFnvzpdvv
QHE8yWi4n67lSyZMxfUlcWV1PBvTFCDKq5EIOzCmBX/fN/xQEZJk73Y88kThd0Wo
hHZJSQUyvd3GsCCcdUb5ig6l53lIY8Dsh8uHQWVfYrCUnvpm3RanCsAz8sZPma0Z
n7fD2o8EEJzfY0LrpnTmAmX2dsyHOdoOGb+e5Yyp5CP+X5Ybp4IocJofL1I43ovj
/2op8K9VeJ/WYq4l4Nqa/fCN4XoBq+oIVRdG82YVkP6tLQOTYRasz6rkSH1G0iQl
PFcsXqMMBDR/ilfIb8eowxKeuKrKQBiJjmxnEzIhLWIMDwZvQd1IdOZn+yodvpDu
MDe77D/czZqhE9u6RIHPbUN2fyxfiO/+cKSia8Jyp4HquPJdHqLDx3M95dMVWQrq
eNlooaBlrdvoo9DQwwqGaCMznBZydU/q+e8RMtRyMmtyknxcdhiEI9+dTLvHlbiH
2RXfoyvfr9QEkcxl18vgR0rm6HzwNYNorFjn1Ii02zMO3WXzQU9dNNlgtPJ7OdDo
rc/hotHqNZTjMiTtICtb86eGvkI7f9qI1gDJukZ4XaOwTyaVJt2rL+DB/9mCFXzO
eOkF142bT8tGSZsJbOOiyK48sSn1jr4J+obttfLAYVHMqKxEKiIoilTFGqCJEXaJ
2R6o9BYGGZXQ53c3SVk/5e8bXy1N5QBdpazVuHlWkVThnKrI9C72DBvwKS0nPpRM
m0/idDgMkc3X6plKV5jcuKy4a+V00cP9x8cp+VrO0MEHkswO7pJCA/kNonLaYzIM
zyp1dtKZZBB0xYdYhptMK3ZfRz924lwpxYoAu5uarLKlK2c2lW1PX/VBuYk788hm
l2Tc/HcxGNQiF+GaqaDT+3A6hemWhWZuGs8HD7c1iR5lyeQpO8s3f4FYwRLQAals
cz6INIBV6HM8QH/eYSbBsa+YnJNxEyf6BneGQKONPwvN+ZfRn0/nTix+MXTsx2PE
3FwPn79k1i5q16WsiCMTVJ9RedcKRH2d0dZQE2WRq/04kmNQUhYmNiy3Q0TD2BTd
w8uvSqO4xJbpWIrFtvddU4iv0mu3Rmj3Z9pKTGxoUeWuPba2LEYzlVGO+nbmwgpt
Lih2H5O93bLD4OnyvJcKR54Ew5W59vyz3V4wrd3yX8Tka1OVLMFNwCqJQWLqPB0l
/ov01Obfw86PUr8vVP2YS+oo5HzqoWoeRRRFdX3imddIvnhDN94zbpPSOXY85FfF
rAkpVl62kIdOAO6l9Eq9BN1vpa9JK7jUZ6PsR+3EblbwfhEvi30q37Mr91545YCU
ddiCr2m88B5NPJvbQjWcBedRPZQp3HmCUm09IYIO534OUMUdEy79UAWqAWlAY9T6
kRGbo8/yPluDL3kb/5epo2y3Yg2w2LmtA6RMg367e99m2i0hlfoiwkdwedKcFG+R
7hzctV0zrtd0kD0plfVxcwmGWlWJiyFqFDPjjGHJWI9h8wh250NpGqYiHFasqFTd
rAfouQwUWEG9XBH+Z2xoP4EuzTJAYCNO09IHrng3Wlp9S69MZ6l6ztw5xhJdB41B
HaSD54FCYjOF0It2/IaRYllBFMYIFxn1MrtW07HVdjC0rt+1OjWGteR20AKOiiaw
f61dtGkB40UDkLajN6K9OcpCiMo3dAVCDd24VOGid9+5DiasZvllykPqs8ElI9oM
x285apMyLZ7MXfdj1b0cRHLUccyd8Q8s3dNEUC71SsTN/qETEFxb/LbgdXDoQptT
fCcQmL009qr7aRDIn7Q2WYW/s97E/4L9GJfmmbu5ZEMoO2Cyln3zR8LVt9hQIAX6
5/w2CJJje0whqB5S0uQMjpbGPC175mgWqAhK0DcfElbMo4KocqX7eExIsFH9OMCP
z7IUkGezYogJLnWfUXMD4juadPfiE9PeDaABzD3OAMYFuQ6GGdd3hDqUsf5eeBsO
uT0Y5j2JcgIiRVyz4mREb+G9oJ7QhP0EMAU4GRvkEebvIciQih+65KngmWM9NqT1
maPPiVvhZTYBXlSwKWhb0sIyxFvWDGDdgzH6edIK+QSfGIDdeJTUIlp+DuYz+yW1
r8PJBZsck3vk5gCP8BRQqcTjBJnBEBsUDR6YPCQp9/XaCUkjwRf/+bspfnGVbAf3
4KhkzxkWtruemQOzPWFbp9ALqeS01eidaRjnqv9l2tEDg01vWjOmopp0WdJfrnvo
wdwQZav63GtKMBvrVdp0piCzhVAboUTPwvnaN++DlBDl5dLvjScIzcZLXuvAIGdz
JMuDamqlZCV4oimUR/OYEkOUB1nAT+LCVkts5fT3zfqDwkwk2qoF3MEDBRZ5BM3S
GM10Wp1sQUgME5U9HOn1etFRJ2YOkbgYCE5/SaVd0z5M3rhxbI67JOqb53L454vI
Rr4daqLxPMdPMBvSmD9M6ryMI/XOjfj2+9UQ+AANycSni+gH6cejig0PTlP0u/Ro
kM7CflmS+L+/X5Y+xFB5krjh2CyQV7tGKlk9ydOLam5b0gd5naclx6z6eJKoJ0TQ
KS0PBW47QiT6h6+Ddzu65d731XOP9N1uhrKBwWmE0acE3Xk5l1F99g9Ff8oSyGWf
UThnxqXmi6LYxdXcrDE7oNf/PVnmafSk95WDCIMa6laVyptzM9ihBP7cmidvULR7
eCU2Kd9QxzY1YoiIUWf9DXOU0mTuhArgYPM81mSkdea95VHxjDFQw3XxWu8VbfJi
fHGiCJvYGob0LeAC48MjoJ9PlIibloDkVYXMhCRHvJLQEZ5o2q4IKB98GRShODt9
j9JB08bj/4VsEKVLhtSvsFaC6f50ytqxtTT+NbcMmMKZU+MYvIhL4wZ79wocNYDC
ZcEMS5R3BAfdW+jv9pC3PZMMkLKGOP5C6/2T/IQdllzbDUS/o1AO7Pg6dGCcBsnp
+/80Bxmf0o2SSLklbKzUw0x7cUvBuYE8vqBSkW4bpx7LwkhF6yQo2Ptpl4OFaAay
C2/MjEbrGQ3kDymibQ62dk8ixIuFu/7B1JkvHtJe7WbDWSAjkeIbRceCf31lrMO8
F8+xpcMlfDTMk35PkokHLK1NQbiqFR4ApMXx1WHk5TJMjZBdQtCnVJpYO7uCxzht
nPO8h9AmLMHmtMZ3XwNbBErC9ZDW1QsYWV9rlTFixE8hhqqu/PxwgD8KfrDgONNv
64oKmHEPgXGtmpqMlr7bJalBe1Wo13IHfvPfcUr1g3Qvc6WiyBhoOSkaxORdy1jw
h9GeouIsh0kxsodpc2rQhuHnSly2lWXdCawvCQ+GJTdu8vUzhuBl5Iyx+VIYktiH
Urq/mi0TVtopduZAEvdabJVl3ILdEcVJPsn+lPoUP59CYlrW3ZlRypnZGib24vnr
qSt6uMCn99QPBGFWE9w7aQReT4NlQFcAZZBFxTpFD2PtbKAKqCA3ZcBJu3aT5sst
SWgSitowzQ4VnGjPDcKeWdL+QRSQ+jVGGGj323n8+OU49RFcCpS+oOdWZMP9cEYk
Hg9futxtcHdLE8srg6HUr+H+rzlatDkd00liYmyVe1PFewbMRI1OGOG9FZEzGbA1
E761Iv4PMiX06/DoyJxukPfHW3X2jHZDExdUM4GeMGPydW5uFWNGGXYuBZDFiN4e
LhxWkyz8ImHIo5fysYo3mV0oB64bbKZAB6cnZKzKbS9jkHGnzOTJWdHqvcpS63hQ
LdxpqTwoYiOLinyLzMITdSGqYtFEuHs3p11g8voeG0AWZylXnEWEc3Fv6ik/RSAz
hKiW7OI7tpPn3Zf8HTSiQm827QOOWmf/4lIYBD585vKWqqlPY1uVNb7IMMhkG5Rr
UAqwpSB4zrLaG1sPYl+ytIk++EFFcVfFwVXTXhQSpJTolBVgzPd79tEMowgIGZtW
p/F+q+PzSXxXfGYpPZNA+BH3X/9Oa3oAr7WNbV/oHTFA+ZMhKPtK/fXqgVcvv1U2
yhiy3f2q2BwIrIq+VI9UhI1AFGQIKsB1+URMr4kgzmVMTrbRRUArbVtITqAk6VA9
OleMFeSCGDQSIpJgnnlAfQ7Wrq2HBlI56AZs/Q5anh5pgx+Y+wiKkX/P4D0medJP
PVcReAZJAoRJMYAb7suzYX40039lK7VIfNpxmB4Mofhl/EztA0IY0my/fc5HjbXE
PBZ3mol3EX7glrvFmhKDmqSr3MFTDZ7riM3BlKY176fuO+i+qJIQVlD6JdaVBlWx
r/+z0IwJ257ux5hbC71LrlkLzNaly4CfSOfAriovpT1qxgTdqZmpvyaCOeixUVft
IR6uxpbtJbtdxPJbK24aanugHKw6Lgc6WK6WSIn9xP06OJOdIcKvy3QqvcPKa4zf
AdDhMzNGpW+7gqyFwwyrjpB1+jDPpG9ssmPonCpJKalZuotJ6Z1Db406NowBZNWN
iuzrMPcPUBbNGNzXo6eHHnWke6qLgELUF1KWfqPhQSe3nbbjwe8CrlIUA9pJR5LN
UJMMuz2M+8tVrF2Qw6KkWyj69HvBL1ivCYRkYk3CBomLSOCVeDy1MA7yNtcs38g6
+KG6PmAQH4M0XZUQG1UBKN8V+tP2fPdwwGfYn09R6tAzBMwd0qXOhpveN/9fPtBu
wa2Z0FGdsTJCdbMv1bX3zHp05NbiR98u7H/uo+VFM15THF2Tz8PO/rpVba82oLbe
nhGFfI4/X2RwmI7m5NjVbQRbLGMSpPvdyJefBMygQv0xzYpL3T+NO29KDCUpGcH/
zrfwKyTjLsxSOrBCZPAc8+/EX5tjzbcTFmclzqK+mcIRUuwAhLsvZwPsG/oY2v9k
cN58quYtlUlOCdk/LAWZXadcJ7NhV5MHwIPGW1OWhyVDBeGAwo42xUJa283RrI6d
19r5/CcK+cwXTTiku78HhXUTIuT3miE/hqiwFxX2HFmpoz/eoIOtbxffsIznOEwq
qmfsB+8EsDZiZGbfLpD899yQUBUVWj2CiVAkX6wuZ2IoXo8L59dXBfkTna8NIkj7
GxhrMa4ouZdcrckuvVv6tsuwEQQqpJZAqhJErA1KsTwgDVGDMI3w1Kq2C0820bZD
qaBClb2w0PhjogBDE2Jg5fVmVGKgrhUJGElrsFQXr9cW6EnqQRZsqGIMWA3GUEpX
wB6t9CUSpTdSUXTtESEFZhQsf/dcbzftdjGF5C/TSf1z+UFaExCBxV7mURQc5iUd
bdTmvEOzkB2IQUKIZuuTFrpl+HU3rNFeEVjEaoayb1pSQCn1Q30c7VoQGekkGEug
/lNfB44DtF2TbICeBPHnR+6imamUSdW7Wdfak7Z6xqcwvQGHMt4Es64LmZ/N+j77
+faMgR8VK/lx6+toALnYlwFX+RX32Mvisd9b88CjN/y0JaVqbR82rKdH3Fg7PCyF
vdylqQMKOfFtfrbssrQz+XIbPN+wVq0weLchzIY0gBqwUE2opbEv3K7y5KArt/Pf
8abulpc7eK6KbnZ7GWXZ5+L0Dl1vP5O3+8ikJffwVZPQOjknxwGlUcsoTrXnCg8f
BjbAJzsWXejFh0tkDogaJVoc/iBhGYPZtuyKKFuklmfvVjV9PUMACaM5vaXMHOTV
fttLK38vkCjif92NjKALUZO6t13FTFUcTZOfpwX7j65WSGbXpvCd0lSkSR32jr6X
PW1p0kg0LiHuCqf5eLzFSL5kX0WExcBxTfy7/Z9ZAoJFqzbSkZVei/m9LdW6wv55
NMtm6N9Z5jpBGzwTBeesvk4wmYwIXslHOQtaK0J9wyDLTbjvhYWQXFhlEGlZvxSh
D6t7fkMdp3ivPy8TTLGu7X/iqV2+JyL6NYy3+VCoNDTo9ILuvVI6yvyyYfXJ3DWI
mvkxteTi8iT9RLJDNqjhEtuUJZmD1qLw7MFJWFzD8doim+8rQjAwkC/Oa9hgFUSa
32mUyXzMNhioW/zPLyxjLjl1rp/6Yo1lK3GkpGuk2LQ67QzKS2+34hH7YoOqhHwR
8HeOC89Owzuu4a/TZg5ygSYQFy/7/Cfzf5NuHWx4htrhZmBDVObgfKs8wFsXoxcU
PeT2rqqAKSRV6uJrQZOqoI9/1B+yegwFpIuXraRgSbJCiqm/qDoka0VuDqhsMmiP
/DMEcEE8OcoxLBRtaIOsY+pyXTJmg4KHH4e56GwY4iGDbiG8iWXHiwHGF34jzZc+
pQ3MJvPA1mi2YC+F8T5CPCL4HmYkEOFdwfiR0eTMb5FAgBKu5z8zHJS2CqvftL8V
cKjvs3gwcdp6Juv9iyQLMq4UtPt3zNldnlqY/LzmMKzsnGgh08nvh+SuP/edERrt
9oN4M/INJOX2uf75TaMXNm+Hse1VNjEjrOZ1znMe2wxVeZCQ5Kka+iXULHI4wli6
MPeiPt43zPuhAT2PNyjDVaQ+aIQVY4d9XvY+R9XziNYMr7d+oSBImxQwcL1hHo+V
h8XBHOqmqDKF148Y0v85SjMf/xtQB+YH/qn+avZ4TVhi2J202+TPLGrh8mZHqT72
7SkfwiUVBc7NaLKlUmCUxBD4hsIRY1z5nS4FajM6p3NWxOdCeHim8wipAuY5mvUM
pI21F/ANeVAeUIMlNywJz0zu2KwWAdzi6eKCgtQRQY6AbXi244NPjTNSxMpSKPF1
ISrQMgAfA9ijbi1DZCT0ByYGk3DnfOHN3rsIrij2vP+DHt6p1iBQ7sAJBYCDZp+9
enLMvUPjRdgQJIvbdhxbiQQkobV6RPzjkDImHGakYo74/Laz92llvWWXnbjlZZQu
6D+n7+D9WXAuZhYjFsUChnI5Odv3aXRDI/vy+642D8tFbozjRACmSG5x4I3Mkh4m
5r1K35hqwoWaiGBluixrhg8ADl/Hjt8UtrH2uvxAVFCdBpgNMSBcMHS0ZsvwU1B9
9JOfcKqD0+uN/JaZ4Vd84TH4pMCYLWMtkuZA08CmYCBnt6NHSZAQrJR68f8SVE4z
KdZgNgrvuMOWhAyLS1Q6+NWOUiPfaYpQArWg8FKhiyC6ddzpPjSlimvEF50aAvKt
vrsCCqms+5HSziwajxugnQEt+2I+3eXQUPzXJICm34DEWa0OsCIe6/tQ3wj3NUo9
g8SU8Ru3CdJO5/H0O5aGqU/xN6RKKHtf2eGJhGdqIWgyIxx/kBMA1PTN6Djg5FE0
CpRmFlDcSdjAT8fwSlbWlmpOVSIAAEaEvVkQHPkBvzc2LnofH/qgjiQewoLWCr02
xlofGZNDT0+rm/4Y2/xIP2yuYa1UOjXbv1D727pGVSq/KumjKx6S5H+CvKVUKr1T
567/JWlSzck7T2uQ73eZuuMFbC6IeEH7X7LmqhKubFxoi72LrD0qh67qi4gs3J5D
Lkgsf0q63yEKPap8pp05+AUfDPYazYAKC/aZ0zdhJGRw/t/O4ohnnA4lgHuah/3/
TniG1hcfu7HomtcHTC76MPdnJ8VCXnESSFeubIz9nOdKtzKKoO62eSNtyVVUoYKF
OV0R7mZu8E539D+DPqC232F3SzyPwo8EnkwK42U8VR/hzEHw6LA5mRff2tEMsX21
llS1jGSpPHLXqiT/WxuawWAi3xxGeMwsvRgTxSPCqiKNnvIXgLgXR/GjRVtt/SoP
0reCdmuwQxQvsjSxp7eu7uboMu5dWlfbBx5cF8FcuFjhTq5OGBRU/c1W33RAeivM
lDwnTqloFEneJU5hmUBLa7+FGzUWxzO7TUQ0iAanXwqWUsAg5WeE1VUEjPoyjwvZ
nLQu4mrSYPpIH5CGtm+eFYEE//kByy2o7wHOeeQ6Mp9nwvW86oQtiyo1fh2n/RFK
0L7xgIEc9QoVp4dNxLX9dctICmR7HKQOBXk47lNtpuwwi+o0KkPDATp7NmBLxH5s
bPTwPP4MIh5Zlp1zEV0jJt7eZpIqcwps26vwFdOVJSfdmyX3YvcgQsJgceZSTtui
QtQjICpoPOkyKmQklw5y/YbBwW3TkJ2dVh5cW5C4p9h9zzA3HVMlhQgZ9tO1PrwY
YlDfWkQuEbCdAvBpVACRlrN84mA1MxBQmieG3PWBcJH30PznkFZtGmPZhQvapqPG
IxNqjK7IKS062qrYwUN58keDOcdsRLsDWR/1spNVHIN5SZeJVKesGj5GdAUwH30k
8e5awNZ2uKXQ6GlWtqNMFPe5BmC4UAzuNgJmBQiGULA7KJyarxNCWC2WaJxl45sI
TvnPA6jkIskrtSDDJiFf/sjW+0rTwFzLZtPV8ryc0zwdv4gU89xeXJDhhtfiYfig
u6Dzyhj0GYvhJXEAxPJwd4gq54sLbxkmBBavdRFFOsk27O36wG0LQJs3GSuDFzkg
AdbuPGrjli0cj9BRWo6E+VkhsQgHLNoj8Gfaj/8wxrni+4uNwK+i6JDjrm/zqptI
SUTwe9z6K9z9RfErNxSws62kAqGIJUUPDYl6/D9dzrgadXPgm/Yqi+QOML+O5HWO
olRT1bZ7ZGa1vNzSlAhHj4ZvZsg2KjvxbcWafSW1dIO0S15J7inNfnLdPqR+++Iu
6et9Rj9TeOIDbnu1orKmMGEMZd1j3j/WAPn48kaSWR7Sj7QAXz3aSt8NiFT2xg/u
evd+jfo5VB9tc4SMfr+ON/nW2dgRh79Fl3yq3FIBCZUhrU5ON4Tdq692j4snCcpi
+ckDZLk5+RXSQBQLn5zWsHedr8zxxTN4NCAt5cxl9v+lVcg1qog3n4EotHO5Nmv1
YGN5CDesKUwuauQ8jhp0SpHryICyMJBmjZmk2FSukNYeyVDRGsk/mFJgVbt7TOhB
cF9z54V8OuuXrucn0baMhIBw+RFYzHcDtYk/08/+25gppVPZ5SgmPTsrdtpGuW5U
u46qenFi8+uU3Umu1UrxBhU9d69Ui8oSigmZkpgMuO79Gleebt3U6Nqss5ZNTxDy
GYRcI5UNg5dlsPtShXgy9iMBM42p/RPfyGI66/v3Y7VjZyukfsfwtfo70YDVunH3
m2as9V0EbxzDlMBxkNsGBHIIC4GXhF+whALPihpAkFTqpLJtCcMSBS6qH6dXunEW
xvS3AEAaNGdxltYs6UTVBO08PAMuK9ZSBUUa3xiqMoZhh7rLZHVGYOrpOhrsbKXZ
Y5wLKmRwPZ/VywpSaFeqHzJLM4aC4/SdsDSMnykmhhgSMdYEy6os8yfHN34QLaap
XscHbe1L1rGdr1yj+/Ncyxeict05Esu9e1sO8uW0ng8CZ0zkqNl0PVbXOuEr37x9
vROgwsNNd5xqCK6DwtjpO4IUBQWw1ZNDMTdbZDTlnzU1CUakii0uNjR4Fmqv2IDO
8giDYQpQcEl9PQqCDrXLCFJfkLhewLJvhcBMYE0dN021U8EH5iVDHmuQ2ZMJ7tfK
4WcMBCqYnrKlek36SarfiVLvyRnqTt0l8HQS+J1jlk1vgYj0qJi1hewewIc/S+9B
b3A5LoqyP9fYtSC6mxmzCbtzo3n+wIM8caPtAW1VmWyLRkEPa3OBw4fjLpLPGtPM
w5Vl/dqrFPzExWgk77TP2Oi+ERk5TSijkHTjoDeIc9EzE3vxLAE6TlcUMX9b/0d1
De7lAgmihVuYt8eBwEOdho4jS4OcmNlsdXXxJhgf0zaPZgde50gP+qjw5pJbteBb
CmbtA3ygkJYvyu779gVro/UVSyTHO0H+zfoPxdODdQEAJ1SpO1BvX/SvDFEg3KTU
rStjQfcJ/j+Z8GKXRrCfUMLta3UuHfC19t4fEYV+dA7MnDIp5oGuKZRsypXpj9x5
s/LSnh3MIEZyeC+OyOdUqVxXLY42vVTT4QHQh7MWKN0jI0AZxOo86kDo9g3/ksxC
X+F4zZaMBUutf1MrMjBqaeoo5OQ19z/xJPFBDtYOjVWxavpFmucyPbn2J7L6UuUh
Jhazq2D7ZtcQ0nZvGuNEkC7QS6BCbk9cRiGRrdSY/SkvdUQ5j7oK599Xr0Wt7mUz
EXU28UK01tGkWmym9n8/p9Te61Qms4Ao0DEcLP0Py8YYd9OkvIm99t10F3AGttpY
/AFNZTDGyOAO7v/KB8mmdpLDiF4G55cdVA5gdrq2su1FzrummR9qh/r40UgxyFsf
Iqxn28GkYz+pub60AXpD6bSKYRABNX1FGSWu0tY4JD4F6TBlsi2r4WRN0wB903zA
jnbmiNtBAuz4vVG4g+0UGVl5X5eNrgAw2qT5rK59N4d9RwVLeZNef257X1kJQwvA
Iz3Z8MJP/pf6AvLRVyGhf3RGxKlv//4/XIKsXwdBpEh6Q5iQbZ78r9q1ZVnmO364
ucz8kTNhgpZ+ILE3rcsIPkekZeyMsOjga3woVxNZzHYnGqFIZ2o1tzj9G55PE5RW
rSffEJm48WOkPO/TwZoKjXN2wIfhw1itGc4ocaViRw6Tgy8yb0fwXAuk1Gi5eTeR
sI5KK/FwDnXejV3yp12t6H/nr61EA70BhI1PmfXK/t6UkoY1bX6af34FXAuggXhg
8dlgiSIpUYcXU8jTDIAe1bDHq92+EwszgWu/HT2BF1JIf2iDrYWCJO7NJRS1LZ++
f96Ne1iNLSyLHm8ePWhdihIQd/awln9BrzisrFuLn2ZTt20PvvLO83x6e3uqbmsC
MLcOtXBwi/+LQkHszGLv/nlpslUKaTX/ygoNGaBzInBe+wtIlTJ6LOQ9adF1NWMC
7Ii23HCpqlvW7jQoqQ/eH1RcdRIzU0YS/lBoE4z314Eqx8fzqWbp0Mb0/TNn7VMd
Nxz/Dgl7XF3m14er3Z7DNe8quGRnqiMFcJ1mjlRLenFA5d7lFME6J0tvx/6MCOCq
DC4aKv7cWqGAYGMUsRWBWutlWUXiWlw/Y89Ncx+6hhVcV3BCrEaM8mOwgjjsEB4c
JKRmdLmJz0JAi8rHeJF0RKfBSYZHXVDjSo4/oLaKFggH6DA4ZLii/5v9Bn1p4Kxf
86bI/803psebAMKLfvb3v1PpJU0zGGF2wUBikX5ZRymlkinWlYRxzKYGh5cUmxmJ
XdMyA5wynu5LoBavY+Tcw3Rw8IXu7ALCJlCZTAGDVsuZfuFkb6QEVY+Zpb1belLV
KtN2xEvg6eajGUJDqf0gn0focqt28gsSGPP5o8Ixam1Cytbih+0zs3SgdLELIUBc
3u5U1jmkB4D0HEpRnOSQWSbCCi+/VwOnPaRxfPHn80z09fc0Hr0OzDrB2x2vz7ti
zr2MlHRl/itTP30XpqyIwJ+0yvAo9EHjTJjDfVTNDE+Wkh4MS4lQ69ls/pyn0YYZ
nbfTgJ4ihQHS7OOZfj5dZmP9FyniCQ0K5g+JXHHOjbJwCbfkz1J4lENTVj0FL1S7
xGmpkvAR+DeOTFlqJ1Ucz5v6Cg8pgUX5Q6meeA23hxJAdZycCvl52aty9p3xcL0E
adXsO0NJvPxPxxMKp1CyHuglqfBcix0K7Xs5TVT+B7oCDDmo5biEo8FuxsZ3g49v
bnWCwXrdvJsCZsg72nSp2zCidzE6x8RWOXOeSo9u7L2/0VdRHbjKd7hUSwvc6v4F
7vJlv8zHwiaRdrnSkankBsaQL6jgxdLVTy8IGKiuY8QBaTX4YlkKQZ7UGnCwsgeo
8Xe0HdVW8D/eKeXkUXQG0M6ofY40Sl4c5ZmVYAOKvjMA7SurGhVtRzquMTiEGZY0
mEraXxS0LLs65pW/bBnBLouT83f+/tHWshsZ1DJuBfgJ8dq+KOmDQ51t9Mxoh5YJ
KfAceUmv0wPl/lOdSR0U4SpthcjmuoP+9M22zqC1RoEQSKJzPUKx+VV+i3ND99p7
vFEqvO9y9GS7oyiA7NFbFpT6dbIp77rCoWtibmFG+6sje9u5PgGLdoQLwGdUzgN8
KTdLrmD0h7d3ZMoJG/srWHondxNSsm30PJ63JIOJKBZvzH2IqYYmOacHLf9XIDo0
1BpYFmgSIU2JMme8MN7gJQvNoKV+YKoCiAJ8L0+9LOrm39p2pUdcSFDJyL3hGsDm
sZOqH1erQujHXAn6WB6+F3CtlMpshJLPuB5AbUDqhFIw6x6Fp4i895aZkPqw1Ihv
wAQVnFTI5E/A5+jx+110GOpK0r7MJ0Zazsid8KoZlzMFvHZgEl6pAOHfrxVHfoBg
Ny18khyOM63uDTuGrbTh65TrVi9+Mwr6oyT7EcBiFFbbRDdifEgpBLxWRC4sQ6Cx
4/VRXPvXhliftuEQ+l+KUl8GJkD2pi92YmvB50DhVkoFcmrVVOr2i4L9i8UycGa/
b6GkpPRw2zrsmYTJSXXtWdqTtmzs6donWQO9KnMSBIM4mJtdXb/1vM3b6YCHRLRu
SvS4SSM8IFdruKSc0MYfa+aI4bCRdgtSy4dUZjusTNzZPNmz0A36YvdqabgkrVKu
83wWZ84hlrU4kh3cgiq0kY6WrZYnxtPMb1dQUSnL48ly6Me7X3aTOoLV4FcjIjX8
NNpQPH93s9lVSqFy5RYfoy064rFn5rcbkL6LQspUfkbINo+o+WCypzBc4t5qaujh
bXp2nYskBBZubXNVe70zs5SOXgFrYxxVmdGmEH8O6VY6aBfNR8RIx7w7BZnVI/Ze
6rXSgqxmC0LOxdR18iwQiewAXWEneM+5Zq4vq1cCHh/QaZ6QRKGsynS2kSqM/pjj
bKleoRXmDj+tN5VSeqOwJ3HdQ6iPu5pBBxdX5++mmTfgyhwyc9cOUpxFfkj+22QF
I6avuPQdsaU1onUxrlcQgo1jlYS8PSR6K3pZngG69XgJ1bgs4L5FKqDX3je1hFCr
6+od0WRQIBOZziC9hS7qjkGVHNQujsVPnlfDMZQJtui75LMkdxMSuhsX0I61e8Xo
JusaCpGeEL6LvBAw+/VgiXhR5boTpDaHykf4HzXGXzURIJgo/cSOENbBsVbdNRhH
KtqPeQvRmYZlpW+m0/8QiijDZkVPXEafSOjE5cks4F+MnYiTgSlpw6jXoHmEy/Do
0dWEsNEdTgLlO9lbUraq3uFjoe0mQmiRLm8goKGu1ypta1F5SCFyZCfBo/I0HVeS
N2JJe+wJUVVVJPlDcPXLZzm+2v7jr9mwMNJwSZZrN2YLbkmM/odaPAPK8y7itVOG
o3xZ+txEtYxwy8pgIsu+//8AtfnU5wvYa0asDrNwG5fi+cMwcL7Mbas/zqOH250T
sd8fPGF34NdAlvqkpEtSbwkaatwCu+2OASGUXtgF8+BqXz2V4XJ0B0rhpIZ2QMAz
SoxjSGE3KL0ZqR2mRJrCwJrJmexdbzEpLeDrJ3GUAernupWKpny4DRT4HC22TmUd
7/eaIDdhhswVOMA4Pgq6Kai4aWrV47KtrWsR8CksZD4rWnRHVp8WUdeCNt5L5qFa
8q4HkazOYYUguZc4tXY1bWM9hbj4JsLWMbs7IppEr/O6j7ZjR+tsePKX6Q7owuWk
Y0RZdAOarCFh1KSbeqmf/lFyiuDPGoGDyjHLFKLiz/Kv3TBikZgzG3JarVcfc4GB
LesEaTUD+7c8JMdPUia9wjenTz/PSbD5sz5Uo+cm5o9GX4DwjFGFgmPawT9kVniq
hbHsCph8KJlqwuHkhaaMP54004WNtfdrFriFHsrCgn6ZEioMyUvY43mTETmJVxAV
sqlu4CW0Z05xayU6n1oiWMQ21kBpvAaVgujhXmwlgKHrnNu+RyGwEBo5WM1GMcGJ
H/WWZmXQklLssa5/WJBmLefiUOnqFfAqSgAjH3hS7bCW52/yDJCWXVLKhaRMKUC9
Y7+iEgLbJPecmBtD2IKp70jcpHW90qQLKeTf2YydbeNbTCLER+ZrGZtEbFtFz9gk
wWYp5D+/V4Vl3yL9LEPV/xD65+pERDyOgsyhDbrVSWsW6sLxYyfASLdeiYRVvfN4
KonijO9Te1p/Sw4JJg4Bmjsz+oZGFI0+YvDSmgCSEf50EYaQdiU9lA38YzOGMvLs
Lkxmx9Z6r0bsZWKNn4eIR5VS4/WKShNuF8US8hi0QPGFSM9EXuYVsPRgRaP6qdDl
9pbrIqe3/NBZFxgA0GGZoF6yIce84qlBcH9U60zBWkNaYlKg8sQ3icgbWtABwoKN
igCVkeED8tBDG2O8M228zox8TNAZSqKcWILUgDlAeaHYdOGW2N0NmaBir2g2PC4x
VGb39vuMBVbXKEekg6F9bz7hGg+c3woPihphNNf0qVfZRtaPDL0e0nekiC+md737
MnmfW8Hu28mb5hL2T+u61W5VLWR/wLom5KzeAjlHef+PVCn5hOulw+8zAU1PF+Nr
/HUWGJaZE7GJ8Oj2usfJ92y7LTFRaDy6mO5Nl4wRWiCeudndFv6pd9MuaQ8LITnE
00zOLDHxUUKY0t47rJ9FD9q3vAHS3YjMd/haHBCSnc93J9zHHc5EBan6qhbfucqP
MmVtw5kbUHMGldNim0tlSIaIH25lVYzt6dlYsHoA49ozhChmh8u8NQGfdCbGWISJ
zfu3p13PoMg8nSgG7Yhufie4fj+c2K/+/3uIn+YTaY4apjAQyo1OKB8AfamxF3qP
k2GgOHgWR5BBQW1vZZM/rszHxTYRtBte+rFfutTDG1cXDz8l2IfoZoOP2ROeX6uQ
55ycK80s0Middw0NeyFpsa4BU2rUM917ckUoDj1ZrdiFT88B6vTXG1YKF4hIrlBb
A8csn9m7O+anioSrdUlqLLBdtgYrkPzUaeIKLwX/SQeL9DENUSJ20NMhcqgNRPs+
hi46+vFU9kQw5LSnBNyDCgU3XKeu9sR7CwEJLqYaTb9gBg/8w73kHisFmEqNVR4J
sXCU3kzdR7L4EvK72zald8hjGQNXE86Sio1UC/EYmR4EZdCQbfwwLHeT1rkkRWsr
oqsb95vEUsQX0TUg6VGLE7PwHf3ZyghD+CDxtTFTSlw4eBUfMiq5aZiD7nOazYBG
ZncLl8kndph418BPxiMrQZN1vwnaacAGdyPEaKTwe3IVOHrgFA3GedrFZJg8MM15
wpTQt+eM1nYIqYkCMXncJ2MrGdLe17OD6Oeq2LQ41weUNMf2Xxk5kenEMSe8wfLo
PTXByyUy6I3rJ9WUp2Z5sSGm9nmOKS+jg9Kaiad7yICE09lxOiZmIrMopv8bDNPk
qNqnqjhSupghGKkks/KD6iZHJ2si4eICwfIT0p1+8cU+tBjcwmMjYtEZf+kyfCak
xpNli8T9rU6shsMg8Hz24YfZXl2+jaGK8gMGG8TLDJ7VSVLf/DUKTwkEJ6TFUedC
0kqvL/5wn+7RLQVyCsb2rXbLsoZe8W2Vvk54iuou50S7+9yVdCtsyK9QHVK+6ylW
xdFwoilqr2v00//3aOgnOTmymuiFni9n4EZscz32/BZnF2TLg02aqXttgVhHawUV
gTo6kKmrHjuvK/gyQuQbhAMKxgoGNJa3pHTT1TkRFJuUggcW4cGVN00mTphCy0Lo
QEmy7xK8sByY5ix0ujIRHjNca64GojjCzlkLsZDENOoXbmHPLCgV4EtLz/ac+XAF
n2LCRkUqKaR8SP3vRdS/mTwW8ULABjVf6VsjHZGNYyGGjlGI50Ph7AZ7IZveDVaR
BhZa1NR+ltc3lm9hStXZUxoaGzKuI6+3NiMDcRwXxORa/dIVg1Zsh3EfmZJHwyUj
Xje7fVl1UHSKCw7usxZCLIEKn4T6WVIBkulMfVnGJunucmhXLK9TIcnl02zBZs1c
Oan09uWheaMScxQGUtR8JI0lm2U7h309nkafXC2Nm4Oc/Bh+csVKDoGcpzdV6eKE
5XEPpom+sJjr+3Jm6KG8y/+oFYyMnbG6oY0VUFGaY+eMN9THKGIylgdJWpV2WDO3
MZWUhxJSx65G8XI8GY9cnlYUUJXv1Xdj2/dFx1/4bkJ61rmHxsQ7lJjbSaqlC2OX
g4u6hbXFkPj1VKmQ+9UE3zilE6p7cMmdZu3+26Ojf/oXAO8qsUvy9ku2vs0BaCII
nerbkfJrBblNmimQeQbFSOfgF0v9ygXS7gVqS2iYHsH1wk/gCgFV6eMFk8yjmt2x
n3NwyjBSMEDmm1cFCsZITY4GVPqmVvld7vWO5IxwYe95Ce6fr2OQu0VmqAfcMrNR
k9sreTwra60qwlDTmcTQUj6IorAKv4wZBKH6ioWNmQc7+jpteK/OsOto3/eorhnD
8Q2sIgWV2Lw8Qt0dR6o49YOAPYRNp++Y0lJN4+Qn66ShD+KjbIM6jwcBX5njDdKq
m/B+oS+f1aUJkxxF0QoUDirGzaV7ysiPgiCow33p/9DM54O5R64SESfXsT4SB1eE
Wg+o9qwf6uYQMVEFkHeKmwsSRiWp51GGDjVoJLEsRqcVcVIFpof4EMMLUujMPQ9R
tSG4ecv9Ad/DMDXF1IoQuXS5R4vq/tDeXuiLu+pUCpltQj18DK1FHGtXpAv0aGsZ
KK3ZUqKD0nF3hWrv+SmoxJy0qF7Iu2Fl4UOWR/Z/3jtfN7HNpP6sCU+fgvqJ7czn
SPds0Dl0msHmblQuZXrtELizLB5kXmrN4jQOGA52gC0zdN0IvzHQI5PvPR06dtHt
ExZ9VgMCtNQVf/OI2R8a1gQHk1TTCqe1kTOgG3iPIK7oHBwYukeFJIO78HRQdM0n
ptLG77MytfhJ5y8n8gyiEuxXONyvinm3o1VNhGOlpbkxtvJRtNuH5p0V/61bbX6w
3EzF3RHJK8jnqwbI9UapAe3zwdz300Qbecf5AS6mo0CpePkGHlhkmMPGygICfK6S
Nd/QYWRlo+4nSGLNZdNKiDMArz3GJMRR0SK3aP1d0l+inAw1MKHAbQtg3RvA6FhL
J/62ppOVlJERhn43j+Ew8XBx7QSARHYCY+397z8ugf/ZGfiO625kbG3URZIUAchy
Q8Mn5GkoHxmZOTaatQO8WE9v8NKKSPeAije21fb3EnaaXYol2c/NwSDlXX8TFPBE
3jl6OtLx3MvrH1DPIml4u2clmJc4lSVZ1G9/xt+RNIrU9XTFF2i/N6KkDzsOLfk1
d9+Y+sHNBNSpdm+Uok7XN+HAtmnNanOcTko61pi7Ti1mSQmGBi+6zPZ7aCPqN7ec
euKAfffpesZUVJ+Sc31TiV+DgiKV8cCcCyTUWC8fE+jX15R/cU8MO/oj/M5MSShH
8xUo7dJcZETJOBMdXBLCWDIAzBL8HS3fcIM0Cv6Dsm1V7xwmlfJ4h2luH6OkQkAt
FJFGxRjEqs11uAxXzSglrTEBDUGvUl3Wo7DALjqP4esuFha5jKB5XM25C0urSUZa
LUb3hIcM+m+YVvNTeJXlMIIpbt5nRMt3oaDClyq2jZLt2QIfy9Y5dPCfDK+49V6s
IxFtroEHpOEQwM0BI+EOL2mp0npDh8RsYLPv/7bfbjRxVisTW8vuHhiwvPkIgSgN
6jg+YO7PMyHZa10w5QUoU4lUCE4JrciKsoI0KYL3e1lqC2heBjsTgo61MTKXMe5H
zcyAYE+M5TlVcbY+/QKvIMyT6xOQVCfN6xs9EdCOaVuT6mzu80esZzyECi/p4W5p
KyHo+6kD52Pg3ehBuoioTTFarmiqcQqlX/HLy73aoCthYHcTR+B5KHfT5CdPrpGE
YNImObQ2yvY7MGdPInbwYH+G9ZEb4cjvl0z5IEyGG1hXBxkzl+UV3gPLkrX/o8gJ
rhbqtfh7B7sfMt+BAmBQF08gjbNqIqnCR/+Caunt7TdaI9ToA64IKuwSOTKMN0UP
U9xE5h7HbOVPDDHjrlJ/JppZB4I5tRfsLB5ofA9cMetY1XWFfmjQ4Ixzr7L2ZwU3
VRKeL2nt8J4MkK+uAh1hV1zuyWb93V7vqYoch6iKcorkPVKcjDXBAplTaQgzDnMH
pJtFhaPdwD1WWPJMDtfanYvpIuNqScUSGAQ2D9CQWpufyNumgDPnIZZ8cJE3H9P3
bDB0DiMQH+rv8bB3diIXAk79S4W/1rsw3IuPN7M3fhsBKXjjo8LD6alTKwIs9vQz
WPKO+bHCB775NRPQ0g163EOQ/0eDS49vx1nKdHngEswxZaV4hCPt0CVpWHeByF6I
oMR/T5K8pgkp39DBfzRNfZ2aO3j+eP+KfxeJVI++1IHqjDGfmtJcHscVXftLrAiH
sBmkszRLzHPhlpWUb6WuuFVPLWwXddpAeVJxxlhVIKq9jzgbXv3YUCZkySVpZE/U
8gJ1z2ZMVmDr9tvOijrXtPv7SIt/NeaQsCXooEH4pamF/HF6Ld6ONgU+GjvEScWE
GygZZBWB0aBIGNI0JrXB9fiiMHdh/mG8B7JQNkSX4b2XdH93EFdiY4GkI9tE6/aZ
xhY3bEiu99jozECpWKpcLbl95E/OdMX8m/Vor4+tLjCM84GYbD66cJiCf8b/Fmk7
qCNcJ7V5aUY/a0dr+NU2omKUBjvmOy8DOH4Knn7HVLMh9uVFM2tSvjTr9P6Ftg52
cS6YDwMTi4bkzPDT8gKsWsnFAlMPyJyzr9WVO1vMN1y9QpIFbBBuWmhVpag+5wmw
pEto4NtUJGYR8lNzmHXIlzbTH9C6WDG6pr96etM4Fc/T2WlySyMD1uL8nQqGzMpV
423DrxCsq6IsZGWaBHBXhy2ddDThFNLRHZ1RlxYUQjex+ZsKj+OlQiH+aJEyZjmC
DKvLcG+/83H3XI4tZ4Tkbroi8QAMRyfFNtU41mv3dsMUSkZ+QM/k64wa4X6dFsH8
bToz5SOjAgeZ0UJuzXPJJeT97M/KEEtfzk3YTOMK0oOBPeVUgaknumUno9qgvCsl
6uBI/MrbbvFuvfe9Gcd1x4aef4uFIOxjVfZNMZeKTzvyfQz9yO0Dls9kU6S8hNzw
KmdjkFSyw5ZAzqYA4AXD7dFijufm6y7Bum4Kqk02A2/HWsZb26kZ+tQHLePOZTjS
j6IzNujK0iibN8G0ggE0PvGWWzt9xLtNwm/jGY9PJIBMa7JQQ0+15glFhd5q3NQs
hPTwNQarB/nZB0W2NKYtt0aonPQmA+m6RNsKVsh6MQfCe6OON0VcDs/R8DsULqga
FxbTbfnQkmWjr+R2g/bJK4dCmQmyAsPtlS8vklhPKEDhS1Gb7X3TxhXRda2EKHIh
axbTVfjiJH9tKOxJN4Pmte6QrKl/Bcde5qUKx9WtDwA022kxUMWeZM59gics84CI
R9PPy297kpF5oz4NULwl5NEvpeqiwBbnx/u3Y6auVgILK047pZwNR2Guw13v/bab
NgOE0Lgg67sOvzF76W4MbwZfy6cWI6fEGsEGgdGIuIIBmDAPaSxHh3rySL5o5KJ/
mzaIBWwrcOlp31pLV+XwiwB90rT3cC8gxKRCpppY0WL8MQa3d7huFR8eILSwjcht
KAjnB+srqsE1Aw5ok1oHFZz7gHPg9F2bUH/SfsiOkwA0yovx4VgG3er+MR0KMJzi
CysN4OSs859vZwWFzkXiBw4VafeOKIvMxQo3yXESyRAP08C7Yqur5rxTbHgIqzGX
KIUs/DYYSwxNm3cSW3dPG+S/MO2sgR18xXyWVNQP//Q=
`protect end_protected
