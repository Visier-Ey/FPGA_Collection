��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���d�v����0�i�=\��A��?��� (��1_B�f�	�Ѻ+|n��y��Q4�]�aY�����*2�y%����>��������K������ �
�D��z�z��C�y�B����
_�U��hkF<�~x�ܕ�c�y�L�-��T��{�-�md�}��M[�xЎ�Y�^�JS�ڣ�mYlY�����n��B�}@�u�н�~�s������r��FA�%E�����������DJ
?�G�%�	��0��O�N�O��0�*������T �ڽWP/��#��uD��ŧ�ɒ��x�?����3�����gѾz*�O�!�$��T���������x���ݭ��~)F��Yh4�0]+��5m� �f̵���CT�y�'�1,p�?0,V�N �|j��XP�����Pk}K�%�MK􁸺�mY��N�|,}a\uZ�>�ԝ��]���ǯl8�[�~ce��H�
xK����1���J]���*l$�	�gDИ����=��u��d�]�7��&���9�^F;War�mX��1;[)lH�����{�/`?�ޅ[�SS��SGM��3�gu���G�+�/�>zݏ��,*+9�E��L���KO� �w�-���3�w�n��m�O~5�/c̥4�!�JWu�����ɭ�B��j!-�GG��bo�zf�gO��$�PK,6X&� n�d�������<���4�==t�ǿ�ӸR^����?^ A7���U���죎`teeQ[�`�V���t7��FZ�oJ�I��6%I�E�2I�[��L>u@R�����ڴ��.е0o��k�l?yF=����}����RO fu{���MBP��E�g�����J�Ȱ��2S�ֿ�y����tH��IV�,X���'s"�у*��$��HUײR��pgm�23x���X��O��/�������/�&�S��S@KIU�E��n\u1�i>���.�;�|/���" ���"��ۑ���=�I��N��4��*]�ܱ�(� �'| ���FLd�l�Ԁ��Gׂ( ��z[��#���ވ+��ܹ�U���\�!C>'�Y�"�/�񼀴:P���N��$�~�COAVH����+�譾2Y�����`^2�F�6G�t1\����K���e&�2I��2��� Q�\&�H��
���ҾcH�7G�!=y��	�	Z�7��� ǫ�zlD�9���'���)}�H���Lr}�q��X��T�b�S�i��EoGC"���U��M�8LQ�o�[��\�aF���@�xUs�%L��Տ1ۜ���HU��s�(l�䥧�'΄�'q� 
��[x[�\WW���?�P��#�1d��4��FՂ[��!�\�V&����2���ZfE���_�sK�~|Q��Ws�6#�@���4��	U��+	�t���%~�%��Œ���eG�Vch�,��l�C��QYx������g �(k�G̕�Tޜȷ��<$��)rE7���J���ʜvk#ZL��La��9d*����Q�&FS0���$E��`�0[��B�fPx4j?��x\0�<���5��)d�n�x;k��)��ܽs�	/*
ý��T���U��F�j���H]�L�}F��5���CS�c]��B�п4���=rX�sxe�4��{�86"�����q
.N�4�Uݷ��WD�ҏ�%�"\������lK�U��)+en"�V��%̷��/���<� ���D�� �너��!�gs��B'~�H�Rk�Ǧ��hxuH�ڋ|���g�aQ��00Ծ#�k����\���^��)*�����n��@a�����q7��+�#��B ~�9+VFѣ��}�Sc���Qz�j����Y�5��9@�ُ��\8��1j`>���gƴ��o�ʧw�.�{�����o Stiy�]6���D �jr|=�Se�g���� �ګu.D)�ڸ[4z���ژG�t��T$3��VX�$�0�Q�*!\eb��dS8A������e
Q_������>.���<!�O��%��R�-��T��N�x�gT�'s=�w@I���T�x�Ri�p�7�P�6��+��sE�QC�٨��ډ���T�0����#]�.ЏT����\��=z��SO���ug־q+���^����N�tWWf�Ŝt�P�L'�2#�ţ"G�aP�+�(�q�÷�q�'=%2/u�?��9�}R�>͵��/��:Ā� �I�#^m��19=��u��^p��P��bn�~�#�˘�y͸��/]+�z��œ�f�����aӈ+D�t #\��INә������1�H�K�0e!̘ŏn�Ӓ���ѧ����t�%�d�X> Tu��w���d�#�^og��In{A��u����@1�>�KQz {��B=�v�$q?svd� h�[v���!-2!�g�X�~�D�<V9*M��~3�Nx����׽�I��)��Ĺ�fv�+o� ���� X����Z��p�
HJ�!�c=a��=��ѯ��կr��voG�j�/6�j�ih5�A�.N�ڗ�%����+Z�<w<K��N��n�w�ğ`��.��-F�+v��Hj�Hw�F����]G���ʹ�,��=�
��`k}J�ny?�Y�n�������bÿH��+y杀 ��rL�΁H�d�*Ɓ��8u��ZER���^�@�%�>aS���&?�P8	��ڷT���%��b��C-3�l?��M�=���#���8f���\
�4��,���<0jkS��>��������WV��02�2�lMB�� �Vb�*���T��"y�Pr�S����m���h $�*A�-�xg�b~&��Wԑ��Q��"�ǧq�=��2UL��<k�DGe����G"1��	���O�t%u)2�T��|Ʒ�X��JS�@�w��p\u�,7~���F�U�7�<(+�'5��Ocqhk�-�Р��Oн3f2(��>�.��{��������-mD\qSA�Ns�7@���&��zX� |�g�[  q��bqn݌��HU%��\����.;s��#����YO��`A-5���Ȧ���!3�r�.J�Ln�>X�s��߆#���^���_���|�d\2�d����2�N�d�cs�z&ɀ��#�q�;�@0���5�\�5�(t�w������� �Jl�YC���"��pb��#�Uc8�#{�����v���X;l&���t��Da0:�ths�d&yS���^#�Hc��	%�ƌ��M�u諔���Avn����`�-s��I��R"0#�VZmzt�77�@����y5$�ca�"f������qV�}�[҉I�?J�-�P��e꤭�}N�����iD������	4�Ӷ� �Ч!MB�|TZYW�� w�44�O24[�{Au�5��T�B=0M=&����I�˃�?w��6�)���o�#3�^�-�h����؏�Iuwvx�5���%*�&I���Ģ�'���2�!�TN��u�ٽ��/;xA�e>��5�d.d��Q�$oV��P�6��t��&H�#ͧ��Rץ�P}����bBd⺊)m.�9hl�=�-r��F�}%>O|�PV�y B)B��ӻv`�,m�����%u�c�xS�"�zpZR��oQ��*mP�n�i���7@�8;�PA^�r����������,�-'�vLL@c9���i�a%~�2u�j�����W���������+��5 J�^�S1�Ӭ:�82���� �t�Ю}��9k^�@ZB���	��Do��|��V��=��DZQ�V���1߫%JLp�XW-��	�RLt�O�L�c'�[����]i�wg�����}L�A  �ᓬX: �U�Bm"�/�E��fFp�M���ޢt�c!��g����l��t��(d?�NG���M�lC�s�����m��o��5!]�~썁�]�-n�u
�L�C����c�i&��v��`Dʉ�TH��%�Y�g�3 ��O��,�Z��Ϗ�?�n��O��F�DG#��'E�0]��]߲nR�g��D�j& x �P�y��t����{-�E\�3�W]F�����q���Zq�կm�n����@ ��m�/����~[�DQޅ�M;�p���vIx4l�L@��9E�Q����6VB�Q��=�_�� ��Ur����슝�v�{���4J��ބ��C����Y3�`����e���j�
g'��je�@�%��%1���	�5X���E°�6w?���!�'n!���h�\d`_����} P�����A����ʡ��wZ՞�ŁM����o;��{:y=��*P�2T�'H鼩p2V��	�N{�MM{�T�S����.�H����3cb8��e@]����m^�"I��Nzw5�
Nb�2�17&��g��]�HoK8���f� ��(���Z��Kzgg��B�R���L��~��e���TJ��d �tU�/a@z&p�Ze��ظ���}�j:�05-��������a<�S �u��W�8q�%��a���4���:6�U,��F�-���w��"�߲3m�����C��ٵ�t��dߔ�>\h���LG¯�G�jX5Aj�cR^��!0�0��}��3��S[>��k���,��`��S�B��,M #��)�s���"���o]�d~�v(�A�eoY�9OۃN��(pj�n�[hE�S�-���n�fgr�b�)�Z2�pv���#�3ƨ	e�w���i�g�y�I(A��D��ߴ7HVӬ�8J��"�Ӂ�DkaN.����Mc��^A��$y����ax���@�͵���^�c��Xc���s��н=��F�|��:�>{�d}t�n�Âh�L����J:�wM�t�������$ɮ��>�K�_���O����a���>4z������%�kp��1��^g��u����@��<�l��z/j���2f���,�)!w5{�)eP�Z+��Cî�].*�0��mp���X�^s���q��K�:o�������+�-�#	 �;$��gۇE�u������3-�������e��1�/�s��1��o"3���׆˖��d����hz�*1�$�V�T%����~�`��AL��"{�ؖR1��
�oư����� ��1Q�1hBr0�u���]������Eg�ŵĪ��4v�~ٙ���v?��K�<Z��`�(�Q�"Kh���F� ��Q��T�c���SB_���9!������֊��w��`�� ?{��:�$oXE�{����]�"w���L-?�V�k�1���zo������'\�clx-���\���4*�kH��W����&V��kbҧh"[xw`ʭ���֕�;ܝ��)�w�k줁��p,?�ػBL0�V�a�<���z>2���ɡ��̔G�X~�1r<��,Β�����嫳z7����uD�Hˋ[�0VH0-�p�p��|Y�=)�d�E���5Z\n�]��i����,�8���1g���I1���?�~$�DKXA�JbI���g�$_akl#����;̽��|����ϒ�h\��D�~Ș~7�ʌ��ܥW�pB��܇�����+�bI�9A^�ɑ���w[k(�]��_�s����C�g�XP�ߏ����Ĺ���qH-�����*��!����=�\=l=�0+��iH_�0Ҡ� h�@��)��/�C٤��b29豯�W�4,�W+%=A�ZϺ~��\n���yಆ"��6�8�y`�7�XQTm11�q����	��g���ҟ� ǲ;�(�*��'��,Q����r5�
X;G�c��6���\�����$��
�n^�Q��P�`~�g�Vt�J�M��f�ޫż)�s�_K-C:�tGP��켔1.��<t~X]����Ċ� �W��w�d�'G���# b;�K	��ۄjZN/T}�b�8 6�����Hl�}�x�8d2�%������Y�Fcᚣ��f�HZr��I�Q|
I4 $j%���U'�u�1��r�zP��B>'�5{��U>�=��1��4A�M�%����jǿ�%�܂UK[Oа�����ɚ>�Pe�Ԃ�\5C+Ĩ��Fѡ3w�!�e�#zi	r���i]WwU�߯���_�	���I6�}��gl���d��B�A�Ϣ�B�5Y���
 �^�Z;ǊQ�b�P��z�s{H���=����c>-׶��6z��4:Q��o��O�<j���"��UM2�@8�}D��@W��E� ��FęcF�Na��bZu�3J���5@+YG���H2{��>6�Vn�B����]�1ru��P����v�N{p�x�V�L�)F���ۙi)F�A��~[[��IQh�8�N����N��L)n	K�R�v�=c�/�`:C��'U#�ϡj"kt|:�h���a�^?�n_	�-�V)˄��%O�NG��������Y\���K���%�Yj-�*X7�45��ǳQ`�Nc���	��}���#��}���r� U,��5����+�.�K��n~L�Ҭə�ZTʿ� �x=W֜��8c�Aŷz���\���(Twøe��Wv��Z�~E4�2R�/�G�d<>�#���}(���.c��/5!>P��S^�[�p� QpЯ�%�>���+\`�9�	p�E�e�LU�� Ϸ�0�x��{�.6xp��c��ި��;�7�Ta�.�Z�7 �.W�O� V���B������[?�3���;�鿕��H�B���e̷�kӛ��� �'9�Xsԡ��p��>u�t,h@��t��j�|[�j��,�᳊ z�k�J>O:R�*�����6�Cj�[b���_�-)z��֪����fʕ2'����R��V�%u�KmrE�MJz�wh��^�@%�U�.d��Y�Lq�/��W~$O?��^��1,��^D�T`B9�	�R(&<6�&q@�_��d2�9��^�L�1MA��v��A��ؤM`��G-D^�2��4pA�6|�
�Q-�-C�a���G.�)�Ԟ�`3�9%4�F��Bt�|'RK��t��iҀ��OLh�F��_�"*e��|�����r��Z�?#�UU�a�� ��M��"�`ŏ�"�O@Y=����O1�'���d��E���T�sG��:(~Ev�yޡ�~�D4��((u�M�xg�x��ny��ǟ�ʰ���u@�!�`(�B���^���0����3F�Ĝ�wvۡt)�a�c戯��IVk�'���f�(��@��"�+Ě>�&ȥ�"F���(�K��@�!�~vY��X�>��D�b>?}�����#G���!6Z�sl��{[�[_���rggXS>[��"��=��)�Z�j7�������~&-�r'll9%�(v��s��":v-7��u�nEA���	��tH~q-��sT\w���o�����B�"�0"')n}��ʮSKj㽊&No�Ԩ�3֨���h�����r��^��h/��=�:kL���b���m<�L�B�nđ߾f������Ʋ��@I:��6h�@e�uU�cC��U� Mr�K�Q�k�~fE��ݹ�V��4�����y,�����1�����6��7�""����"�H��� ���g��҇P�S@��B%�kF�s��j�)O���_�j��I��|B� ���<�z{��Eky�-�#X�
 ��.QQ����ڕ���`�TH0"��f@«��K㗆n��*B�Ii޼fT]$X�,qY��/����|TJlZ9�a��b$"�e�!�%4��qǋhzw쀻䆓�_���Բ䚩i����w ������y-q�aϿ�␲�7K���������wV��R^���(�v��N7̀ƼR6*�@JՏ<I='0�++���P]��'�+OQ/`��p]�Z�\�`J��S�V��a#����-�D~(�,�g�i�h ��d �?�63Ʌ��)�E��~r�?r�z�菸`B@�u�%�H?����#��p0=N����J�"�z�%
�/����7���t��9uj�Xy{���=�C��k'I��>ShE"q��y�0e'�Z0��=$go��a��%�r�{��~`)׊���Px:L��M�A#���̠���D͗���w���;H|Z�m@�5ᡃ0/	h���uB,�P����ds&��d'Fҡ����\�B1�S���ո���f�6F�����M �BP�Sf�,h����RJk2���J�)�n�,O�})�:�EAz��e��a" ���VPo<F*��y��3t�\ūA� fX�]�������'���<L8�һ=����x6�Y��/�tC��g<�����'<�dٸ2we��)<2��\��O��}�.Q]��<���v:��nWl�4��a�\K���l��
T�#��˫�QnR|vEl'J\���������N���͒���{��6��+�R2�p��RG��XY$�j���;߹_�J�X�Nl熐4�Z���RWA��eD����/B#��lG�$��̇�����1���S0�٬����~�r��o�#��l��x/k�x���7Vϱ�K�Zeu�)_���Ó�ا�n�~�)�Kb/|u����I��b!�%��-�����5!�'��d��h��%���Â��~f3i�կ��N�� ��٫��Q��,֑�w)�v�>Ԇ\0��$�V�~8��~um���TX<���*ǐ�u"��P붐Ҫ������"�J�Yie``RH#�e6��R�mqԿ��w�\�C[���z: ��2�#Sz�D��n�ɨZ ��k
�c�b(�)k���upͲ���s���Y���M�wC�e���Gk[>y|�K#��=��c$\.���05 ��:v'��v�>��>>�ep���zRkT���n����M�+�{�X��v oTuQ/�63e
/���t��t3���M92\��vxh"n�r�����h�J��˂��a�@7��B�Y#^^,��{}��m�&���]�N��������po�FG%��#9�0)صȿ�Ʒ|����"�*.[~�9$��%�pd���ל0�B��������:��V|]A@�B�kST�l�rm�X�F_�[)p@N�ڪP�%"sì #����v�E[�5=���
�V!�iG���/@u"��cFl���!-=.�A�9In��������5\���,r5Ȱ��T	{!�$�;�!h�Jx�����9J��e|��߬nM��P��������s7�x��H�� ���$P����DO��B��������J��F�1�����F!�����5]j�{����C ���	�ˀ��g��#�"�c�V1��e�d) Ӧ��R�`i� ^}��WB����e@��M*w&�x�o��n.�
�>�=�����!�HSy7ĤT��^�V��H�������*8>����2O��䬜�e~Q����g.��~N�c��n�sU�(�^y�✬�6Ϭ�%�<�*��-�Иg��R�m\Z?�1�&�*&��Vr�]��a5Sa��#'o����M�����	W�U>7�4V�ʂH������̄��~j�x�`�4ɰ.=�>;f$�<o@ٚV�=Z�9�+,KqU1��x�,��F�N��Uyp�,䎴O�wM[Ef�G0L�������pN��̯*�+��đJ\��ZE̱!���B �/�Yl�{�,4X�&j;a�ƊݯqR��'n:e����G�\���q$��{�F:e�����F����`I3�ʌ��' P�+��BR�\�-W��O��`�
�꦳����{Y���E���;��O��f7aE����k�s��i��u��c�Ӏ�� �/D��S��2�V���#�/��d��T2���u-mU��wDJx��
�]�o��/�ϖ��IYu��4�tE��q��i�L?�%�s�Qϥ�m���4���O��7r$w�Y�xw^� 턹�>�Gz��⻓�s�b3}�m�c���Wx���E�)�R���������x���?�N]�
�6���_���UI?�?��#!������p5���#�}����2����Q��!��6V_1g���0� ��a2ϳ�x�?����������)MP��f`�ԫB�u'L����Nb,��8\���|� �=P���=��z��{�RO�,�����~PbH�\f);���%����`����6&�T^�)ٴ�$@]�ѕ��_�Gk����l�����c2,dPe��S5����Җ� r�4�tk�NZW%��!Iq �H�{�r،����d���#�oR��!��1��Ӹa^j%U�x:뗼�+	M����*��+����o	ܠ�/��5�ȕ/;��N�A!�e �U�D>�����b��.\�>�~�&�L{����'w6.�eNɅ:�g�ƅ6�@�G�u�P�Н����y���g͐��ϡ E���;V`�x+��LJ�s�D���q)3{����ʐ����1B��-kd8�����yV霖��TYA�*��uaD4�|��0t�
�Aj�����v]a�ٻ9	�n��I���������)��\��ܚ�{Q���#�zJk������4(��슝�t�0�Ѿ�w��`8�F��Ԝ̆�<Z�j���4�쥯.:[}��}�|L�2�@�0@�W�����������/,<�\�{�6�0�/��'��{$M%�j��O��7��˅�=�� �_}'q1��[��>�(�νꥄ���3�ĎB�Ii��ʺ|kNމnh�^�sS�zz�36)���8����.�r����v�'K���g�{��%���������͗3!LWBtrWցt\=QFS��Ӛ���2l/#9�Rs�ϩhl!�����c���6�.(�/A�3�#T�wAU�-�=�,R�J���xv���:UZ)��;
����x[�3�>�%{+�i��J:��F�Q ����r��",�ʘ$>/��>�Y��P=?�l[�F�X=��'>Q��9��6�����*_�ԀL���е�EAmI����hy�]Ŀ���wmC2�v	tW,���:���Y[Q��	��6R�8<�D���_Q�5�Q�<�-b�^c�
4�"�dq���n���h�d���������&�c��0�����6��T�~��0���G')�0%�GV (�z��W�ߋ�}�Ė}����˲�H!�pS�	�m`�.���&�-��tp�#�ß��du�&ט��)o�;'�	�|��Yڒb����:�&�Yk�ȓF&1��4���2`�o�]����V���f��F�R�q���`�
7�-�7��L�j+���	�C�5���B�q�5�;z`sC������+���cB~��ܮ.��ݠ��m||�����Q�&qĜXJg���n3���p��t���$2Q栙=Mm��K�Y�2H��8A���h�X?
�R�C�t:�����ܮ��qqI|*���h�Z���K�kN�|�,���~��T�(�}za�(�w��:g��Z����I�Bu!ȕx�~'��λrRs 1C/�Ш�+���Jk���̀��)ʴ-��y�)���}��c-R��V���ջ��H�-����[�N��Dw ���`vv������gA*Da .Ŕ&tC?�?Dvγ	����Z�H��eA��i=�I
'�'~,��o�0(�J��`�]ßF/�����( ���jO�c�b0e�R���ۃ:H��k1��z�p>��?e�|���$�\�����&��"���|�d���AS�(��u.�ޏ�׷$�
�9��]��~�װ�}߼�ԛU?��4@��K"�`+pC܀��y=�J�"��}�,�k%��Їt�X9;�C��ߑSeOYc]1.���D3���OH�������g��	
�|?�M0�>9T���$�A����-:r���&	}-`����!
>��DN�����`�x��g%-V��,FKT���b_׈����ţ��}��-��2�gb�W��NA2�>�I~g�'����kYn��`�a*��U��M0CHCe���L3�Az�~r��dTE�̝YP7VT���Mx��cJ����t��Z��������8c��[C��p0���B�:��PX���r��%�;��J.ߤ�Aoa��Puj���0��څ�z������-H�1�)��V\xHä��4�]/�J���Sv������-S�=㩬ghѧ����z�SIS���o⾫݄w"�u����>� ����Pa~�i��Ѭ�4誽�4.��6kW@�B�}&�]JR�]V �
�X��#(�O�C��
��l�/�e��D��3S�s�'���5혫�\MC������ۯԗ���鬢8-�CD�khm0�-g�{=�3J�J<3/ҝ5���L�a6��&���[�A3XәO�#	�φ`]�)�(�l�[�I�.��[ƵzJ`ic�m���Yg�(�\L���j$����9�aJ G����`����\�!�uW���a���))�����)l��l����댙���@�Ñ`D�� ��b�\�x!)f�f��%%\�q���u���1Q�0��Rۂ��jr�)������}h�$E28�A�>����o5�=c�^�ֽ"��� ��|� ���Sv¸'����H/>#�T
a��K`}~�L��������
� a���鰩1V�}��H'ʙ�����)�_W�R��[��������:L�r��WZ?퀛ByO%B9��q����.�)��O���&n�'b#����h`�������s�J�� ϯѕ�!ؾ����f�������T�s����ҵ*�Ҷ��Tim��B1g��Ƈ�x��:H��%l0��+b��TtJ��o��y5�O+�}CaA�- ��8�	?�a0��_��LUf�^�$7�9(ǐ�f=u�A��Ag ���H+Z��W�+� �O �\�T���c��:�_�}W�mI2��9+� ���;[A����}��'L��g�d$�l������;�<��v���������ڪ�D�x(n%��B.��D6쑢�sPH`~.K$�*Au�_�ԅ7���t���<uu���R�ԍI,�J����ux2���"2Gs��6���Gs@�z=/:R�"�_�m�"M��o���[�36:�m�L���<��#�?����m���M�Q*��-��L�e/���F��f0�E�4����ia�.�Lt+�xq�Uk�z��d���U��y�<�b���o�v�����܀�qǎ����*@��,�3eS�"Z�����S[(ISW�8P7y�{��m�q�=��f2��k�=0������>H<u�2%źe@����4����k	����ϴ�^h:d�a��p�SP���awNz&�"�,L�.�Z�ly��|2�!�=6�F��L���fO��͞�}v��:t����%ҦU��ؙ�-�|Զa�[�`���*��Q�PC�yl�\5��_^�e�Lj����-]J�з�9ES��44���[Ϣ�@�lY�s�B�%�e)��[�t�%�WfA .�b/�񝖒UC�);VmE L�%~�`�iZ�d�أ:dׅ����f��yowvOeJ��,�̪�����V�m��l�Y')����b�#��,A�6�2~B%k|����On��y����8���)�F+���� ��_���Ξ��)J/���{Vd�{��bX=ԇc���D��e�e��=��e"�c��,j�5�5"�lc���1�|,��N�-�YJ��ք$�o�CIp=_vZQ,�薶�θ6gQ��pI�D�����=p�blp���h��'oA5�k29�Y����v֓6,b�)�����P����E$�Ѕ�wY��O�C.q��1�r|>�Xʩ_4O�$�zݶd!}�͘1�k!��6��W��{��d��P�k���9ǋ�S�;���V_� ��M�r��3�,+OK�.ҟx��z�x:tIA�v����s- c�����W_�US>�����d��(�K��-"Q��ߥx�Sx���K7��
�N{��n]�D��bFp�$����۷�cW �/��Z����t���@�P"'�?(< �ӵ�9���G���3�a��q��O��Q����6z�;�w�2�җM&�˻i�G�&�����\[H�-d:�./���)��U�9������Q_�J�s��7�(Y���Z�B�a�"7�4 -=ָĭ��X���M!@m�v؇��ִ�����=��d{S���-��S���]�����-�v���J�D��|�uf:�/��J�t��
���@@��iy��k?k�����,C~
���/nKS	����%��fZ�sr��o���fd��a-��J�J��X����y�@X��BX��_�r�ݰ#�Z�qEY�[�wgA�.#-*�z�҂�a��)���ۂ;���}�U`�����ͦ��A4�7�%��4Z��XZ�r��6ҭ����ɶN�[�c�B-3qp��ueazȁ�J�a�Xǀ.��d��%�Kk�q���=���`���g��>;7D�a\x���2��?�f޵�����梌�����ܞ
�X� <���`�?@�K�~���فb.�������+�)��i7�@ %;o0��8/N��.+Q{!��q����DҶXK_1`Q=���;2Ƥ	��_�؁���-����5����2���x:�E$s�t�ӽ�Ǧ�A��=��U�7��Df#�E�1%A��A��eH5}[��o�(��[(�8m3?_���=2)�&*
������K�lWԉi�\�Tj�L�M�[g����tR�5��^�Ѽ�]�}4����o���n��{Pq�}��:�-��u�������p����xl�4׽�H��p��̈��Z��	6��X��f�(rL:�9<���/��=�%~�ރ]�Pt?D����7���[��U87^��#�C˙s�эE�YU��n\��v��<�p����ݑ�����,Җ�d|�[�O�=����1߳�L�u�A�j8e��9��/PѤm���6}˺W'mF_/��ޖ���V����f�����U��P�����a��G)�S��R.�S��c�ꑛ��>:TـN�5���<�u#�ӏ���[�~hY�Q�Lg�����ĜQ�&�X�Vc�\�=T�'#�t~�O���n��z8�Smh�삤���SAJ�'�!����Hl��mX��<r���Mk:���(���GqJ'�E�y�]���&���,���Fg�M�O6���ȕ����a�����幧�Z�ג�
���n��|2[��j�9����-%E߭U�OxWc!��!�c�r9/��	j�Nh�����N��U	C��Z@aҘ�ܨ���ea�g̱�(��e�u�ؙF��f�����=��a]��{�:�H�#�A��B6�9вEƗ�3��{RAc��\OL/ɬ=�����&5C@tƷ!?�_ő�[g�O2��{0��ŋ̊����G���s���=��Ťf�L-N(B~���t�N8k\QP���6��,�<��W�L0��:��J]C���b��{����].U.μB�Wr.oŐ؞><p�Ô�z�2d����6/��C�ģ�$�]P�顺�v�`�ϴ�5j�"���y����Y�;U�ғ�D���6ܤQ�xܳs7��N��x��-�I>%�M�C0�a+o�qR�!�?����a��H��|��CS�Kc� ֝��g��g[q<5���s��,�ɴtC\���0߇]tZ��E33���y��nGc�����k�ٙ�wѬ\�����a�])��C{��.T�A�9�Q����<�A��-���Q�^l���|������������<)AҶ��V�:���޹۷�
����Epk���J�z[*���װf	s���	�����a�m��h��%-z?��Xå'��\Bu��v�)����hC�ת͏�y��NFX=�6��?I �ro��N����N����"���z��.�r�i����Ae��
��C��S��"�Hfi@�,��z՟%
�X���$x��5ZE[7��h+�4D�w|n�5�4��̂gM�s�9��M��,����:x�.3��*�0�I��qȣ[	�L�Ma���Z����}	�r��zP+�n�9(ݎ!��'����<�G��m���Y��aF�rO�U�"+j�[�OA=/�O�9�Ik��iT����v�dL�����B����F�f!&^Db
��0Ф`���Г�?��,=��
�Y��3����7K�K^�Yh/WlG��|�s�~�k�5�,)�o�]F���P�WO��x2�d�ą7������H�φ��,C��R���)E�o�Z���n�lY����^�F��(��<��Ϊ[��#�%m�x �`^`����'-=G�Ž�B�F��A�uc�%h�z�0�;d��@*PhbCcl� T�)��Ehr�L�*l.{�e�a��Ӌ� ��t��yB��'^��<�!�w�L�O/�/_}[���G��O��O=�E�3/�����Cn���*ۑ�#��J-��(ᗪ+���kԦ3��"�US�Aky
wf��'������:�����G����� \YY��Mہɖ�%��r����G��w�_�[b���0��r7vŮ5g�B�.<J86�4���2��?���׊�w-O�����%�D_�{`N��+��ߩ"l�I�I����",��[����m#p�~�jm8��M�������ΑjLo����+];���E3
���~�4�. ��������Ѧ�+�s.��q-�	��*��2��Z�ͽ������ܰ]g�p򧎶҃R	�k����
��9^Y�Uq���,{qZ��5.(G�CU���Qc��2 ��?��h.��%�(sW�q,+5�F٘�q��k`7���_���xzV�sgB�ua�����)�kT�
���<<���4ŗ*�>  :
U��E�â��x�����o���AO��bt�lo�"*T?��@���b�V�t�si.:j�¦��0�O{�,���s�J�~9\���QK��	a��J�1�-L��(