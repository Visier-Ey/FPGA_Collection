-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
NFX9rlwllI3OUhcl54vmLW6j3fvy9GE5Cp/jHIDVBhljzUeZ/+OacaT55mFywKiEKJqzjtbn7XCD
rLVSLS2hcwUb68oMdxNjcARgPwruU+T+xzXcZ8re20AJJJOq1TZVtEOhZt03oTUn2uUT3nE/kisF
Gk538Wbn57l2JMxPXW26bnSFlcnmcExaOHrd9sQ6SJddTSpD/k2q++7JJFxzKQHWIgpu4vm2OdzN
n1VGTKxIoHUzIBIElQr6/J6CzR4GZ2bzDlIfqdcSSP2wDBS2BLC8XwiKkgpOgF0EXErzgPDIB/xv
oUP2UXdItGhfmiwp7GLqOyjGgatE6CZR/6V/Rg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 16528)
`protect data_block
4WrhGbGHtw8m2k3o15tqK4GUHfOcinCZ4vxmNR+ixO+LC7lVxMlIrgqxyaHBg52hJ7TkoHJ0KCOY
CGCYRPJSu8Bd4k0Wyjw8OSh0yB//6qU0lh8KZV7nkiaIIoMlM2gdLXjMX3A6eE3hgPUYiTH+sIFP
/rERLIMnrRr9HRFVeyBLaiGIspo055PHNV9Z89XGp+r7pGCNbbNL+cH6SnhTcIqeLhkghjlKGKQj
tDspwqQjuwilp70xQ3m50selXCSXLnorh8m5FTWxXwhO1dyBvdDu05TJLlw2hmMuWVxbtLv3bvhk
9BXBTrzvm9NaJ6hVy31YoRCrf9tLHwisefQS8h7x2nEvvFieEB3IyGixHFgQodwiYxkhdBALpnvQ
9p+UMlfs8G2IRhO9ALisH3zek4mIu0cQYKv9YB8SxSCerS2E2RsPMlXXCuYH8KfCTYHyfr6nkFn3
qBcs1/pKIdwK9UWNNcet7ZY26qGdbtFodIZ//9OQ++gAAFcaXd6Sc8E0KhomIpTFV3uSHtjftULb
jKBXYXkJpwntPRyJc5h0l5bOJ4WDM3BTtskPQSAw7JoQMu4/G6O0+OMsi1RyY+kIgL4jNMzaMzVx
TfCLvqo1eN44ztcKMXl0H7nIFR2HhOHAhVja29HdKpzujJOsw+X7kYCUaGdedHWiBSifCaWa0exr
iU43paD0VqCAloOQ4Z2mc1qJS1FLgnzktzf+OWfjLAmIYOWSdXvhXnW5s/ocV44YEeB4U2xbOLOt
6aeNwi8OKgI6pB/CYMX66CdsM8wS8bPJP1Q6pgvqQq31IPe/Q8Fggw92iYHHHPHEP1oSjHCyJZm0
CzN2rvXYLQTSXPAlMe35qCdUybJMn+ail9rZVHMozp9Asa8GqYAY3RWfxfiQwKlnQTKm705SBonH
D6CScOwIcye+avkKyD2YCxNb5zbqKVr5bYKH8+WPIde4CPcuXGaPTVCjq6ZLACrt8wf46gREsf6q
FATOVxXK7fiRA0vnrC1mgqzNXYwQDffGscnEiyOcvzm9iM1B6bvHCjD1XEJtfFch3Mk9MpmiwZpc
3P2bVjpGWg6TncrD7T2Jy0BplIjnqyHSuuz5C+shARWLC+M4JVnQHOwTUYVSHfcFM7s/LWwgrTpw
PFqhTs4uYOkFapemZiE7FTM6V29u7GRuMffKlghfI+b5BiF7qYfM0cgsVqb7m8e5EHz6lzfmMcy3
1Sw2ucWih77WueEQi4ucMp40z5b7qWA7Zz2oNaq1gUV1m+2R3w/ZVYvTMXOe7ALeMzD9g51EElzv
dqm12zuytIUU2Z9RZ6xJrIGBZZhnczuy08VRgIyjwXO+EUj5ikXeh03PWeCEy1MKo6MjBa6qV6QW
d8LLN6gsMYULgxB29OeEt2UNmOq/cvY7cUB3n7OMNJjnJwHXK5Pva+jEjLAb7/pEdw2qjLznTAEZ
Ba4GC3cugIdSvuAMQLYwYSCk5XJGcdwEjPWqCYBrn8wv53Rij5TgKcpYfs87cYyZtHXGNZJnnCt5
wXcNQvOXmIJmsf+WaA/X3epILoNKEQYyuENu6lRQ3On62RfrUbkIojNREdpjqKbJUZcJB7w3DNnE
kqKJaOl8hjzbdpkh1vqUgdcEE6s7U4IHqrzuUiCxbgglWOexOe5gRueZmQ8zQ9JodlZmptQHCPcV
MelDXZZsQSa6nUA2NAZyUZh2efL5viM/PRG+umsH+GsZHG12DU4TXaXWjmg39YA9EzMexjGwOsIS
YR5L9xTC8N62dxfPdtm6klzdK6YDsArpy5BuYY2e94ec1gI///P1vdI8fqJVTFYlE3ZWnneB/Tjl
bU5ogI7xb4F6FfeuJ0YB6NMmVtNYrNlWwPPWA5qY3M8nGUw+S9w6VS9VDQPP1qo96h1un3VEiKWU
e8+8NJwzE+yGUnng9Ht0ratSwcMfR/f/e8ltQc2N+k8jh83/sPvtccX8NEfQ0ZX9wXrQabJlQK3e
ZlXgI4ycL2+uN/A9XI8jy8+glv19Nped/PRuFLjhwGbwVbJXLA2ycahzOHL+/ivu7wQyAo52DC0W
td9DE5oPl+hspFLvPHUPJXrOkw53rOpCekKrCA4sBfRsqu/tNMmS/zwJVpMeAwBvoD4MrlvvtmLp
fVPBQwepSCdOoBmfCSk6iaKThLFrgLzD1/8HgxjISw9KkkRXVYZsdAun2c1n0o46wAF9MFTYZFOT
vaERRMLst1oYegebtR4WgqjNzOC81mvqiCmk6zZ5l4AjFionID1B0KSVjBbRFspjS1p785O9xpBE
+zg4osVQrBhVpVdBp85dNNEFxft0bD6oMAqs+bq8btHy1W11/lpo6Kr51+8hSoJNP1R90gwivxUU
U6DeC8aqNrC2064jkXumHsKUSrggTpvrF4cUUrtAaiz4k/dUauFvue5glZHChPPVl/bwZPvwu99i
zoNmUZjh29fV8+iDnhgMntbeFtCuJxUiJrPtzJzhaN2WuilUc0pT4XrLarXYk9ZzGFXYGyGemaYH
kEDqpSOLCZVwp6ge85Hq5fcx0jI6Hsl9fUiejHZwCOzaUmo5UuTjcbXUqWH1w5EoR+lQ0ai3njtG
P0uGdGd8iBrYC8lUG6YkvMXiTlV1XJq8hHS1VZLVUIl3rtKekyRQ2TgtP55vM15ehxXSOH6JqDaA
up2s3ktCYSrwRF9qVdtfoJL0lKOieiP3psWr+G/fivYe2kzshuZzaPEcn8QmdIlP1xtU3a20Rsyb
Js3EGX3zrIz5ytp/BeUifzJiu3yN+3t6TY1N+B+NaSV2FxkuSPMMql6ztzf8+uJ93VyVrpxVr9CU
MaFbqT7GvUWr5QmMkM3+ykGE4LPN5GjPZCgBRAjLiB7Ik9ZqH0NGvU+96fYBxGdM6HznydoKFWqR
OqmQLpZ02O50bsfq8Iovvqi6kHqISwtWfudNyfrOy5xsqVInoC2zGor7zulXGIE96Dfua9R8vwx8
v1bPdkuMfcLoS0eXZP9DagDettRn/ytPoEzz/7kYWwTq2hyPWlYXWDodjGTl5nghwp9q2bAjmYBn
NI7mevg9esjpe+cZVLAgkUE8WU1JQJQ9uaAe3vmH0QEfC5spL/+DtWx8a8lQSdW7Dk+QBfDPZAPH
e4gAzWV+Ea3ewTAKbQAL/VEVo7hSc3NSIqGkfS0vQNCILZ2u8jBHfuzF8ZKxt8mTkHE1vR1TrODj
AwYATXE7JQC5XkB30BN5kfhM8cwxk0IIwE2HypsL6JaXJwyGfdJYBCMXu/9f6XC2yZ1/qpK5j+tT
8gMRA5cpbk7sn5UjndYuCy+tC8Sk6WTc8hu7Exdbs6fce+N6xKfP3CZpco8n66QeUNFZoKQOzlR8
GxA/XwRVGcvHmBUxI4tGpAgnaQDqKOh/wFR8NYAxQdyKQ7sTYJhp8uEDvStFtINkYuqd8QrrpOZ6
jvohDisQSzoXYREh6J/ZadHmRZxL5r0tF8mHXL/k3rauBoibfDLzSw+HFZiNNhMWVWiPBLqK9ATA
ho+vNFKQ3rALNMyLdnri+fL0DSh4GYWOg7wQUlvtpiOIQKECFalo+5bjBodvc5tYVnRj7Y/FOcW3
NjF4BfuQlsoIIA+6HAft8T6eO1kW0Jd/H8VPJk9wM7i8kRjhtPa8Wac2XSfH17iZDqbdFDlrr5H1
BVF9WPX2LrteSvKxxkM58NyYmPioA1ljCGnhBT0DuX1bLfKR/pujI472fw069o/+YtE1Sc00Ld91
ZlkYiVaXUZBBVSP28sg756leNPaQhVqqWi7PC4Op74/4Vw3FGYVpWLv9EnSDHpS4xEa+rzESZ9A4
go3clMFH2cfIdKyRqJr11Of/CF/EnVlQeW0GF8rnuiOtpvEGy9iMNL5q/UA7FJGKUztr6WGHx70N
j0lUVS92SD4PQhG6MJJE5t9ENQJOT81ZzftcDvnnih4Fx8ZwB6ogSRX6yX0I+IZVoGoKi6TtSdm/
wC+zHmIO7estdCFzmjylSNuGCeTwjPxwqp1ZMdoBOjq9TOjiJkADNhyWNaF99lWkVBkiVk0eq514
WRFfalExwcYB8ABW5AYHCRfFaXYDzz3aPmvwdf8cUe7ukvioeusDpEsDk/EEWxr1fE3GKAMAYtzb
tARXUC+7pTlOiD9hsuLNFSukK8YikBru1DJ8Hfb5nUY7r8bMfCOjg+PG9rO8/bFz5iyZa/hb3fjh
88f9bikIn9JaXbcYCk8CwJof6693Y+tpd5mONEXOtQg6a7DaA0kbEW6Qs7ygluOo9ewrOg1msvaI
+V7tBPhnhGVKtDjTSJHmXKS91qnl/ijshCWgSkKYa9XM+UujOkt0iGHxZV5BMEzLcyoYU0iDucI+
wJErkbZ1T0UvP7lp0V7XKTwGzGM/77b9xvWiI9nCr3R5Lwlex/IxKA47DatmHBCIrYc6i7iWclCX
QJKosgD2/2D9JX127UTY2g9P5abmhc0icl8lbDzHcCELEg7Hdd+jY/vbRJpdv40o9qHG31/9x7Eu
BzVKKUYQsDvjGwKdCTkXttG7Mu48n3kDOBDxigfiuCh6yweWAgdDHvPgCPWLiRSgZL2Ogp6jSl0Z
lf1hQucZK6DxVYeXkg29pfrI2yS83UOe01903+07Knzg/Tq9IFgYQ+hoKMuTZOZq2Qm0e6BIqWLG
7tfiRrAwol3ARwnIBWS7RNmTyYdjghShvMLkHNGwvAmT7veb17jn+5YEmSN4N7eqkaAkKuQ6Y1KC
9VNddjVLin8F9lDRrmIciyQNsDdlJtCc94XROJtFAaiUxyrdgUyyMN446929Z7IeqHXV9RdxV1bn
eb3b/JAeuhKYkx8RphYDYNorQKCs0ODfq1NMod/4WcY0ubKsmj6/txyvzh9sph8RIjLBAIpMz8Zp
kAOrQn6cmX31lrOA060eJbxFJM7rjTLNPozgjVHxBogtZs4DbnbcZJrQS9cdjza1e/MGUwHhv//P
POYCD0t+otQIUROL70hsYdbWKsc2GhkYez0iWAXJg3AxwDxi40rBV6epSgo+rP30ChSxhO4C+7Iz
hjm4im2CAt1of7KQMogppDcZI1jo5MHyaRFBoa+t6CAxmMmi6ST+EZk+ARlp0fOMOItzpoBT+gkb
VeyNTmMj/bBRIIC8SDtOSBwx6Dlkp5oLJLDZXf+bvHG9W4zlhHz1tNeuRvtExfcKOvZU1+vzsaxW
+DkS3hpSHPr/aaiNB66rzd1Dwhe9aVdRW7rifS4nnYfzg5TWG5jnPFV5SSrE1efcNayWxZvESoGP
tlpRfiaZk2Mp+PU7aBFfzoeXgr+JTOcBH1DFZ+v2dTZb/zWGTky8ASVS0b5l7fFtgWP2L3PxdP0b
uRs6IxfaDFW70O7k6XtI1BZcIWCaROYKKkwpP/bFIC0ZHmO98BXwtBdlPV7dziBZnEEeIikR+r17
JakfhjNw7PTrun5eWfvCgyRJxx5dAvOZ/BIAk84xFnHiSE/fVkEWZoXkyFCix9Pqa0xz8jNJ9v3W
Rbe7+6ljF42QBjvtXpCln7Jj0Zs+SmoHfYdwk+BfGpb1oAWX9iAyKsOudhNxOblz79GMJJ5jobtu
V/Cs1hcrLFUdn8SdLtc8k1qWTXZGpa6Yn2mGaOD2YxPKR/qJAZrdGS/XPwQf+ZBLQPACDo86c95k
i4iOPBCd5satYzhaGg21be8OHM/GXOxDb8cep5uyuYlIAFPR/W85W7H1vAnrsRdjkgyuALuxxX7Z
LQjMbmsBA2vsDt2VKDY2nCCc9yBcmiXl0iZHGudLvwG7pSlQMxvz48KoNntN5tMewqgGlrdqzi38
uAHAtEjNiqLA8lj8KZYch446gi2o3fXvZNUGn2/6ZiQbVQbhvQj4PO2hdJwzxzA68lUqsdel+yKU
DlAVAJ0N8Criz4p3X2p5ReS4U6Ag+iPS7/D4RTIj85Qo8kHUZ0GrhEY3mh0ZvwZbA5mg/duCBS5P
5Bwbee8AKfJkC1o75RB9IAkKerUcuNNrLXo0UbBBiGE3UU9RPAfqSt4K4ektxGEU27ZFo2I2wvhX
ezPow7x8vvlnnpxf/J7pI4y77x265bcxL/caNQyMPK5s8sOtnLp4/k7ym4bHs7SQNm2W/tVOXDYv
C7RClXY3Y8l5q+TKCptF/wdC1bWgnr1k5QoaODKI/zr2ieeBNQVhcQdejDwybx/NXSZfPol/eKNf
ZA4IbXuHucxlFVwNf805R0tI7Ftjjxn/wpPAf86HIDe0XNuzvAiXfu44BpofgSSs+2GMOv0BvruP
jfMzs0lOdWjzOQ00MOHxjGFCr4pFn2vegj3O6NPrd+i1yl1uLdjqDVOpud1xPdz3NjrUkCwRVUy9
q6Exf3aB8mkeXOS8+ALmxNF4L8RQRUQOZEdu4K4lfa3WnL86Xxtd9Wvk+MEF8LvQhFSQDbkxJnWa
C+E8bm6Ajl0G554NXMYeJ28vHSB+QgJgcoMkcAYCoRYiDJdIxNOUvVBfyRblMfrMFZODgiDH7Sbm
0YLBWZmQ7mp8ly8rFwud7ELWTRACJJTRiQ08DF8qDs1vYs3XiqPnzpF7QbtGuATSdDJ7aWkULGjM
R4ftVuae4G1AnEUTyiX/ehig+kRHTTHsS0ef4vHpHCAMOsh0XfgsoJef+AbXDVSMKKOAOAV1Xj8k
VSNDDmxR5NS3rXu/fhCaiLXyZrmzq5A2HSTonJeVGsw6EyQMX74y7YPtCO906tjPgmGfccalTupY
kwaBE13snzdF7cw3r8uKc9jezVu/vqo4tlRlS8Q9UMy6BRNaSPDEJYPNXgQfUXBbEJ3AoqQCDoDH
ky4YxOjdvvuFkfYzH2D7fEqOO05XnQS0s+9EMmZeqySwUAQg0gKnzkU55XZIU3oeEhWDPSrnosvP
O2wx1DCH4lWdbN0vnmDpie5cPsWnz8t55mMM7hpSbpBL1qzTqQf1Jo84lSeMVDd3J0sbEwHawFfe
A0ZG0dvw+tKFM/Hm6dpqWPGA1qNgnW0HvFk8fmoAJUIKhn9T/LwqsI6PZfDHYf4XM9Cww1FIr2GO
McPUgzxiv32J0PoFXPkA663Uoo6typSqX6Ma6pfOPk4WtIpl9ENE9/2eO+PTez0TK1zDxey+K7Q9
SwXjbXjpoPPI8duihmTrsd2HCOh5PIO7GIEMTyRfavulTX4yaXFVBNE3tVi/oeAJQSrCcyI2N/uZ
5lD+oLI5A6cBZ12vYUUZ70iJbcwtEaIeaxs0zXyC+3b+QdZNIjto7Qy/UAquy7zGUpzvpfreVXU3
XaXODYmnfce162T90aKpQBI/HLOK0ZyMumfpdx/5hjOcM6bDR9Qcywf438RpBtlgWqUNgH21nYsu
qlFzvx4JSfdH1wPy2bxFRt/j6omx3ig6b/aIkSSbbMQHngYVXVUg1twOBH5So3AuetQX3EvLYqWM
k/O5kXBwHhdqdKaTRrXvnQQAxSO2GVCWpNmyV7t2zur7n6R2vEaJVP8aigaWT7nB7Uyv2I4y438T
/rHnqgzS/EVns/bXa9LuwHOQ5D+hNJtGIVdNI07XnKtIGw5WjSoR8BVown3TYoQ7CIg8yEn1WfET
yvtK8f8H8y534Fi0f6FTai0zHdVONDoJBajoQ+b0UZOVLQOHUyke4ijDVI09vuuvJdYSXW0qc5j+
9hX8isNjMqu93KW+7R88KZtXBj0hPFpB2kqQdSjmtWULVO5feH9TZT6YScf9vjoQT3v+qOwK5vmr
/4p+RXGW5ZhNNegl2PSXbBmVv40/hMUwfGQdEQDLMKKsr58hnJIGlWKgqlHTk3jI/e9zIa5P/Gt4
QOZfgVsBbEhc0WtBaGUD2to4PqE3WhHl5zBJY+/51mO/gBvtZyJ7LzR1qYgtGfm+eoQJxhDGXWDJ
E79JmI8W5+pnyCkeEjPqY5NagTw4oD5CReX61l75EdIb3IdbCDxZcKeW/M9cWciVI5RwPn+F2FGG
nPJAqKtE2yOA7dyBHR5r9HDpxTFn12CsJdHrc2qCH4DlH8/M+wfVs0KpZQKcSlyWrvTOGP+iq3h0
M+9P+7jQ8VMtJAaleNgO01OyM/YxgLMPjugOd44PQT8S/Is81NBshgW201jt/CQPQTurI5t0ute2
TwAhccxTIAoiMkzmaopwFUpTGT2XU4vUpz54gHEbsRIKxSLxOcxJZWzxdapHYcCkmnYNyTrwuglG
//nzwlsDi+HLsouI69mrX1s/WempliUhzgyl5gFSAbB2er02YUdAcGq72C7keZx3b1hBt5MqED2b
0tEz+ckbzqbBCh3PnO8SxzW0Qdc6Bk51gOss9cUrQ8Y9kOv10tB0ZAgA1jfVP/TShV2+vk/dO6mN
gu6ZgQ0oJm1w2jNCgubBPmxkoc4yTJ4kghe+nz6qDRI9QZA/Vo5DmUQg7HgAC+lgZqXtUJ/ikxsB
a7+HdnJs/UItS9JW/uBUSxQ3Y/LOgx0AMayaXDMwFg3V/VrvOFwIAZl5CTxC4EACrlY8oxyfEd56
GqLZJaU7Uykcr4HDPZgFw3AkIQ14gdTvxzps8iYXB7FUao95Ow3/Tl3yybcTbj0kNYhf2wuXktr0
C2wcFuwAt/cJxMLaaNbmM/ZG+Uf51wyroiWv1u1BL6jagkBtToIowmzSIO/Tst8H2HCw8w3CPoa7
zoBPByk6EJp8I7DD5yptZ/wQd75mA4TOV9qCorpb8cFbWMaU6wGJT5hCjFvaHdqEYU76U6yBdNsj
7unBdsxjPAjlo9v8hQ3Pjrrq+R2ahXjTtD7QhA4O1KpigSG3BkjjuWR1/bU+Yki9QQMxRm/gpAKy
QUxfOXRz5peG6IVCywxHS27dGgwu7Ip8iuw63HeyxCatt2/yHlWL5l9wnc9CArnMRsT7Eq8DEZx3
bfXTJUxixUERGDfrCigODS7AtnmDTK/5fMEBiewsMNoNQsoaMCfN7vVfUQrLDRx6KsGPMNqn4fgB
qS6+R8Njj+e/Pwt4a/nfNPrzqmkPD3iizGlZTCYpNkpz6WmsIrgy8T0Q718xi22CRq1oI34Tucva
2UUCJ3mdeiGw1MzNYGXRT+/yp1oNelvgYLPA6b3AcDtTYOD5UMDXZn8VKQBINbmo2qQkdcV9w9Qh
NE9TyihkrF/jYIecHnx8OqfJVoJdwawLCVbFJJg+QffJLJDk/jZWODqR7ToH7Yngt6IoyiPPZFeA
vCdAfhQypH0VDeoLiV9VSOqwLEwG4hn9NeM7lPkTaAGFxt6jzL91U6K6ngXC3ZXSdNAuKCx0QsLX
duudKj3ppJiRZRWBzI7vetaCfBM4FvaOU6luTMJwdGYbJrFBAxDj/aqw2yhYLllWDv164fwrc8oQ
CBtnkxiaNi9XXU7MHelCtJYlhZMYoPpobp0ieQO+DutRPXdGuuNNb2HgSJAqzsOu3KF+fgB2VWAu
r4UHX3CbfpafXXRqfIGrpUJ2L5aGqns3qQfXI899FOJG0cZHRyEJ8TEsiI6rtOL+lA8iPh0J02T0
7Nn1TWzVEW1MCrZA/l7G/onjeNlYlxEuuA1C9Cb4mNqyMHTwwt3LmFAOWYLaFGwlbgtFL010ck+g
P8k+k9TohpNVXTePY3TyG3E2cKIChiSwxBHTDOhXdeWTnzgQ5q36dqnT0rzXc4Ff1u8eYurPWo0S
O4Duo76P295eF7sgZBUAHMD6LT0fngwzjixsZuKRWMM9DhYKkIB82CFMJzhhfmOavVHfIzyJXD7q
M23EDeZoRkbSm5cZT4r9KEo55laLaWoM52+LgFqME/EbbiyDeEcjenNR68qjIs5u2NKwKlFbLeIE
7q+4OcVC/2G5g5w64UtG2gkCUsiacKD8JBRv9OByIISUHcQGIR/t4fxCys8oFL+8Vx2/WYYxnH3o
eEouBGtI48VYsknFkOWp8sr6GX4gUUhMxp+HwQMLMzvZw0JmqvGszbXrm5VIVZMQ2XfRuXxL8hZK
ZeibcnN/1abFqPXCarOmHH6PnQNFamPw+2YkY1rRn9g16Vv4syXfpvUZfCKlXRJG2eZTV2pkZ63x
GdWDvAxCSqlOZixtmeshSs1klLbdFO8tknWO0bi2rx5kQxZGQyS8EvMcQnjoZhUJ2V4b4a/kF/d+
BReocWhJcizObCWRYJlPtODkvBb9nlzVZiBhKgHR/zHeLY+UmBAUv7fEPTHVfWmCnc3vsKh/CBek
HLzFRK+mfD+fNC2wnxUg2T7sE4/6oyAqZEsiCkSJSnOVKQswBcF5PeXkFLGqeM9KvvkIE7ERjFw8
PBLMDOACOqWJcEKkpojCtT2cSU4x3yi4jaKaDKWJUipY5bzTxRzOz0n45hZD/BMsFhV3sKqjEalq
ysKZpqJn58dqKZ3qMx4KgX2eWh2iXldB82Yf8Pp9WpCv1WwGEh4KYAzhrXmjWBlxXRuvAW86Digx
mc0X79D31c2vUI0jnxqjxUBQ1mQIf1cWU93U23KGG4YLcv8fWEqqiNbmz45SfBxZ4rPMiiSnHTMl
JPcBB1g78iYTWsnzpHehZbBNjjBJioULDejV1ZGOsdrkPB/it+PTStPaIGfKN0E4Pmk61bgKOA+2
SSdm5H3M5YzfMdvlI+mtvBZZBwg9DVyGSht/dOx3IO/rAmfPFePeOBjYMoja8RvIayg42F/3Lqjk
Y1NVU3CFGzQ3s/jQIgadA5McSkFVEX+veok2xqwEypfcG+V3RsPwjOJ/0nION+GWX/g5K5SwsOjC
iZ7fhMF/idLpACpgnn7F+b+pDcm5bb514U/qYupUW4NkwNxfJuNNxvwZZcVhgla9MVN4uwM+XMFs
Dnl9zG84bptJRIvSZsILG59b5ihFqlTwZ6T8iE1Jb7eOBU/oRpQi6cNbfEeXrNHsfsQdKm84nCFF
dIlTVOaKR6/rwflZ0LjP395u7Zf2/0lSWbUDUj2CBCaupsoSeSykGHtkTKL1upbOtuJkGAO2PVbk
ZwhHAst4xf3GRY2pYUEUsJynR+WTwS995NoVe3p9XNiSu2UCbawbIXH4jkeIiRurZVG8j03FxHIa
9Yip132EbLU5fTEriI0FcQNbnGcO5p0UwNPDH4DOAUc98YW/7z826uP1GA18PLMHxmBYTjSKbJ5L
gYVQLalXSJo9K0xaIT9hSdSWOk5TcSMK8m1dbL9TxonA7+essUhcKdpHmC+11AtBGEF5ClSI/LAw
19vV3Nbv6+P1rrpRba5rHGYyp5OZXKP9WcyBHK/oqSn9oxKafD0xaMRyAS86Po5ScyyjFOsLHQXc
n70bE9gP2K8Me+UKNJxVg7d4xTTPFlAgqd3081DK1vXdRikAM3MzZY3s0lDf4xMgw4PCzp2mgWEg
Q1Yhpm7fYUVMjM4WPrrs7q741cchez7Z+fxAeupiy4+FxBeyNEejb0LS6RoS+OfWEDGmUoY/Sdgq
0S5MUZG4YWljvE0eSDJxoG+z+KMBG4uWVaGextrvfB6CxNspuKV4XOHltI/kuV5ZycqgVuvczQ6g
gvCH7aN0WbxHEjxp253LSOk6MvyvrMI+DK1aQFYxbctk+qQSIuJdb6v+CBetT5t5JkrSqyEKs7oB
6CTBWRXRfsusZAUY01vVsQH6JOysqYhUFsM4FpqGsfEsDKahuMpeZ6ARd2wPIXYoYwu262mVf2+Q
yVL3Ap4QC+CC+a297bvP1YvW4VfvjgnC6mdcowlAj0ckU8Kek5+8FMUlpavPZJty/P/AWBD2JP8I
aU9PUjdmwc6w981lRxA34fswSmIA+4GXZ6cVVj1+GQyQe+KrOVvr0YsEaARcddT/EXkDHbljEGff
kiVwTWkHwAjQodQiuBbMacLqkyW0uyrOdb334LvW1szX2/5ENW5/PSG8m0UOg2NyWTdLExBmgDGt
GRf3swUx81T9Wq85xVC869BkYnfI1DGu00m3eRIo0bvam96s82Z0x36DLlFQSa1er0ZYytkY1EWc
NEN7ludswMV1Qvd1bXBdkGla8vYwJQMkEGpsYvha6h7Ml4KfHyWZDG08wqjf8Q52XZwUp68Uy3ou
aiCTxrV0FqHy2B2ML5b3B9HkLlwEJPr7HPyl0aRoMRgq9tXyTShTem94EiA9InEjg9VENW6o0crX
G4hg9gRUcTF4OfhMRYmhyQEUuQ0/cdUDkNPilrO6w9FQ+UXDrXaXsU2n7N0YxYJKwp1t88x3fjWZ
/lrc0wi8ylsPUK2AMtd+/P7yq2bPZNZObErT9f1kbJLkis+5P2FQlh6IzwiRxlFpgrioNf31kqfd
0/KBnzNyA3DHGdj9AcvmK9SI9dj6fFYM5XPxcRjKOAxVrqStkLSJ9SWxaoMBBIqFqFSz6vap6qy1
xN9PlOycbpIa3aj7d4xAp9OM944fr8+ny6h3bzaxy4oKIh5L5MgnpLEzbWX1WZJ/StRIEjngfzly
MCKlkcvWqiH1etFmlLWLgrfdDX77cXDzSf4gVIMUKSkKsnEY44h/zxCocBpTU9wYmAHAIszRwofq
cVafr2GbnmR3ZcOjBb5VqZfICh2Y9p8ROmz2nODAKmVYeWpplKShDoXeOUOIprtryPXymTaZoBFX
SN5Btt2iAwpv0SxMZwphxt1VCzD2d1Pz4yM7expLnhbPY3xcZ8jIjyNUEKpBATdLS9tYo033y2cJ
LLbGGedXa/bqH7sYiLju6cJ0nPfjTSCpGaehOhKVCHZJzp3C7UBd76h3Bh7+gRkddsWY0h5iPGKC
IMS8LajlpwP6oIGIiCT4yY5VOR871LnLHJhlBzHL2/PmM20TF4QSkxCf2W25vgXCV1Al2T/CGAlj
hT38FrSzpWR78VG8A5SXQjs2n2f1VBSOqPGw00C3IGcoKJ5Pha3HsyChjn7E4xJQFFAdkmSPvSOP
U9b9GkOSlzJusu76WYmpxXOGcqfAdGX8vlVAQ4Up/ymHcsNQSEvXV5AFrTu5wWfFLmumpvpRFZAr
Qmv+ygYpxu9bEgD6IM7kyTQkhaNqb1c41rh9/hWNMKUp9g/PySE/Lm/FHqShNfDunEt4nHiMXhEx
52kUZ374TC35VTNtWuarqiiLvwbbXKZ7qK/E4ZQ9UGmfLuMlJMj6vLjAQHLVmNUba+0lxFvYnJrV
XHhNk3cduhC+yeG1SayGm8yvtr/w4NCt6xyyJqvxcg7MREoD72iO7ZAexg2ELXloCIrsgPN36+0P
hpuBtqWpv13B/FmnQUohQwDF9oU8kYHG/6qMZTeGM3ZOSFaivGs2frDGoJq2+1+HfTVmzzwNBDNI
+/+PvoMICPU4Kb4puDF8uFksLA/ZwnE5I2lnNLDdj1jGdzNQxn3VqI5HdF7iO+EEzjwOUMSZz5Hn
AaMv3eNTt4vU65+e5iwioDDY2XF3VYgR9nLffzV7VUjDySHG6PyxTOxeUTkroJeXIaeHCpP6NdlM
tlmYlV7oimkowlNpjmgiwdr3GbauiUPMZhhnJqgz926j0Za6DNmdXy1nANcmXxOIOmSCqtfH9lsd
Nk2FCZ/EH1PbtHeci2XVebKm0wgV/+Vb4Wp2cw8fP3t7QWuW21t1AWmTNs5+cJW7DvgCq8k9k3Vh
fmPUH/lB8M8BvbkqLbGynuc3fsbXuybhkAhh2NNzwmyUJ0CgW3JHwv4QhvWXMog+xXh3BJnb7eC0
0xea41Op3uF3tgmCDrO82vb9dD3L1OU2LikqXixR1zAdtDWGkUXocikBf2yEiNBrWqyGcfuosfrI
Cz2aqgVtJklThO/Z28nfx0cyCnksErrf0CwA+K29/6Uxg7CUQeN4plrXuHFqzEG4kuvFv1/dNC5m
EJcyjKDDRb8KVT9MV0pZyfDkpI4qmZA6Yt89TfO0H0NaxstxgIvMERpygxDFBgsJFZHvt5dj5FAF
iZs7PK9gjYQjs+2qYRM5EAW+yFS8SC60AhoKN8wxWJQa5hiYj/QYJcHDGXiLU4d4gZlZVqnGWUOB
sR6MO8BkYm5hLBSUZH4upz2ADtPhFuDWSoA6GdnVgMJya5D75dqAZuGAbrBYL+U2xjqM9PGTDMDk
vtXsfv91ijnpWXokZrBk1oltOmATU0QgRofYjZxf4umZdPkCc8RKwpQpVDCXBxhDpu89WyNo5Qup
J5+eR/KMVJfQMUD8RzdAA6GEtPJZ7J/QZujlkprWdEEA7AEj6jcXtaWzMYpRHF+fHRRZpriW3L0d
amKA27W6xeiYFZoEI1OGChWyT7La8bdz6WjXyN50kQn2eKFWKfouWobBaFDxW0AGiHcPlgOP8vMB
OHmm30xdwUa9ohv24N74ae+zTvWRKAJzpQHjAY0KhX0bqX4arw6zIQvq5D/1m0ZqAunb7wxM/k6K
YEPkE5uxhlQA62U7nvO4gHOfEWtSsfKLMDHUhKO0HlkuYFwm/HkiJ93hfO4lNbsoh8ERaU/pXEJI
0bZk1nhPebDFvfdI8IbgBsbg5v9HUZ0hOh3sEkX/O6WOzLMx0BjhzTh9fqocCjmuu35BqioDq1Ru
D4iAXiACVaYekqKTQ1x/bSHGmGMtepL/JfLu8I6R0vGEelsqLu86j+2Wbk3kt5DpHS6AEK5iv1gz
OkXAo1zCJjIImKxk8RiYikwTcre07YiYkmtfg7lwv9UFy2UCobLfhZpO7ewxSa9HY7Rby9uddGoT
u9gpYqM9AV1E1Ia+owY9Z9DB3NjuEaohTwcIo7/TgDTvTpEmoVZgTvILdn7OctodU9ZgZA6pOnuE
aPAYCgs1CGjkY3GxwMAB4NiS48F8IY9/di3QEi45nEURbgfhg7+r+Cbo2yHFw5tNIzHPKiUsne2W
CUsNjB7/utGMWhFbbSfpXv+ZENrQuNFK15BrMnZOuFOmUvLzEHxjlSqwfTuRo5PjaibjoK7+vUQ8
j3Yo11e7fKJlgGQ9O/IJfaIWvBQbJVP4z4aYDgDIJZJwkJ+QdSzrU2yI7W5sr5jDb2qyg3czY1sB
gNQjokQSltLD97d3T3mEv8TQdTe4dohi7UBo2mXrqIyhvHK6J6jtWvMbSRdeaWi9R3VCBUUBMZQO
bfwB7aOWED3LmW/mbP3JIUwsGdY4O24CqY03mXq2afYZgGgrBAnSPk/G5tfPVsRkxONevZVoXU17
uy6b/2yabUXQ1zRfxjsQhaS34dNOJdkrIOH+Nmd6LuB0s7K5dtN0xvUiAsvKopaUH5Xr0oEVglKF
dJHtZsBmS71Lm0TjUx6X5J5hxPKyszhJa0aPdlqlUUE/Y92KnT1EgATxf/TbRhTjrW6uXVRau5D3
F7TxxApLR1/rWtEp1MfT7VaITv3SPARkLl9wRkuSjk2gh9SEVf3GFUHZb7w1gQlAXg31VYn3dp4i
Knu8XTb6GHJe2KATexmOVcjbn1aa407j/IxmAGcCmdzAn2zQAE8lY784wMOKTYk7XDaC2WCzlK/6
ZnPuHUaAJ4MtYvIWFu3WcHC8jtPEAQesRtAsmYDq6wZv2d9rVeSMEBoLvVu5QOtAQYl1d0kamEV4
DaDsb/tpeb1cad6h9FiiTy0wf7ol+gUmcMXVG9X75vsDdj1YOZSqYAd7FzNBAprgyt5j7Xq+ePX4
wgV9RJBA97/lXSg/23pz50YOiTdat9V95J87JqhX5Y4CuQ/oRJJH8B+wUx0BUD4YRGRSR3dwUg+w
RJDkNyZvLQ2JeG9aBrAtH0kcyi/SA3qoWz/bb7m26BLEFlvsn9UJwSigKFqj0vAO1Z4Ut4BejF3j
oPxZyxqTW/CIjm+F+v4QTmDDbZKdGHLBZEqpMyaEEErmtS4kDTGEBprQ71JHMvkE7zmH6B/q7QuK
OzOLDcdhX2TdvAaIv9T6dakJwuAU91Z8w9b8I1zJousZev0IuyhwuV1jQBbJOBUjigDD7utQ6sXy
WGc2BdSZkKJ/sBzbALVC1SRoD3N4xrO5QAakFl8XruGhAfp98M45joPECr9FVGMtSfEsePseEM+6
ESVggGHQZB55aBs4l7L/XdGEQW5K+4o95NrNPa3eFgllpX4hQXyErRIhVMA0SOMQus+uivKhJnX1
9oc63axod+hSfyXaO+p1EH8EhYtAXtFeXTD0Nj1mj4W5H7gRDT1xF0J79LOhh+K14SXwO9OeVycS
LyK8W28GaineFTJGbngiZlk+6CyUpz5FL+1xcK8NLDQU1ffEkX/3YRdRP6M9G9vZSPnIfzFKYsa1
rfUkTruSGlB9gm3tQt2iEGiDycW5/F2WFbBdB3VRN12HvRFQRCHeNVkwMXrxej92C8QAhA/MYEm5
W7Tchg3PdYS84Loj3j23nWLBKrtFOYydDXm8WoHPf3WmTT4Jn1v/egsnaBFwFWSdbUHGBptAXsOe
LNM1+UY7y48D/G+R72xkYVn12luCUV5lwRaeYSJ5YVhIOTsmMcnZNHg78/kw/ka1pldALCv2OadN
n7z/lu35EtQsqCo3j2VRBDJhUY4F6Gho8T/vfUmXCTa7YDtzGJIda6pxhRt/Ayp+dRRFWG66jphd
sGDvjfP4CgFAWA62t6eHZsXmdTFmkpkMpSDH7cfshqoo5/XXWuKjlDSAwgnXOpX74KwfLRv91gg/
LUlRpTv7Uepb/HmP2Eqqc82z6oj6W78xYbIIO3Vsb/WyMMJXSy7eTCzs9OCun8YQWo6KQ0yajSdm
sbVb1yBbC2TrURlqlid2VhVd6C+5lRfol/SsBjmzv4LHbDJW1Ldbrw8BYKpFQ/pa2Ay/HbdhxJse
N8YOCdJtsovrgD8qptCEWQvuIM+7gAUoZQJhXUWEy/UYPHyJW/O4vyGwv7C4bvrnqrDBd2KIg1gm
XSKcU13Jugh5A9duYvos1h77vndaxkglpSRRtbGLKoy4wciu0U8TDecVBV1FOXgMWmL5xUZ4Y4Jk
Qk1BLk4CRH1kFdnBOl+xqqXKGgzaK29ZglhKzMIRl+DNkenEl9WZI2b1/tnG4nUQVKXnLdVGT26b
q9hzVFI/UkEaMcGHgfrYwlyCe6cCf5ItNJXQygsCRQ1V/HSIc8Q4OaKL0GkJeA+ekEOfxUj9V8pk
NgE5EFv38TCuFfSHn/L8FEyIo1Lx2aXO/1ngeH9TFnBrxVz+K667ydiW7th45FRVfVr1at99w9XM
tsc4VoEOKBuUHWsf2uq0Z1hTaMNxNa9EPf+z0a0Ac01EMI3384s5jABRtxOG0Z54xhnrZcULkpBn
+tYdQJbvjodJFaG3QYWXtq5qO01jWPZGxGQ4yPSJ9v8o+l4IRAAkhDcVzgMMvj0CPDW25aJoZmzv
uTREEIDMl/JbXfioYLNwpYxmMW8Nqixzs6PMINYjWaQrxs76XKAbcphjCyDJyqLVoSfgOQRbNVHx
2DeNCNVlUcX6iEbC3P4PwOZJVFWukZQZMWkujbrq9hjak0EhbhDkDuACPezSFiwgMqrYrypgjZRG
t6FXDLv2aTMi6fmtJk2TJtTh0PP1BH9NoptCJMmSdL0AIdvRliQL/aHsG29vErPi1X3MyHHwsNJV
H4cj4V1PWLbrSxx47dkupkjJAp4L8GR2ZdcX2iQr5Vk7lmmHoz7vB+5mQVrJoKDYHef3RV8lFI0L
Mbmr7YvEmjrufC7t9+Qkfxq5JvovuAAM+0gnNdXK6OwCXnXJW0+TOQsurqvrsWuqhmuxSW9/kM/J
fMgpngR7ixnNFYZW21lDPyhewsecZ3R9ikEamOPTKgfCJE5WIpajSLKW5CD78szHjFfOF1mhE4II
zs7a27ob3faQbLr9Bw7n9krYCorXh+P1y6YibknF6ZH4uqvzb9cvuIpWTSCwiiO8BheKEcA4JpGX
Fu09/zGs72Ivf4T1NNlcANUsOn0aVs1Pk1Js/+EgeQ0Jugmmen8PO7Gca3PeNI5///wWTxz7k4T6
G2oxolPelsQdq7XeAwHpQl5y0RRhxHjDpV25ErGAXTC4RjFflybc2usR+1pNXusyuksYGudnpn8q
6VSAFndvZuRnEwi3OxxeG6MoI7xjG34JRIIF0Hi6Vb/0FXfC6EfvcU0Q8PCDYkmpP4VPBvnROW2z
/s7nyTaAB4Z3KENXGf6+CBZNa7PXxUvM2gaNro7bIicEuzRomfsLIcO8fZYPsaom3cHqgqHbTCBZ
JK7x1bKdsG+ZaOiqHU7IJrzsgJ5T3QH7rGthoVloEKk88RkF6Zp5017H1O1XKUX61nTvaeM06pV5
tU2ih9LMFc3PD7HVpIXUg8O6sqdsAZx4rRjPjwXtX40RvYQE1ygI/C7hYtaSAc9oPezepLdomnDA
R5uI7vwbwaIiNtSfNuE+QOw/A0F59wtsuuR2uDsUBIqK+glmPH6paqxbA19WfJRl1+4z+QVNhp5S
6tSqZzxRRmRtUwM1lBAa7z4eF9lpuz5pU3MMG8GHLd5REawBuzAJHABVIsZj5QD222mMYTekNf5M
JGwcDaLNwAR1tB0N5bRIgdS5axLo+We4vdHKWNLM/dnQ/+kNM4cYWvT1mfaL7BVe8SxJeZMIEZgA
lXfSIsw0zPLYQ0HbvtgD9QOTQ4lrcxBkZwTCMD9OiZ24O3Tx3SBLKtp/rhljttz4vdzgwAzJuGsy
L2ULLie3WwwHYObzuvNzZ/hCBaKpvdRC1QlPANadKwYX3E7oxY26c/D+fP4JcClD7ZkUz8GC8pBH
VoBLGLyudQWABXkbucV/E1jSRzMeQXlvtIUbsobPW0nrGNHZm3XmH+ZDLqPu/UTAJm3vL94nnlOL
iGA2LHem36rSdLqUkbRJZgYkRiG+0kc2uDpxP9eQUEgVlh1sx5RYCNh8CQf2g6slMPZqLW0GAcTa
PAgQWkEK32q1yYHda+g5pnp0wZ5HH1EbA+LRB030GIGOtd6rJidEffL6QnDqHFwI8FhVBTAu07wR
VlcSY/VzCq04PhZc2KoKuV3DUCYHCP6lA9L1Qz7nWtjDyuqIH7MlothdPQAacrOdd3MJyy1MDHRQ
2Ztjj7E4iVLaBOr1/yuKrodNntCWgdkNcRzJStXjqmdgso7GmiBptx//Sw/Gz0YmgxI2AN7EjycU
SLPOA4dJNqp8/DBC+Al28rZtiJhUQGetIRTijVTSdITwqHI2ranjJXHUtqplFM3RQfBn7XhMFswX
5rJJIGRtJEm+s/poqrOQVifwB4nZpI4+HHEVKaiiLw9foHQuuad0f3NuPQ0Rc/vgwuyGwoRYi67W
4+VgpYMv/wSlqR3RY1FG1rFtHEhpXoOdZsw2DIKFgPbfqbLH+98higlNnoULU4QnBkq0cJg18zNI
yilN7vaemSN7usqJHfRYtTEqI2WSetpgrIQvlSP27RhPvrS56hv5hWNWFT/zxFkKTf3wejHPIJ/G
7SIZlaQh/w63p1DyuQiRVD0x0egTnaZYaSaI43jHva0SLfaSf4eX8Ce69sq2TsRrS07q3WF7nmKd
nQJvFrI+Cbc+/LdrMuUo0fizkbTaSrY3DaphIyBwL8EKGuetrrrhlZ/sbqJNitb3+lQ29gdP2/Vo
X0Sec+u4idkRJtUlIqr6XHpwDvcGq/4+xLaJY7QLB9UNfp9G5o0ziDsXsiJkDzRmNN6BWQdvhdzL
NJIySiwyMuVgNMQsCrjsSrKiap2yj73bA7czVSO51IqCywc65IWt7PJi0Y3HHTlNpmDGdrGv9J+f
7DI+qWhH2w53mEFXS9thwQa6AUu/mKddhfMekdJ56mXofpfd7ivIfhtb5IZnoD5kTz8qoJ6L9aBC
bODqpTthU5hgYi1Jo/En/U7aly4tJXavTjCjTQCDBTswsowOdUkjUbuksmGNtLFVopyrsfXNq7+c
KvbOx23tfLiq16FDWwjd5h/MOcoqHiZ5XH2RVURwxHfvU+9nnB6icNOx5R6IllWYI+G5g+GySh2T
54ScP7TePTgf407N20nuXBoTTK/HUnnkFkvRjFhSlz1EfDN6+z6BIYJa1gjPqrpPlQU7hMDgCIjU
F0OKELVd3o2IZhoy/IluLmlMIl/Oh5RjICsAru04MqPjKrLme6dFXjn8xMYkvdiaa6WOiAL+n4++
EdLlHaB1ruQkMwOs0fi9SoUdPh1XHOmuzkYa/Nb1SQCN0vzOngcriFIGJLNJr4nXlFaNHYKBBnhx
cB3kq0PZEzSMt2F568ZvHHzW4O781ZRrNrLXZVEL/ScuWDwqQbp2fGPq1KPFrOU4P5tt1J3LCJyx
fOLWcBP4qD9c7OqNhjB7OlmVRDkgiJok1fhaiqUSDp2+k+TJce0gonR8PxVHvFsdnSE2GncAJbzi
3x1J8OyVv+/pam3jIo+0r/7vQ6lpuN//00dOM5tsWXFgy9W8KgWdaEv4R7H6CWoqSycBMQ9fYHVr
kZvqHwBUkImVXOYcdwwi0QGM1s+5v48pT3lgF2kZ+95grtjRJx72HOzsyV37r/U/0ZXZYUyeA0Of
u1b0rTb06wXmcH029fjBy12ZJo1EqPILHqCW4X1+ZyiqIv0ky/YWg5FH8nba5//m3N0dNV8Ngo4V
BtO7ugimARAVEOHX5rWqw7xKGkV5P7naueE+eiegsfUm8eTc68tF3FkjcQ0K2zraXoUN5xdD6ewJ
ai3h3X4/zEyCP95CJS/kpfWBeA4nT95bVq5SbV84AdiPSPYT1JH2cTioqFnDviX0Tj3tYFxNhNtm
x0ae8LybFV1Lhfxijf2W7PIuJspszWBhJb+ZBr56ZB+72zQnRPV8AflJreiQZeZNIqj+J/oJkL/Y
1ql+8DqSEnbVw1Pim27zGjd5P/dns4DXuGeREMrl0/mWTQodWzxbP8r09r+yNUXdGIdt+QUGN/Ml
79vhKXMFq/eu3Ei9BkU/4DDHAYnQsqZehoyaZ6kR6dff31LCuOK70CNjYeodkGhMN8mBJli56TYv
l7O4Wze0fHjeMBbsq+66dMuR8WPEvNTR3f5NFwmpgy/c474WnaWLNHTsVm2O582eEjZxd00ZJJKu
UGBGfIuwPeIxPWKXOYS8W2HZ5JKTWiJSu5HXAV9CHAVGMoTG3C2URCpPakSWjaUJkp37NdjbOHat
heFrhKA1MozG4McXSwhcoub13lzNshKRRicDDHoEXzQq+9DG3aTHUgWww/NTRAQGWywb+HybiJeg
JmmXDpwvnRykzFvpc4dMWnuTT3Ck5OKrYEDiGGIMcEnMKURFlINME2UTEOyszcS5mfUQNxZPuGGd
6KqyUIEcQdSuyWYX7NpYusC8rAL01ejylxZfGwx5HjtRFXJZOMtmFayiu7M5I4Kba1j6WK1cUURk
XlqMfLYDOauiDuxb1+1/hs/lXHXCzWo1Z+86UoCDhwP22LbMYIKIBot7fxZWup7eYYvYCMBPl2TN
TWxghR0Mhks1xKKHA0L1+f1d2T6HelZLi5MOxvWDMlZwI9k0aE08H3J2HLCZkDaMKql7oGsuTv1Y
B5YF/nag6iS6noPqYZhqb2eiffF8p8uPjorM3a7xeG8GjKTAV2aDqjXVoA/3m2bSUb1FDYUf9RwA
xjmtlHi75q4yTkGKNPf4d9UG7tXVRWcJ95zbYIoZ1Pd5yLRYR8sgZpivXA6EGRuXy81Bt8maCT+p
hX2SBoeNnH78ckKcrJ4V67aAwfqnEi3gdhzs8M8gzknIAJAVUdWrNd12pVdaGZgPAI5VRcUiGh5b
5/kKXh44bDJBYtcgaeTweURQzy14Nw37BI4uHlLa3gFJaijWBOr3D+7mpSX74ilRskev73Y1ZYUG
VbfAD08YAjWun/q0INlAeq/YhUkZJQQCd+dWdsrBVlu/Pybvbyol341pgylAWvkobn/hHr7YwT9x
epPG26qYEB/bgGXYAY5KJc8+SF6Iv8n31W63gAEwhgoWDgYEy6+bnFciMNxmpW+Rb25HAynYHAV1
grsrDlo4su+ZrF+pbZLWQqypBwkXaBKskbS4B5b7rnvjpT9ddV2SN5JddtGps+cYU91BhKYRuBNZ
0MEqEbe9hP0D7XoSYoZNFl/abDuXHzVovJpR0zFnjBgfockKPILVjFfwWqOmk1t7dhGoTvJi782i
8gRgsO6upzF1+IXB1deDBkVMpFynSEnJtLPmPAZ3ujirJk9rMVIfOJH+/IzjChYhNxqLZBfMPVJ0
CkUbJdBvSLQoB8LD+10F0Zpat5Uh0KR1oIx3vzjT+FZ8iQyR1RYM6DsS1cJcKw/dfIqOzWZBZ76q
tZ9HPKfpomATkJgEgkjUrhCMrEkeudYvtIxjHnmoF9CxfG2rt6qvlKanv8P+x2LHoH90ECvnzg==
`protect end_protected
