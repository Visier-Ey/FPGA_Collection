-- (C) 2001-2025 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 24.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
Vp0kCP0fAv4N2f+ia8jwAr6ZIgsHGLlkRiu1mR26MwNX8TRXASz3xsyfxKOIqqul
/nfqCz+Z2ZFnVaGbDp/grq1CVB+CSrcD2ZB3orprv7JxB55hXXM37O2soiQNVodn
20rK9pgrCOtAcHb8WDtlTPLC0OSILqdXNOQE6hnu/cc=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 5561)

`protect DATA_BLOCK
ME0lCoWDeF1Rnl9w+B2PLvNAWb8jjOfr0N+KmQ3ElV67BSxcZWdGvmft+x131ADW
GkvqiX9ZOPMcYBvqlD577+2hNlQrVQ5FpR2fkZODjBrakNKpIkyqUHDJEZYQc0Ys
O7LCkRx3fJNhim1v3KdeaACckWCtkXDnZ7e08iloIxChDN5a3JxkBvCzplz0mhrw
hKf4jMCQqCKfC1d7hmSqI40IatqWZu1A0sbyS4TcgVGunRUoJn6mtRXmtjJdTcCj
k5IjrebjxBAoW1YpkctxwBgaPHK0avH2KMRgM9i0eK9khm4k6Am668RTJVnzJCgs
eIdjoEItwgrYGznJe6LuYjPt3t22yQMhawONtMeyTUbjuOkGKxPeSarlCLm03vZn
yJSenCsg5MroMJylqb9oPymLTLNeYRuznpTP9qF0dwwdWhoiXrpSVngBl4d+Iakv
/duj9GCgoGO0qA7QeUE1X56cIo/N0v53h8F3ad3e5WZ+i38d20cKcLixjAbvjQtn
t78kKaTNX9LN7wMK67Vfh7c7I+zlMC9X4br1cyMplX4LR2TcS+82olj2KexNXUz+
xEOdN8eI2sWZ4Ji0yrZ/TXObDZmo9vGOsUbxeokUN5+RNpfRxNKP5Gxc7AIq1y3K
Zb7z9ir5f3/ielQm1yBOm4lPI1M7UhAgIjmKG3XG2YbCu3moPz+ZWGVGy0xdqfxO
BvLaVd4BPdeF9AXl19y44cNusTQCWFwhJBJE5i97KKpC43hC8N3jOHcBlHIzb7kT
dgTadQWVoOOFr5jYIuNS4SRgf0j/bXOQvXldfe49XNxl+urK50Jfpfia8weESVWH
SKE5vjVnL+2zG0NeoVaVyJbhd5tsnZINGJxsfeGRlZrYUKTbOOe46909BZGeaW7+
5N8IJoNi0hY9dG7V7wGuvJv6ezAMZe2GOYCGKruG/KnHVbvd+CLLJEr+pmZHh7oy
6Vs8wmhgWuKkkMTDarhFVwO2U5DofIno/Rv0KvTd2XmQIYnWC4JKzi27KZNXlJMD
6SIu8ut0utdhbi/v5ikcZfDByAeWcJTMsb/aB+4LbD8v/tDSVIpAbRhJZTpTdqYZ
Psam9odWSZ/UUgyH+FOyqoqvRb6c5ekFQe/+l3W+N3o7UM38ba28+7a5eVy4qzmW
Y8O8U2tKAAwT0SeXWkE3N3O863eSddb2YapmBposdZ86GMFRlUMc/QSc55T/GsBj
05lEhnLpdo0FpcemPbECMYAm1MWL0KtdlVLwUEfu2QW9Wlc/bTFvJXFW4XFMs7Qn
PKYqpnvAtQdUM8L85iw7y7rh1bBT+SuLj66LryqRDUo0P7ox/0eypQQHw5HkMYuE
VIoZD/mQKSZrgJXPUu4VIx77b/AI0hj4Yt9rYkAuOxnHmGqCVH9BnRCmO7jGm8q0
rTVgmf7y08Ywr+gldwKA/SK8oZ4o10QiryVpKkWBu6TJvDu8UkgkIODRMR4cVlF5
lKgOlafQZ8Q11mE4xRtX5LWc5QSEDdBxpbnEsyQoNzt/sX1Kdg6nZ3Z6/+rDtk1v
o95BC3blwmeZqxbCT4PA9mrxU4NmZe2r2ntGgcBByAtFTHyzoynN9ABJoI2rmn+3
RcxQ0cl8R1Mqjt6wXTzRXl9KfG29XT3Gmg8TO7ZST8qNnQqbAHrLwXwbWsm4twsW
dP9kcLBN/nxL/F76TiGvExBN7JIH4p5qjD+xN1/tIWR7N+BbLbBi4ipPHnS2Qzi2
J/AEomEsGW6wbdLQh1rh6EZ7OtJgRAsaQnhvsBkeeh1frV7zFP5AnvtT1ZKgbAb4
0lmxf4UJGRK6KBq8EQ4kAeWjOQJwqHaHOjihUFEeNylGSb3kXWBOLhl8W14WdpsJ
2OvdONbPiyxRVvSKfL4GyhOpZbf8CEFSDHsIbN3bABUA4EiRqn/r1MoCgws2glWr
NjsuycQfz8TgDmW+R/Vkgaxwkc4ShEWW+qmCHkJW1ILP68kBisdSIXTncxuBqajD
Otq7MCuXpzRzt1jHtLAkDHqQOGvWaZNvkBdmsgYOeUKnyfz9nuZ4Wa39D6Nrwzrk
5xFGh++4jjEePzuw0PkV45XXcvLzJQeo0M6CpCs45uPsYma3iw8J9lsiwkK7a8BO
J/vuesURXlFvSEXlV5O6R2kUNDzpfC0P+peaV577i3JOL815XQDzckCMb++qLPzR
5jWUd4eF27IuNabaN+7AF8kbABUMINo4ilWcTBt6g8YHburAfn9x4pG3RseYfR7m
hMVl5mgt2AqomIBlYO3lDA90exX30EtGoJIvVUduRc0UJH1xlVgi2qJg9Z2y6YTm
wSND3ydHLldxXBoZ6Gmi5Du+5wtjTWlpHsMCNcORS1R/zt1g9hO45zLn0ViFzQb7
mP79nbuzwzBlRqvv9DLDQkIFXS5dqBxBpbpbYBTP49zCHvZqxRiVOYNXZrjl1JJE
EKGqjs82nWtBGYvG1/bsSM6u2242giV800qvKaKvu7TdTPJHYtrrMOv+Ghj9Rzcp
w4lwh/o/8LDwSKhrBDXgU231KFCpSNTXwXcTbG9RPmSA0B+S6TNX53ofC7bwSPcl
UzPZx5vTShL7Y0rYOhZFvCMnFMzQKzS7biHTtNuj8pikjljk82dEzHFDoSPHmTXd
NnEfGYhBckjnZFK99QN+f8TPryHg8N5427vM7fGD+ZVNoCy00dBPUZ2nJqkttRg5
wSb2xhL3pPwjzFf3yG4Dc+w/FNjjjx8lCjoOrNb9VxEHlQb4w6ZvwgGCz1X8MDsJ
cFXu9UCUaWJ65FhA+pJxHXqTvTDSfqfAc5EqKjF0stpE9kPGbFjHu/Auf9VEXfYI
PCEx5WPOb0lQNo+D3DGqy2Zt7hq+xQQFW39WcoqYRtgFKAtaGEOecTu3gR3MfTlT
GV9QO/9ZYik2UBnI7MnlA453ihpALLQ1YaWIi8rrDLzrTS+qc3ZdPVyyY3viSt3D
ZjuFuhvwvF3ejKol3fizlXLO48T6YvDKD6oVnHSvd20st7g9XZRD9e1rsz5IRvyz
hKkw1ZDEftfHV2O9U7wizDXYabq55+sqAfL+tCpiHeMGaKHsK5osc12c1DFIVJRH
skHr5HgJ+W3GMQ69T7XDcE+C++8x3gyFba6DsnYSkh0Ho7+z+Ln7osHseThWFJPb
y3x/jgZl53PUKKf1o9ux5EGyK3H34izOo+pp5pAPuCYgiW3zROeZV1kYabo1hCWx
tC4sllf/dy4B5+X79S1UhU5zc+/lhDTjedGIc91g9s5KmnVk314j4mpBMRxLxAJk
0mYziXZRMVxL9OAdxxxCI1k0pAIEEgnOEJMx7giCMD+bvStyYarTAQFRBwhLnvgE
5YNI8rs1Hi23iPYEmQMpoKJOhAsH0T51UM3xgbyHFcbZxECv7GKWow2+dBB3pwmb
r+RRvWVwh1RFgh9g1rDYZwvS0sWNERbckU/oPGHMJUZ6M0X5RaYp61uDd5c0aRoR
pHmqJHEGejyqWRbmqJRlZRvfuJ33tnX0FGKxmlttWdJlZ/htqY8dhhKTQi/rOvco
jVyBnY/a8wjhHUNLyCE6vqU6iz7CDYm/68U72wBxG/8iyMPeDIZ0tAdK5uHDScX9
+zwPxEw+sk3/8HcVnzIm8aNe2cxwI3l4k4uTDCeKrAODJlBPO1Tm6O3GGWw/CHcC
/+zx+UBm345YkEXwTL/0PNl3U7oXgmmJHBWjL10MEkTJhvEzAl2RCuC+7UhNf2w1
9srZDP5OkWnnvdY8iBDUPJL+9Mcps2ExHDKv8xy5Q8VD3tnJ8WG7tqeJakpwzKHE
l4qbjh3uSMLUDUqz5dK1smr0fw+kYsfO2X1BkkkU20hPwRtGUrIAV9EpM++Z7K4k
a/hmOqgZxXWwzJB0nWGlPxt1cGACO/w1aIQa9NVcCMzni1x4IT1UwXX+pGKlH/kE
vE2CAOR1mGug2UGuALkm9xLgS6w4C4wTZjytwOu/ZodVNxQpEFoxGXqzEkm3+JUu
HO4KKxGWyCGqeYU7aoRmInrpJFnbmheeEHjrQUw65cgcm3gU4wjg6j5VZjgGq6Eu
DPcAgkQtjftvBOGlCp+tphDFjQeRKBUqm1eASBuaMxA/EjQAyq89ohgxTyXr7Dfe
w/s5/nCG829uxnEwu3yGdyatQr92pVqdWHL5RDwWarcMcFQ4K7C2gJAjAzJ2zrek
jn/1faN42YJlFHs+sdnIwmgUiPZTd2p8vGl/rjoJI8Put/yroDB2+RHJp2wclBVh
bA1BjLcaxqm4sNcDBMGiYZfEcRN1SKs3s4xTNaDflTlqrglz/he810J15js2MGAd
UCsZAjBv5or0X1KG4Px7Rm4purGAbQytgS5ju3c1x1zjfUir3QtBhMEfGKBxh0iO
qgasp5FSvzSjximkUrFVqRBTYy4NE/xcK1qHuPJdsAhBx0qARFZo57c4As35L0wP
SUu0pIK1cv0uaVU6AEvE8kWrOJetNpOKRFl4xv21Q4mO1H6KD+9gDzPvqbfMk0ws
UVys7HhoWnXD73iU9gN81rcnc80i8CxhetvJXdSvGDoLkB+8bs+/XGEdXvvWmxgx
LWE8zelde/WVmc9PTZJgOiHelrQK2BOuC162XFUW2mlszHIOYlfadHYgFpOv9I2h
pMrX8iWnY9LHP4Tk+vsXIjHWKY9jkMDtnUvUtkx1axSGkIlkJkUd8KRNizuWjaOg
g+6g+S9rsQe2GybRoi/0Geay8FBvoVIRVZAAYaRtBvX2XHnU9Dcc1U2nb0eFGktg
kvj9yZerKstvWrWJdvONC9VgieeLxog6ZoL9NBn3ySCJXkNxq9c89dV+NEbvOgWn
rDi26cEBAAy6wGzNkWC4WXCuBNdB3tnJF/KRszYNwZKpPENRX7ONU6CsoRhPQXck
diKo0uk+O9hVsR6DguGKos6VdEHvqkdgEkJPTffoQQ2hToI/PNcCtH6TZ4OjZxa+
svHbR1ZnAurcCxwzB4lkzQM64iygNtZt/NEeGFY5OxoqjQf14kjTpjhDcOQIJ48X
v/cBar5c54rQLcKUYnw2lkW2WyibgR2TReeAx+BL4FRITkIAJO4MIBHrnAnCgCET
Eqi/t7eKxRjU//Md+F+H6PdPBq+x5HjlldKr77km8AjsfYuWT+qtDPsP+xnxnM6v
MtRE1IMMqOQgXsIjgc71lYXpdLEsyA9+3GaCIcKcppkgV53YYPoFIgQ+DMyNa1Hb
Ck8CaJQ+ym2PHyxLsF9ghWf6o4eloSD22ECjl78ygZdtG7RHxTM2TYwqczIjjH6S
BBFM2Q0ez5wB/wZ3ztYWsNvZKjuukOFwCVzSb0Wn3LrfUhHCh6CfEWf1TccuVSfX
9d82M8mUne3pUHOXgYUUy5LaDHdw9iPWwIl27qLvkNPbHqBe4BAITO1ct995VXbN
+cQycocJraHVLmTJuBAU+kpUILih+ujmLxKF8hIycr4QV1mwOmpIRsSYHPwZNhma
JGIhlOifu00JiBYmHdTnPX+JsInz5lODxXXvOLu/536UZDJ7VzugHlV/E3JshDpj
Jy8xphA+1RetIByIqcaq/OA0RFuc+tHGuS0p4E28XJ6QOPzN4ZHvWpusleqzQPxd
Jgp+QVQVwuvBkgsOr0m+96aH/kzhpc76FEivUmYKdFRRzz04L2EuSWDJ69wDCkyN
iVNjty5sLxSqChE/GNAdIdgWu5HuSmE3N8sNNXdlS59UwLttzzyqN8TcK6uWRMzs
DIu1OfxjCklq3lxmxVE8PIuChBMs4uo3fWDWs9YU/6HFYF7OZuE1nAAorcQefgWr
sFjPOc2CUdnClE5lO9EDBt/IQkpmccgFIbAhmZMVcNVcpMeKkZ3XjEi2zw7SoqsQ
Xglra9Zh5n50YNtypkBiHR3L97iyOkhBt99CjWCT+r/wQA3SOaQnqpi6S2Euq/Fy
0gB7xpOv/jaV5Tyq8xHFfemDebQfE1EbP7ztDwo0lz/3U8yaX9dE9ontZJyCVqch
Ix+ezoV91v/hdJP5f3sDMhDktStOAZqqTmS8H4RTrMWD/ubDPmQid5Lif9y4P95V
8rlJ8F0pQzuxe4uI/8PaghBQ1ObyA2I3VyV6ShH9sEH0Qp9zjYT/UTMTmSRTHRmI
BEkXkapmmP5c6LuCW42aoEKqlb+8T4wJ/XJI2WxM06GB/JNkctEqdmsEkxYnXkSq
KSSWax/OG3UJVVD/Cunqa/xQRx87HgFgzslRH931TFIypb3eXYm7lVQU7/P+/Iul
ISbm2Q91Qo3bEBWl6ljRJwGWKpJlKEUDIP8KElGMwz/KegKYHYPNN6jFu0Q5wWbE
9ui8abcxLq4gonpmNWvdH+gb+RI+SZt1y9MzaruZ+51RLWLbYSgI9SA67+uvDAm1
OS/jO+9NLFGjg/x7yT+TRK72vC/wmweiIfJXOkOAV4p2a9eshwwH46AqWBxkkxrj
Fg1zKY1zT/irUXPV6p3iu82wm0MGbLET5EOx58dVmH5r4yUHEdrveNBr1c7eDOia
snnT+P1W7UkoMI3pSYoSNjMc6WkfUWLaZEZ6vnBVwFrAgbrZ8EbBskY6zoipTWd8
+o41FLX2WbdfatIMfZpErOywkdFRpA6JVrxOphYdXZJ5LAak5WkXNStjsbTb+4lc
Msb7Hk++I0I9kdLMK4VO/HokZXvyNQ3A19BbZQkJ0f7FVLGXhSLcxruDZvzpcjUj
8PAyQ9zwftUS3hXn7GpC+h7HYZGEzNRuS2ZcgXjaThczSxon1VnJzWVxkt1toolp
paTq7NcGMEEd46MJN5WkwhzWY+g+Mz9pWLXoeSeMg0qar/fHmEnFTw/WfYngFU5P
Dr6350LYgJGN68bmG2LHOldwbgk+PwvmW32UJ/RpKY69ghZ+8bPBGZdnzjUf0zYy
w2ZP1gx1ojE52IMcvVyF8FUTgdgmdgtT/9SNa/BGDT1pKjQakJ7PBWJndjtU3vRJ
8nqqohwO2xbRU2grJ7YME7ORqOSr01sABXqZH+02CiLycGShvR73z1dpVpd1sWSW
4DwHUv0oD/T8qafURvTxzWehIq5TpA4rK2KqJn7KtRMRF6TFTw6rOsNP1KLs54xA
y9wp7sFH/nkMUombvEPYKhDJLQQzsTMQdTBzj/DEZmnhDWfxM9gTyPm8INp3TNi2
iWvmQqbG6BoaAityCphN7llbTYsxt6ixqzWFC6fKB/25dJDNeBRojnhOnaaGr//j
W3aJxwcndvyIt+iXj38NlijCbpks+2pq4cEm6CDfI0upo0SkUa7/8fQfFiAWdzH8
u4SHzHOHmYxX8PHSsCqbGj7+wLGKBzlw+oLdJLP4AwNMF2SwaFxtCJVDwRoigAfR
ZFmdqjhf83dYyD/9rophoiEpTEzVsAC59afw6oHnbJ6gV1DopFZqYG2BSCl81OD8
AZcOYa213eCSJef7PM+YFNsAeSI9B29+uOywX8MyfzMxvQN2n43QnFNPCnVwIJ/F
OsqzxNIaNsxV+M4AE0Mz+w==
`protect END_PROTECTED